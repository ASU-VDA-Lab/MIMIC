module fake_netlist_5_1571_n_13034 (n_924, n_1263, n_977, n_1378, n_2253, n_2417, n_611, n_2756, n_1126, n_1423, n_1729, n_2739, n_1166, n_2380, n_1751, n_469, n_1508, n_82, n_2771, n_785, n_549, n_2617, n_2200, n_532, n_1161, n_1859, n_2746, n_1677, n_1150, n_2327, n_226, n_1780, n_1488, n_667, n_790, n_1055, n_2386, n_1501, n_111, n_2395, n_880, n_544, n_1007, n_2369, n_155, n_552, n_1528, n_2683, n_1370, n_1292, n_2347, n_2520, n_1198, n_1360, n_2388, n_1099, n_2568, n_956, n_564, n_423, n_1738, n_2021, n_21, n_2134, n_2391, n_105, n_1021, n_1960, n_2185, n_4, n_551, n_2143, n_2059, n_1323, n_1466, n_688, n_1695, n_2487, n_1353, n_800, n_1347, n_2495, n_1535, n_1789, n_1666, n_2389, n_671, n_819, n_1451, n_1022, n_2302, n_915, n_1545, n_2374, n_864, n_173, n_859, n_951, n_1947, n_1264, n_2114, n_447, n_247, n_2001, n_1494, n_292, n_625, n_854, n_1462, n_1799, n_2069, n_2396, n_1580, n_674, n_417, n_1939, n_2486, n_1806, n_516, n_933, n_2244, n_2257, n_1152, n_497, n_1869, n_1607, n_1563, n_606, n_275, n_2011, n_2096, n_26, n_877, n_2105, n_2538, n_2024, n_2, n_2530, n_1696, n_2483, n_755, n_1118, n_6, n_1686, n_947, n_1285, n_373, n_307, n_1860, n_2543, n_1359, n_530, n_87, n_150, n_1107, n_1728, n_556, n_2031, n_2076, n_2482, n_2677, n_1230, n_668, n_375, n_301, n_1896, n_2165, n_2147, n_929, n_2770, n_1124, n_1818, n_2127, n_902, n_1576, n_191, n_1104, n_1294, n_659, n_51, n_1705, n_2584, n_1257, n_2639, n_171, n_1182, n_579, n_1698, n_1261, n_2329, n_938, n_1098, n_2142, n_320, n_1154, n_2189, n_1242, n_1135, n_24, n_406, n_519, n_2323, n_2203, n_2597, n_1016, n_1243, n_546, n_101, n_2047, n_1280, n_1845, n_281, n_240, n_2052, n_2193, n_2058, n_2458, n_2478, n_291, n_231, n_257, n_2761, n_731, n_371, n_1483, n_1314, n_1512, n_709, n_1490, n_317, n_1236, n_1633, n_2537, n_569, n_2669, n_2144, n_1778, n_227, n_2306, n_920, n_2515, n_1289, n_1517, n_2091, n_2466, n_2635, n_2652, n_94, n_335, n_2715, n_2085, n_1669, n_2566, n_370, n_976, n_1949, n_343, n_1449, n_308, n_1946, n_1566, n_2032, n_297, n_2587, n_156, n_2149, n_1078, n_2782, n_1670, n_2672, n_775, n_219, n_157, n_2651, n_600, n_1484, n_2071, n_2561, n_1374, n_1328, n_2643, n_223, n_2141, n_1948, n_1984, n_2099, n_2408, n_264, n_1877, n_1831, n_1598, n_1723, n_955, n_1850, n_163, n_339, n_1146, n_882, n_183, n_243, n_2384, n_1036, n_1097, n_1749, n_347, n_59, n_550, n_696, n_897, n_215, n_350, n_196, n_798, n_646, n_1428, n_2663, n_436, n_1394, n_2659, n_1414, n_1216, n_290, n_580, n_2693, n_1040, n_2202, n_2648, n_1872, n_1852, n_2159, n_578, n_926, n_2180, n_2249, n_344, n_2353, n_1218, n_1931, n_2439, n_2632, n_2276, n_422, n_475, n_777, n_1070, n_1547, n_2089, n_1030, n_72, n_2470, n_1755, n_415, n_1071, n_485, n_1165, n_1267, n_1561, n_496, n_1801, n_1391, n_958, n_1034, n_670, n_1513, n_1600, n_48, n_521, n_663, n_845, n_2235, n_1862, n_673, n_837, n_1239, n_528, n_2300, n_2791, n_1796, n_2551, n_680, n_1473, n_1587, n_2682, n_395, n_164, n_553, n_901, n_2432, n_813, n_1521, n_1284, n_1590, n_214, n_2174, n_2714, n_1748, n_1672, n_2506, n_675, n_2699, n_888, n_1880, n_2769, n_2337, n_1167, n_1626, n_637, n_2615, n_1384, n_1556, n_184, n_446, n_1863, n_1064, n_144, n_858, n_2079, n_2238, n_114, n_96, n_923, n_2118, n_691, n_1151, n_881, n_1405, n_2407, n_1706, n_468, n_213, n_129, n_342, n_2753, n_464, n_363, n_1582, n_197, n_1069, n_1784, n_1075, n_1836, n_1450, n_1322, n_2101, n_1471, n_1986, n_2072, n_2738, n_1750, n_1459, n_460, n_889, n_2358, n_973, n_1700, n_477, n_571, n_1585, n_461, n_2684, n_2712, n_1971, n_1599, n_2275, n_2713, n_2644, n_2700, n_1211, n_1197, n_1523, n_2730, n_1950, n_907, n_1447, n_2251, n_1377, n_2370, n_190, n_989, n_2544, n_1039, n_2214, n_34, n_2055, n_228, n_283, n_1403, n_2248, n_2356, n_488, n_736, n_892, n_2688, n_1000, n_1202, n_2750, n_2620, n_1278, n_2622, n_2062, n_2668, n_1002, n_1463, n_1581, n_2100, n_49, n_310, n_54, n_593, n_2258, n_12, n_748, n_586, n_1058, n_1667, n_838, n_2784, n_332, n_1053, n_1224, n_349, n_2557, n_1926, n_2706, n_1248, n_230, n_1331, n_953, n_279, n_1014, n_1241, n_70, n_2150, n_2241, n_2757, n_2152, n_289, n_963, n_1052, n_954, n_627, n_1385, n_440, n_793, n_478, n_2590, n_2776, n_2140, n_2385, n_1819, n_2330, n_2139, n_476, n_1527, n_2042, n_534, n_1882, n_884, n_345, n_944, n_1754, n_1623, n_2175, n_2720, n_2324, n_1854, n_91, n_2606, n_2674, n_1565, n_1809, n_1856, n_182, n_143, n_647, n_237, n_407, n_1072, n_2218, n_2267, n_832, n_857, n_2305, n_2636, n_2450, n_207, n_561, n_1319, n_2379, n_2616, n_2154, n_1825, n_1951, n_1883, n_1906, n_2759, n_1712, n_1387, n_2262, n_2462, n_2514, n_1532, n_2322, n_2271, n_2625, n_18, n_1027, n_971, n_1156, n_117, n_326, n_794, n_404, n_2798, n_2331, n_2293, n_686, n_847, n_1393, n_2319, n_596, n_1775, n_2028, n_1368, n_2762, n_558, n_2808, n_702, n_1276, n_2548, n_822, n_1412, n_2676, n_1709, n_2679, n_2108, n_728, n_266, n_1162, n_272, n_1538, n_1838, n_1199, n_1847, n_1779, n_2767, n_2777, n_2603, n_352, n_1884, n_2434, n_2660, n_53, n_1038, n_520, n_1369, n_409, n_2611, n_1841, n_1660, n_887, n_1905, n_2553, n_154, n_2581, n_71, n_2195, n_2529, n_300, n_2698, n_809, n_870, n_931, n_599, n_1711, n_1662, n_1891, n_1481, n_2626, n_1942, n_434, n_1978, n_1544, n_2510, n_868, n_2454, n_639, n_2804, n_914, n_2120, n_411, n_414, n_2546, n_1629, n_1293, n_2801, n_965, n_1876, n_1743, n_935, n_121, n_1175, n_817, n_2763, n_360, n_36, n_1479, n_1810, n_2350, n_2813, n_64, n_1888, n_2009, n_759, n_2222, n_1892, n_28, n_806, n_1997, n_2667, n_1766, n_1477, n_324, n_1635, n_1963, n_2226, n_1571, n_187, n_1189, n_2690, n_103, n_97, n_11, n_2215, n_7, n_1259, n_1690, n_706, n_746, n_1649, n_747, n_2064, n_52, n_784, n_110, n_2449, n_1733, n_1244, n_2413, n_431, n_1194, n_1925, n_2297, n_1815, n_2621, n_615, n_851, n_1759, n_843, n_1788, n_2177, n_2491, n_523, n_913, n_1537, n_705, n_865, n_61, n_2227, n_678, n_2671, n_697, n_127, n_1222, n_75, n_1679, n_2190, n_776, n_1798, n_2022, n_1790, n_2518, n_1415, n_367, n_2629, n_2592, n_452, n_525, n_1260, n_1746, n_1647, n_2181, n_2479, n_1829, n_1464, n_649, n_547, n_2563, n_43, n_1444, n_1191, n_2387, n_1674, n_1833, n_116, n_1830, n_2517, n_2073, n_1710, n_284, n_1128, n_139, n_1734, n_744, n_590, n_629, n_2631, n_1308, n_2178, n_1767, n_2336, n_254, n_1680, n_1233, n_2607, n_23, n_1615, n_1529, n_2005, n_526, n_1916, n_293, n_372, n_677, n_244, n_47, n_1333, n_2469, n_1121, n_2723, n_314, n_368, n_433, n_604, n_2007, n_8, n_949, n_2539, n_100, n_2582, n_1443, n_1008, n_946, n_1539, n_2736, n_1001, n_1503, n_2054, n_498, n_1468, n_1559, n_1765, n_1866, n_689, n_738, n_1624, n_640, n_1510, n_252, n_624, n_1380, n_1744, n_2623, n_1617, n_295, n_133, n_1010, n_1994, n_1231, n_739, n_1279, n_1406, n_2718, n_1195, n_1837, n_1839, n_610, n_2577, n_1760, n_936, n_568, n_1500, n_39, n_1090, n_2796, n_757, n_2342, n_633, n_439, n_106, n_1832, n_259, n_448, n_1851, n_758, n_999, n_2046, n_2741, n_1933, n_2290, n_93, n_1656, n_1158, n_2045, n_1509, n_1874, n_2040, n_563, n_2060, n_2613, n_1987, n_2805, n_1145, n_878, n_524, n_204, n_394, n_1678, n_1049, n_1153, n_2145, n_741, n_1639, n_1306, n_1068, n_1871, n_2580, n_2545, n_2787, n_1964, n_122, n_331, n_10, n_906, n_1163, n_2039, n_1207, n_919, n_908, n_2412, n_2406, n_90, n_724, n_1781, n_2084, n_2035, n_658, n_2061, n_2378, n_2509, n_1740, n_2398, n_1362, n_1586, n_456, n_959, n_2459, n_535, n_152, n_940, n_1445, n_9, n_1492, n_2155, n_2516, n_1923, n_1773, n_592, n_1169, n_45, n_1596, n_1692, n_2666, n_1017, n_2481, n_2171, n_123, n_978, n_2768, n_2116, n_2314, n_1434, n_1054, n_2507, n_1474, n_1665, n_1269, n_2420, n_1095, n_1828, n_1614, n_267, n_514, n_457, n_1079, n_1045, n_1208, n_2093, n_2038, n_2320, n_2339, n_2473, n_2137, n_603, n_1431, n_2583, n_484, n_1593, n_1033, n_442, n_2299, n_131, n_2540, n_636, n_660, n_2087, n_1640, n_2162, n_1732, n_1009, n_1148, n_2051, n_109, n_742, n_750, n_2029, n_995, n_454, n_2168, n_2790, n_1609, n_374, n_1989, n_185, n_2359, n_396, n_1887, n_2523, n_1383, n_1073, n_255, n_2346, n_2457, n_662, n_459, n_2312, n_218, n_962, n_1215, n_1171, n_1578, n_723, n_1920, n_1065, n_1592, n_2536, n_1336, n_1721, n_1959, n_1758, n_2338, n_2737, n_1574, n_2399, n_2812, n_473, n_2048, n_2355, n_2133, n_1921, n_2721, n_1309, n_1878, n_1426, n_1043, n_2585, n_355, n_486, n_1800, n_1548, n_2725, n_614, n_337, n_1421, n_88, n_2571, n_1286, n_1177, n_1355, n_168, n_974, n_2565, n_727, n_1159, n_957, n_773, n_208, n_142, n_2124, n_743, n_2081, n_299, n_303, n_296, n_613, n_1119, n_2156, n_1240, n_2261, n_1820, n_2729, n_2418, n_65, n_829, n_2519, n_2724, n_1612, n_2179, n_1416, n_2077, n_1724, n_2111, n_2521, n_361, n_700, n_1237, n_573, n_69, n_1420, n_1132, n_388, n_1366, n_1300, n_2595, n_1127, n_2277, n_761, n_2477, n_1785, n_1568, n_1006, n_2110, n_329, n_274, n_1270, n_1664, n_1486, n_582, n_1332, n_2231, n_1390, n_2017, n_73, n_2474, n_2604, n_19, n_2090, n_1870, n_309, n_30, n_512, n_2367, n_1591, n_2033, n_84, n_130, n_322, n_1682, n_1980, n_2390, n_2628, n_1249, n_652, n_1111, n_1365, n_1927, n_25, n_2132, n_1349, n_1093, n_288, n_2400, n_1031, n_263, n_609, n_1041, n_1265, n_1909, n_44, n_224, n_2681, n_1562, n_383, n_834, n_112, n_765, n_2255, n_2424, n_2272, n_893, n_1015, n_1140, n_891, n_1651, n_1965, n_239, n_630, n_1902, n_2151, n_1941, n_55, n_2106, n_2775, n_2716, n_1913, n_504, n_1823, n_511, n_874, n_2464, n_358, n_1101, n_77, n_102, n_1106, n_1456, n_2230, n_2015, n_2365, n_1875, n_1982, n_1304, n_2803, n_1324, n_987, n_1846, n_261, n_174, n_2066, n_1885, n_1455, n_767, n_993, n_1903, n_2490, n_1407, n_2452, n_1551, n_545, n_441, n_860, n_450, n_1805, n_2176, n_2204, n_1816, n_429, n_948, n_1217, n_2220, n_2455, n_628, n_365, n_1849, n_2410, n_729, n_1131, n_1084, n_1961, n_970, n_1935, n_911, n_1430, n_83, n_2645, n_2467, n_513, n_2727, n_1094, n_1354, n_560, n_1534, n_340, n_2288, n_1351, n_2240, n_2696, n_1044, n_1205, n_2436, n_346, n_1209, n_1552, n_2508, n_495, n_602, n_574, n_2593, n_1435, n_879, n_16, n_2416, n_58, n_2405, n_623, n_2088, n_405, n_824, n_359, n_1645, n_2461, n_490, n_1327, n_2243, n_996, n_921, n_1684, n_233, n_2658, n_1717, n_572, n_366, n_815, n_1795, n_2128, n_2578, n_128, n_1821, n_120, n_327, n_135, n_1381, n_2555, n_2662, n_2740, n_1611, n_1037, n_2368, n_2656, n_1080, n_2301, n_1274, n_2554, n_1316, n_1708, n_2419, n_426, n_1438, n_1082, n_1840, n_589, n_716, n_1630, n_2122, n_2512, n_562, n_1436, n_62, n_1691, n_952, n_2786, n_2534, n_2092, n_1229, n_391, n_701, n_1437, n_1023, n_2075, n_645, n_539, n_803, n_1092, n_2694, n_238, n_1776, n_2198, n_2610, n_2661, n_2572, n_2281, n_2131, n_2789, n_2216, n_531, n_1757, n_890, n_1897, n_764, n_1919, n_1056, n_1424, n_162, n_960, n_2308, n_1893, n_222, n_1290, n_1123, n_1467, n_1047, n_2053, n_2163, n_634, n_2328, n_199, n_1958, n_32, n_2254, n_1252, n_348, n_1382, n_1029, n_925, n_1206, n_424, n_2647, n_1311, n_2191, n_1519, n_256, n_950, n_2428, n_1553, n_2664, n_1811, n_2443, n_2624, n_380, n_419, n_1346, n_444, n_1299, n_2158, n_1808, n_1060, n_1141, n_316, n_2266, n_389, n_2465, n_2650, n_418, n_248, n_136, n_86, n_146, n_912, n_315, n_968, n_451, n_619, n_408, n_2440, n_1386, n_1699, n_376, n_967, n_1442, n_2541, n_74, n_1139, n_2731, n_515, n_2333, n_57, n_351, n_885, n_397, n_1432, n_1357, n_483, n_2125, n_683, n_1632, n_1057, n_1051, n_1085, n_1066, n_721, n_2402, n_1157, n_2403, n_841, n_1050, n_22, n_802, n_1954, n_2265, n_46, n_1608, n_983, n_1844, n_2760, n_2792, n_38, n_280, n_1305, n_873, n_1826, n_378, n_1112, n_2304, n_762, n_1283, n_1644, n_17, n_2334, n_2637, n_690, n_33, n_1974, n_2463, n_583, n_2086, n_2289, n_302, n_1343, n_2701, n_2783, n_2263, n_1203, n_1631, n_2472, n_821, n_1763, n_2341, n_1966, n_1768, n_321, n_2294, n_1179, n_621, n_753, n_2475, n_2733, n_455, n_1048, n_1719, n_1288, n_212, n_385, n_2785, n_2556, n_507, n_2269, n_2732, n_2309, n_2415, n_2646, n_1560, n_1605, n_2236, n_330, n_1228, n_2123, n_972, n_692, n_2037, n_2685, n_1953, n_1938, n_820, n_1200, n_2499, n_1911, n_2460, n_2589, n_1301, n_1363, n_1668, n_1185, n_991, n_828, n_1967, n_779, n_576, n_1143, n_1579, n_2233, n_1329, n_2743, n_2675, n_1312, n_1439, n_804, n_537, n_1688, n_945, n_492, n_153, n_1504, n_943, n_341, n_250, n_992, n_1932, n_2755, n_543, n_260, n_842, n_650, n_984, n_694, n_2082, n_286, n_1992, n_2429, n_1643, n_883, n_1983, n_470, n_325, n_449, n_1594, n_132, n_1214, n_1342, n_1400, n_900, n_2362, n_856, n_2609, n_1793, n_1976, n_2223, n_918, n_942, n_2169, n_1804, n_189, n_1147, n_1557, n_1977, n_2153, n_2468, n_1610, n_13, n_1077, n_1422, n_2364, n_2533, n_540, n_618, n_896, n_2310, n_2780, n_323, n_2287, n_195, n_356, n_2291, n_2596, n_894, n_1636, n_2056, n_1730, n_831, n_2280, n_2192, n_964, n_1373, n_1350, n_1511, n_1865, n_1470, n_1096, n_2094, n_2670, n_234, n_1575, n_1697, n_1735, n_833, n_2318, n_2393, n_2020, n_5, n_1646, n_2502, n_225, n_2504, n_1307, n_1881, n_988, n_2749, n_2043, n_1940, n_814, n_2707, n_2751, n_2793, n_192, n_1549, n_1934, n_2311, n_1201, n_1114, n_655, n_2025, n_1616, n_1446, n_2285, n_2758, n_669, n_472, n_1458, n_1176, n_1472, n_2298, n_2471, n_1807, n_387, n_1149, n_2618, n_398, n_1671, n_635, n_2559, n_763, n_1020, n_1062, n_211, n_2303, n_1824, n_1917, n_2295, n_1219, n_3, n_1204, n_2810, n_2325, n_178, n_2747, n_2446, n_1814, n_1035, n_287, n_555, n_783, n_1848, n_1928, n_2126, n_1188, n_2588, n_1722, n_661, n_2441, n_41, n_1802, n_2600, n_849, n_2795, n_15, n_336, n_584, n_681, n_1638, n_1786, n_50, n_430, n_2002, n_2282, n_510, n_2800, n_216, n_2371, n_311, n_830, n_2098, n_1296, n_2627, n_2352, n_1413, n_801, n_2207, n_2080, n_2377, n_2619, n_2340, n_2444, n_2068, n_241, n_875, n_357, n_1110, n_1655, n_445, n_2641, n_749, n_1895, n_2574, n_1134, n_1358, n_717, n_165, n_939, n_482, n_2361, n_1088, n_588, n_1173, n_789, n_1232, n_1603, n_734, n_638, n_2638, n_866, n_107, n_969, n_1401, n_2492, n_1019, n_1105, n_249, n_1998, n_304, n_1338, n_577, n_2016, n_1522, n_1687, n_1637, n_2034, n_1419, n_2711, n_338, n_149, n_1653, n_693, n_2270, n_1506, n_2653, n_14, n_836, n_990, n_2496, n_1886, n_1389, n_1894, n_975, n_1908, n_1256, n_1702, n_2259, n_2794, n_567, n_1465, n_778, n_1122, n_151, n_2608, n_306, n_2657, n_458, n_770, n_1375, n_2494, n_2649, n_1102, n_2392, n_1843, n_711, n_1499, n_85, n_1187, n_2633, n_1441, n_2522, n_2435, n_1392, n_1597, n_1929, n_2807, n_1164, n_1659, n_1834, n_2097, n_2313, n_2542, n_489, n_1174, n_2431, n_2558, n_1371, n_617, n_1303, n_2206, n_2063, n_1572, n_1968, n_2564, n_2252, n_876, n_1516, n_1190, n_1736, n_1685, n_118, n_2409, n_601, n_917, n_1714, n_966, n_253, n_1116, n_2000, n_1661, n_1212, n_2074, n_1541, n_2576, n_172, n_206, n_217, n_726, n_982, n_2575, n_1573, n_1453, n_1731, n_2217, n_818, n_2373, n_1970, n_861, n_1713, n_1183, n_2307, n_2766, n_1658, n_899, n_1253, n_210, n_1737, n_2201, n_2722, n_2117, n_2745, n_1904, n_2640, n_1993, n_774, n_1628, n_2493, n_2205, n_1335, n_1514, n_1777, n_1957, n_1059, n_1345, n_176, n_1133, n_1771, n_1912, n_1899, n_557, n_1410, n_1005, n_607, n_1003, n_679, n_710, n_2067, n_527, n_1168, n_707, n_2219, n_2437, n_2148, n_937, n_2445, n_1427, n_2779, n_393, n_108, n_487, n_1584, n_665, n_1726, n_1835, n_66, n_1440, n_177, n_2164, n_421, n_1988, n_2115, n_1853, n_1356, n_1787, n_2634, n_910, n_2232, n_2212, n_2602, n_1657, n_768, n_1475, n_1302, n_1774, n_1725, n_205, n_1136, n_1313, n_1491, n_754, n_2811, n_1496, n_179, n_1125, n_125, n_410, n_2547, n_708, n_529, n_1812, n_735, n_2501, n_232, n_1915, n_1109, n_126, n_895, n_2532, n_1310, n_2605, n_2121, n_1803, n_202, n_2665, n_427, n_1399, n_1543, n_1991, n_1979, n_791, n_732, n_1533, n_2224, n_193, n_808, n_2484, n_797, n_1025, n_1930, n_1955, n_2765, n_500, n_1067, n_1720, n_148, n_2401, n_435, n_2003, n_159, n_766, n_1457, n_541, n_2692, n_538, n_2354, n_2246, n_2008, n_1117, n_799, n_2264, n_2754, n_687, n_715, n_1742, n_1480, n_1482, n_1213, n_2489, n_1266, n_536, n_872, n_2012, n_594, n_200, n_1291, n_1297, n_1753, n_2283, n_1782, n_2245, n_1155, n_1418, n_89, n_1972, n_1524, n_1689, n_1485, n_2806, n_115, n_1011, n_1184, n_2184, n_985, n_1855, n_2425, n_869, n_810, n_416, n_827, n_401, n_1703, n_1352, n_626, n_2197, n_2199, n_1650, n_1144, n_1137, n_1570, n_1170, n_305, n_2023, n_2213, n_2351, n_2211, n_2095, n_137, n_676, n_294, n_318, n_2103, n_653, n_2160, n_642, n_2228, n_2527, n_1602, n_2498, n_194, n_855, n_1178, n_1461, n_2697, n_850, n_684, n_124, n_268, n_2421, n_2286, n_664, n_1999, n_503, n_2372, n_2065, n_2136, n_2480, n_235, n_1372, n_605, n_2630, n_1273, n_1822, n_353, n_620, n_643, n_2363, n_2430, n_916, n_1081, n_2549, n_493, n_2705, n_2332, n_1235, n_703, n_698, n_980, n_1115, n_2433, n_1282, n_1318, n_1783, n_780, n_2601, n_998, n_2375, n_2550, n_1454, n_467, n_1227, n_1531, n_840, n_1334, n_1907, n_501, n_823, n_245, n_2686, n_2528, n_725, n_2344, n_1388, n_1417, n_1295, n_2316, n_672, n_1985, n_1898, n_2107, n_581, n_382, n_554, n_1625, n_2130, n_2187, n_2284, n_898, n_2773, n_2598, n_1762, n_1013, n_1452, n_718, n_2687, n_265, n_1120, n_719, n_443, n_1791, n_198, n_1890, n_1747, n_714, n_1683, n_1817, n_909, n_1944, n_1497, n_1530, n_2654, n_997, n_932, n_612, n_2078, n_1409, n_788, n_1326, n_119, n_1268, n_559, n_825, n_1981, n_508, n_2186, n_506, n_1320, n_1663, n_737, n_1718, n_986, n_2315, n_509, n_1317, n_147, n_1518, n_1715, n_2102, n_2562, n_1281, n_67, n_1952, n_1192, n_2221, n_1024, n_1063, n_1889, n_209, n_1792, n_1564, n_1868, n_1613, n_733, n_1489, n_1922, n_1376, n_941, n_2326, n_981, n_2560, n_1569, n_2188, n_68, n_867, n_186, n_2348, n_2422, n_134, n_2239, n_587, n_63, n_792, n_756, n_1429, n_399, n_1238, n_2448, n_548, n_812, n_298, n_2104, n_2748, n_518, n_505, n_2057, n_1772, n_282, n_752, n_905, n_1476, n_1108, n_782, n_2717, n_1100, n_1861, n_2129, n_1395, n_862, n_1425, n_760, n_1901, n_1900, n_1620, n_381, n_220, n_390, n_1330, n_1867, n_31, n_1945, n_2772, n_481, n_1675, n_1924, n_2573, n_1727, n_2710, n_1554, n_1745, n_2735, n_769, n_2497, n_2006, n_42, n_1995, n_2411, n_2138, n_1046, n_271, n_934, n_1618, n_2260, n_826, n_2343, n_1813, n_2447, n_886, n_2014, n_1221, n_2345, n_654, n_1172, n_167, n_2535, n_379, n_428, n_1341, n_2726, n_570, n_2774, n_1641, n_1361, n_2382, n_1707, n_853, n_377, n_2317, n_751, n_2799, n_2172, n_1973, n_786, n_1083, n_1142, n_2376, n_2488, n_1129, n_392, n_2579, n_158, n_2476, n_704, n_787, n_1770, n_138, n_2781, n_2456, n_961, n_2250, n_2678, n_1756, n_771, n_2778, n_276, n_95, n_1716, n_2788, n_1225, n_1520, n_2451, n_169, n_522, n_1287, n_1262, n_2691, n_400, n_930, n_181, n_1873, n_1411, n_221, n_622, n_1962, n_1577, n_2423, n_1087, n_2526, n_386, n_994, n_1701, n_2194, n_848, n_1550, n_2764, n_2703, n_1498, n_2167, n_1223, n_1272, n_2680, n_104, n_682, n_1567, n_56, n_141, n_2567, n_1247, n_2709, n_922, n_816, n_1648, n_591, n_145, n_1536, n_1857, n_1344, n_2041, n_313, n_631, n_479, n_1246, n_1339, n_1478, n_1797, n_432, n_1769, n_839, n_1210, n_1364, n_2357, n_2183, n_2673, n_2742, n_2360, n_328, n_140, n_2292, n_1250, n_2173, n_369, n_1842, n_871, n_2442, n_598, n_685, n_928, n_608, n_1367, n_78, n_1943, n_1460, n_772, n_2018, n_1555, n_499, n_2531, n_1589, n_517, n_98, n_402, n_413, n_1086, n_2570, n_2702, n_796, n_1858, n_1619, n_236, n_2119, n_1502, n_2157, n_2552, n_1469, n_1012, n_1, n_1396, n_2744, n_1348, n_2030, n_903, n_2453, n_1525, n_1752, n_2397, n_740, n_203, n_384, n_2208, n_1404, n_80, n_1794, n_2182, n_35, n_1315, n_2234, n_277, n_1061, n_92, n_1910, n_333, n_1298, n_1652, n_2209, n_462, n_2050, n_2809, n_1193, n_2797, n_1676, n_1255, n_258, n_1113, n_29, n_79, n_2321, n_1226, n_722, n_1277, n_2591, n_188, n_2146, n_844, n_201, n_471, n_852, n_1487, n_40, n_1864, n_1028, n_1601, n_781, n_474, n_542, n_463, n_1546, n_595, n_502, n_466, n_2612, n_420, n_1337, n_1495, n_632, n_699, n_979, n_1515, n_1627, n_1245, n_846, n_2427, n_2438, n_2505, n_1673, n_465, n_76, n_362, n_1321, n_170, n_1975, n_27, n_2296, n_2070, n_161, n_273, n_1937, n_585, n_2112, n_1739, n_270, n_616, n_2278, n_81, n_2594, n_2394, n_1914, n_2135, n_2335, n_745, n_2381, n_1654, n_2569, n_2349, n_1103, n_648, n_1379, n_2734, n_312, n_2196, n_2170, n_1076, n_1091, n_1408, n_494, n_1761, n_641, n_730, n_2036, n_1325, n_1595, n_2161, n_354, n_575, n_480, n_425, n_795, n_2404, n_2083, n_695, n_180, n_656, n_1606, n_2503, n_1220, n_37, n_1694, n_1540, n_2485, n_229, n_1936, n_1956, n_437, n_1642, n_2279, n_2655, n_2027, n_60, n_403, n_453, n_2642, n_1130, n_720, n_0, n_2500, n_2366, n_1918, n_1526, n_863, n_2210, n_805, n_1604, n_1275, n_2513, n_2525, n_2695, n_1764, n_113, n_712, n_2414, n_246, n_1583, n_2426, n_1042, n_1402, n_269, n_2049, n_2273, n_285, n_412, n_2719, n_1493, n_657, n_644, n_1741, n_2229, n_1160, n_1397, n_491, n_1258, n_1074, n_2004, n_1621, n_2708, n_2113, n_251, n_160, n_566, n_565, n_2586, n_1448, n_2225, n_1507, n_1398, n_2383, n_1879, n_597, n_1996, n_1181, n_1505, n_1634, n_1196, n_2019, n_651, n_1340, n_2274, n_334, n_811, n_1558, n_807, n_2166, n_835, n_175, n_666, n_262, n_1433, n_1704, n_2256, n_99, n_1254, n_1026, n_2026, n_1969, n_1234, n_2109, n_319, n_364, n_1138, n_927, n_20, n_1089, n_2013, n_1990, n_2044, n_2689, n_1004, n_1186, n_1032, n_242, n_2614, n_2511, n_1681, n_2010, n_1018, n_2242, n_2247, n_2752, n_1693, n_438, n_2599, n_713, n_2704, n_904, n_1588, n_1622, n_2237, n_166, n_1180, n_1827, n_2524, n_1271, n_2802, n_533, n_1542, n_1251, n_278, n_2728, n_2268, n_13034);

input n_924;
input n_1263;
input n_977;
input n_1378;
input n_2253;
input n_2417;
input n_611;
input n_2756;
input n_1126;
input n_1423;
input n_1729;
input n_2739;
input n_1166;
input n_2380;
input n_1751;
input n_469;
input n_1508;
input n_82;
input n_2771;
input n_785;
input n_549;
input n_2617;
input n_2200;
input n_532;
input n_1161;
input n_1859;
input n_2746;
input n_1677;
input n_1150;
input n_2327;
input n_226;
input n_1780;
input n_1488;
input n_667;
input n_790;
input n_1055;
input n_2386;
input n_1501;
input n_111;
input n_2395;
input n_880;
input n_544;
input n_1007;
input n_2369;
input n_155;
input n_552;
input n_1528;
input n_2683;
input n_1370;
input n_1292;
input n_2347;
input n_2520;
input n_1198;
input n_1360;
input n_2388;
input n_1099;
input n_2568;
input n_956;
input n_564;
input n_423;
input n_1738;
input n_2021;
input n_21;
input n_2134;
input n_2391;
input n_105;
input n_1021;
input n_1960;
input n_2185;
input n_4;
input n_551;
input n_2143;
input n_2059;
input n_1323;
input n_1466;
input n_688;
input n_1695;
input n_2487;
input n_1353;
input n_800;
input n_1347;
input n_2495;
input n_1535;
input n_1789;
input n_1666;
input n_2389;
input n_671;
input n_819;
input n_1451;
input n_1022;
input n_2302;
input n_915;
input n_1545;
input n_2374;
input n_864;
input n_173;
input n_859;
input n_951;
input n_1947;
input n_1264;
input n_2114;
input n_447;
input n_247;
input n_2001;
input n_1494;
input n_292;
input n_625;
input n_854;
input n_1462;
input n_1799;
input n_2069;
input n_2396;
input n_1580;
input n_674;
input n_417;
input n_1939;
input n_2486;
input n_1806;
input n_516;
input n_933;
input n_2244;
input n_2257;
input n_1152;
input n_497;
input n_1869;
input n_1607;
input n_1563;
input n_606;
input n_275;
input n_2011;
input n_2096;
input n_26;
input n_877;
input n_2105;
input n_2538;
input n_2024;
input n_2;
input n_2530;
input n_1696;
input n_2483;
input n_755;
input n_1118;
input n_6;
input n_1686;
input n_947;
input n_1285;
input n_373;
input n_307;
input n_1860;
input n_2543;
input n_1359;
input n_530;
input n_87;
input n_150;
input n_1107;
input n_1728;
input n_556;
input n_2031;
input n_2076;
input n_2482;
input n_2677;
input n_1230;
input n_668;
input n_375;
input n_301;
input n_1896;
input n_2165;
input n_2147;
input n_929;
input n_2770;
input n_1124;
input n_1818;
input n_2127;
input n_902;
input n_1576;
input n_191;
input n_1104;
input n_1294;
input n_659;
input n_51;
input n_1705;
input n_2584;
input n_1257;
input n_2639;
input n_171;
input n_1182;
input n_579;
input n_1698;
input n_1261;
input n_2329;
input n_938;
input n_1098;
input n_2142;
input n_320;
input n_1154;
input n_2189;
input n_1242;
input n_1135;
input n_24;
input n_406;
input n_519;
input n_2323;
input n_2203;
input n_2597;
input n_1016;
input n_1243;
input n_546;
input n_101;
input n_2047;
input n_1280;
input n_1845;
input n_281;
input n_240;
input n_2052;
input n_2193;
input n_2058;
input n_2458;
input n_2478;
input n_291;
input n_231;
input n_257;
input n_2761;
input n_731;
input n_371;
input n_1483;
input n_1314;
input n_1512;
input n_709;
input n_1490;
input n_317;
input n_1236;
input n_1633;
input n_2537;
input n_569;
input n_2669;
input n_2144;
input n_1778;
input n_227;
input n_2306;
input n_920;
input n_2515;
input n_1289;
input n_1517;
input n_2091;
input n_2466;
input n_2635;
input n_2652;
input n_94;
input n_335;
input n_2715;
input n_2085;
input n_1669;
input n_2566;
input n_370;
input n_976;
input n_1949;
input n_343;
input n_1449;
input n_308;
input n_1946;
input n_1566;
input n_2032;
input n_297;
input n_2587;
input n_156;
input n_2149;
input n_1078;
input n_2782;
input n_1670;
input n_2672;
input n_775;
input n_219;
input n_157;
input n_2651;
input n_600;
input n_1484;
input n_2071;
input n_2561;
input n_1374;
input n_1328;
input n_2643;
input n_223;
input n_2141;
input n_1948;
input n_1984;
input n_2099;
input n_2408;
input n_264;
input n_1877;
input n_1831;
input n_1598;
input n_1723;
input n_955;
input n_1850;
input n_163;
input n_339;
input n_1146;
input n_882;
input n_183;
input n_243;
input n_2384;
input n_1036;
input n_1097;
input n_1749;
input n_347;
input n_59;
input n_550;
input n_696;
input n_897;
input n_215;
input n_350;
input n_196;
input n_798;
input n_646;
input n_1428;
input n_2663;
input n_436;
input n_1394;
input n_2659;
input n_1414;
input n_1216;
input n_290;
input n_580;
input n_2693;
input n_1040;
input n_2202;
input n_2648;
input n_1872;
input n_1852;
input n_2159;
input n_578;
input n_926;
input n_2180;
input n_2249;
input n_344;
input n_2353;
input n_1218;
input n_1931;
input n_2439;
input n_2632;
input n_2276;
input n_422;
input n_475;
input n_777;
input n_1070;
input n_1547;
input n_2089;
input n_1030;
input n_72;
input n_2470;
input n_1755;
input n_415;
input n_1071;
input n_485;
input n_1165;
input n_1267;
input n_1561;
input n_496;
input n_1801;
input n_1391;
input n_958;
input n_1034;
input n_670;
input n_1513;
input n_1600;
input n_48;
input n_521;
input n_663;
input n_845;
input n_2235;
input n_1862;
input n_673;
input n_837;
input n_1239;
input n_528;
input n_2300;
input n_2791;
input n_1796;
input n_2551;
input n_680;
input n_1473;
input n_1587;
input n_2682;
input n_395;
input n_164;
input n_553;
input n_901;
input n_2432;
input n_813;
input n_1521;
input n_1284;
input n_1590;
input n_214;
input n_2174;
input n_2714;
input n_1748;
input n_1672;
input n_2506;
input n_675;
input n_2699;
input n_888;
input n_1880;
input n_2769;
input n_2337;
input n_1167;
input n_1626;
input n_637;
input n_2615;
input n_1384;
input n_1556;
input n_184;
input n_446;
input n_1863;
input n_1064;
input n_144;
input n_858;
input n_2079;
input n_2238;
input n_114;
input n_96;
input n_923;
input n_2118;
input n_691;
input n_1151;
input n_881;
input n_1405;
input n_2407;
input n_1706;
input n_468;
input n_213;
input n_129;
input n_342;
input n_2753;
input n_464;
input n_363;
input n_1582;
input n_197;
input n_1069;
input n_1784;
input n_1075;
input n_1836;
input n_1450;
input n_1322;
input n_2101;
input n_1471;
input n_1986;
input n_2072;
input n_2738;
input n_1750;
input n_1459;
input n_460;
input n_889;
input n_2358;
input n_973;
input n_1700;
input n_477;
input n_571;
input n_1585;
input n_461;
input n_2684;
input n_2712;
input n_1971;
input n_1599;
input n_2275;
input n_2713;
input n_2644;
input n_2700;
input n_1211;
input n_1197;
input n_1523;
input n_2730;
input n_1950;
input n_907;
input n_1447;
input n_2251;
input n_1377;
input n_2370;
input n_190;
input n_989;
input n_2544;
input n_1039;
input n_2214;
input n_34;
input n_2055;
input n_228;
input n_283;
input n_1403;
input n_2248;
input n_2356;
input n_488;
input n_736;
input n_892;
input n_2688;
input n_1000;
input n_1202;
input n_2750;
input n_2620;
input n_1278;
input n_2622;
input n_2062;
input n_2668;
input n_1002;
input n_1463;
input n_1581;
input n_2100;
input n_49;
input n_310;
input n_54;
input n_593;
input n_2258;
input n_12;
input n_748;
input n_586;
input n_1058;
input n_1667;
input n_838;
input n_2784;
input n_332;
input n_1053;
input n_1224;
input n_349;
input n_2557;
input n_1926;
input n_2706;
input n_1248;
input n_230;
input n_1331;
input n_953;
input n_279;
input n_1014;
input n_1241;
input n_70;
input n_2150;
input n_2241;
input n_2757;
input n_2152;
input n_289;
input n_963;
input n_1052;
input n_954;
input n_627;
input n_1385;
input n_440;
input n_793;
input n_478;
input n_2590;
input n_2776;
input n_2140;
input n_2385;
input n_1819;
input n_2330;
input n_2139;
input n_476;
input n_1527;
input n_2042;
input n_534;
input n_1882;
input n_884;
input n_345;
input n_944;
input n_1754;
input n_1623;
input n_2175;
input n_2720;
input n_2324;
input n_1854;
input n_91;
input n_2606;
input n_2674;
input n_1565;
input n_1809;
input n_1856;
input n_182;
input n_143;
input n_647;
input n_237;
input n_407;
input n_1072;
input n_2218;
input n_2267;
input n_832;
input n_857;
input n_2305;
input n_2636;
input n_2450;
input n_207;
input n_561;
input n_1319;
input n_2379;
input n_2616;
input n_2154;
input n_1825;
input n_1951;
input n_1883;
input n_1906;
input n_2759;
input n_1712;
input n_1387;
input n_2262;
input n_2462;
input n_2514;
input n_1532;
input n_2322;
input n_2271;
input n_2625;
input n_18;
input n_1027;
input n_971;
input n_1156;
input n_117;
input n_326;
input n_794;
input n_404;
input n_2798;
input n_2331;
input n_2293;
input n_686;
input n_847;
input n_1393;
input n_2319;
input n_596;
input n_1775;
input n_2028;
input n_1368;
input n_2762;
input n_558;
input n_2808;
input n_702;
input n_1276;
input n_2548;
input n_822;
input n_1412;
input n_2676;
input n_1709;
input n_2679;
input n_2108;
input n_728;
input n_266;
input n_1162;
input n_272;
input n_1538;
input n_1838;
input n_1199;
input n_1847;
input n_1779;
input n_2767;
input n_2777;
input n_2603;
input n_352;
input n_1884;
input n_2434;
input n_2660;
input n_53;
input n_1038;
input n_520;
input n_1369;
input n_409;
input n_2611;
input n_1841;
input n_1660;
input n_887;
input n_1905;
input n_2553;
input n_154;
input n_2581;
input n_71;
input n_2195;
input n_2529;
input n_300;
input n_2698;
input n_809;
input n_870;
input n_931;
input n_599;
input n_1711;
input n_1662;
input n_1891;
input n_1481;
input n_2626;
input n_1942;
input n_434;
input n_1978;
input n_1544;
input n_2510;
input n_868;
input n_2454;
input n_639;
input n_2804;
input n_914;
input n_2120;
input n_411;
input n_414;
input n_2546;
input n_1629;
input n_1293;
input n_2801;
input n_965;
input n_1876;
input n_1743;
input n_935;
input n_121;
input n_1175;
input n_817;
input n_2763;
input n_360;
input n_36;
input n_1479;
input n_1810;
input n_2350;
input n_2813;
input n_64;
input n_1888;
input n_2009;
input n_759;
input n_2222;
input n_1892;
input n_28;
input n_806;
input n_1997;
input n_2667;
input n_1766;
input n_1477;
input n_324;
input n_1635;
input n_1963;
input n_2226;
input n_1571;
input n_187;
input n_1189;
input n_2690;
input n_103;
input n_97;
input n_11;
input n_2215;
input n_7;
input n_1259;
input n_1690;
input n_706;
input n_746;
input n_1649;
input n_747;
input n_2064;
input n_52;
input n_784;
input n_110;
input n_2449;
input n_1733;
input n_1244;
input n_2413;
input n_431;
input n_1194;
input n_1925;
input n_2297;
input n_1815;
input n_2621;
input n_615;
input n_851;
input n_1759;
input n_843;
input n_1788;
input n_2177;
input n_2491;
input n_523;
input n_913;
input n_1537;
input n_705;
input n_865;
input n_61;
input n_2227;
input n_678;
input n_2671;
input n_697;
input n_127;
input n_1222;
input n_75;
input n_1679;
input n_2190;
input n_776;
input n_1798;
input n_2022;
input n_1790;
input n_2518;
input n_1415;
input n_367;
input n_2629;
input n_2592;
input n_452;
input n_525;
input n_1260;
input n_1746;
input n_1647;
input n_2181;
input n_2479;
input n_1829;
input n_1464;
input n_649;
input n_547;
input n_2563;
input n_43;
input n_1444;
input n_1191;
input n_2387;
input n_1674;
input n_1833;
input n_116;
input n_1830;
input n_2517;
input n_2073;
input n_1710;
input n_284;
input n_1128;
input n_139;
input n_1734;
input n_744;
input n_590;
input n_629;
input n_2631;
input n_1308;
input n_2178;
input n_1767;
input n_2336;
input n_254;
input n_1680;
input n_1233;
input n_2607;
input n_23;
input n_1615;
input n_1529;
input n_2005;
input n_526;
input n_1916;
input n_293;
input n_372;
input n_677;
input n_244;
input n_47;
input n_1333;
input n_2469;
input n_1121;
input n_2723;
input n_314;
input n_368;
input n_433;
input n_604;
input n_2007;
input n_8;
input n_949;
input n_2539;
input n_100;
input n_2582;
input n_1443;
input n_1008;
input n_946;
input n_1539;
input n_2736;
input n_1001;
input n_1503;
input n_2054;
input n_498;
input n_1468;
input n_1559;
input n_1765;
input n_1866;
input n_689;
input n_738;
input n_1624;
input n_640;
input n_1510;
input n_252;
input n_624;
input n_1380;
input n_1744;
input n_2623;
input n_1617;
input n_295;
input n_133;
input n_1010;
input n_1994;
input n_1231;
input n_739;
input n_1279;
input n_1406;
input n_2718;
input n_1195;
input n_1837;
input n_1839;
input n_610;
input n_2577;
input n_1760;
input n_936;
input n_568;
input n_1500;
input n_39;
input n_1090;
input n_2796;
input n_757;
input n_2342;
input n_633;
input n_439;
input n_106;
input n_1832;
input n_259;
input n_448;
input n_1851;
input n_758;
input n_999;
input n_2046;
input n_2741;
input n_1933;
input n_2290;
input n_93;
input n_1656;
input n_1158;
input n_2045;
input n_1509;
input n_1874;
input n_2040;
input n_563;
input n_2060;
input n_2613;
input n_1987;
input n_2805;
input n_1145;
input n_878;
input n_524;
input n_204;
input n_394;
input n_1678;
input n_1049;
input n_1153;
input n_2145;
input n_741;
input n_1639;
input n_1306;
input n_1068;
input n_1871;
input n_2580;
input n_2545;
input n_2787;
input n_1964;
input n_122;
input n_331;
input n_10;
input n_906;
input n_1163;
input n_2039;
input n_1207;
input n_919;
input n_908;
input n_2412;
input n_2406;
input n_90;
input n_724;
input n_1781;
input n_2084;
input n_2035;
input n_658;
input n_2061;
input n_2378;
input n_2509;
input n_1740;
input n_2398;
input n_1362;
input n_1586;
input n_456;
input n_959;
input n_2459;
input n_535;
input n_152;
input n_940;
input n_1445;
input n_9;
input n_1492;
input n_2155;
input n_2516;
input n_1923;
input n_1773;
input n_592;
input n_1169;
input n_45;
input n_1596;
input n_1692;
input n_2666;
input n_1017;
input n_2481;
input n_2171;
input n_123;
input n_978;
input n_2768;
input n_2116;
input n_2314;
input n_1434;
input n_1054;
input n_2507;
input n_1474;
input n_1665;
input n_1269;
input n_2420;
input n_1095;
input n_1828;
input n_1614;
input n_267;
input n_514;
input n_457;
input n_1079;
input n_1045;
input n_1208;
input n_2093;
input n_2038;
input n_2320;
input n_2339;
input n_2473;
input n_2137;
input n_603;
input n_1431;
input n_2583;
input n_484;
input n_1593;
input n_1033;
input n_442;
input n_2299;
input n_131;
input n_2540;
input n_636;
input n_660;
input n_2087;
input n_1640;
input n_2162;
input n_1732;
input n_1009;
input n_1148;
input n_2051;
input n_109;
input n_742;
input n_750;
input n_2029;
input n_995;
input n_454;
input n_2168;
input n_2790;
input n_1609;
input n_374;
input n_1989;
input n_185;
input n_2359;
input n_396;
input n_1887;
input n_2523;
input n_1383;
input n_1073;
input n_255;
input n_2346;
input n_2457;
input n_662;
input n_459;
input n_2312;
input n_218;
input n_962;
input n_1215;
input n_1171;
input n_1578;
input n_723;
input n_1920;
input n_1065;
input n_1592;
input n_2536;
input n_1336;
input n_1721;
input n_1959;
input n_1758;
input n_2338;
input n_2737;
input n_1574;
input n_2399;
input n_2812;
input n_473;
input n_2048;
input n_2355;
input n_2133;
input n_1921;
input n_2721;
input n_1309;
input n_1878;
input n_1426;
input n_1043;
input n_2585;
input n_355;
input n_486;
input n_1800;
input n_1548;
input n_2725;
input n_614;
input n_337;
input n_1421;
input n_88;
input n_2571;
input n_1286;
input n_1177;
input n_1355;
input n_168;
input n_974;
input n_2565;
input n_727;
input n_1159;
input n_957;
input n_773;
input n_208;
input n_142;
input n_2124;
input n_743;
input n_2081;
input n_299;
input n_303;
input n_296;
input n_613;
input n_1119;
input n_2156;
input n_1240;
input n_2261;
input n_1820;
input n_2729;
input n_2418;
input n_65;
input n_829;
input n_2519;
input n_2724;
input n_1612;
input n_2179;
input n_1416;
input n_2077;
input n_1724;
input n_2111;
input n_2521;
input n_361;
input n_700;
input n_1237;
input n_573;
input n_69;
input n_1420;
input n_1132;
input n_388;
input n_1366;
input n_1300;
input n_2595;
input n_1127;
input n_2277;
input n_761;
input n_2477;
input n_1785;
input n_1568;
input n_1006;
input n_2110;
input n_329;
input n_274;
input n_1270;
input n_1664;
input n_1486;
input n_582;
input n_1332;
input n_2231;
input n_1390;
input n_2017;
input n_73;
input n_2474;
input n_2604;
input n_19;
input n_2090;
input n_1870;
input n_309;
input n_30;
input n_512;
input n_2367;
input n_1591;
input n_2033;
input n_84;
input n_130;
input n_322;
input n_1682;
input n_1980;
input n_2390;
input n_2628;
input n_1249;
input n_652;
input n_1111;
input n_1365;
input n_1927;
input n_25;
input n_2132;
input n_1349;
input n_1093;
input n_288;
input n_2400;
input n_1031;
input n_263;
input n_609;
input n_1041;
input n_1265;
input n_1909;
input n_44;
input n_224;
input n_2681;
input n_1562;
input n_383;
input n_834;
input n_112;
input n_765;
input n_2255;
input n_2424;
input n_2272;
input n_893;
input n_1015;
input n_1140;
input n_891;
input n_1651;
input n_1965;
input n_239;
input n_630;
input n_1902;
input n_2151;
input n_1941;
input n_55;
input n_2106;
input n_2775;
input n_2716;
input n_1913;
input n_504;
input n_1823;
input n_511;
input n_874;
input n_2464;
input n_358;
input n_1101;
input n_77;
input n_102;
input n_1106;
input n_1456;
input n_2230;
input n_2015;
input n_2365;
input n_1875;
input n_1982;
input n_1304;
input n_2803;
input n_1324;
input n_987;
input n_1846;
input n_261;
input n_174;
input n_2066;
input n_1885;
input n_1455;
input n_767;
input n_993;
input n_1903;
input n_2490;
input n_1407;
input n_2452;
input n_1551;
input n_545;
input n_441;
input n_860;
input n_450;
input n_1805;
input n_2176;
input n_2204;
input n_1816;
input n_429;
input n_948;
input n_1217;
input n_2220;
input n_2455;
input n_628;
input n_365;
input n_1849;
input n_2410;
input n_729;
input n_1131;
input n_1084;
input n_1961;
input n_970;
input n_1935;
input n_911;
input n_1430;
input n_83;
input n_2645;
input n_2467;
input n_513;
input n_2727;
input n_1094;
input n_1354;
input n_560;
input n_1534;
input n_340;
input n_2288;
input n_1351;
input n_2240;
input n_2696;
input n_1044;
input n_1205;
input n_2436;
input n_346;
input n_1209;
input n_1552;
input n_2508;
input n_495;
input n_602;
input n_574;
input n_2593;
input n_1435;
input n_879;
input n_16;
input n_2416;
input n_58;
input n_2405;
input n_623;
input n_2088;
input n_405;
input n_824;
input n_359;
input n_1645;
input n_2461;
input n_490;
input n_1327;
input n_2243;
input n_996;
input n_921;
input n_1684;
input n_233;
input n_2658;
input n_1717;
input n_572;
input n_366;
input n_815;
input n_1795;
input n_2128;
input n_2578;
input n_128;
input n_1821;
input n_120;
input n_327;
input n_135;
input n_1381;
input n_2555;
input n_2662;
input n_2740;
input n_1611;
input n_1037;
input n_2368;
input n_2656;
input n_1080;
input n_2301;
input n_1274;
input n_2554;
input n_1316;
input n_1708;
input n_2419;
input n_426;
input n_1438;
input n_1082;
input n_1840;
input n_589;
input n_716;
input n_1630;
input n_2122;
input n_2512;
input n_562;
input n_1436;
input n_62;
input n_1691;
input n_952;
input n_2786;
input n_2534;
input n_2092;
input n_1229;
input n_391;
input n_701;
input n_1437;
input n_1023;
input n_2075;
input n_645;
input n_539;
input n_803;
input n_1092;
input n_2694;
input n_238;
input n_1776;
input n_2198;
input n_2610;
input n_2661;
input n_2572;
input n_2281;
input n_2131;
input n_2789;
input n_2216;
input n_531;
input n_1757;
input n_890;
input n_1897;
input n_764;
input n_1919;
input n_1056;
input n_1424;
input n_162;
input n_960;
input n_2308;
input n_1893;
input n_222;
input n_1290;
input n_1123;
input n_1467;
input n_1047;
input n_2053;
input n_2163;
input n_634;
input n_2328;
input n_199;
input n_1958;
input n_32;
input n_2254;
input n_1252;
input n_348;
input n_1382;
input n_1029;
input n_925;
input n_1206;
input n_424;
input n_2647;
input n_1311;
input n_2191;
input n_1519;
input n_256;
input n_950;
input n_2428;
input n_1553;
input n_2664;
input n_1811;
input n_2443;
input n_2624;
input n_380;
input n_419;
input n_1346;
input n_444;
input n_1299;
input n_2158;
input n_1808;
input n_1060;
input n_1141;
input n_316;
input n_2266;
input n_389;
input n_2465;
input n_2650;
input n_418;
input n_248;
input n_136;
input n_86;
input n_146;
input n_912;
input n_315;
input n_968;
input n_451;
input n_619;
input n_408;
input n_2440;
input n_1386;
input n_1699;
input n_376;
input n_967;
input n_1442;
input n_2541;
input n_74;
input n_1139;
input n_2731;
input n_515;
input n_2333;
input n_57;
input n_351;
input n_885;
input n_397;
input n_1432;
input n_1357;
input n_483;
input n_2125;
input n_683;
input n_1632;
input n_1057;
input n_1051;
input n_1085;
input n_1066;
input n_721;
input n_2402;
input n_1157;
input n_2403;
input n_841;
input n_1050;
input n_22;
input n_802;
input n_1954;
input n_2265;
input n_46;
input n_1608;
input n_983;
input n_1844;
input n_2760;
input n_2792;
input n_38;
input n_280;
input n_1305;
input n_873;
input n_1826;
input n_378;
input n_1112;
input n_2304;
input n_762;
input n_1283;
input n_1644;
input n_17;
input n_2334;
input n_2637;
input n_690;
input n_33;
input n_1974;
input n_2463;
input n_583;
input n_2086;
input n_2289;
input n_302;
input n_1343;
input n_2701;
input n_2783;
input n_2263;
input n_1203;
input n_1631;
input n_2472;
input n_821;
input n_1763;
input n_2341;
input n_1966;
input n_1768;
input n_321;
input n_2294;
input n_1179;
input n_621;
input n_753;
input n_2475;
input n_2733;
input n_455;
input n_1048;
input n_1719;
input n_1288;
input n_212;
input n_385;
input n_2785;
input n_2556;
input n_507;
input n_2269;
input n_2732;
input n_2309;
input n_2415;
input n_2646;
input n_1560;
input n_1605;
input n_2236;
input n_330;
input n_1228;
input n_2123;
input n_972;
input n_692;
input n_2037;
input n_2685;
input n_1953;
input n_1938;
input n_820;
input n_1200;
input n_2499;
input n_1911;
input n_2460;
input n_2589;
input n_1301;
input n_1363;
input n_1668;
input n_1185;
input n_991;
input n_828;
input n_1967;
input n_779;
input n_576;
input n_1143;
input n_1579;
input n_2233;
input n_1329;
input n_2743;
input n_2675;
input n_1312;
input n_1439;
input n_804;
input n_537;
input n_1688;
input n_945;
input n_492;
input n_153;
input n_1504;
input n_943;
input n_341;
input n_250;
input n_992;
input n_1932;
input n_2755;
input n_543;
input n_260;
input n_842;
input n_650;
input n_984;
input n_694;
input n_2082;
input n_286;
input n_1992;
input n_2429;
input n_1643;
input n_883;
input n_1983;
input n_470;
input n_325;
input n_449;
input n_1594;
input n_132;
input n_1214;
input n_1342;
input n_1400;
input n_900;
input n_2362;
input n_856;
input n_2609;
input n_1793;
input n_1976;
input n_2223;
input n_918;
input n_942;
input n_2169;
input n_1804;
input n_189;
input n_1147;
input n_1557;
input n_1977;
input n_2153;
input n_2468;
input n_1610;
input n_13;
input n_1077;
input n_1422;
input n_2364;
input n_2533;
input n_540;
input n_618;
input n_896;
input n_2310;
input n_2780;
input n_323;
input n_2287;
input n_195;
input n_356;
input n_2291;
input n_2596;
input n_894;
input n_1636;
input n_2056;
input n_1730;
input n_831;
input n_2280;
input n_2192;
input n_964;
input n_1373;
input n_1350;
input n_1511;
input n_1865;
input n_1470;
input n_1096;
input n_2094;
input n_2670;
input n_234;
input n_1575;
input n_1697;
input n_1735;
input n_833;
input n_2318;
input n_2393;
input n_2020;
input n_5;
input n_1646;
input n_2502;
input n_225;
input n_2504;
input n_1307;
input n_1881;
input n_988;
input n_2749;
input n_2043;
input n_1940;
input n_814;
input n_2707;
input n_2751;
input n_2793;
input n_192;
input n_1549;
input n_1934;
input n_2311;
input n_1201;
input n_1114;
input n_655;
input n_2025;
input n_1616;
input n_1446;
input n_2285;
input n_2758;
input n_669;
input n_472;
input n_1458;
input n_1176;
input n_1472;
input n_2298;
input n_2471;
input n_1807;
input n_387;
input n_1149;
input n_2618;
input n_398;
input n_1671;
input n_635;
input n_2559;
input n_763;
input n_1020;
input n_1062;
input n_211;
input n_2303;
input n_1824;
input n_1917;
input n_2295;
input n_1219;
input n_3;
input n_1204;
input n_2810;
input n_2325;
input n_178;
input n_2747;
input n_2446;
input n_1814;
input n_1035;
input n_287;
input n_555;
input n_783;
input n_1848;
input n_1928;
input n_2126;
input n_1188;
input n_2588;
input n_1722;
input n_661;
input n_2441;
input n_41;
input n_1802;
input n_2600;
input n_849;
input n_2795;
input n_15;
input n_336;
input n_584;
input n_681;
input n_1638;
input n_1786;
input n_50;
input n_430;
input n_2002;
input n_2282;
input n_510;
input n_2800;
input n_216;
input n_2371;
input n_311;
input n_830;
input n_2098;
input n_1296;
input n_2627;
input n_2352;
input n_1413;
input n_801;
input n_2207;
input n_2080;
input n_2377;
input n_2619;
input n_2340;
input n_2444;
input n_2068;
input n_241;
input n_875;
input n_357;
input n_1110;
input n_1655;
input n_445;
input n_2641;
input n_749;
input n_1895;
input n_2574;
input n_1134;
input n_1358;
input n_717;
input n_165;
input n_939;
input n_482;
input n_2361;
input n_1088;
input n_588;
input n_1173;
input n_789;
input n_1232;
input n_1603;
input n_734;
input n_638;
input n_2638;
input n_866;
input n_107;
input n_969;
input n_1401;
input n_2492;
input n_1019;
input n_1105;
input n_249;
input n_1998;
input n_304;
input n_1338;
input n_577;
input n_2016;
input n_1522;
input n_1687;
input n_1637;
input n_2034;
input n_1419;
input n_2711;
input n_338;
input n_149;
input n_1653;
input n_693;
input n_2270;
input n_1506;
input n_2653;
input n_14;
input n_836;
input n_990;
input n_2496;
input n_1886;
input n_1389;
input n_1894;
input n_975;
input n_1908;
input n_1256;
input n_1702;
input n_2259;
input n_2794;
input n_567;
input n_1465;
input n_778;
input n_1122;
input n_151;
input n_2608;
input n_306;
input n_2657;
input n_458;
input n_770;
input n_1375;
input n_2494;
input n_2649;
input n_1102;
input n_2392;
input n_1843;
input n_711;
input n_1499;
input n_85;
input n_1187;
input n_2633;
input n_1441;
input n_2522;
input n_2435;
input n_1392;
input n_1597;
input n_1929;
input n_2807;
input n_1164;
input n_1659;
input n_1834;
input n_2097;
input n_2313;
input n_2542;
input n_489;
input n_1174;
input n_2431;
input n_2558;
input n_1371;
input n_617;
input n_1303;
input n_2206;
input n_2063;
input n_1572;
input n_1968;
input n_2564;
input n_2252;
input n_876;
input n_1516;
input n_1190;
input n_1736;
input n_1685;
input n_118;
input n_2409;
input n_601;
input n_917;
input n_1714;
input n_966;
input n_253;
input n_1116;
input n_2000;
input n_1661;
input n_1212;
input n_2074;
input n_1541;
input n_2576;
input n_172;
input n_206;
input n_217;
input n_726;
input n_982;
input n_2575;
input n_1573;
input n_1453;
input n_1731;
input n_2217;
input n_818;
input n_2373;
input n_1970;
input n_861;
input n_1713;
input n_1183;
input n_2307;
input n_2766;
input n_1658;
input n_899;
input n_1253;
input n_210;
input n_1737;
input n_2201;
input n_2722;
input n_2117;
input n_2745;
input n_1904;
input n_2640;
input n_1993;
input n_774;
input n_1628;
input n_2493;
input n_2205;
input n_1335;
input n_1514;
input n_1777;
input n_1957;
input n_1059;
input n_1345;
input n_176;
input n_1133;
input n_1771;
input n_1912;
input n_1899;
input n_557;
input n_1410;
input n_1005;
input n_607;
input n_1003;
input n_679;
input n_710;
input n_2067;
input n_527;
input n_1168;
input n_707;
input n_2219;
input n_2437;
input n_2148;
input n_937;
input n_2445;
input n_1427;
input n_2779;
input n_393;
input n_108;
input n_487;
input n_1584;
input n_665;
input n_1726;
input n_1835;
input n_66;
input n_1440;
input n_177;
input n_2164;
input n_421;
input n_1988;
input n_2115;
input n_1853;
input n_1356;
input n_1787;
input n_2634;
input n_910;
input n_2232;
input n_2212;
input n_2602;
input n_1657;
input n_768;
input n_1475;
input n_1302;
input n_1774;
input n_1725;
input n_205;
input n_1136;
input n_1313;
input n_1491;
input n_754;
input n_2811;
input n_1496;
input n_179;
input n_1125;
input n_125;
input n_410;
input n_2547;
input n_708;
input n_529;
input n_1812;
input n_735;
input n_2501;
input n_232;
input n_1915;
input n_1109;
input n_126;
input n_895;
input n_2532;
input n_1310;
input n_2605;
input n_2121;
input n_1803;
input n_202;
input n_2665;
input n_427;
input n_1399;
input n_1543;
input n_1991;
input n_1979;
input n_791;
input n_732;
input n_1533;
input n_2224;
input n_193;
input n_808;
input n_2484;
input n_797;
input n_1025;
input n_1930;
input n_1955;
input n_2765;
input n_500;
input n_1067;
input n_1720;
input n_148;
input n_2401;
input n_435;
input n_2003;
input n_159;
input n_766;
input n_1457;
input n_541;
input n_2692;
input n_538;
input n_2354;
input n_2246;
input n_2008;
input n_1117;
input n_799;
input n_2264;
input n_2754;
input n_687;
input n_715;
input n_1742;
input n_1480;
input n_1482;
input n_1213;
input n_2489;
input n_1266;
input n_536;
input n_872;
input n_2012;
input n_594;
input n_200;
input n_1291;
input n_1297;
input n_1753;
input n_2283;
input n_1782;
input n_2245;
input n_1155;
input n_1418;
input n_89;
input n_1972;
input n_1524;
input n_1689;
input n_1485;
input n_2806;
input n_115;
input n_1011;
input n_1184;
input n_2184;
input n_985;
input n_1855;
input n_2425;
input n_869;
input n_810;
input n_416;
input n_827;
input n_401;
input n_1703;
input n_1352;
input n_626;
input n_2197;
input n_2199;
input n_1650;
input n_1144;
input n_1137;
input n_1570;
input n_1170;
input n_305;
input n_2023;
input n_2213;
input n_2351;
input n_2211;
input n_2095;
input n_137;
input n_676;
input n_294;
input n_318;
input n_2103;
input n_653;
input n_2160;
input n_642;
input n_2228;
input n_2527;
input n_1602;
input n_2498;
input n_194;
input n_855;
input n_1178;
input n_1461;
input n_2697;
input n_850;
input n_684;
input n_124;
input n_268;
input n_2421;
input n_2286;
input n_664;
input n_1999;
input n_503;
input n_2372;
input n_2065;
input n_2136;
input n_2480;
input n_235;
input n_1372;
input n_605;
input n_2630;
input n_1273;
input n_1822;
input n_353;
input n_620;
input n_643;
input n_2363;
input n_2430;
input n_916;
input n_1081;
input n_2549;
input n_493;
input n_2705;
input n_2332;
input n_1235;
input n_703;
input n_698;
input n_980;
input n_1115;
input n_2433;
input n_1282;
input n_1318;
input n_1783;
input n_780;
input n_2601;
input n_998;
input n_2375;
input n_2550;
input n_1454;
input n_467;
input n_1227;
input n_1531;
input n_840;
input n_1334;
input n_1907;
input n_501;
input n_823;
input n_245;
input n_2686;
input n_2528;
input n_725;
input n_2344;
input n_1388;
input n_1417;
input n_1295;
input n_2316;
input n_672;
input n_1985;
input n_1898;
input n_2107;
input n_581;
input n_382;
input n_554;
input n_1625;
input n_2130;
input n_2187;
input n_2284;
input n_898;
input n_2773;
input n_2598;
input n_1762;
input n_1013;
input n_1452;
input n_718;
input n_2687;
input n_265;
input n_1120;
input n_719;
input n_443;
input n_1791;
input n_198;
input n_1890;
input n_1747;
input n_714;
input n_1683;
input n_1817;
input n_909;
input n_1944;
input n_1497;
input n_1530;
input n_2654;
input n_997;
input n_932;
input n_612;
input n_2078;
input n_1409;
input n_788;
input n_1326;
input n_119;
input n_1268;
input n_559;
input n_825;
input n_1981;
input n_508;
input n_2186;
input n_506;
input n_1320;
input n_1663;
input n_737;
input n_1718;
input n_986;
input n_2315;
input n_509;
input n_1317;
input n_147;
input n_1518;
input n_1715;
input n_2102;
input n_2562;
input n_1281;
input n_67;
input n_1952;
input n_1192;
input n_2221;
input n_1024;
input n_1063;
input n_1889;
input n_209;
input n_1792;
input n_1564;
input n_1868;
input n_1613;
input n_733;
input n_1489;
input n_1922;
input n_1376;
input n_941;
input n_2326;
input n_981;
input n_2560;
input n_1569;
input n_2188;
input n_68;
input n_867;
input n_186;
input n_2348;
input n_2422;
input n_134;
input n_2239;
input n_587;
input n_63;
input n_792;
input n_756;
input n_1429;
input n_399;
input n_1238;
input n_2448;
input n_548;
input n_812;
input n_298;
input n_2104;
input n_2748;
input n_518;
input n_505;
input n_2057;
input n_1772;
input n_282;
input n_752;
input n_905;
input n_1476;
input n_1108;
input n_782;
input n_2717;
input n_1100;
input n_1861;
input n_2129;
input n_1395;
input n_862;
input n_1425;
input n_760;
input n_1901;
input n_1900;
input n_1620;
input n_381;
input n_220;
input n_390;
input n_1330;
input n_1867;
input n_31;
input n_1945;
input n_2772;
input n_481;
input n_1675;
input n_1924;
input n_2573;
input n_1727;
input n_2710;
input n_1554;
input n_1745;
input n_2735;
input n_769;
input n_2497;
input n_2006;
input n_42;
input n_1995;
input n_2411;
input n_2138;
input n_1046;
input n_271;
input n_934;
input n_1618;
input n_2260;
input n_826;
input n_2343;
input n_1813;
input n_2447;
input n_886;
input n_2014;
input n_1221;
input n_2345;
input n_654;
input n_1172;
input n_167;
input n_2535;
input n_379;
input n_428;
input n_1341;
input n_2726;
input n_570;
input n_2774;
input n_1641;
input n_1361;
input n_2382;
input n_1707;
input n_853;
input n_377;
input n_2317;
input n_751;
input n_2799;
input n_2172;
input n_1973;
input n_786;
input n_1083;
input n_1142;
input n_2376;
input n_2488;
input n_1129;
input n_392;
input n_2579;
input n_158;
input n_2476;
input n_704;
input n_787;
input n_1770;
input n_138;
input n_2781;
input n_2456;
input n_961;
input n_2250;
input n_2678;
input n_1756;
input n_771;
input n_2778;
input n_276;
input n_95;
input n_1716;
input n_2788;
input n_1225;
input n_1520;
input n_2451;
input n_169;
input n_522;
input n_1287;
input n_1262;
input n_2691;
input n_400;
input n_930;
input n_181;
input n_1873;
input n_1411;
input n_221;
input n_622;
input n_1962;
input n_1577;
input n_2423;
input n_1087;
input n_2526;
input n_386;
input n_994;
input n_1701;
input n_2194;
input n_848;
input n_1550;
input n_2764;
input n_2703;
input n_1498;
input n_2167;
input n_1223;
input n_1272;
input n_2680;
input n_104;
input n_682;
input n_1567;
input n_56;
input n_141;
input n_2567;
input n_1247;
input n_2709;
input n_922;
input n_816;
input n_1648;
input n_591;
input n_145;
input n_1536;
input n_1857;
input n_1344;
input n_2041;
input n_313;
input n_631;
input n_479;
input n_1246;
input n_1339;
input n_1478;
input n_1797;
input n_432;
input n_1769;
input n_839;
input n_1210;
input n_1364;
input n_2357;
input n_2183;
input n_2673;
input n_2742;
input n_2360;
input n_328;
input n_140;
input n_2292;
input n_1250;
input n_2173;
input n_369;
input n_1842;
input n_871;
input n_2442;
input n_598;
input n_685;
input n_928;
input n_608;
input n_1367;
input n_78;
input n_1943;
input n_1460;
input n_772;
input n_2018;
input n_1555;
input n_499;
input n_2531;
input n_1589;
input n_517;
input n_98;
input n_402;
input n_413;
input n_1086;
input n_2570;
input n_2702;
input n_796;
input n_1858;
input n_1619;
input n_236;
input n_2119;
input n_1502;
input n_2157;
input n_2552;
input n_1469;
input n_1012;
input n_1;
input n_1396;
input n_2744;
input n_1348;
input n_2030;
input n_903;
input n_2453;
input n_1525;
input n_1752;
input n_2397;
input n_740;
input n_203;
input n_384;
input n_2208;
input n_1404;
input n_80;
input n_1794;
input n_2182;
input n_35;
input n_1315;
input n_2234;
input n_277;
input n_1061;
input n_92;
input n_1910;
input n_333;
input n_1298;
input n_1652;
input n_2209;
input n_462;
input n_2050;
input n_2809;
input n_1193;
input n_2797;
input n_1676;
input n_1255;
input n_258;
input n_1113;
input n_29;
input n_79;
input n_2321;
input n_1226;
input n_722;
input n_1277;
input n_2591;
input n_188;
input n_2146;
input n_844;
input n_201;
input n_471;
input n_852;
input n_1487;
input n_40;
input n_1864;
input n_1028;
input n_1601;
input n_781;
input n_474;
input n_542;
input n_463;
input n_1546;
input n_595;
input n_502;
input n_466;
input n_2612;
input n_420;
input n_1337;
input n_1495;
input n_632;
input n_699;
input n_979;
input n_1515;
input n_1627;
input n_1245;
input n_846;
input n_2427;
input n_2438;
input n_2505;
input n_1673;
input n_465;
input n_76;
input n_362;
input n_1321;
input n_170;
input n_1975;
input n_27;
input n_2296;
input n_2070;
input n_161;
input n_273;
input n_1937;
input n_585;
input n_2112;
input n_1739;
input n_270;
input n_616;
input n_2278;
input n_81;
input n_2594;
input n_2394;
input n_1914;
input n_2135;
input n_2335;
input n_745;
input n_2381;
input n_1654;
input n_2569;
input n_2349;
input n_1103;
input n_648;
input n_1379;
input n_2734;
input n_312;
input n_2196;
input n_2170;
input n_1076;
input n_1091;
input n_1408;
input n_494;
input n_1761;
input n_641;
input n_730;
input n_2036;
input n_1325;
input n_1595;
input n_2161;
input n_354;
input n_575;
input n_480;
input n_425;
input n_795;
input n_2404;
input n_2083;
input n_695;
input n_180;
input n_656;
input n_1606;
input n_2503;
input n_1220;
input n_37;
input n_1694;
input n_1540;
input n_2485;
input n_229;
input n_1936;
input n_1956;
input n_437;
input n_1642;
input n_2279;
input n_2655;
input n_2027;
input n_60;
input n_403;
input n_453;
input n_2642;
input n_1130;
input n_720;
input n_0;
input n_2500;
input n_2366;
input n_1918;
input n_1526;
input n_863;
input n_2210;
input n_805;
input n_1604;
input n_1275;
input n_2513;
input n_2525;
input n_2695;
input n_1764;
input n_113;
input n_712;
input n_2414;
input n_246;
input n_1583;
input n_2426;
input n_1042;
input n_1402;
input n_269;
input n_2049;
input n_2273;
input n_285;
input n_412;
input n_2719;
input n_1493;
input n_657;
input n_644;
input n_1741;
input n_2229;
input n_1160;
input n_1397;
input n_491;
input n_1258;
input n_1074;
input n_2004;
input n_1621;
input n_2708;
input n_2113;
input n_251;
input n_160;
input n_566;
input n_565;
input n_2586;
input n_1448;
input n_2225;
input n_1507;
input n_1398;
input n_2383;
input n_1879;
input n_597;
input n_1996;
input n_1181;
input n_1505;
input n_1634;
input n_1196;
input n_2019;
input n_651;
input n_1340;
input n_2274;
input n_334;
input n_811;
input n_1558;
input n_807;
input n_2166;
input n_835;
input n_175;
input n_666;
input n_262;
input n_1433;
input n_1704;
input n_2256;
input n_99;
input n_1254;
input n_1026;
input n_2026;
input n_1969;
input n_1234;
input n_2109;
input n_319;
input n_364;
input n_1138;
input n_927;
input n_20;
input n_1089;
input n_2013;
input n_1990;
input n_2044;
input n_2689;
input n_1004;
input n_1186;
input n_1032;
input n_242;
input n_2614;
input n_2511;
input n_1681;
input n_2010;
input n_1018;
input n_2242;
input n_2247;
input n_2752;
input n_1693;
input n_438;
input n_2599;
input n_713;
input n_2704;
input n_904;
input n_1588;
input n_1622;
input n_2237;
input n_166;
input n_1180;
input n_1827;
input n_2524;
input n_1271;
input n_2802;
input n_533;
input n_1542;
input n_1251;
input n_278;
input n_2728;
input n_2268;

output n_13034;

wire n_6643;
wire n_6122;
wire n_10564;
wire n_7981;
wire n_9936;
wire n_4706;
wire n_5567;
wire n_12148;
wire n_9194;
wire n_3241;
wire n_3006;
wire n_12407;
wire n_6579;
wire n_9325;
wire n_7164;
wire n_10794;
wire n_5287;
wire n_6546;
wire n_12872;
wire n_9655;
wire n_2899;
wire n_5484;
wire n_3619;
wire n_10515;
wire n_3541;
wire n_3622;
wire n_11207;
wire n_11326;
wire n_5978;
wire n_8174;
wire n_5161;
wire n_5776;
wire n_6551;
wire n_5512;
wire n_10793;
wire n_5207;
wire n_12853;
wire n_9044;
wire n_6786;
wire n_12327;
wire n_7206;
wire n_7303;
wire n_10552;
wire n_9083;
wire n_12215;
wire n_4963;
wire n_4240;
wire n_4508;
wire n_8363;
wire n_9408;
wire n_12975;
wire n_11802;
wire n_7710;
wire n_8383;
wire n_5035;
wire n_5282;
wire n_10885;
wire n_2843;
wire n_11583;
wire n_11349;
wire n_3615;
wire n_8328;
wire n_7461;
wire n_12641;
wire n_9331;
wire n_6649;
wire n_8060;
wire n_7154;
wire n_8551;
wire n_3202;
wire n_8002;
wire n_12924;
wire n_4977;
wire n_3813;
wire n_10108;
wire n_8594;
wire n_6810;
wire n_7660;
wire n_12071;
wire n_6276;
wire n_11016;
wire n_6072;
wire n_3341;
wire n_12738;
wire n_3587;
wire n_4128;
wire n_8976;
wire n_3445;
wire n_4145;
wire n_8617;
wire n_5033;
wire n_3785;
wire n_10883;
wire n_7686;
wire n_4211;
wire n_10117;
wire n_12139;
wire n_9846;
wire n_12328;
wire n_8603;
wire n_7024;
wire n_12493;
wire n_3448;
wire n_7205;
wire n_9204;
wire n_6742;
wire n_9769;
wire n_3019;
wire n_11342;
wire n_9312;
wire n_10363;
wire n_8319;
wire n_6694;
wire n_3776;
wire n_9610;
wire n_7616;
wire n_4517;
wire n_7486;
wire n_4425;
wire n_4950;
wire n_4988;
wire n_11450;
wire n_8244;
wire n_12028;
wire n_9273;
wire n_12357;
wire n_4615;
wire n_6580;
wire n_6090;
wire n_12515;
wire n_7010;
wire n_11678;
wire n_5480;
wire n_6549;
wire n_8105;
wire n_6913;
wire n_7867;
wire n_10756;
wire n_3010;
wire n_7315;
wire n_11801;
wire n_11653;
wire n_7004;
wire n_8961;
wire n_4131;
wire n_7772;
wire n_10761;
wire n_11299;
wire n_5402;
wire n_5851;
wire n_3188;
wire n_5509;
wire n_9773;
wire n_8574;
wire n_3403;
wire n_11089;
wire n_11077;
wire n_3624;
wire n_8864;
wire n_3461;
wire n_12861;
wire n_9173;
wire n_12709;
wire n_3082;
wire n_7641;
wire n_11296;
wire n_3796;
wire n_5154;
wire n_3283;
wire n_9363;
wire n_8681;
wire n_7468;
wire n_9796;
wire n_5469;
wire n_6431;
wire n_11800;
wire n_12012;
wire n_12462;
wire n_5744;
wire n_12266;
wire n_9049;
wire n_3340;
wire n_11947;
wire n_3277;
wire n_5453;
wire n_11917;
wire n_7861;
wire n_9907;
wire n_4499;
wire n_4927;
wire n_8413;
wire n_9738;
wire n_5202;
wire n_5648;
wire n_10745;
wire n_7667;
wire n_6931;
wire n_9539;
wire n_8114;
wire n_9811;
wire n_12970;
wire n_6618;
wire n_6408;
wire n_9993;
wire n_9208;
wire n_3214;
wire n_10421;
wire n_7523;
wire n_4311;
wire n_3631;
wire n_8706;
wire n_3806;
wire n_4691;
wire n_13000;
wire n_5922;
wire n_8158;
wire n_11594;
wire n_12100;
wire n_6698;
wire n_4678;
wire n_9500;
wire n_8104;
wire n_10399;
wire n_5848;
wire n_10420;
wire n_12575;
wire n_11635;
wire n_5406;
wire n_12501;
wire n_6085;
wire n_3947;
wire n_3490;
wire n_12819;
wire n_7421;
wire n_7306;
wire n_11505;
wire n_8819;
wire n_10535;
wire n_6214;
wire n_7493;
wire n_10360;
wire n_3868;
wire n_12027;
wire n_3183;
wire n_3437;
wire n_9420;
wire n_7804;
wire n_8089;
wire n_12111;
wire n_12075;
wire n_12078;
wire n_9557;
wire n_3353;
wire n_4203;
wire n_3687;
wire n_9382;
wire n_5241;
wire n_12175;
wire n_6939;
wire n_12604;
wire n_7528;
wire n_11615;
wire n_10307;
wire n_10781;
wire n_3156;
wire n_8290;
wire n_8262;
wire n_9206;
wire n_11507;
wire n_3376;
wire n_7562;
wire n_12626;
wire n_11497;
wire n_5037;
wire n_9388;
wire n_10193;
wire n_11541;
wire n_4468;
wire n_5661;
wire n_6991;
wire n_3653;
wire n_5562;
wire n_8885;
wire n_9772;
wire n_10437;
wire n_12142;
wire n_10430;
wire n_3702;
wire n_8147;
wire n_4976;
wire n_6586;
wire n_11111;
wire n_11354;
wire n_5008;
wire n_10177;
wire n_2976;
wire n_3876;
wire n_8310;
wire n_11052;
wire n_4811;
wire n_5398;
wire n_6096;
wire n_6707;
wire n_10175;
wire n_5852;
wire n_12767;
wire n_3420;
wire n_6920;
wire n_6868;
wire n_9311;
wire n_12754;
wire n_5144;
wire n_9422;
wire n_4758;
wire n_3361;
wire n_10672;
wire n_9040;
wire n_9795;
wire n_8380;
wire n_9027;
wire n_8962;
wire n_12225;
wire n_7402;
wire n_4255;
wire n_5577;
wire n_10626;
wire n_7592;
wire n_4484;
wire n_3668;
wire n_11316;
wire n_7152;
wire n_6512;
wire n_9966;
wire n_11272;
wire n_4237;
wire n_2934;
wire n_3550;
wire n_8126;
wire n_5689;
wire n_10392;
wire n_5894;
wire n_12670;
wire n_12152;
wire n_7801;
wire n_7992;
wire n_11588;
wire n_11689;
wire n_9161;
wire n_10231;
wire n_7463;
wire n_12101;
wire n_3418;
wire n_8556;
wire n_10316;
wire n_9369;
wire n_4901;
wire n_9033;
wire n_8305;
wire n_10683;
wire n_6725;
wire n_7613;
wire n_2859;
wire n_9429;
wire n_3395;
wire n_12576;
wire n_7083;
wire n_4917;
wire n_7086;
wire n_7349;
wire n_10514;
wire n_6464;
wire n_2863;
wire n_8317;
wire n_10730;
wire n_10958;
wire n_10562;
wire n_11273;
wire n_11962;
wire n_8653;
wire n_7647;
wire n_5825;
wire n_7779;
wire n_7712;
wire n_2968;
wire n_11303;
wire n_7316;
wire n_6820;
wire n_12224;
wire n_3593;
wire n_5343;
wire n_9780;
wire n_10252;
wire n_4421;
wire n_10438;
wire n_9824;
wire n_6098;
wire n_12237;
wire n_7019;
wire n_12751;
wire n_6686;
wire n_11664;
wire n_10523;
wire n_4836;
wire n_11720;
wire n_5062;
wire n_4020;
wire n_10202;
wire n_11398;
wire n_11659;
wire n_3915;
wire n_4469;
wire n_4414;
wire n_6561;
wire n_6584;
wire n_7452;
wire n_5184;
wire n_7956;
wire n_8939;
wire n_4532;
wire n_12824;
wire n_3339;
wire n_9489;
wire n_8604;
wire n_3735;
wire n_3349;
wire n_7323;
wire n_11365;
wire n_12269;
wire n_7195;
wire n_6701;
wire n_10988;
wire n_7478;
wire n_3007;
wire n_11836;
wire n_6769;
wire n_7683;
wire n_6592;
wire n_11150;
wire n_5686;
wire n_12298;
wire n_12019;
wire n_5463;
wire n_5236;
wire n_3310;
wire n_3487;
wire n_6191;
wire n_6062;
wire n_7903;
wire n_11003;
wire n_12299;
wire n_9625;
wire n_8440;
wire n_3983;
wire n_10980;
wire n_4405;
wire n_5433;
wire n_10367;
wire n_8525;
wire n_4195;
wire n_8416;
wire n_4969;
wire n_4504;
wire n_9570;
wire n_12232;
wire n_9368;
wire n_8064;
wire n_5909;
wire n_7575;
wire n_8879;
wire n_10664;
wire n_4408;
wire n_9115;
wire n_9694;
wire n_9367;
wire n_4531;
wire n_6043;
wire n_11520;
wire n_12812;
wire n_2987;
wire n_6271;
wire n_7171;
wire n_4567;
wire n_11099;
wire n_7701;
wire n_4164;
wire n_5315;
wire n_4234;
wire n_4130;
wire n_11859;
wire n_8931;
wire n_3611;
wire n_2862;
wire n_5348;
wire n_5055;
wire n_8214;
wire n_9072;
wire n_6793;
wire n_7873;
wire n_9612;
wire n_3187;
wire n_12777;
wire n_2828;
wire n_9971;
wire n_8729;
wire n_7127;
wire n_5397;
wire n_4471;
wire n_6550;
wire n_5031;
wire n_10575;
wire n_11746;
wire n_3392;
wire n_3975;
wire n_4444;
wire n_5709;
wire n_3430;
wire n_7568;
wire n_10803;
wire n_3208;
wire n_6021;
wire n_9720;
wire n_3331;
wire n_4983;
wire n_5695;
wire n_7814;
wire n_9213;
wire n_2911;
wire n_10187;
wire n_10400;
wire n_11330;
wire n_10778;
wire n_4916;
wire n_5860;
wire n_6926;
wire n_11121;
wire n_3649;
wire n_9607;
wire n_4302;
wire n_7589;
wire n_6928;
wire n_7965;
wire n_5862;
wire n_6304;
wire n_8228;
wire n_8210;
wire n_5189;
wire n_10586;
wire n_6956;
wire n_10040;
wire n_5381;
wire n_4786;
wire n_3257;
wire n_7026;
wire n_4160;
wire n_6782;
wire n_5854;
wire n_11911;
wire n_5516;
wire n_4051;
wire n_9554;
wire n_9262;
wire n_11599;
wire n_12412;
wire n_3009;
wire n_8387;
wire n_7002;
wire n_12782;
wire n_3981;
wire n_8898;
wire n_8410;
wire n_7141;
wire n_10935;
wire n_5936;
wire n_6126;
wire n_9761;
wire n_12284;
wire n_12612;
wire n_11102;
wire n_8795;
wire n_9649;
wire n_10164;
wire n_10269;
wire n_11039;
wire n_8501;
wire n_12567;
wire n_10401;
wire n_6027;
wire n_6598;
wire n_9254;
wire n_9529;
wire n_11535;
wire n_3224;
wire n_4647;
wire n_3752;
wire n_6342;
wire n_6638;
wire n_10651;
wire n_7308;
wire n_5254;
wire n_12180;
wire n_3526;
wire n_6900;
wire n_8953;
wire n_12731;
wire n_9726;
wire n_11686;
wire n_8823;
wire n_12153;
wire n_3790;
wire n_10851;
wire n_7264;
wire n_3491;
wire n_11730;
wire n_12608;
wire n_7457;
wire n_4613;
wire n_12383;
wire n_7718;
wire n_10918;
wire n_4649;
wire n_7617;
wire n_9197;
wire n_6269;
wire n_8843;
wire n_11942;
wire n_5615;
wire n_4795;
wire n_12057;
wire n_2891;
wire n_5902;
wire n_4028;
wire n_7768;
wire n_5479;
wire n_10964;
wire n_3819;
wire n_7974;
wire n_12902;
wire n_9106;
wire n_6013;
wire n_7357;
wire n_5083;
wire n_8247;
wire n_9564;
wire n_6927;
wire n_9627;
wire n_7975;
wire n_10864;
wire n_6503;
wire n_5888;
wire n_8172;
wire n_4186;
wire n_8941;
wire n_8940;
wire n_9739;
wire n_7310;
wire n_10598;
wire n_11835;
wire n_12070;
wire n_13021;
wire n_4731;
wire n_11444;
wire n_3747;
wire n_5698;
wire n_5592;
wire n_7521;
wire n_12430;
wire n_4618;
wire n_3346;
wire n_7593;
wire n_4742;
wire n_6256;
wire n_7716;
wire n_2876;
wire n_4099;
wire n_7406;
wire n_7600;
wire n_3484;
wire n_3620;
wire n_10223;
wire n_11353;
wire n_5870;
wire n_9812;
wire n_4295;
wire n_11823;
wire n_9646;
wire n_5303;
wire n_10451;
wire n_10553;
wire n_12718;
wire n_12393;
wire n_10201;
wire n_12249;
wire n_7076;
wire n_11814;
wire n_12719;
wire n_8780;
wire n_10215;
wire n_11205;
wire n_9465;
wire n_12932;
wire n_9928;
wire n_4694;
wire n_8456;
wire n_9970;
wire n_4533;
wire n_3038;
wire n_11138;
wire n_5081;
wire n_9894;
wire n_10100;
wire n_10278;
wire n_5124;
wire n_10436;
wire n_3068;
wire n_2871;
wire n_5807;
wire n_5863;
wire n_5943;
wire n_4244;
wire n_4603;
wire n_2943;
wire n_11048;
wire n_4254;
wire n_3143;
wire n_9129;
wire n_3168;
wire n_6982;
wire n_4697;
wire n_7286;
wire n_7137;
wire n_12625;
wire n_9957;
wire n_10915;
wire n_4190;
wire n_3994;
wire n_9558;
wire n_11292;
wire n_11487;
wire n_11753;
wire n_4810;
wire n_7848;
wire n_6727;
wire n_3317;
wire n_11782;
wire n_8218;
wire n_10689;
wire n_9267;
wire n_12371;
wire n_7539;
wire n_8769;
wire n_7229;
wire n_4391;
wire n_10538;
wire n_8514;
wire n_5954;
wire n_3263;
wire n_11865;
wire n_4157;
wire n_4283;
wire n_8368;
wire n_4681;
wire n_12163;
wire n_8334;
wire n_12258;
wire n_9918;
wire n_4638;
wire n_8159;
wire n_3455;
wire n_6097;
wire n_10773;
wire n_11397;
wire n_8639;
wire n_10621;
wire n_5047;
wire n_3452;
wire n_11600;
wire n_12516;
wire n_5346;
wire n_5517;
wire n_7125;
wire n_6677;
wire n_7797;
wire n_4707;
wire n_8216;
wire n_4527;
wire n_5109;
wire n_6624;
wire n_7121;
wire n_10924;
wire n_11844;
wire n_10874;
wire n_7869;
wire n_6466;
wire n_12871;
wire n_10942;
wire n_12602;
wire n_12295;
wire n_4156;
wire n_9956;
wire n_4848;
wire n_9095;
wire n_9715;
wire n_2937;
wire n_6008;
wire n_12198;
wire n_3095;
wire n_8337;
wire n_11201;
wire n_8257;
wire n_11781;
wire n_10292;
wire n_7983;
wire n_11550;
wire n_12077;
wire n_7781;
wire n_8125;
wire n_12166;
wire n_12786;
wire n_5624;
wire n_4918;
wire n_5714;
wire n_5806;
wire n_3856;
wire n_9246;
wire n_7624;
wire n_10653;
wire n_9683;
wire n_11945;
wire n_12117;
wire n_12110;
wire n_2914;
wire n_4898;
wire n_12216;
wire n_2869;
wire n_6221;
wire n_7160;
wire n_4002;
wire n_8063;
wire n_9931;
wire n_6805;
wire n_12098;
wire n_6185;
wire n_5010;
wire n_7762;
wire n_8731;
wire n_3623;
wire n_2846;
wire n_12102;
wire n_13009;
wire n_2925;
wire n_3773;
wire n_8950;
wire n_3918;
wire n_10624;
wire n_12802;
wire n_6568;
wire n_2857;
wire n_9011;
wire n_5358;
wire n_9899;
wire n_4528;
wire n_3932;
wire n_8295;
wire n_12570;
wire n_4619;
wire n_4673;
wire n_6004;
wire n_6351;
wire n_7552;
wire n_8059;
wire n_4822;
wire n_3516;
wire n_8995;
wire n_8146;
wire n_3797;
wire n_11502;
wire n_6901;
wire n_8082;
wire n_11965;
wire n_2947;
wire n_11997;
wire n_9094;
wire n_5580;
wire n_4299;
wire n_5937;
wire n_4801;
wire n_7183;
wire n_12456;
wire n_11424;
wire n_6411;
wire n_3515;
wire n_8339;
wire n_2886;
wire n_3287;
wire n_11816;
wire n_9195;
wire n_3378;
wire n_7746;
wire n_5435;
wire n_12768;
wire n_10867;
wire n_11361;
wire n_10701;
wire n_11062;
wire n_6873;
wire n_4279;
wire n_4769;
wire n_4632;
wire n_10741;
wire n_5373;
wire n_5745;
wire n_8032;
wire n_7139;
wire n_12710;
wire n_12483;
wire n_8640;
wire n_4294;
wire n_9332;
wire n_10016;
wire n_10070;
wire n_5279;
wire n_4232;
wire n_4125;
wire n_8351;
wire n_4949;
wire n_10190;
wire n_2941;
wire n_11499;
wire n_8196;
wire n_11580;
wire n_12128;
wire n_6594;
wire n_5493;
wire n_4790;
wire n_7857;
wire n_9054;
wire n_10812;
wire n_10150;
wire n_9460;
wire n_9638;
wire n_12682;
wire n_13028;
wire n_6387;
wire n_12389;
wire n_7223;
wire n_7890;
wire n_2952;
wire n_12464;
wire n_4847;
wire n_6179;
wire n_9281;
wire n_7338;
wire n_5321;
wire n_3058;
wire n_10134;
wire n_11379;
wire n_7964;
wire n_5096;
wire n_9740;
wire n_4365;
wire n_9475;
wire n_8865;
wire n_9661;
wire n_10861;
wire n_6019;
wire n_12313;
wire n_12147;
wire n_11070;
wire n_9190;
wire n_6222;
wire n_7165;
wire n_8110;
wire n_3505;
wire n_11245;
wire n_10635;
wire n_12874;
wire n_6223;
wire n_8838;
wire n_8475;
wire n_4610;
wire n_6435;
wire n_12909;
wire n_9143;
wire n_3730;
wire n_4489;
wire n_12990;
wire n_7235;
wire n_5210;
wire n_6976;
wire n_4967;
wire n_6486;
wire n_8488;
wire n_11286;
wire n_5657;
wire n_6889;
wire n_6083;
wire n_4992;
wire n_8766;
wire n_6844;
wire n_3001;
wire n_7795;
wire n_8969;
wire n_12240;
wire n_11631;
wire n_7404;
wire n_3945;
wire n_9891;
wire n_10555;
wire n_4542;
wire n_6295;
wire n_10897;
wire n_11147;
wire n_3597;
wire n_9087;
wire n_11700;
wire n_9804;
wire n_10287;
wire n_8087;
wire n_8119;
wire n_10135;
wire n_9321;
wire n_7885;
wire n_12468;
wire n_4198;
wire n_2897;
wire n_2909;
wire n_5857;
wire n_10983;
wire n_8173;
wire n_4534;
wire n_4500;
wire n_11833;
wire n_9800;
wire n_7437;
wire n_5014;
wire n_11053;
wire n_6241;
wire n_8420;
wire n_3185;
wire n_6087;
wire n_8019;
wire n_9186;
wire n_3523;
wire n_9951;
wire n_2829;
wire n_4597;
wire n_6846;
wire n_4329;
wire n_4087;
wire n_9243;
wire n_11335;
wire n_3811;
wire n_3200;
wire n_5756;
wire n_12294;
wire n_11336;
wire n_11057;
wire n_11247;
wire n_6041;
wire n_7822;
wire n_12186;
wire n_8851;
wire n_6994;
wire n_10987;
wire n_4257;
wire n_3453;
wire n_7449;
wire n_11262;
wire n_7329;
wire n_9359;
wire n_5708;
wire n_10402;
wire n_3213;
wire n_8687;
wire n_6790;
wire n_12860;
wire n_10001;
wire n_10666;
wire n_3077;
wire n_7194;
wire n_11363;
wire n_6273;
wire n_3474;
wire n_11783;
wire n_8740;
wire n_11661;
wire n_11026;
wire n_3984;
wire n_6807;
wire n_11889;
wire n_5927;
wire n_10189;
wire n_12939;
wire n_9879;
wire n_4665;
wire n_8221;
wire n_8468;
wire n_7708;
wire n_7696;
wire n_11756;
wire n_3679;
wire n_11232;
wire n_11419;
wire n_3422;
wire n_3888;
wire n_5638;
wire n_9975;
wire n_10997;
wire n_7115;
wire n_9335;
wire n_4189;
wire n_5670;
wire n_9171;
wire n_12778;
wire n_8815;
wire n_9942;
wire n_11081;
wire n_3707;
wire n_12813;
wire n_11407;
wire n_5584;
wire n_8952;
wire n_3429;
wire n_11654;
wire n_3849;
wire n_3946;
wire n_9247;
wire n_9933;
wire n_5965;
wire n_12907;
wire n_3229;
wire n_4463;
wire n_7958;
wire n_10209;
wire n_8128;
wire n_11519;
wire n_4687;
wire n_5751;
wire n_10434;
wire n_5664;
wire n_12011;
wire n_9441;
wire n_11668;
wire n_11913;
wire n_4670;
wire n_11978;
wire n_4084;
wire n_4703;
wire n_10829;
wire n_5641;
wire n_8667;
wire n_6218;
wire n_4037;
wire n_8863;
wire n_7281;
wire n_10233;
wire n_2922;
wire n_11810;
wire n_3275;
wire n_3499;
wire n_8106;
wire n_9362;
wire n_10690;
wire n_10311;
wire n_3421;
wire n_6824;
wire n_11198;
wire n_11767;
wire n_8717;
wire n_6189;
wire n_3618;
wire n_11595;
wire n_9216;
wire n_11168;
wire n_8299;
wire n_5262;
wire n_9200;
wire n_6993;
wire n_6037;
wire n_3683;
wire n_7245;
wire n_3642;
wire n_11872;
wire n_5963;
wire n_3286;
wire n_3808;
wire n_5980;
wire n_8892;
wire n_11235;
wire n_12007;
wire n_10146;
wire n_4763;
wire n_3590;
wire n_9067;
wire n_12712;
wire n_5310;
wire n_9152;
wire n_12846;
wire n_8287;
wire n_11906;
wire n_4594;
wire n_6153;
wire n_9074;
wire n_7989;
wire n_10790;
wire n_3424;
wire n_5970;
wire n_6418;
wire n_12908;
wire n_6564;
wire n_3583;
wire n_8657;
wire n_12505;
wire n_12747;
wire n_3560;
wire n_12577;
wire n_4076;
wire n_4714;
wire n_12426;
wire n_3215;
wire n_5146;
wire n_4776;
wire n_11122;
wire n_9287;
wire n_4102;
wire n_8197;
wire n_9511;
wire n_10052;
wire n_8081;
wire n_7192;
wire n_3171;
wire n_12309;
wire n_6671;
wire n_10407;
wire n_10449;
wire n_11324;
wire n_12164;
wire n_6591;
wire n_6266;
wire n_10950;
wire n_7161;
wire n_11566;
wire n_7580;
wire n_7153;
wire n_9880;
wire n_10072;
wire n_9843;
wire n_5213;
wire n_3020;
wire n_3677;
wire n_8609;
wire n_11869;
wire n_5441;
wire n_3462;
wire n_6517;
wire n_3468;
wire n_2910;
wire n_11579;
wire n_8559;
wire n_7350;
wire n_10838;
wire n_5690;
wire n_12140;
wire n_10369;
wire n_6967;
wire n_5885;
wire n_10920;
wire n_9248;
wire n_6433;
wire n_10321;
wire n_12178;
wire n_3546;
wire n_7535;
wire n_6893;
wire n_9128;
wire n_13003;
wire n_8452;
wire n_10506;
wire n_4443;
wire n_5461;
wire n_11082;
wire n_4507;
wire n_7178;
wire n_7480;
wire n_10224;
wire n_7632;
wire n_4575;
wire n_3012;
wire n_12554;
wire n_10671;
wire n_8771;
wire n_8140;
wire n_8476;
wire n_9528;
wire n_3244;
wire n_12912;
wire n_6501;
wire n_8981;
wire n_10157;
wire n_12200;
wire n_11529;
wire n_9507;
wire n_6028;
wire n_3130;
wire n_3822;
wire n_3569;
wire n_5629;
wire n_4452;
wire n_4348;
wire n_5634;
wire n_5430;
wire n_9533;
wire n_12611;
wire n_5362;
wire n_8137;
wire n_6709;
wire n_4355;
wire n_3494;
wire n_12322;
wire n_8469;
wire n_10808;
wire n_6798;
wire n_12303;
wire n_12507;
wire n_5702;
wire n_5050;
wire n_5063;
wire n_5229;
wire n_7844;
wire n_5199;
wire n_3771;
wire n_11430;
wire n_3110;
wire n_11882;
wire n_12023;
wire n_9665;
wire n_4572;
wire n_3073;
wire n_8423;
wire n_12171;
wire n_12395;
wire n_12472;
wire n_12815;
wire n_5527;
wire n_6986;
wire n_11146;
wire n_8090;
wire n_5609;
wire n_12239;
wire n_5416;
wire n_10504;
wire n_4026;
wire n_11279;
wire n_4104;
wire n_10975;
wire n_4512;
wire n_3554;
wire n_4377;
wire n_5266;
wire n_7471;
wire n_3178;
wire n_9436;
wire n_5355;
wire n_9562;
wire n_6745;
wire n_11516;
wire n_11005;
wire n_8260;
wire n_4521;
wire n_8481;
wire n_4488;
wire n_5977;
wire n_6811;
wire n_3051;
wire n_6209;
wire n_6875;
wire n_10566;
wire n_3750;
wire n_3632;
wire n_11451;
wire n_4588;
wire n_11980;
wire n_11076;
wire n_7905;
wire n_3299;
wire n_6853;
wire n_4519;
wire n_12121;
wire n_5551;
wire n_7766;
wire n_7594;
wire n_3715;
wire n_7803;
wire n_7340;
wire n_10837;
wire n_6699;
wire n_7747;
wire n_6073;
wire n_8205;
wire n_5767;
wire n_8401;
wire n_6324;
wire n_3040;
wire n_12116;
wire n_8651;
wire n_5640;
wire n_10199;
wire n_13020;
wire n_8284;
wire n_10688;
wire n_12261;
wire n_3568;
wire n_9255;
wire n_10039;
wire n_8828;
wire n_5655;
wire n_5475;
wire n_11239;
wire n_12259;
wire n_12338;
wire n_3737;
wire n_6138;
wire n_7603;
wire n_8510;
wire n_8810;
wire n_9034;
wire n_3255;
wire n_9203;
wire n_9601;
wire n_5692;
wire n_4856;
wire n_7726;
wire n_10443;
wire n_11623;
wire n_12825;
wire n_7494;
wire n_2997;
wire n_5921;
wire n_12222;
wire n_8024;
wire n_9946;
wire n_4400;
wire n_5168;
wire n_3326;
wire n_10887;
wire n_9967;
wire n_6477;
wire n_10735;
wire n_10274;
wire n_8739;
wire n_3734;
wire n_8133;
wire n_8373;
wire n_8919;
wire n_11740;
wire n_4778;
wire n_10482;
wire n_6159;
wire n_11012;
wire n_9647;
wire n_6283;
wire n_7396;
wire n_9912;
wire n_5322;
wire n_11698;
wire n_7116;
wire n_12779;
wire n_4352;
wire n_7519;
wire n_10485;
wire n_4441;
wire n_6943;
wire n_9329;
wire n_4761;
wire n_6827;
wire n_10652;
wire n_12465;
wire n_6173;
wire n_8318;
wire n_8542;
wire n_11059;
wire n_4347;
wire n_4095;
wire n_3196;
wire n_8543;
wire n_8846;
wire n_10791;
wire n_4593;
wire n_6312;
wire n_3492;
wire n_11236;
wire n_4727;
wire n_4568;
wire n_12852;
wire n_5371;
wire n_12334;
wire n_4043;
wire n_3601;
wire n_6997;
wire n_5418;
wire n_11196;
wire n_11629;
wire n_10411;
wire n_12847;
wire n_7770;
wire n_10286;
wire n_12511;
wire n_11643;
wire n_2973;
wire n_7664;
wire n_10913;
wire n_5316;
wire n_9890;
wire n_3831;
wire n_10273;
wire n_3801;
wire n_6300;
wire n_9609;
wire n_9883;
wire n_10172;
wire n_7815;
wire n_12014;
wire n_9046;
wire n_9361;
wire n_8163;
wire n_11609;
wire n_6131;
wire n_4893;
wire n_5032;
wire n_10806;
wire n_6537;
wire n_5933;
wire n_12305;
wire n_4948;
wire n_4000;
wire n_9864;
wire n_3240;
wire n_4406;
wire n_12485;
wire n_7023;
wire n_8972;
wire n_9300;
wire n_12408;
wire n_12238;
wire n_7428;
wire n_5112;
wire n_10694;
wire n_5386;
wire n_11509;
wire n_6783;
wire n_11351;
wire n_9353;
wire n_4748;
wire n_9766;
wire n_7465;
wire n_3931;
wire n_4010;
wire n_11271;
wire n_8293;
wire n_2840;
wire n_5017;
wire n_9832;
wire n_10754;
wire n_2822;
wire n_4710;
wire n_12409;
wire n_11307;
wire n_4607;
wire n_5123;
wire n_9954;
wire n_4117;
wire n_8737;
wire n_3636;
wire n_7961;
wire n_10953;
wire n_11761;
wire n_7847;
wire n_9997;
wire n_10703;
wire n_11973;
wire n_3083;
wire n_4487;
wire n_5001;
wire n_9334;
wire n_7149;
wire n_8252;
wire n_6459;
wire n_9622;
wire n_10847;
wire n_11565;
wire n_2981;
wire n_11252;
wire n_8450;
wire n_4817;
wire n_7700;
wire n_9284;
wire n_3380;
wire n_5644;
wire n_3460;
wire n_3409;
wire n_9147;
wire n_8367;
wire n_3538;
wire n_12454;
wire n_10103;
wire n_8834;
wire n_6869;
wire n_8078;
wire n_10922;
wire n_10413;
wire n_11571;
wire n_4849;
wire n_10738;
wire n_12587;
wire n_4867;
wire n_5424;
wire n_7914;
wire n_3198;
wire n_10995;
wire n_7967;
wire n_9794;
wire n_11858;
wire n_4728;
wire n_7117;
wire n_9354;
wire n_8471;
wire n_11904;
wire n_12324;
wire n_4247;
wire n_4933;
wire n_12130;
wire n_6977;
wire n_4018;
wire n_8474;
wire n_12643;
wire n_3900;
wire n_7984;
wire n_10185;
wire n_11131;
wire n_4902;
wire n_11478;
wire n_4518;
wire n_10591;
wire n_11656;
wire n_12955;
wire n_4409;
wire n_4411;
wire n_11673;
wire n_11821;
wire n_8361;
wire n_6313;
wire n_3872;
wire n_11701;
wire n_10856;
wire n_4336;
wire n_6569;
wire n_4777;
wire n_9494;
wire n_6555;
wire n_9614;
wire n_11283;
wire n_12948;
wire n_9551;
wire n_3877;
wire n_6639;
wire n_7516;
wire n_2995;
wire n_5496;
wire n_3977;
wire n_3547;
wire n_9154;
wire n_10677;
wire n_7596;
wire n_4052;
wire n_5864;
wire n_6536;
wire n_3459;
wire n_4398;
wire n_3155;
wire n_8553;
wire n_6490;
wire n_8301;
wire n_10610;
wire n_6961;
wire n_4954;
wire n_12574;
wire n_12697;
wire n_9437;
wire n_5460;
wire n_7628;
wire n_9276;
wire n_4304;
wire n_6761;
wire n_9346;
wire n_11229;
wire n_3911;
wire n_5333;
wire n_6294;
wire n_11636;
wire n_6767;
wire n_8518;
wire n_4431;
wire n_7427;
wire n_4192;
wire n_6802;
wire n_7527;
wire n_12162;
wire n_5570;
wire n_3736;
wire n_6326;
wire n_9514;
wire n_4805;
wire n_11919;
wire n_9402;
wire n_10456;
wire n_12634;
wire n_11675;
wire n_10343;
wire n_4885;
wire n_7838;
wire n_8364;
wire n_7786;
wire n_5983;
wire n_9580;
wire n_9005;
wire n_5804;
wire n_12236;
wire n_7979;
wire n_6376;
wire n_3565;
wire n_6167;
wire n_8621;
wire n_8993;
wire n_7926;
wire n_4701;
wire n_5910;
wire n_7411;
wire n_12632;
wire n_7101;
wire n_12398;
wire n_5040;
wire n_6730;
wire n_6948;
wire n_10979;
wire n_10487;
wire n_10332;
wire n_9162;
wire n_9921;
wire n_9443;
wire n_6582;
wire n_8910;
wire n_7752;
wire n_9897;
wire n_11570;
wire n_10807;
wire n_6996;
wire n_11855;
wire n_9817;
wire n_11667;
wire n_9301;
wire n_6974;
wire n_7731;
wire n_8753;
wire n_6765;
wire n_7577;
wire n_8388;
wire n_9401;
wire n_8321;
wire n_6921;
wire n_11290;
wire n_8044;
wire n_8091;
wire n_8486;
wire n_7845;
wire n_3533;
wire n_10750;
wire n_2877;
wire n_12292;
wire n_7709;
wire n_9689;
wire n_4631;
wire n_3035;
wire n_11592;
wire n_11466;
wire n_5194;
wire n_9982;
wire n_6898;
wire n_12056;
wire n_6710;
wire n_5717;
wire n_7162;
wire n_5464;
wire n_6565;
wire n_8508;
wire n_12679;
wire n_8261;
wire n_12811;
wire n_12581;
wire n_5886;
wire n_7080;
wire n_9886;
wire n_7744;
wire n_12897;
wire n_8034;
wire n_8841;
wire n_10970;
wire n_3639;
wire n_7302;
wire n_6533;
wire n_12837;
wire n_4965;
wire n_3079;
wire n_10264;
wire n_6960;
wire n_8201;
wire n_6426;
wire n_6634;
wire n_7180;
wire n_5610;
wire n_5239;
wire n_6836;
wire n_11983;
wire n_12605;
wire n_11043;
wire n_4747;
wire n_5197;
wire n_8947;
wire n_9671;
wire n_6972;
wire n_2924;
wire n_9297;
wire n_8788;
wire n_10472;
wire n_7111;
wire n_7549;
wire n_4111;
wire n_5785;
wire n_4587;
wire n_3731;
wire n_11415;
wire n_2946;
wire n_6344;
wire n_5305;
wire n_5994;
wire n_4538;
wire n_6093;
wire n_10499;
wire n_8093;
wire n_11680;
wire n_6010;
wire n_7247;
wire n_11446;
wire n_9225;
wire n_8061;
wire n_6833;
wire n_11972;
wire n_5376;
wire n_11103;
wire n_7481;
wire n_10435;
wire n_12220;
wire n_10066;
wire n_5204;
wire n_7292;
wire n_10341;
wire n_12230;
wire n_4094;
wire n_3503;
wire n_8811;
wire n_12995;
wire n_7150;
wire n_2866;
wire n_3561;
wire n_7687;
wire n_10184;
wire n_10498;
wire n_12867;
wire n_8507;
wire n_9662;
wire n_10508;
wire n_2917;
wire n_9057;
wire n_3661;
wire n_3536;
wire n_12497;
wire n_4150;
wire n_4878;
wire n_12406;
wire n_6265;
wire n_8861;
wire n_11749;
wire n_6821;
wire n_8661;
wire n_11417;
wire n_3934;
wire n_8545;
wire n_12725;
wire n_4985;
wire n_6373;
wire n_6988;
wire n_8755;
wire n_5788;
wire n_11490;
wire n_12401;
wire n_8573;
wire n_8191;
wire n_11704;
wire n_3922;
wire n_3846;
wire n_7692;
wire n_5897;
wire n_6887;
wire n_10865;
wire n_11343;
wire n_9809;
wire n_12185;
wire n_3074;
wire n_8683;
wire n_10081;
wire n_8836;
wire n_6676;
wire n_3673;
wire n_6347;
wire n_6492;
wire n_7016;
wire n_12161;
wire n_3768;
wire n_2861;
wire n_9448;
wire n_3943;
wire n_8136;
wire n_8446;
wire n_9799;
wire n_7742;
wire n_10577;
wire n_9313;
wire n_8916;
wire n_3293;
wire n_7955;
wire n_5795;
wire n_7072;
wire n_5508;
wire n_10037;
wire n_12424;
wire n_5582;
wire n_10234;
wire n_4022;
wire n_7374;
wire n_7440;
wire n_9989;
wire n_11766;
wire n_4852;
wire n_7758;
wire n_11639;
wire n_7547;
wire n_12114;
wire n_11967;
wire n_4869;
wire n_9438;
wire n_4700;
wire n_7201;
wire n_4035;
wire n_11457;
wire n_3294;
wire n_4426;
wire n_10832;
wire n_12490;
wire n_10036;
wire n_12571;
wire n_11932;
wire n_3415;
wire n_5746;
wire n_2817;
wire n_5292;
wire n_3139;
wire n_10853;
wire n_12508;
wire n_12582;
wire n_6648;
wire n_7880;
wire n_12052;
wire n_4601;
wire n_8075;
wire n_8857;
wire n_11275;
wire n_4220;
wire n_8587;
wire n_12337;
wire n_9675;
wire n_10030;
wire n_5630;
wire n_9667;
wire n_10676;
wire n_11819;
wire n_8071;
wire n_3431;
wire n_10815;
wire n_12928;
wire n_3169;
wire n_3151;
wire n_11589;
wire n_11309;
wire n_12927;
wire n_3284;
wire n_3070;
wire n_4066;
wire n_2884;
wire n_11803;
wire n_7513;
wire n_11067;
wire n_12321;
wire n_4515;
wire n_4351;
wire n_11274;
wire n_5264;
wire n_9537;
wire n_11174;
wire n_3126;
wire n_7413;
wire n_4403;
wire n_10833;
wire n_11770;
wire n_7540;
wire n_8646;
wire n_4858;
wire n_4509;
wire n_3700;
wire n_9866;
wire n_5504;
wire n_8630;
wire n_7622;
wire n_9602;
wire n_7005;
wire n_11266;
wire n_11151;
wire n_4223;
wire n_7353;
wire n_6219;
wire n_10071;
wire n_9885;
wire n_12592;
wire n_12698;
wire n_8315;
wire n_6965;
wire n_9260;
wire n_5025;
wire n_2966;
wire n_8314;
wire n_6720;
wire n_12048;
wire n_8149;
wire n_6032;
wire n_11413;
wire n_8581;
wire n_7174;
wire n_8565;
wire n_6205;
wire n_6362;
wire n_6402;
wire n_4644;
wire n_7166;
wire n_4456;
wire n_5060;
wire n_7607;
wire n_8209;
wire n_9159;
wire n_5334;
wire n_4346;
wire n_7816;
wire n_9654;
wire n_3170;
wire n_8560;
wire n_7591;
wire n_5775;
wire n_8141;
wire n_3311;
wire n_7830;
wire n_3272;
wire n_7282;
wire n_6491;
wire n_8302;
wire n_10015;
wire n_9306;
wire n_2898;
wire n_7151;
wire n_11652;
wire n_11682;
wire n_12801;
wire n_6229;
wire n_11091;
wire n_11929;
wire n_9978;
wire n_5731;
wire n_8612;
wire n_5581;
wire n_3628;
wire n_3691;
wire n_6668;
wire n_7446;
wire n_10362;
wire n_4235;
wire n_7053;
wire n_3018;
wire n_8724;
wire n_11331;
wire n_11640;
wire n_5831;
wire n_10171;
wire n_12552;
wire n_7473;
wire n_4435;
wire n_10183;
wire n_10471;
wire n_2939;
wire n_8070;
wire n_6835;
wire n_6419;
wire n_6039;
wire n_12704;
wire n_11237;
wire n_3807;
wire n_11601;
wire n_11741;
wire n_5884;
wire n_9279;
wire n_8457;
wire n_4764;
wire n_5653;
wire n_8922;
wire n_8248;
wire n_7966;
wire n_9509;
wire n_6258;
wire n_10095;
wire n_10549;
wire n_7070;
wire n_5394;
wire n_11721;
wire n_6755;
wire n_9563;
wire n_7276;
wire n_7351;
wire n_12256;
wire n_7942;
wire n_10057;
wire n_4655;
wire n_12477;
wire n_3161;
wire n_4581;
wire n_12184;
wire n_11093;
wire n_12245;
wire n_6084;
wire n_10301;
wire n_4827;
wire n_9496;
wire n_8411;
wire n_12657;
wire n_12740;
wire n_9644;
wire n_7412;
wire n_7157;
wire n_6436;
wire n_7666;
wire n_12089;
wire n_6472;
wire n_3477;
wire n_5421;
wire n_8527;
wire n_7211;
wire n_10394;
wire n_10154;
wire n_4399;
wire n_11097;
wire n_11681;
wire n_6531;
wire n_5309;
wire n_7901;
wire n_8689;
wire n_11522;
wire n_9750;
wire n_4782;
wire n_9980;
wire n_10818;
wire n_12145;
wire n_8988;
wire n_11105;
wire n_4363;
wire n_2887;
wire n_12377;
wire n_12647;
wire n_12721;
wire n_4864;
wire n_9251;
wire n_10141;
wire n_7368;
wire n_8549;
wire n_12541;
wire n_3054;
wire n_4335;
wire n_6567;
wire n_5889;
wire n_12316;
wire n_11849;
wire n_6771;
wire n_11578;
wire n_10916;
wire n_10208;
wire n_6389;
wire n_10182;
wire n_9616;
wire n_12399;
wire n_8004;
wire n_10929;
wire n_8658;
wire n_9959;
wire n_8375;
wire n_10403;
wire n_5764;
wire n_10260;
wire n_5428;
wire n_6910;
wire n_9291;
wire n_9092;
wire n_10261;
wire n_6442;
wire n_12285;
wire n_3391;
wire n_6102;
wire n_8908;
wire n_4259;
wire n_5541;
wire n_10384;
wire n_6441;
wire n_5543;
wire n_10372;
wire n_9818;
wire n_10237;
wire n_9283;
wire n_5678;
wire n_5935;
wire n_4865;
wire n_11219;
wire n_4056;
wire n_4564;
wire n_3840;
wire n_7677;
wire n_5085;
wire n_3518;
wire n_8569;
wire n_2956;
wire n_3733;
wire n_8676;
wire n_10118;
wire n_5950;
wire n_12379;
wire n_7929;
wire n_10028;
wire n_12257;
wire n_3738;
wire n_10691;
wire n_8399;
wire n_5995;
wire n_12246;
wire n_11069;
wire n_6162;
wire n_5116;
wire n_4526;
wire n_3464;
wire n_6331;
wire n_6006;
wire n_8421;
wire n_3245;
wire n_4417;
wire n_6109;
wire n_11268;
wire n_6278;
wire n_9304;
wire n_12655;
wire n_6787;
wire n_10777;
wire n_11066;
wire n_6872;
wire n_4899;
wire n_6208;
wire n_6632;
wire n_9310;
wire n_5411;
wire n_7754;
wire n_4798;
wire n_9830;
wire n_9913;
wire n_11728;
wire n_7027;
wire n_3509;
wire n_3352;
wire n_8001;
wire n_5671;
wire n_3076;
wire n_8322;
wire n_12272;
wire n_6990;
wire n_12862;
wire n_8403;
wire n_3535;
wire n_6349;
wire n_3251;
wire n_11796;
wire n_2931;
wire n_7631;
wire n_6830;
wire n_8999;
wire n_12662;
wire n_8754;
wire n_5185;
wire n_7939;
wire n_8675;
wire n_7898;
wire n_10715;
wire n_12136;
wire n_6359;
wire n_9375;
wire n_3118;
wire n_8596;
wire n_10665;
wire n_10073;
wire n_10291;
wire n_3511;
wire n_8858;
wire n_8666;
wire n_11873;
wire n_3443;
wire n_8313;
wire n_7763;
wire n_10296;
wire n_7498;
wire n_3644;
wire n_5076;
wire n_3336;
wire n_3935;
wire n_7377;
wire n_11228;
wire n_3521;
wire n_8555;
wire n_5379;
wire n_3562;
wire n_3948;
wire n_4750;
wire n_12517;
wire n_6301;
wire n_12031;
wire n_11743;
wire n_2918;
wire n_3232;
wire n_10512;
wire n_8610;
wire n_12993;
wire n_10324;
wire n_12663;
wire n_7945;
wire n_5945;
wire n_11261;
wire n_9323;
wire n_6744;
wire n_2958;
wire n_4981;
wire n_3125;
wire n_3114;
wire n_9985;
wire n_10765;
wire n_12039;
wire n_3612;
wire n_11023;
wire n_2954;
wire n_8615;
wire n_11382;
wire n_4835;
wire n_5811;
wire n_4430;
wire n_6439;
wire n_10026;
wire n_8677;
wire n_9355;
wire n_8602;
wire n_9714;
wire n_12938;
wire n_7381;
wire n_10041;
wire n_5565;
wire n_4081;
wire n_7948;
wire n_4407;
wire n_3132;
wire n_7291;
wire n_8102;
wire n_9540;
wire n_3951;
wire n_4894;
wire n_13033;
wire n_9753;
wire n_5780;
wire n_8460;
wire n_9105;
wire n_5643;
wire n_3238;
wire n_11305;
wire n_3210;
wire n_10149;
wire n_12680;
wire n_13017;
wire n_11137;
wire n_11607;
wire n_5846;
wire n_7430;
wire n_9700;
wire n_3267;
wire n_12930;
wire n_4995;
wire n_8871;
wire n_10649;
wire n_9476;
wire n_12722;
wire n_7870;
wire n_9875;
wire n_11265;
wire n_10593;
wire n_12042;
wire n_5524;
wire n_8824;
wire n_3964;
wire n_3772;
wire n_10597;
wire n_9963;
wire n_6104;
wire n_4446;
wire n_3373;
wire n_6475;
wire n_3884;
wire n_12469;
wire n_8470;
wire n_9582;
wire n_12172;
wire n_11739;
wire n_10817;
wire n_6465;
wire n_10060;
wire n_9574;
wire n_12049;
wire n_3726;
wire n_6496;
wire n_11687;
wire n_9732;
wire n_11050;
wire n_2892;
wire n_12666;
wire n_2907;
wire n_8238;
wire n_9882;
wire n_12205;
wire n_6998;
wire n_10779;
wire n_6145;
wire n_3577;
wire n_11789;
wire n_8699;
wire n_2820;
wire n_7305;
wire n_10242;
wire n_10086;
wire n_9992;
wire n_12885;
wire n_11347;
wire n_4057;
wire n_4332;
wire n_4314;
wire n_3347;
wire n_7980;
wire n_3216;
wire n_3809;
wire n_11617;
wire n_7075;
wire n_7545;
wire n_11581;
wire n_7846;
wire n_10981;
wire n_6076;
wire n_4288;
wire n_3567;
wire n_8438;
wire n_6194;
wire n_10673;
wire n_10869;
wire n_7695;
wire n_5066;
wire n_12917;
wire n_3939;
wire n_6092;
wire n_7275;
wire n_5401;
wire n_6357;
wire n_5843;
wire n_4241;
wire n_3321;
wire n_8095;
wire n_12616;
wire n_7537;
wire n_3212;
wire n_3152;
wire n_10128;
wire n_10746;
wire n_12217;
wire n_12287;
wire n_12950;
wire n_7489;
wire n_5106;
wire n_10339;
wire n_11559;
wire n_5468;
wire n_11867;
wire n_2920;
wire n_4265;
wire n_6335;
wire n_8112;
wire n_12835;
wire n_5883;
wire n_6985;
wire n_8642;
wire n_5319;
wire n_7451;
wire n_8624;
wire n_6238;
wire n_9090;
wire n_11989;
wire n_12800;
wire n_10684;
wire n_10441;
wire n_12036;
wire n_12177;
wire n_9149;
wire n_10590;
wire n_9174;
wire n_12850;
wire n_11175;
wire n_12962;
wire n_3705;
wire n_6548;
wire n_4705;
wire n_3159;
wire n_5455;
wire n_8894;
wire n_9226;
wire n_6366;
wire n_3778;
wire n_5337;
wire n_5706;
wire n_9018;
wire n_3304;
wire n_12336;
wire n_10949;
wire n_3912;
wire n_7236;
wire n_9835;
wire n_12044;
wire n_11727;
wire n_12905;
wire n_4604;
wire n_7269;
wire n_8878;
wire n_5223;
wire n_10934;
wire n_5962;
wire n_3795;
wire n_5020;
wire n_6602;
wire n_4419;
wire n_4477;
wire n_6620;
wire n_3179;
wire n_6502;
wire n_9702;
wire n_3256;
wire n_7560;
wire n_11725;
wire n_10279;
wire n_11291;
wire n_7326;
wire n_7060;
wire n_7572;
wire n_3086;
wire n_6885;
wire n_12495;
wire n_2927;
wire n_4217;
wire n_4395;
wire n_8807;
wire n_12565;
wire n_2821;
wire n_9968;
wire n_5074;
wire n_5364;
wire n_9924;
wire n_6529;
wire n_8732;
wire n_8169;
wire n_11958;
wire n_3728;
wire n_8803;
wire n_3064;
wire n_9515;
wire n_3088;
wire n_8017;
wire n_10527;
wire n_5895;
wire n_4639;
wire n_6951;
wire n_3713;
wire n_8801;
wire n_3663;
wire n_12584;
wire n_5649;
wire n_5046;
wire n_5166;
wire n_7169;
wire n_12654;
wire n_6423;
wire n_9252;
wire n_3246;
wire n_10785;
wire n_7140;
wire n_7233;
wire n_10228;
wire n_11311;
wire n_12999;
wire n_5088;
wire n_6558;
wire n_8522;
wire n_5457;
wire n_7352;
wire n_7986;
wire n_9948;
wire n_7134;
wire n_5532;
wire n_12823;
wire n_11528;
wire n_12422;
wire n_6950;
wire n_7246;
wire n_12234;
wire n_6525;
wire n_7650;
wire n_3434;
wire n_9871;
wire n_11807;
wire n_6631;
wire n_6892;
wire n_11705;
wire n_8203;
wire n_7663;
wire n_9423;
wire n_11378;
wire n_11521;
wire n_11998;
wire n_4227;
wire n_4033;
wire n_4289;
wire n_9660;
wire n_9108;
wire n_11222;
wire n_4780;
wire n_8680;
wire n_9631;
wire n_10643;
wire n_7056;
wire n_4243;
wire n_4982;
wire n_12293;
wire n_10427;
wire n_3695;
wire n_4330;
wire n_6683;
wire n_8727;
wire n_10389;
wire n_10423;
wire n_6292;
wire n_5544;
wire n_3832;
wire n_9900;
wire n_11080;
wire n_7729;
wire n_3987;
wire n_7339;
wire n_5987;
wire n_7740;
wire n_6180;
wire n_5352;
wire n_5824;
wire n_4991;
wire n_11533;
wire n_12572;
wire n_5538;
wire n_8138;
wire n_6658;
wire n_10863;
wire n_6264;
wire n_9608;
wire n_9137;
wire n_6925;
wire n_8990;
wire n_5919;
wire n_10077;
wire n_12988;
wire n_8206;
wire n_9144;
wire n_12512;
wire n_7767;
wire n_11940;
wire n_8190;
wire n_6176;
wire n_9778;
wire n_8622;
wire n_5410;
wire n_11808;
wire n_3332;
wire n_7146;
wire n_8092;
wire n_3048;
wire n_3937;
wire n_10250;
wire n_6124;
wire n_7672;
wire n_8242;
wire n_4525;
wire n_12118;
wire n_12609;
wire n_3782;
wire n_7482;
wire n_12176;
wire n_9850;
wire n_6864;
wire n_9531;
wire n_7893;
wire n_2978;
wire n_4208;
wire n_8331;
wire n_7090;
wire n_3786;
wire n_11549;
wire n_7158;
wire n_7156;
wire n_2888;
wire n_5742;
wire n_5992;
wire n_3638;
wire n_8649;
wire n_8684;
wire n_6494;
wire n_5503;
wire n_8323;
wire n_10828;
wire n_4177;
wire n_12353;
wire n_6199;
wire n_11139;
wire n_8296;
wire n_3763;
wire n_9139;
wire n_11584;
wire n_9430;
wire n_10417;
wire n_5958;
wire n_6614;
wire n_7749;
wire n_3022;
wire n_11695;
wire n_7839;
wire n_4264;
wire n_8882;
wire n_10310;
wire n_12053;
wire n_7504;
wire n_10333;
wire n_3087;
wire n_10996;
wire n_12795;
wire n_9272;
wire n_3489;
wire n_8708;
wire n_10880;
wire n_12045;
wire n_7360;
wire n_10810;
wire n_12274;
wire n_7681;
wire n_10636;
wire n_12348;
wire n_8448;
wire n_8076;
wire n_7301;
wire n_9041;
wire n_11360;
wire n_5129;
wire n_11886;
wire n_9643;
wire n_8904;
wire n_7375;
wire n_7102;
wire n_5500;
wire n_8277;
wire n_3060;
wire n_11920;
wire n_4276;
wire n_7794;
wire n_11479;
wire n_12006;
wire n_7366;
wire n_8184;
wire n_5219;
wire n_5605;
wire n_3013;
wire n_9944;
wire n_5170;
wire n_5654;
wire n_7025;
wire n_8304;
wire n_5320;
wire n_10258;
wire n_3049;
wire n_6947;
wire n_11534;
wire n_8586;
wire n_5107;
wire n_9648;
wire n_5999;
wire n_4485;
wire n_8557;
wire n_9376;
wire n_10507;
wire n_8636;
wire n_7309;
wire n_4626;
wire n_6863;
wire n_9288;
wire n_10835;
wire n_6637;
wire n_6100;
wire n_7860;
wire n_6735;
wire n_9541;
wire n_9521;
wire n_8212;
wire n_4975;
wire n_6358;
wire n_9759;
wire n_12500;
wire n_12781;
wire n_7911;
wire n_11848;
wire n_8530;
wire n_9278;
wire n_9378;
wire n_11227;
wire n_8665;
wire n_5602;
wire n_9456;
wire n_9086;
wire n_3089;
wire n_7876;
wire n_6050;
wire n_11401;
wire n_9711;
wire n_8933;
wire n_7244;
wire n_7960;
wire n_5405;
wire n_12922;
wire n_5253;
wire n_3985;
wire n_9485;
wire n_4760;
wire n_11375;
wire n_4652;
wire n_4624;
wire n_9555;
wire n_10959;
wire n_7610;
wire n_12842;
wire n_9999;
wire n_11813;
wire n_9994;
wire n_10814;
wire n_5903;
wire n_6371;
wire n_8690;
wire n_8538;
wire n_7043;
wire n_12753;
wire n_3440;
wire n_10859;
wire n_6171;
wire n_7751;
wire n_8643;
wire n_6510;
wire n_4569;
wire n_6468;
wire n_9142;
wire n_9613;
wire n_4897;
wire n_11134;
wire n_9440;
wire n_3542;
wire n_3436;
wire n_5491;
wire n_8825;
wire n_11716;
wire n_12366;
wire n_3940;
wire n_7788;
wire n_5842;
wire n_6352;
wire n_8300;
wire n_2985;
wire n_10531;
wire n_5722;
wire n_7534;
wire n_9462;
wire n_5636;
wire n_7719;
wire n_11357;
wire n_9202;
wire n_5065;
wire n_7287;
wire n_10699;
wire n_12208;
wire n_7032;
wire n_8451;
wire n_11386;
wire n_3637;
wire n_2842;
wire n_4523;
wire n_2868;
wire n_5492;
wire n_9237;
wire n_10941;
wire n_3141;
wire n_11448;
wire n_5084;
wire n_10567;
wire n_6850;
wire n_8435;
wire n_5667;
wire n_3164;
wire n_12122;
wire n_10770;
wire n_3570;
wire n_5260;
wire n_11693;
wire n_7119;
wire n_8835;
wire n_4919;
wire n_10714;
wire n_9788;
wire n_4025;
wire n_5328;
wire n_3936;
wire n_6354;
wire n_5918;
wire n_7634;
wire n_11755;
wire n_4503;
wire n_3507;
wire n_6959;
wire n_3821;
wire n_6909;
wire n_11221;
wire n_7851;
wire n_6332;
wire n_9807;
wire n_3367;
wire n_4464;
wire n_7006;
wire n_9573;
wire n_5877;
wire n_8963;
wire n_12351;
wire n_3096;
wire n_6306;
wire n_7682;
wire n_3496;
wire n_4114;
wire n_6434;
wire n_12040;
wire n_12443;
wire n_8713;
wire n_6751;
wire n_7068;
wire n_9392;
wire n_12133;
wire n_4556;
wire n_11084;
wire n_6322;
wire n_8668;
wire n_8353;
wire n_5454;
wire n_9390;
wire n_7704;
wire n_10326;
wire n_7773;
wire n_9416;
wire n_6667;
wire n_7526;
wire n_8817;
wire n_6530;
wire n_9518;
wire n_4089;
wire n_12491;
wire n_7376;
wire n_6156;
wire n_5913;
wire n_7268;
wire n_7044;
wire n_12452;
wire n_5621;
wire n_2919;
wire n_8213;
wire n_12233;
wire n_4327;
wire n_8591;
wire n_7973;
wire n_11885;
wire n_4218;
wire n_6429;
wire n_3146;
wire n_10966;
wire n_5165;
wire n_7239;
wire n_10047;
wire n_12633;
wire n_5573;
wire n_11253;
wire n_6405;
wire n_11551;
wire n_8532;
wire n_11380;
wire n_12936;
wire n_12035;
wire n_6613;
wire n_4353;
wire n_8043;
wire n_9196;
wire n_11172;
wire n_7969;
wire n_6248;
wire n_2921;
wire n_12915;
wire n_7821;
wire n_4990;
wire n_6088;
wire n_12275;
wire n_10784;
wire n_5529;
wire n_10248;
wire n_6894;
wire n_12947;
wire n_7267;
wire n_4959;
wire n_9589;
wire n_4161;
wire n_5800;
wire n_11539;
wire n_9898;
wire n_9373;
wire n_3992;
wire n_11976;
wire n_12308;
wire n_8606;
wire n_4103;
wire n_4466;
wire n_6204;
wire n_10351;
wire n_7915;
wire n_3625;
wire n_8121;
wire n_8868;
wire n_10408;
wire n_10921;
wire n_7387;
wire n_7431;
wire n_11731;
wire n_7654;
wire n_10551;
wire n_12760;
wire n_2945;
wire n_10656;
wire n_2837;
wire n_4844;
wire n_6296;
wire n_11531;
wire n_12318;
wire n_10313;
wire n_10639;
wire n_2979;
wire n_5257;
wire n_9983;
wire n_6290;
wire n_6288;
wire n_3655;
wire n_12700;
wire n_4688;
wire n_4765;
wire n_8276;
wire n_8718;
wire n_12364;
wire n_8182;
wire n_5645;
wire n_11392;
wire n_5180;
wire n_11204;
wire n_3640;
wire n_13025;
wire n_12985;
wire n_5779;
wire n_11627;
wire n_4388;
wire n_4206;
wire n_12340;
wire n_12478;
wire n_6140;
wire n_9039;
wire n_8359;
wire n_7441;
wire n_9849;
wire n_8597;
wire n_4738;
wire n_6211;
wire n_12788;
wire n_8562;
wire n_3909;
wire n_11485;
wire n_8211;
wire n_9962;
wire n_12826;
wire n_8430;
wire n_6307;
wire n_8007;
wire n_10871;
wire n_6164;
wire n_3207;
wire n_3944;
wire n_12752;
wire n_7394;
wire n_8600;
wire n_8311;
wire n_8943;
wire n_8441;
wire n_12194;
wire n_4434;
wire n_4837;
wire n_10747;
wire n_7022;
wire n_3042;
wire n_9829;
wire n_6860;
wire n_4219;
wire n_10459;
wire n_3659;
wire n_8978;
wire n_5012;
wire n_10121;
wire n_4620;
wire n_11387;
wire n_8198;
wire n_9988;
wire n_5697;
wire n_7188;
wire n_8526;
wire n_10705;
wire n_7573;
wire n_7879;
wire n_4438;
wire n_9848;
wire n_7087;
wire n_3510;
wire n_6147;
wire n_3218;
wire n_7985;
wire n_10334;
wire n_12689;
wire n_11691;
wire n_11358;
wire n_9045;
wire n_9466;
wire n_6515;
wire n_9348;
wire n_6011;
wire n_8278;
wire n_7722;
wire n_7935;
wire n_8592;
wire n_6645;
wire n_11128;
wire n_12271;
wire n_8226;
wire n_3150;
wire n_6984;
wire n_4325;
wire n_12843;
wire n_10716;
wire n_12273;
wire n_10235;
wire n_10090;
wire n_10153;
wire n_11649;
wire n_10937;
wire n_7193;
wire n_10018;
wire n_8987;
wire n_4133;
wire n_3775;
wire n_11489;
wire n_6897;
wire n_7256;
wire n_12391;
wire n_4184;
wire n_5203;
wire n_12420;
wire n_9071;
wire n_10568;
wire n_9356;
wire n_9464;
wire n_4481;
wire n_12314;
wire n_3416;
wire n_6460;
wire n_4379;
wire n_7128;
wire n_7595;
wire n_9239;
wire n_10053;
wire n_6183;
wire n_10051;
wire n_11373;
wire n_7522;
wire n_5882;
wire n_9606;
wire n_4030;
wire n_10359;
wire n_7881;
wire n_7436;
wire n_4490;
wire n_3138;
wire n_7380;
wire n_7012;
wire n_11216;
wire n_4397;
wire n_12356;
wire n_10998;
wire n_7502;
wire n_9492;
wire n_2928;
wire n_8960;
wire n_7335;
wire n_7103;
wire n_4820;
wire n_10648;
wire n_10151;
wire n_6246;
wire n_11194;
wire n_11804;
wire n_3770;
wire n_8025;
wire n_5094;
wire n_6383;
wire n_9031;
wire n_11107;
wire n_4938;
wire n_9717;
wire n_11434;
wire n_9516;
wire n_11645;
wire n_12073;
wire n_7020;
wire n_8434;
wire n_4179;
wire n_11244;
wire n_3469;
wire n_12848;
wire n_8175;
wire n_9693;
wire n_9991;
wire n_5336;
wire n_12155;
wire n_8850;
wire n_9103;
wire n_11254;
wire n_9477;
wire n_5672;
wire n_4641;
wire n_3220;
wire n_5548;
wire n_10253;
wire n_10822;
wire n_5601;
wire n_7248;
wire n_7662;
wire n_8895;
wire n_3855;
wire n_10589;
wire n_12390;
wire n_12160;
wire n_11297;
wire n_10349;
wire n_11991;
wire n_5339;
wire n_4931;
wire n_6099;
wire n_3158;
wire n_10946;
wire n_12150;
wire n_5693;
wire n_8046;
wire n_3113;
wire n_11173;
wire n_6904;
wire n_11183;
wire n_3760;
wire n_4078;
wire n_11922;
wire n_8867;
wire n_2856;
wire n_10473;
wire n_8239;
wire n_9599;
wire n_4146;
wire n_4360;
wire n_3666;
wire n_7825;
wire n_8183;
wire n_8924;
wire n_9001;
wire n_12840;
wire n_10893;
wire n_3828;
wire n_10218;
wire n_12964;
wire n_3288;
wire n_5514;
wire n_4404;
wire n_5091;
wire n_7533;
wire n_8578;
wire n_11548;
wire n_9777;
wire n_4787;
wire n_8848;
wire n_10903;
wire n_3667;
wire n_10458;
wire n_11868;
wire n_9222;
wire n_10148;
wire n_6626;
wire n_6563;
wire n_5486;
wire n_9366;
wire n_6611;
wire n_10775;
wire n_11248;
wire n_10543;
wire n_9449;
wire n_3703;
wire n_4903;
wire n_3558;
wire n_11114;
wire n_11260;
wire n_11901;
wire n_12994;
wire n_5599;
wire n_6116;
wire n_7186;
wire n_10337;
wire n_4356;
wire n_8230;
wire n_9869;
wire n_10478;
wire n_12252;
wire n_11981;
wire n_6819;
wire n_8725;
wire n_4432;
wire n_5251;
wire n_7936;
wire n_6473;
wire n_12951;
wire n_9741;
wire n_4291;
wire n_11956;
wire n_10956;
wire n_10637;
wire n_11805;
wire n_5403;
wire n_4386;
wire n_12131;
wire n_12280;
wire n_4149;
wire n_8391;
wire n_6310;
wire n_7840;
wire n_10698;
wire n_11381;
wire n_9397;
wire n_2982;
wire n_8202;
wire n_11775;
wire n_11797;
wire n_12453;
wire n_10834;
wire n_7429;
wire n_3545;
wire n_6688;
wire n_12557;
wire n_7906;
wire n_8948;
wire n_8678;
wire n_9754;
wire n_4019;
wire n_10783;
wire n_2900;
wire n_9179;
wire n_7148;
wire n_5782;
wire n_6714;
wire n_4637;
wire n_7017;
wire n_7250;
wire n_7462;
wire n_7658;
wire n_7828;
wire n_8340;
wire n_8905;
wire n_12020;
wire n_4935;
wire n_8691;
wire n_12051;
wire n_6365;
wire n_10619;
wire n_4785;
wire n_3426;
wire n_3454;
wire n_3820;
wire n_5608;
wire n_3741;
wire n_11322;
wire n_3410;
wire n_12455;
wire n_10136;
wire n_7401;
wire n_8812;
wire n_12920;
wire n_9169;
wire n_6828;
wire n_12785;
wire n_11758;
wire n_5298;
wire n_8704;
wire n_6355;
wire n_5596;
wire n_7887;
wire n_11162;
wire n_8058;
wire n_4413;
wire n_12559;
wire n_9177;
wire n_10078;
wire n_6777;
wire n_5728;
wire n_11987;
wire n_8394;
wire n_9269;
wire n_3990;
wire n_4493;
wire n_7835;
wire n_10719;
wire n_12614;
wire n_3475;
wire n_11106;
wire n_9289;
wire n_8181;
wire n_10463;
wire n_12797;
wire n_8722;
wire n_10827;
wire n_12429;
wire n_6420;
wire n_6945;
wire n_11218;
wire n_2882;
wire n_9350;
wire n_7356;
wire n_5726;
wire n_7288;
wire n_7637;
wire n_11467;
wire n_7124;
wire n_10454;
wire n_11795;
wire n_12384;
wire n_3672;
wire n_7294;
wire n_12629;
wire n_12668;
wire n_12123;
wire n_5290;
wire n_12972;
wire n_3197;
wire n_7018;
wire n_3109;
wire n_10312;
wire n_11374;
wire n_11167;
wire n_12146;
wire n_7321;
wire n_9166;
wire n_10663;
wire n_10501;
wire n_5095;
wire n_10265;
wire n_10452;
wire n_8707;
wire n_3002;
wire n_6754;
wire n_10766;
wire n_12435;
wire n_11999;
wire n_6583;
wire n_6622;
wire n_6936;
wire n_8747;
wire n_5324;
wire n_3897;
wire n_7691;
wire n_5928;
wire n_3845;
wire n_8742;
wire n_10470;
wire n_10563;
wire n_12921;
wire n_7108;
wire n_6882;
wire n_11455;
wire n_7585;
wire n_9125;
wire n_4570;
wire n_7386;
wire n_8552;
wire n_10288;
wire n_5101;
wire n_4296;
wire n_5019;
wire n_5911;
wire n_7362;
wire n_7888;
wire n_7417;
wire n_12029;
wire n_12548;
wire n_9641;
wire n_9960;
wire n_7187;
wire n_11884;
wire n_5589;
wire n_5841;
wire n_12727;
wire n_10776;
wire n_11611;
wire n_9785;
wire n_9923;
wire n_8224;
wire n_10771;
wire n_7544;
wire n_3458;
wire n_11087;
wire n_5712;
wire n_3330;
wire n_11960;
wire n_4606;
wire n_6166;
wire n_8628;
wire n_4774;
wire n_11422;
wire n_6966;
wire n_3887;
wire n_7542;
wire n_6781;
wire n_9228;
wire n_7255;
wire n_4093;
wire n_12227;
wire n_8037;
wire n_8084;
wire n_7120;
wire n_7218;
wire n_12597;
wire n_4672;
wire n_7147;
wire n_3519;
wire n_7221;
wire n_10967;
wire n_4174;
wire n_8289;
wire n_9801;
wire n_3374;
wire n_3045;
wire n_10249;
wire n_11029;
wire n_9645;
wire n_4766;
wire n_8045;
wire n_11199;
wire n_5633;
wire n_8697;
wire n_13029;
wire n_2896;
wire n_8077;
wire n_4074;
wire n_4600;
wire n_6980;
wire n_12674;
wire n_5583;
wire n_11826;
wire n_9457;
wire n_4460;
wire n_8026;
wire n_11317;
wire n_3645;
wire n_7889;
wire n_3223;
wire n_3929;
wire n_6064;
wire n_6110;
wire n_10742;
wire n_6237;
wire n_7196;
wire n_12913;
wire n_10390;
wire n_9330;
wire n_6341;
wire n_10012;
wire n_9365;
wire n_6590;
wire n_5501;
wire n_8444;
wire n_9178;
wire n_8654;
wire n_10035;
wire n_10753;
wire n_9181;
wire n_12112;
wire n_7923;
wire n_3938;
wire n_5377;
wire n_11033;
wire n_2878;
wire n_6697;
wire n_5652;
wire n_6453;
wire n_6135;
wire n_7559;
wire n_11798;
wire n_3498;
wire n_12346;
wire n_4110;
wire n_11853;
wire n_7081;
wire n_9307;
wire n_3189;
wire n_10795;
wire n_10300;
wire n_10257;
wire n_6449;
wire n_7832;
wire n_7968;
wire n_3154;
wire n_9238;
wire n_12714;
wire n_11079;
wire n_11166;
wire n_6141;
wire n_2905;
wire n_10099;
wire n_8449;
wire n_11217;
wire n_12732;
wire n_3965;
wire n_3566;
wire n_10985;
wire n_4349;
wire n_8493;
wire n_7584;
wire n_9224;
wire n_3788;
wire n_10244;
wire n_12400;
wire n_4313;
wire n_6983;
wire n_12671;
wire n_7843;
wire n_10377;
wire n_6036;
wire n_11469;
wire n_10984;
wire n_3366;
wire n_12863;
wire n_12347;
wire n_8958;
wire n_10801;
wire n_11898;
wire n_8443;
wire n_4863;
wire n_12041;
wire n_9756;
wire n_7222;
wire n_3242;
wire n_9624;
wire n_6071;
wire n_3525;
wire n_8161;
wire n_11710;
wire n_3486;
wire n_6808;
wire n_8734;
wire n_9547;
wire n_11341;
wire n_8271;
wire n_9594;
wire n_9901;
wire n_11619;
wire n_11238;
wire n_9895;
wire n_10878;
wire n_6724;
wire n_3995;
wire n_2953;
wire n_9277;
wire n_11608;
wire n_4036;
wire n_12756;
wire n_6571;
wire n_5100;
wire n_7470;
wire n_9189;
wire n_5849;
wire n_8495;
wire n_6251;
wire n_7400;
wire n_9548;
wire n_12088;
wire n_12218;
wire n_3483;
wire n_6635;
wire n_10000;
wire n_3894;
wire n_9472;
wire n_3478;
wire n_11553;
wire n_4015;
wire n_3890;
wire n_5367;
wire n_8994;
wire n_8901;
wire n_8056;
wire n_10725;
wire n_12323;
wire n_9538;
wire n_7623;
wire n_12387;
wire n_10627;
wire n_8954;
wire n_3524;
wire n_5616;
wire n_7597;
wire n_11996;
wire n_5034;
wire n_6733;
wire n_7071;
wire n_8840;
wire n_5988;
wire n_6467;
wire n_6035;
wire n_7859;
wire n_8900;
wire n_10477;
wire n_12798;
wire n_3549;
wire n_11032;
wire n_6522;
wire n_7109;
wire n_11834;
wire n_9434;
wire n_10604;
wire n_11110;
wire n_5959;
wire n_9052;
wire n_7645;
wire n_3658;
wire n_6732;
wire n_4807;
wire n_6562;
wire n_12780;
wire n_6150;
wire n_9176;
wire n_10461;
wire n_12772;
wire n_10559;
wire n_3026;
wire n_11141;
wire n_8157;
wire n_12539;
wire n_13007;
wire n_8346;
wire n_9697;
wire n_4230;
wire n_7882;
wire n_8827;
wire n_3419;
wire n_8309;
wire n_8344;
wire n_5917;
wire n_12589;
wire n_9060;
wire n_5754;
wire n_6016;
wire n_12775;
wire n_8096;
wire n_8100;
wire n_8822;
wire n_3784;
wire n_3941;
wire n_2969;
wire n_2864;
wire n_12043;
wire n_3195;
wire n_9758;
wire n_3190;
wire n_7212;
wire n_3678;
wire n_7908;
wire n_8222;
wire n_3456;
wire n_10479;
wire n_9876;
wire n_5628;
wire n_10572;
wire n_11971;
wire n_6726;
wire n_8406;
wire n_10277;
wire n_11320;
wire n_4428;
wire n_5003;
wire n_11028;
wire n_5252;
wire n_7009;
wire n_6554;
wire n_10230;
wire n_10139;
wire n_6689;
wire n_12476;
wire n_8866;
wire n_6143;
wire n_5614;
wire n_8693;
wire n_5134;
wire n_3953;
wire n_3166;
wire n_10207;
wire n_12536;
wire n_4122;
wire n_3976;
wire n_11368;
wire n_11144;
wire n_7355;
wire n_3979;
wire n_7365;
wire n_4582;
wire n_7777;
wire n_8794;
wire n_2998;
wire n_6277;
wire n_9653;
wire n_4684;
wire n_7395;
wire n_5981;
wire n_11404;
wire n_12896;
wire n_6095;
wire n_7671;
wire n_10429;
wire n_8020;
wire n_12957;
wire n_6247;
wire n_4840;
wire n_10255;
wire n_9257;
wire n_13014;
wire n_3162;
wire n_9270;
wire n_6880;
wire n_3377;
wire n_10901;
wire n_3749;
wire n_10101;
wire n_5720;
wire n_3962;
wire n_13022;
wire n_5325;
wire n_5696;
wire n_12549;
wire n_5375;
wire n_4384;
wire n_8736;
wire n_6499;
wire n_12362;
wire n_6837;
wire n_4423;
wire n_10063;
wire n_4096;
wire n_12030;
wire n_7393;
wire n_2881;
wire n_8400;
wire n_6616;
wire n_9686;
wire n_3282;
wire n_3231;
wire n_7871;
wire n_12018;
wire n_10846;
wire n_6946;
wire n_4996;
wire n_8333;
wire n_8055;
wire n_10195;
wire n_11593;
wire n_11847;
wire n_9718;
wire n_11773;
wire n_4598;
wire n_5064;
wire n_9215;
wire n_5759;
wire n_12060;
wire n_4478;
wire n_5753;
wire n_10628;
wire n_8909;
wire n_5536;
wire n_7484;
wire n_5173;
wire n_11968;
wire n_6305;
wire n_6317;
wire n_3920;
wire n_9762;
wire n_9407;
wire n_10819;
wire n_12315;
wire n_12903;
wire n_4890;
wire n_5691;
wire n_5794;
wire n_11896;
wire n_5027;
wire n_5647;
wire n_7231;
wire n_11897;
wire n_3203;
wire n_10368;
wire n_12484;
wire n_3866;
wire n_2903;
wire n_3921;
wire n_7272;
wire n_9964;
wire n_4106;
wire n_3717;
wire n_13031;
wire n_5738;
wire n_7649;
wire n_9953;
wire n_10356;
wire n_3052;
wire n_5215;
wire n_7324;
wire n_9153;
wire n_6693;
wire n_8786;
wire n_10931;
wire n_8541;
wire n_11711;
wire n_3743;
wire n_12673;
wire n_6734;
wire n_12000;
wire n_10173;
wire n_9571;
wire n_7135;
wire n_11554;
wire n_7014;
wire n_8263;
wire n_10644;
wire n_11159;
wire n_8884;
wire n_4721;
wire n_5597;
wire n_5635;
wire n_10323;
wire n_11350;
wire n_6382;
wire n_9019;
wire n_11310;
wire n_13001;
wire n_7328;
wire n_7635;
wire n_6404;
wire n_12063;
wire n_10229;
wire n_10693;
wire n_5975;
wire n_9737;
wire n_4029;
wire n_11688;
wire n_10493;
wire n_11125;
wire n_8494;
wire n_10554;
wire n_3870;
wire n_6379;
wire n_10382;
wire n_11083;
wire n_7703;
wire n_7066;
wire n_4496;
wire n_3529;
wire n_7358;
wire n_9468;
wire n_10622;
wire n_12449;
wire n_11939;
wire n_6235;
wire n_9870;
wire n_4338;
wire n_7277;
wire n_6504;
wire n_9026;
wire n_3094;
wire n_9710;
wire n_3952;
wire n_7265;
wire n_8638;
wire n_2860;
wire n_11126;
wire n_8710;
wire n_10019;
wire n_6789;
wire n_7184;
wire n_11090;
wire n_6440;
wire n_9725;
wire n_11953;
wire n_6417;
wire n_12845;
wire n_8177;
wire n_12062;
wire n_12636;
wire n_4495;
wire n_4762;
wire n_7491;
wire n_5942;
wire n_2974;
wire n_2901;
wire n_9084;
wire n_7728;
wire n_3442;
wire n_10488;
wire n_10767;
wire n_7690;
wire n_7219;
wire n_7479;
wire n_11040;
wire n_3998;
wire n_11751;
wire n_9419;
wire n_12793;
wire n_3147;
wire n_4141;
wire n_11158;
wire n_7270;
wire n_5940;
wire n_8170;
wire n_12367;
wire n_10579;
wire n_8893;
wire n_12317;
wire n_7390;
wire n_7805;
wire n_10474;
wire n_7807;
wire n_5121;
wire n_9479;
wire n_3386;
wire n_8589;
wire n_4107;
wire n_9973;
wire n_9820;
wire n_12724;
wire n_12954;
wire n_4667;
wire n_11094;
wire n_8320;
wire n_5555;
wire n_6914;
wire n_7978;
wire n_12157;
wire n_3488;
wire n_11161;
wire n_11182;
wire n_10587;
wire n_7182;
wire n_12195;
wire n_4547;
wire n_11839;
wire n_2893;
wire n_11815;
wire n_4004;
wire n_2962;
wire n_5784;
wire n_10843;
wire n_12773;
wire n_6272;
wire n_8153;
wire n_7699;
wire n_6484;
wire n_7674;
wire n_12556;
wire n_6236;
wire n_8620;
wire n_10755;
wire n_5576;
wire n_4668;
wire n_8298;
wire n_11614;
wire n_4953;
wire n_5466;
wire n_6958;
wire n_6840;
wire n_3898;
wire n_6871;
wire n_12789;
wire n_10270;
wire n_11590;
wire n_12649;
wire n_8235;
wire n_11845;
wire n_5284;
wire n_9294;
wire n_9126;
wire n_8370;
wire n_11263;
wire n_11908;
wire n_4997;
wire n_5308;
wire n_4274;
wire n_10573;
wire n_6768;
wire n_4759;
wire n_7951;
wire n_10992;
wire n_4467;
wire n_7506;
wire n_3552;
wire n_12696;
wire n_6717;
wire n_11257;
wire n_3684;
wire n_4735;
wire n_3137;
wire n_7048;
wire n_11142;
wire n_11136;
wire n_10428;
wire n_12664;
wire n_5578;
wire n_8395;
wire n_10989;
wire n_11145;
wire n_12206;
wire n_11745;
wire n_13010;
wire n_11017;
wire n_4113;
wire n_10805;
wire n_8906;
wire n_4686;
wire n_10682;
wire n_5530;
wire n_11414;
wire n_8097;
wire n_10327;
wire n_12940;
wire n_3759;
wire n_6196;
wire n_7416;
wire n_4321;
wire n_4342;
wire n_10528;
wire n_5741;
wire n_8570;
wire n_8902;
wire n_12404;
wire n_5991;
wire n_3933;
wire n_10365;
wire n_7330;
wire n_3206;
wire n_7928;
wire n_12201;
wire n_5506;
wire n_3966;
wire n_5243;
wire n_9819;
wire n_8477;
wire n_5449;
wire n_10236;
wire n_5221;
wire n_6992;
wire n_10433;
wire n_4183;
wire n_12312;
wire n_4068;
wire n_4872;
wire n_10625;
wire n_6000;
wire n_10303;
wire n_9545;
wire n_4233;
wire n_7283;
wire n_3192;
wire n_7099;
wire n_3764;
wire n_11452;
wire n_10557;
wire n_4709;
wire n_5038;
wire n_5311;
wire n_6448;
wire n_11323;
wire n_13002;
wire n_6655;
wire n_12982;
wire n_7892;
wire n_9165;
wire n_11558;
wire n_7304;
wire n_10143;
wire n_13018;
wire n_5792;
wire n_12002;
wire n_6657;
wire n_7756;
wire n_8129;
wire n_5575;
wire n_8580;
wire n_11543;
wire n_7990;
wire n_3324;
wire n_4625;
wire n_3914;
wire n_8122;
wire n_11883;
wire n_10796;
wire n_8259;
wire n_3803;
wire n_8536;
wire n_7626;
wire n_3742;
wire n_7474;
wire n_10855;
wire n_8748;
wire n_7612;
wire n_6113;
wire n_7789;
wire n_4819;
wire n_9056;
wire n_8094;
wire n_9341;
wire n_11429;
wire n_6242;
wire n_7902;
wire n_7088;
wire n_6519;
wire n_10357;
wire n_8572;
wire n_4900;
wire n_10681;
wire n_8120;
wire n_12598;
wire n_6842;
wire n_12942;
wire n_12750;
wire n_12729;
wire n_7588;
wire n_3390;
wire n_12033;
wire n_6206;
wire n_6414;
wire n_3746;
wire n_11241;
wire n_9172;
wire n_3817;
wire n_12441;
wire n_9145;
wire n_6801;
wire n_8099;
wire n_9996;
wire n_11348;
wire n_10059;
wire n_10284;
wire n_4930;
wire n_7680;
wire n_8770;
wire n_5276;
wire n_6308;
wire n_7398;
wire n_6906;
wire n_5078;
wire n_11169;
wire n_4537;
wire n_11041;
wire n_7230;
wire n_8700;
wire n_11160;
wire n_2885;
wire n_9906;
wire n_6629;
wire n_5011;
wire n_10957;
wire n_12827;
wire n_3318;
wire n_4070;
wire n_11124;
wire n_6968;
wire n_9920;
wire n_4282;
wire n_9504;
wire n_6615;
wire n_3485;
wire n_4180;
wire n_7378;
wire n_3839;
wire n_12734;
wire n_12181;
wire n_9482;
wire n_5205;
wire n_9138;
wire n_11152;
wire n_3333;
wire n_9384;
wire n_8637;
wire n_5651;
wire n_2845;
wire n_6144;
wire n_8757;
wire n_4143;
wire n_4659;
wire n_6188;
wire n_5819;
wire n_10147;
wire n_4579;
wire n_4616;
wire n_8903;
wire n_9193;
wire n_3014;
wire n_5998;
wire n_6398;
wire n_11586;
wire n_5023;
wire n_12069;
wire n_11990;
wire n_4105;
wire n_5721;
wire n_5673;
wire n_9527;
wire n_3791;
wire n_5351;
wire n_3905;
wire n_10889;
wire n_12363;
wire n_3368;
wire n_11019;
wire n_8585;
wire n_9064;
wire n_3530;
wire n_8982;
wire n_3329;
wire n_6415;
wire n_10816;
wire n_2994;
wire n_10032;
wire n_6857;
wire n_10489;
wire n_3135;
wire n_5476;
wire n_10200;
wire n_12442;
wire n_7842;
wire n_10898;
wire n_5856;
wire n_12499;
wire n_8709;
wire n_5446;
wire n_9383;
wire n_10825;
wire n_4895;
wire n_6722;
wire n_3573;
wire n_3148;
wire n_9943;
wire n_9735;
wire n_10290;
wire n_6428;
wire n_5944;
wire n_7618;
wire n_3534;
wire n_12818;
wire n_6413;
wire n_7679;
wire n_11132;
wire n_4275;
wire n_6361;
wire n_3970;
wire n_9357;
wire n_11677;
wire n_3438;
wire n_10680;
wire n_12531;
wire n_6231;
wire n_7783;
wire n_4098;
wire n_11036;
wire n_5684;
wire n_5861;
wire n_11927;
wire n_8108;
wire n_10306;
wire n_5976;
wire n_4789;
wire n_11827;
wire n_7862;
wire n_5312;
wire n_10675;
wire n_5850;
wire n_10014;
wire n_3217;
wire n_3404;
wire n_3425;
wire n_5111;
wire n_5890;
wire n_4055;
wire n_2926;
wire n_9986;
wire n_3540;
wire n_10355;
wire n_3670;
wire n_3973;
wire n_10830;
wire n_7820;
wire n_7167;
wire n_8692;
wire n_7833;
wire n_11118;
wire n_8820;
wire n_3249;
wire n_12496;
wire n_7643;
wire n_12460;
wire n_8490;
wire n_10380;
wire n_5113;
wire n_4442;
wire n_9491;
wire n_4698;
wire n_12821;
wire n_9922;
wire n_6712;
wire n_5687;
wire n_12479;
wire n_10530;
wire n_4779;
wire n_8062;
wire n_8781;
wire n_10999;
wire n_10203;
wire n_4966;
wire n_8000;
wire n_10061;
wire n_10899;
wire n_10961;
wire n_4017;
wire n_8808;
wire n_8233;
wire n_5839;
wire n_3397;
wire n_3740;
wire n_9747;
wire n_11811;
wire n_6953;
wire n_4418;
wire n_8685;
wire n_9061;
wire n_9168;
wire n_12361;
wire n_11561;
wire n_12345;
wire n_8575;
wire n_8701;
wire n_11690;
wire n_2977;
wire n_11212;
wire n_6303;
wire n_12593;
wire n_6474;
wire n_6182;
wire n_3723;
wire n_11155;
wire n_5674;
wire n_3600;
wire n_8670;
wire n_6573;
wire n_4134;
wire n_6053;
wire n_7234;
wire n_10425;
wire n_8352;
wire n_7993;
wire n_7930;
wire n_2836;
wire n_5682;
wire n_12984;
wire n_8385;
wire n_8875;
wire n_6392;
wire n_8166;
wire n_11433;
wire n_5167;
wire n_3239;
wire n_8934;
wire n_5117;
wire n_9073;
wire n_3365;
wire n_3476;
wire n_3686;
wire n_4913;
wire n_11312;
wire n_11477;
wire n_7999;
wire n_5612;
wire n_11988;
wire n_6125;
wire n_7963;
wire n_6599;
wire n_6685;
wire n_12311;
wire n_12914;
wire n_2850;
wire n_11964;
wire n_12086;
wire n_4251;
wire n_8389;
wire n_9068;
wire n_3982;
wire n_10537;
wire n_4621;
wire n_10158;
wire n_6560;
wire n_12787;
wire n_10711;
wire n_3176;
wire n_11933;
wire n_8659;
wire n_8804;
wire n_10043;
wire n_4559;
wire n_12703;
wire n_4368;
wire n_6253;
wire n_12411;
wire n_4740;
wire n_7382;
wire n_8439;
wire n_9544;
wire n_8814;
wire n_8369;
wire n_5301;
wire n_11574;
wire n_7800;
wire n_5007;
wire n_3581;
wire n_4077;
wire n_4642;
wire n_7615;
wire n_5898;
wire n_9286;
wire n_10930;
wire n_11313;
wire n_3576;
wire n_11206;
wire n_12263;
wire n_7298;
wire n_12959;
wire n_10131;
wire n_7581;
wire n_4049;
wire n_6641;
wire n_5214;
wire n_3862;
wire n_5563;
wire n_5487;
wire n_6593;
wire n_3495;
wire n_3879;
wire n_6673;
wire n_10696;
wire n_12461;
wire n_12893;
wire n_8789;
wire n_7172;
wire n_7074;
wire n_10685;
wire n_5497;
wire n_8790;
wire n_11223;
wire n_8234;
wire n_11624;
wire n_4724;
wire n_5832;
wire n_7190;
wire n_11515;
wire n_7112;
wire n_7678;
wire n_10082;
wire n_9265;
wire n_11560;
wire n_9080;
wire n_5526;
wire n_8989;
wire n_10152;
wire n_2818;
wire n_3646;
wire n_12645;
wire n_6367;
wire n_6195;
wire n_3345;
wire n_4546;
wire n_6356;
wire n_3584;
wire n_8927;
wire n_11055;
wire n_3756;
wire n_11616;
wire n_9770;
wire n_2889;
wire n_9463;
wire n_7001;
wire n_12090;
wire n_5593;
wire n_5021;
wire n_6514;
wire n_7369;
wire n_5444;
wire n_10580;
wire n_7829;
wire n_4382;
wire n_9939;
wire n_10159;
wire n_3999;
wire n_11390;
wire n_8534;
wire n_2844;
wire n_9911;
wire n_9210;
wire n_5211;
wire n_6559;
wire n_5230;
wire n_10122;
wire n_10302;
wire n_7359;
wire n_5389;
wire n_7144;
wire n_10462;
wire n_4833;
wire n_8756;
wire n_6841;
wire n_11597;
wire n_3056;
wire n_11002;
wire n_9691;
wire n_5110;
wire n_6653;
wire n_12165;
wire n_3295;
wire n_4719;
wire n_4178;
wire n_3062;
wire n_7450;
wire n_5425;
wire n_3289;
wire n_10532;
wire n_8832;
wire n_5737;
wire n_9340;
wire n_10350;
wire n_9351;
wire n_8461;
wire n_8042;
wire n_10977;
wire n_11179;
wire n_6825;
wire n_6923;
wire n_11708;
wire n_9950;
wire n_10418;
wire n_11474;
wire n_10336;
wire n_4228;
wire n_4401;
wire n_8021;
wire n_8839;
wire n_12092;
wire n_11369;
wire n_6112;
wire n_11738;
wire n_6547;
wire n_11240;
wire n_2984;
wire n_6198;
wire n_7439;
wire n_3364;
wire n_5560;
wire n_12074;
wire n_9155;
wire n_11931;
wire n_10925;
wire n_6399;
wire n_8623;
wire n_12109;
wire n_3201;
wire n_11438;
wire n_8758;
wire n_6275;
wire n_5666;
wire n_6575;
wire n_10609;
wire n_3472;
wire n_7924;
wire n_7732;
wire n_6151;
wire n_2874;
wire n_5179;
wire n_7227;
wire n_7040;
wire n_4605;
wire n_4877;
wire n_8511;
wire n_3235;
wire n_7325;
wire n_4968;
wire n_6469;
wire n_6756;
wire n_8595;
wire n_12900;
wire n_8873;
wire n_11376;
wire n_5030;
wire n_3949;
wire n_5961;
wire n_3543;
wire n_7191;
wire n_7459;
wire n_9201;
wire n_9823;
wire n_11051;
wire n_11812;
wire n_9688;
wire n_12330;
wire n_7096;
wire n_12519;
wire n_3050;
wire n_8455;
wire n_11838;
wire n_12717;
wire n_8280;
wire n_3903;
wire n_10102;
wire n_4834;
wire n_10908;
wire n_11333;
wire n_9595;
wire n_5272;
wire n_9530;
wire n_3314;
wire n_4158;
wire n_6826;
wire n_9227;
wire n_6015;
wire n_3254;
wire n_8372;
wire n_5361;
wire n_8598;
wire n_5683;
wire n_10939;
wire n_4171;
wire n_11178;
wire n_12595;
wire n_5847;
wire n_7551;
wire n_9400;
wire n_4045;
wire n_6678;
wire n_11188;
wire n_4562;
wire n_5068;
wire n_3634;
wire n_9025;
wire n_5740;
wire n_2834;
wire n_8282;
wire n_7750;
wire n_10936;
wire n_11840;
wire n_5015;
wire n_12525;
wire n_7697;
wire n_5729;
wire n_7485;
wire n_11685;
wire n_10955;
wire n_10824;
wire n_6748;
wire n_12084;
wire n_8616;
wire n_3115;
wire n_4749;
wire n_10440;
wire n_10630;
wire n_8336;
wire n_4390;
wire n_5302;
wire n_4979;
wire n_11472;
wire n_6752;
wire n_9749;
wire n_4804;
wire n_5545;
wire n_6553;
wire n_9285;
wire n_12997;
wire n_11295;
wire n_9972;
wire n_10058;
wire n_7652;
wire n_8847;
wire n_7808;
wire n_11171;
wire n_6500;
wire n_4270;
wire n_8135;
wire n_9214;
wire n_7051;
wire n_9859;
wire n_11030;
wire n_10295;
wire n_5152;
wire n_9003;
wire n_11443;
wire n_9271;
wire n_9258;
wire n_3680;
wire n_6628;
wire n_12661;
wire n_12693;
wire n_6297;
wire n_5905;
wire n_3497;
wire n_12203;
wire n_6975;
wire n_5409;
wire n_6329;
wire n_2940;
wire n_7536;
wire n_8979;
wire n_12080;
wire n_8529;
wire n_10658;
wire n_5688;
wire n_9763;
wire n_5128;
wire n_10894;
wire n_4566;
wire n_9597;
wire n_2841;
wire n_6293;
wire n_8417;
wire n_9965;
wire n_9076;
wire n_10912;
wire n_7952;
wire n_3322;
wire n_4576;
wire n_9393;
wire n_8498;
wire n_7991;
wire n_7676;
wire n_11769;
wire n_4061;
wire n_12486;
wire n_3250;
wire n_7553;
wire n_6905;
wire n_12623;
wire n_7425;
wire n_5798;
wire n_6381;
wire n_6521;
wire n_2904;
wire n_5307;
wire n_12933;
wire n_12489;
wire n_8967;
wire n_8355;
wire n_9736;
wire n_4767;
wire n_7998;
wire n_4328;
wire n_3004;
wire n_5986;
wire n_8719;
wire n_3112;
wire n_6581;
wire n_10160;
wire n_10678;
wire n_3874;
wire n_6215;
wire n_7095;
wire n_11794;
wire n_5415;
wire n_4676;
wire n_10241;
wire n_5770;
wire n_11495;
wire n_7064;
wire n_5892;
wire n_8762;
wire n_12480;
wire n_4544;
wire n_10180;
wire n_8516;
wire n_8880;
wire n_6577;
wire n_6899;
wire n_8784;
wire n_12335;
wire n_5676;
wire n_7307;
wire n_6545;
wire n_10631;
wire n_8237;
wire n_5802;
wire n_3175;
wire n_3522;
wire n_10852;
wire n_9803;
wire n_4429;
wire n_8977;
wire n_11406;
wire n_8171;
wire n_4591;
wire n_10978;
wire n_10500;
wire n_6370;
wire n_9755;
wire n_3266;
wire n_9805;
wire n_7210;
wire n_4646;
wire n_7899;
wire n_10370;
wire n_9728;
wire n_5769;
wire n_6065;
wire n_7039;
wire n_9659;
wire n_6987;
wire n_12624;
wire n_4563;
wire n_4725;
wire n_9107;
wire n_11428;
wire n_6190;
wire n_5331;
wire n_4169;
wire n_6859;
wire n_3247;
wire n_3091;
wire n_12410;
wire n_9917;
wire n_3066;
wire n_6309;
wire n_11149;
wire n_9520;
wire n_6623;
wire n_12055;
wire n_12925;
wire n_7723;
wire n_12771;
wire n_6527;
wire n_7443;
wire n_11707;
wire n_10550;
wire n_9583;
wire n_7811;
wire n_12413;
wire n_11086;
wire n_5341;
wire n_4320;
wire n_12182;
wire n_5930;
wire n_5814;
wire n_12803;
wire n_4881;
wire n_9036;
wire n_9522;
wire n_5979;
wire n_5271;
wire n_5089;
wire n_10571;
wire n_7015;
wire n_5263;
wire n_3613;
wire n_11772;
wire n_12547;
wire n_3444;
wire n_6929;
wire n_11225;
wire n_11764;
wire n_12544;
wire n_11339;
wire n_4012;
wire n_5518;
wire n_10125;
wire n_4636;
wire n_5637;
wire n_12370;
wire n_4584;
wire n_12931;
wire n_8279;
wire n_5622;
wire n_3910;
wire n_4711;
wire n_11112;
wire n_9723;
wire n_12986;
wire n_3319;
wire n_7348;
wire n_10254;
wire n_5240;
wire n_3335;
wire n_5813;
wire n_3413;
wire n_5495;
wire n_4680;
wire n_5546;
wire n_8912;
wire n_3259;
wire n_9488;
wire n_7143;
wire n_5482;
wire n_7312;
wire n_4191;
wire n_5224;
wire n_4293;
wire n_7155;
wire n_8227;
wire n_3688;
wire n_9231;
wire n_8938;
wire n_6865;
wire n_3016;
wire n_8787;
wire n_5393;
wire n_10017;
wire n_6535;
wire n_3338;
wire n_7213;
wire n_10866;
wire n_3414;
wire n_9047;
wire n_10348;
wire n_12991;
wire n_4671;
wire n_8270;
wire n_4209;
wire n_5966;
wire n_11072;
wire n_7456;
wire n_8335;
wire n_11359;
wire n_10657;
wire n_5041;
wire n_7420;
wire n_11605;
wire n_9798;
wire n_9681;
wire n_8054;
wire n_9414;
wire n_12419;
wire n_8607;
wire n_5431;
wire n_9979;
wire n_9093;
wire n_3261;
wire n_11959;
wire n_6482;
wire n_5026;
wire n_3863;
wire n_11318;
wire n_3027;
wire n_11830;
wire n_10842;
wire n_13012;
wire n_12865;
wire n_8150;
wire n_5059;
wire n_9379;
wire n_5505;
wire n_3127;
wire n_7715;
wire n_9486;
wire n_3732;
wire n_11881;
wire n_6605;
wire n_4250;
wire n_9134;
wire n_5329;
wire n_12481;
wire n_3596;
wire n_4699;
wire n_7007;
wire n_8358;
wire n_9410;
wire n_3906;
wire n_4127;
wire n_10045;
wire n_3297;
wire n_7909;
wire n_9151;
wire n_12278;
wire n_4292;
wire n_3641;
wire n_4577;
wire n_11863;
wire n_4854;
wire n_8281;
wire n_12562;
wire n_11494;
wire n_9182;
wire n_6018;
wire n_5908;
wire n_12744;
wire n_4202;
wire n_7168;
wire n_11850;
wire n_5212;
wire n_9976;
wire n_7736;
wire n_5000;
wire n_8396;
wire n_9591;
wire n_10322;
wire n_2853;
wire n_9838;
wire n_5939;
wire n_7177;
wire n_10033;
wire n_3766;
wire n_12615;
wire n_13027;
wire n_11258;
wire n_9568;
wire n_7780;
wire n_10886;
wire n_2880;
wire n_9261;
wire n_9701;
wire n_7379;
wire n_3350;
wire n_4165;
wire n_4866;
wire n_7444;
wire n_8223;
wire n_5931;
wire n_11468;
wire n_7435;
wire n_4038;
wire n_4109;
wire n_5297;
wire n_7813;
wire n_7030;
wire n_8459;
wire n_5420;
wire n_6311;
wire n_11192;
wire n_12580;
wire n_11569;
wire n_4412;
wire n_3407;
wire n_6654;
wire n_6424;
wire n_3599;
wire n_6816;
wire n_6220;
wire n_3621;
wire n_9752;
wire n_12769;
wire n_5234;
wire n_6740;
wire n_7122;
wire n_12540;
wire n_5835;
wire n_7049;
wire n_7567;
wire n_3815;
wire n_6029;
wire n_8379;
wire n_11563;
wire n_6879;
wire n_5259;
wire n_5440;
wire n_3163;
wire n_5679;
wire n_5938;
wire n_3710;
wire n_9079;
wire n_6702;
wire n_4155;
wire n_11846;
wire n_3891;
wire n_5891;
wire n_10383;
wire n_4144;
wire n_5724;
wire n_10064;
wire n_10876;
wire n_5774;
wire n_8793;
wire n_11852;
wire n_6452;
wire n_4374;
wire n_3379;
wire n_12619;
wire n_8975;
wire n_6791;
wire n_3532;
wire n_9170;
wire n_11679;
wire n_8792;
wire n_5131;
wire n_7280;
wire n_8671;
wire n_6915;
wire n_7110;
wire n_8489;
wire n_7511;
wire n_10831;
wire n_6856;
wire n_7941;
wire n_7791;
wire n_9385;
wire n_3531;
wire n_11186;
wire n_11870;
wire n_12960;
wire n_8484;
wire n_3834;
wire n_2963;
wire n_8454;
wire n_11492;
wire n_10536;
wire n_10238;
wire n_7232;
wire n_8759;
wire n_12268;
wire n_11544;
wire n_4548;
wire n_7345;
wire n_5923;
wire n_8703;
wire n_11233;
wire n_12656;
wire n_5790;
wire n_3258;
wire n_12678;
wire n_10206;
wire n_4989;
wire n_4622;
wire n_4315;
wire n_12880;
wire n_2959;
wire n_9670;
wire n_12876;
wire n_6451;
wire n_6364;
wire n_12711;
wire n_6552;
wire n_10786;
wire n_8325;
wire n_5140;
wire n_6328;
wire n_9598;
wire n_4816;
wire n_8382;
wire n_7827;
wire n_8971;
wire n_6363;
wire n_11646;
wire n_10602;
wire n_10620;
wire n_2983;
wire n_7159;
wire n_8127;
wire n_11878;
wire n_10079;
wire n_10188;
wire n_3810;
wire n_8721;
wire n_9391;
wire n_12458;
wire n_6132;
wire n_6578;
wire n_8889;
wire n_6406;
wire n_10319;
wire n_5598;
wire n_11900;
wire n_9470;
wire n_12132;
wire n_5306;
wire n_6978;
wire n_12104;
wire n_12037;
wire n_9328;
wire n_12467;
wire n_4483;
wire n_12870;
wire n_5342;
wire n_9245;
wire n_10739;
wire n_12911;
wire n_8232;
wire n_4358;
wire n_7477;
wire n_5147;
wire n_3656;
wire n_6918;
wire n_7363;
wire n_4793;
wire n_9833;
wire n_12386;
wire n_11837;
wire n_10213;
wire n_6612;
wire n_10107;
wire n_8664;
wire n_5677;
wire n_4168;
wire n_10872;
wire n_3446;
wire n_5997;
wire n_9455;
wire n_12651;
wire n_5511;
wire n_7863;
wire n_5680;
wire n_9719;
wire n_4806;
wire n_3028;
wire n_4350;
wire n_7295;
wire n_8633;
wire n_9744;
wire n_8842;
wire n_5533;
wire n_5838;
wire n_6058;
wire n_11871;
wire n_8956;
wire n_5280;
wire n_10969;
wire n_6375;
wire n_6479;
wire n_6866;
wire n_12563;
wire n_7831;
wire n_11674;
wire n_12621;
wire n_5235;
wire n_3836;
wire n_3963;
wire n_3389;
wire n_12331;
wire n_12304;
wire n_9698;
wire n_12339;
wire n_6170;
wire n_12270;
wire n_9124;
wire n_10718;
wire n_10669;
wire n_9695;
wire n_4187;
wire n_6447;
wire n_4166;
wire n_6263;
wire n_7093;
wire n_9497;
wire n_5206;
wire n_10895;
wire n_8641;
wire n_8479;
wire n_3222;
wire n_11610;
wire n_11187;
wire n_12210;
wire n_7466;
wire n_5419;
wire n_6130;
wire n_12858;
wire n_2970;
wire n_12382;
wire n_11280;
wire n_10757;
wire n_7651;
wire n_4937;
wire n_3980;
wire n_10513;
wire n_5103;
wire n_3755;
wire n_11148;
wire n_8179;
wire n_5803;
wire n_4258;
wire n_6014;
wire n_4498;
wire n_11396;
wire n_8973;
wire n_6935;
wire n_10194;
wire n_9775;
wire n_7530;
wire n_5285;
wire n_11426;
wire n_3563;
wire n_4064;
wire n_9038;
wire n_8308;
wire n_4936;
wire n_5387;
wire n_9630;
wire n_10692;
wire n_8378;
wire n_3841;
wire n_8733;
wire n_12107;
wire n_8809;
wire n_4770;
wire n_5985;
wire n_2944;
wire n_11723;
wire n_11009;
wire n_4907;
wire n_9652;
wire n_10021;
wire n_5058;
wire n_12381;
wire n_6907;
wire n_11706;
wire n_8500;
wire n_12653;
wire n_6158;
wire n_7661;
wire n_10782;
wire n_9709;
wire n_6541;
wire n_3262;
wire n_6119;
wire n_8447;
wire n_5018;
wire n_11949;
wire n_4006;
wire n_5896;
wire n_4861;
wire n_10457;
wire n_9324;
wire n_3690;
wire n_9934;
wire n_11957;
wire n_5192;
wire n_8548;
wire n_11538;
wire n_5141;
wire n_3716;
wire n_5133;
wire n_8412;
wire n_4712;
wire n_2833;
wire n_6226;
wire n_3191;
wire n_11264;
wire n_3837;
wire n_11211;
wire n_12774;
wire n_3193;
wire n_11880;
wire n_9668;
wire n_3252;
wire n_7145;
wire n_2855;
wire n_3273;
wire n_10385;
wire n_3544;
wire n_11377;
wire n_12064;
wire n_9877;
wire n_4310;
wire n_12503;
wire n_9657;
wire n_10111;
wire n_11302;
wire n_6338;
wire n_12425;
wire n_11921;
wire n_5159;
wire n_9352;
wire n_3954;
wire n_9395;
wire n_12807;
wire n_8425;
wire n_10809;
wire n_9349;
wire n_4674;
wire n_3025;
wire n_4908;
wire n_8241;
wire n_7823;
wire n_9209;
wire n_7467;
wire n_5097;
wire n_10113;
wire n_11267;
wire n_10990;
wire n_7932;
wire n_11626;
wire n_5730;
wire n_3899;
wire n_7550;
wire n_11694;
wire n_4159;
wire n_3714;
wire n_11618;
wire n_9969;
wire n_3071;
wire n_3739;
wire n_9937;
wire n_5816;
wire n_4069;
wire n_7541;
wire n_3718;
wire n_10545;
wire n_12715;
wire n_3092;
wire n_4862;
wire n_3470;
wire n_7241;
wire n_7717;
wire n_5300;
wire n_10595;
wire n_10973;
wire n_11011;
wire n_12015;
wire n_12968;
wire n_9618;
wire n_10732;
wire n_10009;
wire n_11776;
wire n_4850;
wire n_6625;
wire n_11165;
wire n_4813;
wire n_4912;
wire n_3781;
wire n_12135;
wire n_7464;
wire n_9082;
wire n_11366;
wire n_6302;
wire n_9424;
wire n_8274;
wire n_9453;
wire n_5748;
wire n_2942;
wire n_6759;
wire n_5525;
wire n_3106;
wire n_9637;
wire n_8152;
wire n_3328;
wire n_6706;
wire n_10526;
wire n_8550;
wire n_3889;
wire n_6139;
wire n_4256;
wire n_8264;
wire n_7434;
wire n_7636;
wire n_6999;
wire n_7054;
wire n_12817;
wire n_4224;
wire n_6403;
wire n_3508;
wire n_6483;
wire n_8829;
wire n_9183;
wire n_9205;
wire n_12869;
wire n_9009;
wire n_4024;
wire n_6228;
wire n_11315;
wire n_5650;
wire n_10044;
wire n_12059;
wire n_11098;
wire n_12586;
wire n_5400;
wire n_4415;
wire n_5552;
wire n_7299;
wire n_10221;
wire n_4702;
wire n_6888;
wire n_8266;
wire n_8515;
wire n_10109;
wire n_10169;
wire n_4252;
wire n_4457;
wire n_8648;
wire n_6063;
wire n_10329;
wire n_10928;
wire n_9024;
wire n_9030;
wire n_9523;
wire n_9377;
wire n_10891;
wire n_8946;
wire n_10839;
wire n_11875;
wire n_6800;
wire n_5139;
wire n_9716;
wire n_6922;
wire n_9380;
wire n_3481;
wire n_5481;
wire n_6890;
wire n_8744;
wire n_9000;
wire n_9679;
wire n_9116;
wire n_9742;
wire n_9016;
wire n_7503;
wire n_6070;
wire n_9006;
wire n_12514;
wire n_11524;
wire n_10091;
wire n_6651;
wire n_5821;
wire n_7091;
wire n_4491;
wire n_7296;
wire n_6647;
wire n_7273;
wire n_2930;
wire n_5733;
wire n_10029;
wire n_9690;
wire n_3514;
wire n_8765;
wire n_4132;
wire n_5871;
wire n_9852;
wire n_7543;
wire n_4261;
wire n_10600;
wire n_9914;
wire n_11056;
wire n_11514;
wire n_12438;
wire n_6184;
wire n_4886;
wire n_11774;
wire n_8627;
wire n_4090;
wire n_7507;
wire n_9451;
wire n_10849;
wire n_5043;
wire n_11108;
wire n_9760;
wire n_7555;
wire n_5707;
wire n_10947;
wire n_4001;
wire n_3047;
wire n_10272;
wire n_12099;
wire n_9035;
wire n_12009;
wire n_12806;
wire n_4371;
wire n_5836;
wire n_9211;
wire n_5281;
wire n_6716;
wire n_6422;
wire n_12887;
wire n_12776;
wire n_4473;
wire n_3120;
wire n_4007;
wire n_12898;
wire n_4268;
wire n_9677;
wire n_5048;
wire n_11954;
wire n_5521;
wire n_12191;
wire n_7578;
wire n_5028;
wire n_4480;
wire n_3895;
wire n_7475;
wire n_4194;
wire n_8195;
wire n_9070;
wire n_5585;
wire n_6397;
wire n_12578;
wire n_4824;
wire n_4120;
wire n_4427;
wire n_11864;
wire n_3745;
wire n_2990;
wire n_7033;
wire n_9881;
wire n_6121;
wire n_3119;
wire n_9669;
wire n_7531;
wire n_4142;
wire n_9958;
wire n_4082;
wire n_9858;
wire n_8462;
wire n_5561;
wire n_3479;
wire n_9981;
wire n_4085;
wire n_10391;
wire n_4260;
wire n_4073;
wire n_8377;
wire n_11157;
wire n_4163;
wire n_4439;
wire n_12509;
wire n_12235;
wire n_6981;
wire n_3867;
wire n_4372;
wire n_3500;
wire n_9588;
wire n_6954;
wire n_11733;
wire n_3279;
wire n_5799;
wire n_5073;
wire n_5024;
wire n_12471;
wire n_12365;
wire n_5875;
wire n_8428;
wire n_8103;
wire n_4262;
wire n_9021;
wire n_6646;
wire n_8936;
wire n_8414;
wire n_8362;
wire n_12083;
wire n_9682;
wire n_10137;
wire n_10344;
wire n_7131;
wire n_4720;
wire n_7769;
wire n_10882;
wire n_11540;
wire n_11861;
wire n_6903;
wire n_9050;
wire n_11724;
wire n_9303;
wire n_12065;
wire n_9495;
wire n_12167;
wire n_11220;
wire n_4685;
wire n_6101;
wire n_9415;
wire n_5968;
wire n_10196;
wire n_8491;
wire n_9058;
wire n_4334;
wire n_6941;
wire n_9845;
wire n_8831;
wire n_4511;
wire n_5812;
wire n_6148;
wire n_5515;
wire n_8324;
wire n_11459;
wire n_11355;
wire n_6106;
wire n_9822;
wire n_12087;
wire n_6604;
wire n_12243;
wire n_4014;
wire n_7418;
wire n_12267;
wire n_5250;
wire n_3144;
wire n_12569;
wire n_4757;
wire n_7688;
wire n_2913;
wire n_10518;
wire n_11101;
wire n_9640;
wire n_11899;
wire n_8348;
wire n_5607;
wire n_4175;
wire n_8288;
wire n_10613;
wire n_10583;
wire n_4648;
wire n_11481;
wire n_11712;
wire n_11612;
wire n_8269;
wire n_5006;
wire n_7806;
wire n_10335;
wire n_10085;
wire n_10840;
wire n_6566;
wire n_12599;
wire n_8625;
wire n_5734;
wire n_6081;
wire n_8458;
wire n_4892;
wire n_8806;
wire n_7204;
wire n_10560;
wire n_3823;
wire n_8180;
wire n_4173;
wire n_8499;
wire n_8601;
wire n_4970;
wire n_9062;
wire n_3816;
wire n_5404;
wire n_4486;
wire n_4108;
wire n_8306;
wire n_12375;
wire n_12091;
wire n_9722;
wire n_12513;
wire n_6047;
wire n_2960;
wire n_8167;
wire n_5438;
wire n_9791;
wire n_10486;
wire n_12307;
wire n_9229;
wire n_11603;
wire n_11890;
wire n_4627;
wire n_8613;
wire n_9603;
wire n_11790;
wire n_8913;
wire n_11060;
wire n_7354;
wire n_7448;
wire n_8800;
wire n_6244;
wire n_12684;
wire n_8768;
wire n_6861;
wire n_9099;
wire n_3369;
wire n_3783;
wire n_10919;
wire n_3199;
wire n_3843;
wire n_12288;
wire n_9309;
wire n_12418;
wire n_7852;
wire n_10952;
wire n_5725;
wire n_12566;
wire n_7925;
wire n_12415;
wire n_3030;
wire n_9432;
wire n_9454;
wire n_3685;
wire n_4249;
wire n_7571;
wire n_11744;
wire n_9065;
wire n_11650;
wire n_5163;
wire n_11518;
wire n_7748;
wire n_5768;
wire n_12949;
wire n_4961;
wire n_7556;
wire n_3753;
wire n_7640;
wire n_8187;
wire n_10352;
wire n_8881;
wire n_9704;
wire n_4718;
wire n_3555;
wire n_3579;
wire n_11663;
wire n_5190;
wire n_7422;
wire n_7920;
wire n_8433;
wire n_9837;
wire n_10991;
wire n_4317;
wire n_3236;
wire n_4855;
wire n_9431;
wire n_10167;
wire n_3969;
wire n_12681;
wire n_12859;
wire n_9160;
wire n_10911;
wire n_4154;
wire n_9433;
wire n_6588;
wire n_3396;
wire n_9256;
wire n_10442;
wire n_12829;
wire n_11282;
wire n_9706;
wire n_12448;
wire n_7900;
wire n_7050;
wire n_4023;
wire n_9808;
wire n_9915;
wire n_10534;
wire n_4420;
wire n_5685;
wire n_11726;
wire n_5773;
wire n_7136;
wire n_10406;
wire n_10465;
wire n_12188;
wire n_12943;
wire n_8316;
wire n_7318;
wire n_12149;
wire n_6055;
wire n_5138;
wire n_12783;
wire n_8397;
wire n_9184;
wire n_5374;
wire n_10373;
wire n_9133;
wire n_6108;
wire n_8115;
wire n_12129;
wire n_12631;
wire n_6165;
wire n_10965;
wire n_6621;
wire n_7175;
wire n_5349;
wire n_4973;
wire n_7810;
wire n_9109;
wire n_4640;
wire n_6323;
wire n_10517;
wire n_12588;
wire n_12652;
wire n_8523;
wire n_9207;
wire n_11458;
wire n_4396;
wire n_5127;
wire n_6587;
wire n_4367;
wire n_6480;
wire n_7733;
wire n_6731;
wire n_5485;
wire n_10484;
wire n_5766;
wire n_11255;
wire n_5216;
wire n_6597;
wire n_10561;
wire n_9673;
wire n_8891;
wire n_12523;
wire n_7817;
wire n_3818;
wire n_8294;
wire n_11856;
wire n_6933;
wire n_4387;
wire n_7878;
wire n_8338;
wire n_4951;
wire n_12579;
wire n_9010;
wire n_8915;
wire n_4453;
wire n_4170;
wire n_6881;
wire n_11442;
wire n_7289;
wire n_5805;
wire n_7665;
wire n_8131;
wire n_11747;
wire n_9552;
wire n_3719;
wire n_7855;
wire n_11008;
wire n_3681;
wire n_10371;
wire n_11243;
wire n_9841;
wire n_12675;
wire n_13006;
wire n_9230;
wire n_12174;
wire n_7764;
wire n_4308;
wire n_12113;
wire n_12831;
wire n_10198;
wire n_8027;
wire n_6216;
wire n_10096;
wire n_3830;
wire n_10582;
wire n_11425;
wire n_10638;
wire n_8162;
wire n_6817;
wire n_7170;
wire n_7314;
wire n_9132;
wire n_11992;
wire n_6949;
wire n_6509;
wire n_5175;
wire n_3883;
wire n_7260;
wire n_8855;
wire n_10483;
wire n_11657;
wire n_4152;
wire n_12470;
wire n_8546;
wire n_9878;
wire n_11536;
wire n_11717;
wire n_9069;
wire n_8966;
wire n_12154;
wire n_7263;
wire n_8844;
wire n_8487;
wire n_5948;
wire n_4392;
wire n_4660;
wire n_3149;
wire n_5611;
wire n_10662;
wire n_6911;
wire n_3268;
wire n_9674;
wire n_11512;
wire n_11327;
wire n_8533;
wire n_4281;
wire n_4661;
wire n_12799;
wire n_4200;
wire n_3614;
wire n_3301;
wire n_8869;
wire n_5900;
wire n_3466;
wire n_4962;
wire n_9786;
wire n_6327;
wire n_8584;
wire n_11140;
wire n_8932;
wire n_9063;
wire n_8998;
wire n_6607;
wire n_9188;
wire n_9467;
wire n_9372;
wire n_3411;
wire n_10960;
wire n_11078;
wire n_4958;
wire n_9743;
wire n_4271;
wire n_7850;
wire n_7509;
wire n_11620;
wire n_7209;
wire n_5171;
wire n_3586;
wire n_12617;
wire n_6401;
wire n_5554;
wire n_6227;
wire n_12919;
wire n_8480;
wire n_9926;
wire n_7240;
wire n_10094;
wire n_12095;
wire n_10749;
wire n_11907;
wire n_4071;
wire n_4921;
wire n_12432;
wire n_12796;
wire n_8911;
wire n_11352;
wire n_5427;
wire n_5639;
wire n_7725;
wire n_8398;
wire n_3065;
wire n_4361;
wire n_10585;
wire n_5417;
wire n_8772;
wire n_12008;
wire n_4614;
wire n_12279;
wire n_9480;
wire n_8307;
wire n_10896;
wire n_8767;
wire n_9113;
wire n_9158;
wire n_12156;
wire n_3103;
wire n_11851;
wire n_4945;
wire n_4922;
wire n_4732;
wire n_7609;
wire n_8010;
wire n_7278;
wire n_11986;
wire n_12637;
wire n_12301;
wire n_9263;
wire n_8347;
wire n_11734;
wire n_7630;
wire n_11517;
wire n_11022;
wire n_11831;
wire n_10162;
wire n_12302;
wire n_8466;
wire n_6416;
wire n_4693;
wire n_5488;
wire n_12190;
wire n_9632;
wire n_10353;
wire n_8813;
wire n_8354;
wire n_4326;
wire n_6695;
wire n_8204;
wire n_3557;
wire n_7741;
wire n_5447;
wire n_5383;
wire n_4744;
wire n_6127;
wire n_7565;
wire n_11259;
wire n_11197;
wire n_11504;
wire n_9282;
wire n_2851;
wire n_4305;
wire n_5781;
wire n_7883;
wire n_6600;
wire n_10933;
wire n_12192;
wire n_7410;
wire n_12010;
wire n_12977;
wire n_4213;
wire n_2849;
wire n_10546;
wire n_7097;
wire n_12864;
wire n_3692;
wire n_9503;
wire n_6421;
wire n_10724;
wire n_5747;
wire n_7414;
wire n_11427;
wire n_10660;
wire n_7495;
wire n_9782;
wire n_5969;
wire n_9114;
wire n_8312;
wire n_9855;
wire n_4929;
wire n_8040;
wire n_11153;
wire n_9347;
wire n_4964;
wire n_9469;
wire n_9680;
wire n_9746;
wire n_10923;
wire n_6079;
wire n_4802;
wire n_6192;
wire n_9633;
wire n_12746;
wire n_10836;
wire n_6458;
wire n_10884;
wire n_4139;
wire n_3029;
wire n_6746;
wire n_8132;
wire n_12436;
wire n_4031;
wire n_7586;
wire n_10780;
wire n_9501;
wire n_12528;
wire n_7720;
wire n_6719;
wire n_12792;
wire n_5437;
wire n_9148;
wire n_11475;
wire n_5826;
wire n_7659;
wire n_3881;
wire n_12973;
wire n_11385;
wire n_6506;
wire n_4583;
wire n_6287;
wire n_6662;
wire n_8650;
wire n_12916;
wire n_10870;
wire n_12923;
wire n_9585;
wire n_10267;
wire n_8974;
wire n_10379;
wire n_4210;
wire n_5245;
wire n_7189;
wire n_8688;
wire n_4666;
wire n_2929;
wire n_3751;
wire n_10821;
wire n_10740;
wire n_8983;
wire n_10558;
wire n_6851;
wire n_8116;
wire n_12144;
wire n_9338;
wire n_12716;
wire n_6687;
wire n_10297;
wire n_2890;
wire n_6884;
wire n_8356;
wire n_8013;
wire n_9075;
wire n_3698;
wire n_3927;
wire n_4540;
wire n_3961;
wire n_6780;
wire n_6513;
wire n_12463;
wire n_12524;
wire n_4891;
wire n_8519;
wire n_7841;
wire n_10497;
wire n_6619;
wire n_10354;
wire n_11456;
wire n_8193;
wire n_5603;
wire n_10888;
wire n_6804;
wire n_3559;
wire n_9370;
wire n_11647;
wire n_12392;
wire n_12173;
wire n_9409;
wire n_5716;
wire n_3993;
wire n_10138;
wire n_4940;
wire n_6516;
wire n_10358;
wire n_5208;
wire n_7490;
wire n_3588;
wire n_7792;
wire n_10578;
wire n_6924;
wire n_4590;
wire n_7492;
wire n_12168;
wire n_12349;
wire n_10948;
wire n_5606;
wire n_4830;
wire n_12665;
wire n_5231;
wire n_8329;
wire n_5237;
wire n_7809;
wire n_11736;
wire n_4664;
wire n_9626;
wire n_3860;
wire n_8154;
wire n_12067;
wire n_5456;
wire n_3160;
wire n_12546;
wire n_7073;
wire n_11393;
wire n_10007;
wire n_5093;
wire n_10904;
wire n_10386;
wire n_6040;
wire n_3847;
wire n_4946;
wire n_9961;
wire n_4906;
wire n_5727;
wire n_3290;
wire n_9098;
wire n_4663;
wire n_5390;
wire n_7114;
wire n_5347;
wire n_11325;
wire n_9861;
wire n_2824;
wire n_3033;
wire n_3298;
wire n_6788;
wire n_4883;
wire n_11660;
wire n_2923;
wire n_4162;
wire n_10448;
wire n_3665;
wire n_5115;
wire n_12963;
wire n_3264;
wire n_6393;
wire n_9536;
wire n_8566;
wire n_12282;
wire n_8086;
wire n_12620;
wire n_2916;
wire n_8746;
wire n_11411;
wire n_6249;
wire n_4297;
wire n_5833;
wire n_6849;
wire n_12431;
wire n_3800;
wire n_9593;
wire n_9017;
wire n_5407;
wire n_11281;
wire n_11841;
wire n_4608;
wire n_11658;
wire n_5232;
wire n_9703;
wire n_2870;
wire n_7271;
wire n_3991;
wire n_12830;
wire n_3134;
wire n_11025;
wire n_6572;
wire n_12213;
wire n_4172;
wire n_4791;
wire n_6739;
wire n_11372;
wire n_4536;
wire n_10450;
wire n_12397;
wire n_5149;
wire n_5967;
wire n_7569;
wire n_5151;
wire n_7003;
wire n_9565;
wire n_7897;
wire n_4773;
wire n_7962;
wire n_8942;
wire n_5345;
wire n_5357;
wire n_4497;
wire n_6666;
wire n_10320;
wire n_4611;
wire n_8113;
wire n_6812;
wire n_4755;
wire n_5982;
wire n_4960;
wire n_10308;
wire n_2993;
wire n_8652;
wire n_3864;
wire n_4658;
wire n_5135;
wire n_2948;
wire n_7419;
wire n_11545;
wire n_12974;
wire n_5827;
wire n_9337;
wire n_5494;
wire n_11465;
wire n_4362;
wire n_4306;
wire n_6200;
wire n_11437;
wire n_3209;
wire n_3504;
wire n_10304;
wire n_7784;
wire n_11436;
wire n_4422;
wire n_10902;
wire n_8714;
wire n_6123;
wire n_10607;
wire n_6934;
wire n_7094;
wire n_7500;
wire n_11463;
wire n_10605;
wire n_3482;
wire n_11394;
wire n_6082;
wire n_10668;
wire n_8944;
wire n_12487;
wire n_9232;
wire n_12385;
wire n_9320;
wire n_10713;
wire n_4555;
wire n_11191;
wire n_2827;
wire n_9167;
wire n_10464;
wire n_5136;
wire n_7864;
wire n_5228;
wire n_10596;
wire n_10034;
wire n_11068;
wire n_7129;
wire n_3956;
wire n_5758;
wire n_5323;
wire n_7790;
wire n_3572;
wire n_4215;
wire n_6952;
wire n_4280;
wire n_7062;
wire n_3375;
wire n_10875;
wire n_4047;
wire n_12735;
wire n_9526;
wire n_5471;
wire n_8107;
wire n_7642;
wire n_5434;
wire n_12475;
wire n_9077;
wire n_5941;
wire n_7045;
wire n_12646;
wire n_5879;
wire n_11277;
wire n_3167;
wire n_11665;
wire n_5558;
wire n_11061;
wire n_9692;
wire n_5350;
wire n_3423;
wire n_9141;
wire n_5338;
wire n_7238;
wire n_11483;
wire n_3044;
wire n_12733;
wire n_7126;
wire n_9745;
wire n_5669;
wire n_9787;
wire n_3854;
wire n_8674;
wire n_11073;
wire n_12944;
wire n_7931;
wire n_10309;
wire n_12061;
wire n_12265;
wire n_3078;
wire n_12380;
wire n_8482;
wire n_11462;
wire n_8992;
wire n_13032;
wire n_6979;
wire n_11224;
wire n_10024;
wire n_9892;
wire n_6203;
wire n_7405;
wire n_10762;
wire n_7739;
wire n_10490;
wire n_3253;
wire n_8761;
wire n_7207;
wire n_9078;
wire n_8899;
wire n_11127;
wire n_4027;
wire n_7934;
wire n_9015;
wire n_7454;
wire n_9012;
wire n_4599;
wire n_12794;
wire n_5830;
wire n_6796;
wire n_3363;
wire n_4812;
wire n_9233;
wire n_12890;
wire n_9217;
wire n_5760;
wire n_6368;
wire n_3689;
wire n_6556;
wire n_4628;
wire n_11632;
wire n_10974;
wire n_9435;
wire n_5668;
wire n_3451;
wire n_4873;
wire n_5878;
wire n_8926;
wire n_5588;
wire n_4657;
wire n_2971;
wire n_11692;
wire n_11762;
wire n_5765;
wire n_11843;
wire n_3950;
wire n_9389;
wire n_11344;
wire n_4458;
wire n_11403;
wire n_6596;
wire n_12926;
wire n_4121;
wire n_5090;
wire n_6870;
wire n_10520;
wire n_7639;
wire n_12247;
wire n_12881;
wire n_4476;
wire n_5613;
wire n_10914;
wire n_10129;
wire n_4756;
wire n_3869;
wire n_4307;
wire n_5104;
wire n_5042;
wire n_4860;
wire n_4359;
wire n_11510;
wire n_10084;
wire n_7251;
wire n_10519;
wire n_7776;
wire n_12966;
wire n_6080;
wire n_10318;
wire n_7059;
wire n_8561;
wire n_10877;
wire n_8255;
wire n_7035;
wire n_10468;
wire n_5571;
wire n_11854;
wire n_8029;
wire n_12894;
wire n_10906;
wire n_4573;
wire n_5289;
wire n_6713;
wire n_4118;
wire n_5513;
wire n_6747;
wire n_12276;
wire n_6281;
wire n_4803;
wire n_5972;
wire n_10289;
wire n_9381;
wire n_4079;
wire n_4091;
wire n_9873;
wire n_11925;
wire n_12594;
wire n_10905;
wire n_5916;
wire n_5984;
wire n_7029;
wire n_7317;
wire n_13030;
wire n_9575;
wire n_5145;
wire n_12529;
wire n_11817;
wire n_3712;
wire n_6094;
wire n_2935;
wire n_6444;
wire n_11961;
wire n_12001;
wire n_5132;
wire n_5191;
wire n_10298;
wire n_12433;
wire n_6333;
wire n_10940;
wire n_6262;
wire n_12765;
wire n_3085;
wire n_5869;
wire n_8130;
wire n_5925;
wire n_9023;
wire n_12097;
wire n_6240;
wire n_10723;
wire n_5359;
wire n_6412;
wire n_9412;
wire n_5293;
wire n_7782;
wire n_7220;
wire n_10293;
wire n_11824;
wire n_4316;
wire n_3697;
wire n_10361;
wire n_7438;
wire n_11269;
wire n_11270;
wire n_9955;
wire n_10161;
wire n_10432;
wire n_7515;
wire n_11532;
wire n_7574;
wire n_12402;
wire n_4044;
wire n_12728;
wire n_4062;
wire n_6684;
wire n_4524;
wire n_4843;
wire n_8921;
wire n_3971;
wire n_10640;
wire n_11546;
wire n_7065;
wire n_10271;
wire n_11314;
wire n_5510;
wire n_6046;
wire n_7894;
wire n_7868;
wire n_9418;
wire n_6973;
wire n_2949;
wire n_9733;
wire n_5363;
wire n_7285;
wire n_8286;
wire n_5200;
wire n_9502;
wire n_5659;
wire n_5618;
wire n_6325;
wire n_2867;
wire n_9765;
wire n_9029;
wire n_11130;
wire n_3145;
wire n_10163;
wire n_3124;
wire n_6737;
wire n_12262;
wire n_6454;
wire n_4253;
wire n_5356;
wire n_6721;
wire n_8178;
wire n_5369;
wire n_11935;
wire n_5258;
wire n_12708;
wire n_5255;
wire n_10576;
wire n_2852;
wire n_9623;
wire n_11822;
wire n_10424;
wire n_12805;
wire n_7008;
wire n_11035;
wire n_8925;
wire n_10404;
wire n_3517;
wire n_3100;
wire n_8432;
wire n_6111;
wire n_10130;
wire n_12901;
wire n_7505;
wire n_3758;
wire n_3356;
wire n_2835;
wire n_8047;
wire n_6260;
wire n_7501;
wire n_10214;
wire n_3269;
wire n_12971;
wire n_5080;
wire n_11389;
wire n_6665;
wire n_9783;
wire n_7566;
wire n_7937;
wire n_12658;
wire n_7055;
wire n_3506;
wire n_3605;
wire n_12372;
wire n_8268;
wire n_11501;
wire n_12564;
wire n_8053;
wire n_11015;
wire n_5858;
wire n_5817;
wire n_10317;
wire n_6690;
wire n_9840;
wire n_3402;
wire n_5723;
wire n_10491;
wire n_5295;
wire n_6137;
wire n_10712;
wire n_4679;
wire n_4115;
wire n_6201;
wire n_9909;
wire n_10192;
wire n_7113;
wire n_12204;
wire n_4998;
wire n_2988;
wire n_10453;
wire n_11034;
wire n_8735;
wire n_11895;
wire n_7872;
wire n_12543;
wire n_10219;
wire n_5627;
wire n_12888;
wire n_4167;
wire n_8845;
wire n_7242;
wire n_5155;
wire n_3835;
wire n_6461;
wire n_8830;
wire n_12013;
wire n_11662;
wire n_5016;
wire n_3967;
wire n_7954;
wire n_6212;
wire n_3401;
wire n_6908;
wire n_3226;
wire n_7819;
wire n_6570;
wire n_12741;
wire n_8022;
wire n_9532;
wire n_8415;
wire n_9112;
wire n_6498;
wire n_3902;
wire n_10062;
wire n_4730;
wire n_7228;
wire n_9561;
wire n_6692;
wire n_8547;
wire n_10788;
wire n_11500;
wire n_6074;
wire n_10910;
wire n_7561;
wire n_6380;
wire n_3654;
wire n_10892;
wire n_10216;
wire n_9091;
wire n_5996;
wire n_8386;
wire n_8426;
wire n_9326;
wire n_8672;
wire n_11977;
wire n_10049;
wire n_5327;
wire n_7994;
wire n_9180;
wire n_10431;
wire n_11215;
wire n_8540;
wire n_6045;
wire n_9932;
wire n_4713;
wire n_5137;
wire n_6505;
wire n_9220;
wire n_9834;
wire n_3348;
wire n_7415;
wire n_9474;
wire n_7793;
wire n_5796;
wire n_7702;
wire n_9542;
wire n_11530;
wire n_7598;
wire n_6320;
wire n_6489;
wire n_6068;
wire n_12889;
wire n_3358;
wire n_8192;
wire n_5791;
wire n_8791;
wire n_9458;
wire n_10608;
wire n_4204;
wire n_9642;
wire n_5098;
wire n_6772;
wire n_6877;
wire n_9020;
wire n_9910;
wire n_6823;
wire n_6806;
wire n_7426;
wire n_11014;
wire n_5906;
wire n_8350;
wire n_11439;
wire n_12526;
wire n_9100;
wire n_11119;
wire n_11752;
wire n_4743;
wire n_8816;
wire n_3805;
wire n_7957;
wire n_3825;
wire n_8712;
wire n_8048;
wire n_6831;
wire n_3657;
wire n_10395;
wire n_4924;
wire n_3928;
wire n_12255;
wire n_9781;
wire n_8663;
wire n_4859;
wire n_7217;
wire n_9940;
wire n_12068;
wire n_10802;
wire n_6284;
wire n_7058;
wire n_4654;
wire n_6157;
wire n_5423;
wire n_7497;
wire n_8503;
wire n_6785;
wire n_8254;
wire n_6374;
wire n_8959;
wire n_9117;
wire n_6930;
wire n_12784;
wire n_9198;
wire n_4733;
wire n_6017;
wire n_3792;
wire n_11729;
wire n_8506;
wire n_4272;
wire n_11289;
wire n_3974;
wire n_3871;
wire n_11699;
wire n_7735;
wire n_3278;
wire n_8265;
wire n_8465;
wire n_8049;
wire n_12277;
wire n_4269;
wire n_4695;
wire n_6838;
wire n_11902;
wire n_12212;
wire n_12126;
wire n_5736;
wire n_6937;
wire n_12686;
wire n_6443;
wire n_3312;
wire n_6105;
wire n_10080;
wire n_7558;
wire n_12344;
wire n_12250;
wire n_8937;
wire n_12961;
wire n_5069;
wire n_7442;
wire n_10574;
wire n_8272;
wire n_5700;
wire n_6543;
wire n_3285;
wire n_9249;
wire n_11628;
wire n_10594;
wire n_11784;
wire n_12193;
wire n_3968;
wire n_9398;
wire n_5099;
wire n_11622;
wire n_4704;
wire n_4551;
wire n_11763;
wire n_5052;
wire n_6091;
wire n_11606;
wire n_2902;
wire n_12749;
wire n_4957;
wire n_6674;
wire n_10155;
wire n_6034;
wire n_7499;
wire n_4072;
wire n_9751;
wire n_5579;
wire n_8381;
wire n_7085;
wire n_12079;
wire n_4781;
wire n_9579;
wire n_3606;
wire n_11006;
wire n_10879;
wire n_6652;
wire n_7098;
wire n_5004;
wire n_6762;
wire n_7341;
wire n_7895;
wire n_4424;
wire n_11321;
wire n_8366;
wire n_10792;
wire n_8101;
wire n_7611;
wire n_9925;
wire n_10655;
wire n_7391;
wire n_3055;
wire n_3711;
wire n_10890;
wire n_12187;
wire n_12093;
wire n_3315;
wire n_5837;
wire n_3172;
wire n_3292;
wire n_4436;
wire n_6895;
wire n_3878;
wire n_7646;
wire n_4450;
wire n_8384;
wire n_9889;
wire n_5642;
wire n_12705;
wire n_3553;
wire n_7224;
wire n_5880;
wire n_8728;
wire n_6169;
wire n_11133;
wire n_4746;
wire n_12241;
wire n_12211;
wire n_7524;
wire n_5713;
wire n_6005;
wire n_10212;
wire n_8023;
wire n_8052;
wire n_11001;
wire n_7627;
wire n_9998;
wire n_11143;
wire n_10654;
wire n_3131;
wire n_5118;
wire n_5105;
wire n_9729;
wire n_3850;
wire n_4459;
wire n_11757;
wire n_8614;
wire n_2996;
wire n_5793;
wire n_5591;
wire n_7856;
wire n_4050;
wire n_9081;
wire n_7496;
wire n_12446;
wire n_12640;
wire n_3228;
wire n_12699;
wire n_9784;
wire n_5623;
wire n_12856;
wire n_10005;
wire n_10544;
wire n_10217;
wire n_12231;
wire n_5681;
wire n_4853;
wire n_11421;
wire n_11780;
wire n_12745;
wire n_9856;
wire n_9101;
wire n_7399;
wire n_12841;
wire n_6213;
wire n_8656;
wire n_10393;
wire n_6118;
wire n_5256;
wire n_2950;
wire n_11793;
wire n_12527;
wire n_7605;
wire n_11400;
wire n_5220;
wire n_12814;
wire n_5732;
wire n_8897;
wire n_3852;
wire n_9696;
wire n_12545;
wire n_5178;
wire n_11621;
wire n_4520;
wire n_6814;
wire n_7342;
wire n_12354;
wire n_4008;
wire n_8014;
wire n_9825;
wire n_5507;
wire n_10093;
wire n_8564;
wire n_11969;
wire n_7214;
wire n_7472;
wire n_12685;
wire n_5077;
wire n_10850;
wire n_12886;
wire n_8371;
wire n_10945;
wire n_5872;
wire n_11791;
wire n_3858;
wire n_7408;
wire n_8231;
wire n_9250;
wire n_10541;
wire n_6115;
wire n_4502;
wire n_9572;
wire n_6858;
wire n_12196;
wire n_10375;
wire n_11910;
wire n_11948;
wire n_8558;
wire n_3032;
wire n_4851;
wire n_5735;
wire n_9483;
wire n_10275;
wire n_9816;
wire n_12119;
wire n_9253;
wire n_8164;
wire n_7254;
wire n_6944;
wire n_7384;
wire n_9136;
wire n_3072;
wire n_3313;
wire n_3081;
wire n_7837;
wire n_8357;
wire n_10726;
wire n_9426;
wire n_3924;
wire n_8870;
wire n_9831;
wire n_4571;
wire n_8143;
wire n_11064;
wire n_6430;
wire n_6193;
wire n_10614;
wire n_5314;
wire n_6462;
wire n_8422;
wire n_12094;
wire n_12096;
wire n_3439;
wire n_9896;
wire n_9650;
wire n_12730;
wire n_10002;
wire n_5049;
wire n_6757;
wire n_6822;
wire n_4205;
wire n_5953;
wire n_7599;
wire n_5277;
wire n_4723;
wire n_5176;
wire n_11974;
wire n_12202;
wire n_6779;
wire n_6518;
wire n_9767;
wire n_6797;
wire n_11367;
wire n_4454;
wire n_7938;
wire n_8253;
wire n_4229;
wire n_5952;
wire n_4739;
wire n_12534;
wire n_5820;
wire n_5483;
wire n_12120;
wire n_3017;
wire n_9028;
wire n_9055;
wire n_5718;
wire n_10251;
wire n_11562;
wire n_11866;
wire n_6916;
wire n_3904;
wire n_5150;
wire n_11383;
wire n_12854;
wire n_8563;
wire n_9949;
wire n_4838;
wire n_2872;
wire n_5075;
wire n_11655;
wire n_12553;
wire n_7812;
wire n_12816;
wire n_4879;
wire n_5051;
wire n_11552;
wire n_9684;
wire n_3926;
wire n_6152;
wire n_10010;
wire n_9724;
wire n_3996;
wire n_4221;
wire n_8243;
wire n_10226;
wire n_11117;
wire n_8236;
wire n_11046;
wire n_8292;
wire n_2854;
wire n_11547;
wire n_12676;
wire n_4181;
wire n_5777;
wire n_7949;
wire n_8611;
wire n_7046;
wire n_12720;
wire n_4225;
wire n_10475;
wire n_10020;
wire n_9826;
wire n_5142;
wire n_3102;
wire n_10467;
wire n_4153;
wire n_5156;
wire n_5926;
wire n_3627;
wire n_8011;
wire n_9839;
wire n_4300;
wire n_9399;
wire n_3551;
wire n_4783;
wire n_12535;
wire n_2964;
wire n_3769;
wire n_12283;
wire n_12506;
wire n_6589;
wire n_7579;
wire n_4530;
wire n_4267;
wire n_8139;
wire n_12046;
wire n_8123;
wire n_3865;
wire n_3859;
wire n_3722;
wire n_7173;
wire n_10720;
wire n_7917;
wire n_5951;
wire n_7092;
wire n_10907;
wire n_6197;
wire n_6971;
wire n_9938;
wire n_8424;
wire n_9776;
wire n_8859;
wire n_11256;
wire n_7460;
wire n_9658;
wire n_11914;
wire n_3117;
wire n_9605;
wire n_11934;
wire n_12124;
wire n_10868;
wire n_11047;
wire n_3428;
wire n_9013;
wire n_2961;
wire n_8730;
wire n_9417;
wire n_8156;
wire n_9290;
wire n_9212;
wire n_3351;
wire n_3527;
wire n_9721;
wire n_12189;
wire n_10615;
wire n_7698;
wire n_12884;
wire n_7886;
wire n_6154;
wire n_7344;
wire n_6020;
wire n_2883;
wire n_9586;
wire n_7904;
wire n_12310;
wire n_11004;
wire n_4182;
wire n_10751;
wire n_12683;
wire n_2912;
wire n_11287;
wire n_4825;
wire n_5701;
wire n_10706;
wire n_4440;
wire n_10774;
wire n_11208;
wire n_4549;
wire n_12108;
wire n_12502;
wire n_3955;
wire n_9104;
wire n_7079;
wire n_10225;
wire n_11963;
wire n_10570;
wire n_9293;
wire n_11860;
wire n_5120;
wire n_8645;
wire n_10744;
wire n_11625;
wire n_5470;
wire n_4565;
wire n_7675;
wire n_4039;
wire n_10416;
wire n_3227;
wire n_3300;
wire n_4303;
wire n_4574;
wire n_7774;
wire n_5797;
wire n_7922;
wire n_8189;
wire n_8618;
wire n_6696;
wire n_11181;
wire n_11787;
wire n_4839;
wire n_5222;
wire n_8285;
wire n_5743;
wire n_4016;
wire n_9919;
wire n_10396;
wire n_8826;
wire n_6210;
wire n_10123;
wire n_5772;
wire n_12899;
wire n_3435;
wire n_8715;
wire n_3575;
wire n_12761;
wire n_8782;
wire n_6964;
wire n_10083;
wire n_5801;
wire n_6117;
wire n_4231;
wire n_8117;
wire n_12918;
wire n_11825;
wire n_6202;
wire n_7279;
wire n_3165;
wire n_7670;
wire n_11364;
wire n_4923;
wire n_12713;
wire n_3652;
wire n_12522;
wire n_12822;
wire n_9445;
wire n_4097;
wire n_6681;
wire n_5971;
wire n_4083;
wire n_11420;
wire n_12223;
wire n_11470;
wire n_4461;
wire n_3234;
wire n_5392;
wire n_8497;
wire n_12082;
wire n_9930;
wire n_6661;
wire n_8018;
wire n_3303;
wire n_6640;
wire n_12151;
wire n_3916;
wire n_7940;
wire n_11230;
wire n_12757;
wire n_3556;
wire n_7371;
wire n_6962;
wire n_4101;
wire n_10731;
wire n_11074;
wire n_10347;
wire n_11063;
wire n_6455;
wire n_3591;
wire n_7721;
wire n_9727;
wire n_4273;
wire n_3024;
wire n_7606;
wire n_5443;
wire n_12025;
wire n_3512;
wire n_5600;
wire n_4939;
wire n_5169;
wire n_6963;
wire n_10926;
wire n_6644;
wire n_4389;
wire n_6896;
wire n_3930;
wire n_12183;
wire n_4448;
wire n_11669;
wire n_10734;
wire n_6832;
wire n_8798;
wire n_7836;
wire n_12143;
wire n_6160;
wire n_7564;
wire n_11493;
wire n_12158;
wire n_7884;
wire n_8673;
wire n_10281;
wire n_6718;
wire n_9685;
wire n_11486;
wire n_8502;
wire n_6542;
wire n_10126;
wire n_10759;
wire n_11786;
wire n_10650;
wire n_11777;
wire n_6031;
wire n_5502;
wire n_5568;
wire n_9421;
wire n_8577;
wire n_11722;
wire n_7653;
wire n_10092;
wire n_10445;
wire n_5656;
wire n_8531;
wire n_8635;
wire n_6763;
wire n_4831;
wire n_5974;
wire n_9567;
wire n_3480;
wire n_3057;
wire n_3194;
wire n_6280;
wire n_9298;
wire n_11941;
wire n_10116;
wire n_6438;
wire n_10048;
wire n_9059;
wire n_12937;
wire n_8485;
wire n_3662;
wire n_6316;
wire n_7383;
wire n_4319;
wire n_5474;
wire n_8872;
wire n_8752;
wire n_9396;
wire n_4596;
wire n_5413;
wire n_6758;
wire n_12459;
wire n_7976;
wire n_9234;
wire n_9425;
wire n_12648;
wire n_10364;
wire n_5412;
wire n_9620;
wire n_3694;
wire n_6069;
wire n_10963;
wire n_5752;
wire n_10191;
wire n_6874;
wire n_4726;
wire n_4751;
wire n_4222;
wire n_8341;
wire n_12638;
wire n_2972;
wire n_6030;
wire n_3225;
wire n_8521;
wire n_8199;
wire n_11209;
wire n_12976;
wire n_6077;
wire n_8005;
wire n_11718;
wire n_4119;
wire n_3799;
wire n_7743;
wire n_4298;
wire n_5201;
wire n_6299;
wire n_9280;
wire n_9517;
wire n_4474;
wire n_6386;
wire n_9639;
wire n_9192;
wire n_12762;
wire n_9102;
wire n_5217;
wire n_10003;
wire n_10025;
wire n_8016;
wire n_10156;
wire n_8669;
wire n_5957;
wire n_12066;
wire n_11234;
wire n_3383;
wire n_12021;
wire n_8283;
wire n_13016;
wire n_10502;
wire n_3585;
wire n_2975;
wire n_7655;
wire n_5490;
wire n_5029;
wire n_8291;
wire n_4214;
wire n_8176;
wire n_10674;
wire n_5158;
wire n_4884;
wire n_6708;
wire n_7737;
wire n_10179;
wire n_7433;
wire n_11000;
wire n_12447;
wire n_11702;
wire n_4366;
wire n_10466;
wire n_12667;
wire n_4009;
wire n_12221;
wire n_7347;
wire n_8145;
wire n_9487;
wire n_10268;
wire n_4580;
wire n_6792;
wire n_12906;
wire n_7633;
wire n_12851;
wire n_6177;
wire n_5912;
wire n_11431;
wire n_10679;
wire n_12691;
wire n_7798;
wire n_10492;
wire n_11177;
wire n_12980;
wire n_4129;
wire n_4871;
wire n_12416;
wire n_4999;
wire n_13023;
wire n_11454;
wire n_6033;
wire n_9221;
wire n_12989;
wire n_11418;
wire n_5557;
wire n_7397;
wire n_12739;
wire n_7389;
wire n_12791;
wire n_5472;
wire n_7602;
wire n_2955;
wire n_4112;
wire n_8069;
wire n_6002;
wire n_4337;
wire n_5711;
wire n_4138;
wire n_7554;
wire n_5396;
wire n_7693;
wire n_5335;
wire n_8888;
wire n_12650;
wire n_12319;
wire n_6557;
wire n_7300;
wire n_9566;
wire n_12692;
wire n_12403;
wire n_9578;
wire n_8483;
wire n_8797;
wire n_5960;
wire n_8605;
wire n_8041;
wire n_4236;
wire n_9868;
wire n_3270;
wire n_5002;
wire n_11750;
wire n_3595;
wire n_11572;
wire n_7532;
wire n_11038;
wire n_11049;
wire n_9292;
wire n_10460;
wire n_5143;
wire n_7724;
wire n_4238;
wire n_12669;
wire n_11491;
wire n_6142;
wire n_6917;
wire n_7510;
wire n_11109;
wire n_5859;
wire n_10968;
wire n_3571;
wire n_8760;
wire n_4734;
wire n_8928;
wire n_10004;
wire n_10729;
wire n_11894;
wire n_8374;
wire n_8917;
wire n_6163;
wire n_4635;
wire n_10811;
wire n_3501;
wire n_7118;
wire n_8006;
wire n_11806;
wire n_4013;
wire n_3039;
wire n_9884;
wire n_6778;
wire n_6285;
wire n_7946;
wire n_8723;
wire n_9857;
wire n_11737;
wire n_12127;
wire n_11637;
wire n_6025;
wire n_8957;
wire n_12058;
wire n_7257;
wire n_4242;
wire n_11799;
wire n_10944;
wire n_11788;
wire n_6862;
wire n_6319;
wire n_7067;
wire n_4984;
wire n_3851;
wire n_10140;
wire n_3036;
wire n_12868;
wire n_12642;
wire n_10013;
wire n_12600;
wire n_7933;
wire n_3180;
wire n_5283;
wire n_8409;
wire n_9815;
wire n_9110;
wire n_7669;
wire n_5268;
wire n_10110;
wire n_6318;
wire n_10133;
wire n_8215;
wire n_11453;
wire n_11184;
wire n_8220;
wire n_9471;
wire n_9048;
wire n_4561;
wire n_7927;
wire n_11356;
wire n_6089;
wire n_3325;
wire n_3107;
wire n_4021;
wire n_8629;
wire n_3880;
wire n_5122;
wire n_7910;
wire n_11955;
wire n_12005;
wire n_6315;
wire n_10592;
wire n_3186;
wire n_7970;
wire n_4955;
wire n_10476;
wire n_8407;
wire n_5556;
wire n_5462;
wire n_4501;
wire n_3696;
wire n_12953;
wire n_11488;
wire n_12369;
wire n_9394;
wire n_3650;
wire n_8991;
wire n_12300;
wire n_5840;
wire n_13015;
wire n_6343;
wire n_10186;
wire n_11938;
wire n_3157;
wire n_11946;
wire n_9191;
wire n_11918;
wire n_9004;
wire n_12832;
wire n_6049;
wire n_6919;
wire n_7423;
wire n_7865;
wire n_6052;
wire n_11412;
wire n_10700;
wire n_5330;
wire n_4197;
wire n_4829;
wire n_7069;
wire n_12290;
wire n_6886;
wire n_2936;
wire n_12169;
wire n_8783;
wire n_6912;
wire n_8326;
wire n_10496;
wire n_11249;
wire n_10521;
wire n_12838;
wire n_5914;
wire n_11464;
wire n_12325;
wire n_8504;
wire n_10695;
wire n_8445;
wire n_11950;
wire n_11648;
wire n_8250;
wire n_10994;
wire n_11576;
wire n_4715;
wire n_5039;
wire n_9118;
wire n_6061;
wire n_4369;
wire n_12969;
wire n_5378;
wire n_10758;
wire n_8408;
wire n_4543;
wire n_10120;
wire n_11410;
wire n_4941;
wire n_11251;
wire n_7252;
wire n_5542;
wire n_4394;
wire n_9051;
wire n_7133;
wire n_6883;
wire n_10345;
wire n_5519;
wire n_12809;
wire n_9908;
wire n_12748;
wire n_3101;
wire n_3669;
wire n_6009;
wire n_7061;
wire n_8155;
wire n_5278;
wire n_8818;
wire n_11641;
wire n_11633;
wire n_12264;
wire n_7518;
wire n_9123;
wire n_12352;
wire n_5586;
wire n_10232;
wire n_3798;
wire n_4065;
wire n_6378;
wire n_8660;
wire n_5187;
wire n_4944;
wire n_12054;
wire n_5675;
wire n_4135;
wire n_8275;
wire n_9327;
wire n_6601;
wire n_5771;
wire n_7216;
wire n_6407;
wire n_11555;
wire n_9687;
wire n_8297;
wire n_9828;
wire n_6749;
wire n_11984;
wire n_6839;
wire n_10533;
wire n_9519;
wire n_10611;
wire n_7711;
wire n_12368;
wire n_2908;
wire n_10089;
wire n_12137;
wire n_3744;
wire n_4263;
wire n_11651;
wire n_7705;
wire n_2915;
wire n_10455;
wire n_8590;
wire n_3291;
wire n_6051;
wire n_4716;
wire n_12538;
wire n_4942;
wire n_6217;
wire n_6680;
wire n_5844;
wire n_12016;
wire n_7972;
wire n_6532;
wire n_3405;
wire n_4745;
wire n_6155;
wire n_6446;
wire n_8072;
wire n_12644;
wire n_6738;
wire n_6250;
wire n_7458;
wire n_7614;
wire n_7854;
wire n_12017;
wire n_7707;
wire n_10632;
wire n_11672;
wire n_11696;
wire n_3907;
wire n_8050;
wire n_6736;
wire n_5344;
wire n_6526;
wire n_8142;
wire n_10820;
wire n_10601;
wire n_4629;
wire n_6339;
wire n_2932;
wire n_12197;
wire n_2980;
wire n_5225;
wire n_8151;
wire n_6350;
wire n_7013;
wire n_12892;
wire n_3306;
wire n_5662;
wire n_4857;
wire n_3136;
wire n_9802;
wire n_9315;
wire n_9296;
wire n_8599;
wire n_10447;
wire n_4080;
wire n_12373;
wire n_12660;
wire n_4226;
wire n_4741;
wire n_10022;
wire n_5265;
wire n_4752;
wire n_11567;
wire n_10305;
wire n_12855;
wire n_3986;
wire n_4376;
wire n_10031;
wire n_12877;
wire n_5705;
wire n_4753;
wire n_12350;
wire n_10798;
wire n_12388;
wire n_4552;
wire n_7656;
wire n_10760;
wire n_11202;
wire n_3885;
wire n_6845;
wire n_9405;
wire n_12891;
wire n_9302;
wire n_7105;
wire n_5196;
wire n_12836;
wire n_5181;
wire n_11779;
wire n_11888;
wire n_10166;
wire n_2951;
wire n_3008;
wire n_3709;
wire n_6829;
wire n_11684;
wire n_11879;
wire n_5574;
wire n_11054;
wire n_5126;
wire n_6508;
wire n_9977;
wire n_9842;
wire n_3427;
wire n_9887;
wire n_4067;
wire n_5553;
wire n_4042;
wire n_4176;
wire n_7570;
wire n_8246;
wire n_11116;
wire n_9524;
wire n_11129;
wire n_7771;
wire n_4385;
wire n_3320;
wire n_7052;
wire n_5009;
wire n_7262;
wire n_5368;
wire n_9322;
wire n_11937;
wire n_10098;
wire n_10510;
wire n_10848;
wire n_10042;
wire n_8057;
wire n_9122;
wire n_8349;
wire n_5626;
wire n_9333;
wire n_8743;
wire n_6603;
wire n_6114;
wire n_9590;
wire n_6576;
wire n_3651;
wire n_7943;
wire n_4333;
wire n_7364;
wire n_3359;
wire n_8473;
wire n_10993;
wire n_10342;
wire n_7208;
wire n_12286;
wire n_6245;
wire n_12992;
wire n_2865;
wire n_10439;
wire n_11923;
wire n_12844;
wire n_5499;
wire n_6703;
wire n_4375;
wire n_3676;
wire n_4788;
wire n_4717;
wire n_4986;
wire n_5604;
wire n_9676;
wire n_3789;
wire n_3598;
wire n_10444;
wire n_7714;
wire n_9902;
wire n_10054;
wire n_12759;
wire n_8535;
wire n_10728;
wire n_4815;
wire n_9621;
wire n_7202;
wire n_9140;
wire n_4246;
wire n_3580;
wire n_9604;
wire n_7011;
wire n_4609;
wire n_7621;
wire n_5291;
wire n_8068;
wire n_10565;
wire n_10540;
wire n_12935;
wire n_9821;
wire n_11943;
wire n_10748;
wire n_5876;
wire n_10178;
wire n_11995;
wire n_11058;
wire n_6970;
wire n_11842;
wire n_12076;
wire n_12790;
wire n_12979;
wire n_5114;
wire n_6409;
wire n_6704;
wire n_6876;
wire n_4088;
wire n_12659;
wire n_7778;
wire n_3682;
wire n_4357;
wire n_3371;
wire n_9343;
wire n_7028;
wire n_12532;
wire n_4462;
wire n_4472;
wire n_3433;
wire n_7320;
wire n_6255;
wire n_7313;
wire n_7343;
wire n_5288;
wire n_5540;
wire n_5699;
wire n_11473;
wire n_7525;
wire n_7875;
wire n_3447;
wire n_5810;
wire n_11568;
wire n_3305;
wire n_4148;
wire n_4151;
wire n_12702;
wire n_3528;
wire n_6938;
wire n_12050;
wire n_4373;
wire n_12138;
wire n_5762;
wire n_4934;
wire n_5218;
wire n_8785;
wire n_9952;
wire n_12473;
wire n_13013;
wire n_10686;
wire n_8327;
wire n_12606;
wire n_9219;
wire n_7337;
wire n_6989;
wire n_8512;
wire n_4630;
wire n_5408;
wire n_10971;
wire n_4643;
wire n_4331;
wire n_6427;
wire n_4475;
wire n_3989;
wire n_7753;
wire n_10076;
wire n_4846;
wire n_3804;
wire n_4344;
wire n_11924;
wire n_12374;
wire n_8168;
wire n_3296;
wire n_8392;
wire n_7038;
wire n_12967;
wire n_4683;
wire n_5366;
wire n_10132;
wire n_10282;
wire n_9872;
wire n_12956;
wire n_6360;
wire n_11203;
wire n_3116;
wire n_13026;
wire n_9553;
wire n_10900;
wire n_3602;
wire n_2967;
wire n_6146;
wire n_10616;
wire n_9447;
wire n_6270;
wire n_11585;
wire n_9150;
wire n_3706;
wire n_5477;
wire n_9592;
wire n_5451;
wire n_9984;
wire n_12695;
wire n_3923;
wire n_11416;
wire n_4696;
wire n_11526;
wire n_3441;
wire n_11742;
wire n_12179;
wire n_8419;
wire n_11809;
wire n_5086;
wire n_9814;
wire n_10858;
wire n_12038;
wire n_5901;
wire n_6353;
wire n_4011;
wire n_10769;
wire n_9446;
wire n_4905;
wire n_10023;
wire n_10211;
wire n_11877;
wire n_2825;
wire n_3643;
wire n_4876;
wire n_6345;
wire n_12105;
wire n_9461;
wire n_10772;
wire n_9793;
wire n_6691;
wire n_3748;
wire n_8997;
wire n_4278;
wire n_3142;
wire n_4623;
wire n_4910;
wire n_12360;
wire n_12297;
wire n_4410;
wire n_3370;
wire n_12952;
wire n_9874;
wire n_7392;
wire n_5053;
wire n_7912;
wire n_8245;
wire n_6239;
wire n_4553;
wire n_6803;
wire n_10446;
wire n_11735;
wire n_7919;
wire n_3978;
wire n_6340;
wire n_7583;
wire n_4809;
wire n_8109;
wire n_5226;
wire n_7657;
wire n_3660;
wire n_7995;
wire n_11405;
wire n_6048;
wire n_5867;
wire n_8985;
wire n_5079;
wire n_5590;
wire n_10331;
wire n_12103;
wire n_6773;
wire n_9403;
wire n_3833;
wire n_5632;
wire n_8390;
wire n_11480;
wire n_11874;
wire n_4841;
wire n_12115;
wire n_6336;
wire n_3814;
wire n_8463;
wire n_7041;
wire n_7802;
wire n_2838;
wire n_4842;
wire n_4911;
wire n_4340;
wire n_7370;
wire n_3513;
wire n_3133;
wire n_10181;
wire n_10074;
wire n_9731;
wire n_5660;
wire n_11104;
wire n_4645;
wire n_7557;
wire n_11862;
wire n_2992;
wire n_11952;
wire n_6174;
wire n_3725;
wire n_4920;
wire n_12828;
wire n_4972;
wire n_6023;
wire n_6776;
wire n_3128;
wire n_5426;
wire n_9947;
wire n_6463;
wire n_7896;
wire n_9699;
wire n_6372;
wire n_10962;
wire n_11037;
wire n_9305;
wire n_10481;
wire n_7176;
wire n_12003;
wire n_10220;
wire n_10381;
wire n_8517;
wire n_12332;
wire n_5625;
wire n_5778;
wire n_6396;
wire n_3355;
wire n_9218;
wire n_10642;
wire n_11556;
wire n_6669;
wire n_3917;
wire n_9096;
wire n_10634;
wire n_3942;
wire n_10170;
wire n_10142;
wire n_10569;
wire n_12326;
wire n_3765;
wire n_5531;
wire n_9534;
wire n_7826;
wire n_3000;
wire n_5429;
wire n_11044;
wire n_3108;
wire n_3111;
wire n_5818;
wire n_5646;
wire n_6940;
wire n_4557;
wire n_5248;
wire n_11042;
wire n_12141;
wire n_4451;
wire n_6394;
wire n_2875;
wire n_9164;
wire n_9546;
wire n_3844;
wire n_3280;
wire n_12622;
wire n_11226;
wire n_4054;
wire n_5448;
wire n_3471;
wire n_5432;
wire n_7590;
wire n_9358;
wire n_3205;
wire n_11985;
wire n_2848;
wire n_5160;
wire n_11328;
wire n_3003;
wire n_3610;
wire n_8208;
wire n_6995;
wire n_7185;
wire n_10127;
wire n_3564;
wire n_11525;
wire n_3988;
wire n_9730;
wire n_6254;
wire n_6161;
wire n_9066;
wire n_10800;
wire n_11020;
wire n_3457;
wire n_9185;
wire n_9318;
wire n_10374;
wire n_7987;
wire n_8134;
wire n_4324;
wire n_4821;
wire n_10328;
wire n_8631;
wire n_5445;
wire n_3630;
wire n_8694;
wire n_11892;
wire n_8965;
wire n_8647;
wire n_11013;
wire n_3271;
wire n_12343;
wire n_7332;
wire n_6660;
wire n_4771;
wire n_5719;
wire n_7225;
wire n_10529;
wire n_12396;
wire n_6128;
wire n_4086;
wire n_7037;
wire n_11820;
wire n_11587;
wire n_4814;
wire n_12081;
wire n_10314;
wire n_3648;
wire n_5749;
wire n_11697;
wire n_12296;
wire n_8427;
wire n_3075;
wire n_3173;
wire n_9339;
wire n_5332;
wire n_9596;
wire n_5108;
wire n_7409;
wire n_4692;
wire n_3031;
wire n_10006;
wire n_10667;
wire n_7258;
wire n_7432;
wire n_9156;
wire n_11242;
wire n_11441;
wire n_3701;
wire n_11916;
wire n_11435;
wire n_12804;
wire n_11471;
wire n_3243;
wire n_6334;
wire n_3385;
wire n_10346;
wire n_8984;
wire n_6848;
wire n_10539;
wire n_8345;
wire n_10414;
wire n_4708;
wire n_6321;
wire n_7765;
wire n_9708;
wire n_9268;
wire n_8764;
wire n_6794;
wire n_10340;
wire n_4826;
wire n_3343;
wire n_10245;
wire n_11644;
wire n_7761;
wire n_7197;
wire n_12466;
wire n_12701;
wire n_5489;
wire n_12106;
wire n_6400;
wire n_3767;
wire n_12560;
wire n_2873;
wire n_4589;
wire n_9097;
wire n_5057;
wire n_10280;
wire n_12895;
wire n_11432;
wire n_4578;
wire n_12342;
wire n_6705;
wire n_7775;
wire n_9636;
wire n_10256;
wire n_7619;
wire n_12125;
wire n_2847;
wire n_3221;
wire n_5436;
wire n_5907;
wire n_11120;
wire n_5072;
wire n_11391;
wire n_3629;
wire n_3021;
wire n_6044;
wire n_11164;
wire n_11527;
wire n_3674;
wire n_5286;
wire n_8083;
wire n_3502;
wire n_8853;
wire n_3098;
wire n_11371;
wire n_6495;
wire n_5013;
wire n_10917;
wire n_7403;
wire n_6902;
wire n_6470;
wire n_9473;
wire n_3015;
wire n_10727;
wire n_11591;
wire n_10145;
wire n_12341;
wire n_9560;
wire n_5569;
wire n_8038;
wire n_10938;
wire n_9175;
wire n_8711;
wire n_10976;
wire n_5439;
wire n_8229;
wire n_8949;
wire n_10612;
wire n_5619;
wire n_4147;
wire n_6481;
wire n_9810;
wire n_3607;
wire n_4925;
wire n_7548;
wire n_9244;
wire n_9584;
wire n_12047;
wire n_6534;
wire n_11460;
wire n_4974;
wire n_8567;
wire n_10797;
wire n_9439;
wire n_11915;
wire n_4932;
wire n_4510;
wire n_8655;
wire n_9235;
wire n_6181;
wire n_3276;
wire n_6728;
wire n_8705;
wire n_11642;
wire n_9043;
wire n_9768;
wire n_11306;
wire n_3787;
wire n_5119;
wire n_9037;
wire n_5715;
wire n_9085;
wire n_12434;
wire n_8085;
wire n_8777;
wire n_6133;
wire n_11891;
wire n_8852;
wire n_9264;
wire n_6528;
wire n_10114;
wire n_7604;
wire n_7407;
wire n_8185;
wire n_3827;
wire n_12998;
wire n_3354;
wire n_10845;
wire n_4447;
wire n_8513;
wire n_6670;
wire n_12248;
wire n_6774;
wire n_8365;
wire n_11007;
wire n_4285;
wire n_5887;
wire n_4651;
wire n_6741;
wire n_7424;
wire n_11557;
wire n_12405;
wire n_6038;
wire n_4818;
wire n_7727;
wire n_4514;
wire n_4800;
wire n_10599;
wire n_11231;
wire n_3960;
wire n_9550;
wire n_9836;
wire n_3248;
wire n_6282;
wire n_9929;
wire n_12134;
wire n_8035;
wire n_8505;
wire n_11399;
wire n_11092;
wire n_4433;
wire n_11163;
wire n_8874;
wire n_11542;
wire n_2879;
wire n_10008;
wire n_3153;
wire n_6700;
wire n_7334;
wire n_7684;
wire n_7755;
wire n_8098;
wire n_4341;
wire n_10623;
wire n_9187;
wire n_11276;
wire n_4312;
wire n_3399;
wire n_10511;
wire n_5932;
wire n_12770;
wire n_13011;
wire n_6178;
wire n_11575;
wire n_10503;
wire n_6234;
wire n_11732;
wire n_6012;
wire n_4633;
wire n_9406;
wire n_3838;
wire n_10857;
wire n_9342;
wire n_4277;
wire n_7787;
wire n_4140;
wire n_8067;
wire n_3675;
wire n_12421;
wire n_5092;
wire n_10708;
wire n_3387;
wire n_7849;
wire n_5186;
wire n_12550;
wire n_11045;
wire n_7367;
wire n_8619;
wire n_9851;
wire n_9559;
wire n_11993;
wire n_11508;
wire n_12755;
wire n_8679;
wire n_9806;
wire n_8644;
wire n_12306;
wire n_12965;
wire n_11982;
wire n_10516;
wire n_4662;
wire n_3779;
wire n_6715;
wire n_11395;
wire n_5828;
wire n_2831;
wire n_11634;
wire n_7200;
wire n_9860;
wire n_4882;
wire n_4993;
wire n_11887;
wire n_11301;
wire n_7582;
wire n_4832;
wire n_4207;
wire n_4545;
wire n_3037;
wire n_6337;
wire n_4868;
wire n_8923;
wire n_8970;
wire n_10119;
wire n_8332;
wire n_10548;
wire n_11010;
wire n_11408;
wire n_8632;
wire n_6770;
wire n_7745;
wire n_6743;
wire n_8876;
wire n_3925;
wire n_10733;
wire n_10547;
wire n_11670;
wire n_5238;
wire n_10067;
wire n_4059;
wire n_8856;
wire n_12603;
wire n_11604;
wire n_9240;
wire n_4595;
wire n_7877;
wire n_11506;
wire n_11666;
wire n_8945;
wire n_11503;
wire n_8918;
wire n_7799;
wire n_6682;
wire n_5054;
wire n_7673;
wire n_11857;
wire n_5631;
wire n_8028;
wire n_6539;
wire n_7243;
wire n_7179;
wire n_9345;
wire n_4063;
wire n_5399;
wire n_6617;
wire n_6314;
wire n_10222;
wire n_11193;
wire n_11293;
wire n_12439;
wire n_3592;
wire n_5694;
wire n_4650;
wire n_4888;
wire n_7274;
wire n_8774;
wire n_5326;
wire n_12072;
wire n_8779;
wire n_3394;
wire n_8968;
wire n_4874;
wire n_7608;
wire n_3793;
wire n_8404;
wire n_4669;
wire n_4339;
wire n_6595;
wire n_12558;
wire n_12244;
wire n_12199;
wire n_11214;
wire n_4041;
wire n_5459;
wire n_2858;
wire n_7738;
wire n_4060;
wire n_9223;
wire n_9499;
wire n_10647;
wire n_2895;
wire n_11362;
wire n_11288;
wire n_11409;
wire n_5528;
wire n_3097;
wire n_11027;
wire n_12996;
wire n_5391;
wire n_12873;
wire n_8073;
wire n_4541;
wire n_3824;
wire n_5422;
wire n_7785;
wire n_6385;
wire n_6289;
wire n_3388;
wire n_12591;
wire n_5267;
wire n_4494;
wire n_3059;
wire n_10581;
wire n_5523;
wire n_3465;
wire n_4796;
wire n_7373;
wire n_9576;
wire n_9120;
wire n_3589;
wire n_10097;
wire n_10405;
wire n_6186;
wire n_4799;
wire n_5153;
wire n_12726;
wire n_9651;
wire n_12833;
wire n_6257;
wire n_12690;
wire n_3449;
wire n_11031;
wire n_9386;
wire n_2989;
wire n_11285;
wire n_10813;
wire n_6852;
wire n_6346;
wire n_11346;
wire n_12618;
wire n_4775;
wire n_9779;
wire n_5044;
wire n_5809;
wire n_12414;
wire n_11513;
wire n_5365;
wire n_2933;
wire n_7587;
wire n_5045;
wire n_4381;
wire n_4266;
wire n_11250;
wire n_7874;
wire n_3886;
wire n_11340;
wire n_5354;
wire n_4455;
wire n_6274;
wire n_7372;
wire n_7760;
wire n_10588;
wire n_4248;
wire n_9635;
wire n_5915;
wire n_6818;
wire n_9444;
wire n_10943;
wire n_11190;
wire n_5452;
wire n_7226;
wire n_8930;
wire n_4754;
wire n_7057;
wire n_12736;
wire n_7685;
wire n_8031;
wire n_11818;
wire n_8750;
wire n_4554;
wire n_5595;
wire n_6609;
wire n_4845;
wire n_6753;
wire n_6815;
wire n_9364;
wire n_9512;
wire n_9581;
wire n_3053;
wire n_9317;
wire n_3893;
wire n_8593;
wire n_3548;
wire n_4585;
wire n_7730;
wire n_8509;
wire n_9314;
wire n_9459;
wire n_8405;
wire n_3334;
wire n_9549;
wire n_11564;
wire n_10641;
wire n_7913;
wire n_4383;
wire n_11719;
wire n_8492;
wire n_6764;
wire n_5535;
wire n_9275;
wire n_3875;
wire n_10210;
wire n_5370;
wire n_11944;
wire n_7706;
wire n_7891;
wire n_6391;
wire n_4003;
wire n_11785;
wire n_8088;
wire n_5372;
wire n_5299;
wire n_5594;
wire n_4301;
wire n_11754;
wire n_4586;
wire n_4048;
wire n_9865;
wire n_6471;
wire n_11075;
wire n_11511;
wire n_12981;
wire n_6627;
wire n_3777;
wire n_10027;
wire n_5761;
wire n_10263;
wire n_10722;
wire n_13005;
wire n_11771;
wire n_4784;
wire n_7203;
wire n_8429;
wire n_8854;
wire n_9757;
wire n_2999;
wire n_7512;
wire n_5550;
wire n_12333;
wire n_11912;
wire n_5082;
wire n_4046;
wire n_9656;
wire n_10426;
wire n_11284;
wire n_5209;
wire n_3537;
wire n_7215;
wire n_10246;
wire n_3080;
wire n_6636;
wire n_4199;
wire n_13004;
wire n_10617;
wire n_5929;
wire n_3362;
wire n_10909;
wire n_5559;
wire n_3105;
wire n_12694;
wire n_5478;
wire n_11298;
wire n_7388;
wire n_7694;
wire n_6243;
wire n_6488;
wire n_4286;
wire n_9629;
wire n_11185;
wire n_5102;
wire n_3274;
wire n_3041;
wire n_11498;
wire n_6022;
wire n_8686;
wire n_6457;
wire n_10299;
wire n_4470;
wire n_2816;
wire n_12904;
wire n_7982;
wire n_11384;
wire n_10763;
wire n_3616;
wire n_10494;
wire n_4058;
wire n_3664;
wire n_8773;
wire n_10743;
wire n_8225;
wire n_8583;
wire n_4188;
wire n_6867;
wire n_3913;
wire n_8887;
wire n_9556;
wire n_3417;
wire n_5868;
wire n_6230;
wire n_4034;
wire n_6538;
wire n_12810;
wire n_9259;
wire n_9995;
wire n_12820;
wire n_6633;
wire n_9371;
wire n_8080;
wire n_11496;
wire n_6187;
wire n_3327;
wire n_6172;
wire n_10050;
wire n_5275;
wire n_10702;
wire n_4689;
wire n_5071;
wire n_3067;
wire n_7311;
wire n_5989;
wire n_8964;
wire n_11768;
wire n_12085;
wire n_3237;
wire n_9008;
wire n_6574;
wire n_11388;
wire n_11683;
wire n_8929;
wire n_8539;
wire n_6395;
wire n_4402;
wire n_9484;
wire n_8745;
wire n_4239;
wire n_6854;
wire n_3400;
wire n_7996;
wire n_6233;
wire n_4550;
wire n_6456;
wire n_8776;
wire n_8588;
wire n_8554;
wire n_9319;
wire n_3382;
wire n_11748;
wire n_7488;
wire n_3574;
wire n_5227;
wire n_9442;
wire n_10165;
wire n_7198;
wire n_4201;
wire n_10366;
wire n_12207;
wire n_8802;
wire n_9587;
wire n_6784;
wire n_6168;
wire n_9904;
wire n_9157;
wire n_8431;
wire n_8453;
wire n_3316;
wire n_6766;
wire n_5242;
wire n_3099;
wire n_8955;
wire n_3704;
wire n_12510;
wire n_8634;
wire n_3603;
wire n_4123;
wire n_6330;
wire n_5520;
wire n_8896;
wire n_3633;
wire n_4479;
wire n_7950;
wire n_7249;
wire n_9713;
wire n_11210;
wire n_9452;
wire n_10104;
wire n_5947;
wire n_7336;
wire n_4416;
wire n_8837;
wire n_3372;
wire n_7031;
wire n_4539;
wire n_8907;
wire n_6799;
wire n_10115;
wire n_8015;
wire n_10397;
wire n_9974;
wire n_10398;
wire n_5920;
wire n_6672;
wire n_6149;
wire n_8256;
wire n_10065;
wire n_11156;
wire n_10243;
wire n_10087;
wire n_12628;
wire n_7142;
wire n_3230;
wire n_11598;
wire n_5808;
wire n_3342;
wire n_6054;
wire n_7089;
wire n_11176;
wire n_12687;
wire n_4682;
wire n_7916;
wire n_12260;
wire n_5353;
wire n_3708;
wire n_5294;
wire n_6450;
wire n_12445;
wire n_3729;
wire n_8074;
wire n_12878;
wire n_4978;
wire n_4690;
wire n_10174;
wire n_12281;
wire n_10266;
wire n_12879;
wire n_10509;
wire n_12355;
wire n_4437;
wire n_5458;
wire n_3861;
wire n_5617;
wire n_4736;
wire n_7042;
wire n_3780;
wire n_8778;
wire n_8039;
wire n_5244;
wire n_10415;
wire n_6523;
wire n_5382;
wire n_8065;
wire n_6107;
wire n_9634;
wire n_3957;
wire n_12601;
wire n_11893;
wire n_12004;
wire n_11828;
wire n_6775;
wire n_5274;
wire n_10873;
wire n_3848;
wire n_8194;
wire n_12291;
wire n_4284;
wire n_11582;
wire n_8207;
wire n_3919;
wire n_10106;
wire n_12474;
wire n_9241;
wire n_6232;
wire n_6445;
wire n_10422;
wire n_10736;
wire n_7181;
wire n_6134;
wire n_5384;
wire n_9903;
wire n_3608;
wire n_8582;
wire n_10378;
wire n_6056;
wire n_8537;
wire n_6932;
wire n_7036;
wire n_4513;
wire n_3233;
wire n_3829;
wire n_9615;
wire n_3177;
wire n_4053;
wire n_8951;
wire n_7759;
wire n_9600;
wire n_11095;
wire n_7818;
wire n_11180;
wire n_9748;
wire n_9945;
wire n_5125;
wire n_12024;
wire n_4040;
wire n_9927;
wire n_5587;
wire n_6855;
wire n_11876;
wire n_5789;
wire n_8217;
wire n_10046;
wire n_3123;
wire n_5787;
wire n_6585;
wire n_6369;
wire n_5056;
wire n_10954;
wire n_10388;
wire n_8437;
wire n_5249;
wire n_3393;
wire n_8849;
wire n_7447;
wire n_10659;
wire n_7944;
wire n_5198;
wire n_11709;
wire n_5360;
wire n_10804;
wire n_7455;
wire n_5233;
wire n_4887;
wire n_5829;
wire n_4617;
wire n_9295;
wire n_5269;
wire n_3520;
wire n_11602;
wire n_11304;
wire n_6252;
wire n_12934;
wire n_5866;
wire n_6493;
wire n_8568;
wire n_10239;
wire n_12723;
wire n_7947;
wire n_12428;
wire n_4005;
wire n_10841;
wire n_12857;
wire n_9916;
wire n_4904;
wire n_8980;
wire n_5899;
wire n_11630;
wire n_7629;
wire n_8051;
wire n_4792;
wire n_7104;
wire n_3578;
wire n_8716;
wire n_11461;
wire n_3812;
wire n_9844;
wire n_7601;
wire n_4980;
wire n_11135;
wire n_12520;
wire n_11994;
wire n_12457;
wire n_12743;
wire n_6026;
wire n_4290;
wire n_5247;
wire n_7757;
wire n_8030;
wire n_9316;
wire n_9663;
wire n_10168;
wire n_5865;
wire n_13019;
wire n_10075;
wire n_3727;
wire n_5317;
wire n_6544;
wire n_3774;
wire n_10068;
wire n_11596;
wire n_10276;
wire n_3093;
wire n_12533;
wire n_8749;
wire n_3061;
wire n_11024;
wire n_7138;
wire n_7290;
wire n_8544;
wire n_8249;
wire n_12555;
wire n_9628;
wire n_6679;
wire n_8496;
wire n_9789;
wire n_4956;
wire n_5380;
wire n_5924;
wire n_3182;
wire n_12839;
wire n_7625;
wire n_5822;
wire n_10495;
wire n_9299;
wire n_6259;
wire n_12251;
wire n_4947;
wire n_7284;
wire n_11246;
wire n_11715;
wire n_4656;
wire n_12766;
wire n_12983;
wire n_3896;
wire n_6390;
wire n_3958;
wire n_12573;
wire n_12945;
wire n_3450;
wire n_11970;
wire n_4729;
wire n_5786;
wire n_4987;
wire n_5182;
wire n_4971;
wire n_11113;
wire n_12451;
wire n_7971;
wire n_3174;
wire n_12542;
wire n_12376;
wire n_9022;
wire n_10927;
wire n_6630;
wire n_12585;
wire n_10704;
wire n_3398;
wire n_5658;
wire n_3408;
wire n_11613;
wire n_5388;
wire n_4823;
wire n_9427;
wire n_4875;
wire n_3432;
wire n_6279;
wire n_8698;
wire n_8695;
wire n_9344;
wire n_12530;
wire n_8751;
wire n_10603;
wire n_12875;
wire n_3090;
wire n_11085;
wire n_3762;
wire n_6813;
wire n_9764;
wire n_12808;
wire n_5564;
wire n_11294;
wire n_13024;
wire n_8273;
wire n_11021;
wire n_9242;
wire n_9498;
wire n_8442;
wire n_7106;
wire n_8472;
wire n_9535;
wire n_6042;
wire n_7644;
wire n_12494;
wire n_10011;
wire n_6057;
wire n_4137;
wire n_7529;
wire n_8986;
wire n_6675;
wire n_11905;
wire n_12488;
wire n_4529;
wire n_4323;
wire n_3034;
wire n_12229;
wire n_6476;
wire n_8200;
wire n_3972;
wire n_10055;
wire n_7907;
wire n_10982;
wire n_8188;
wire n_11926;
wire n_11951;
wire n_8528;
wire n_12219;
wire n_6207;
wire n_5539;
wire n_10764;
wire n_6268;
wire n_6878;
wire n_6286;
wire n_9088;
wire n_3308;
wire n_12630;
wire n_6524;
wire n_10787;
wire n_5036;
wire n_12910;
wire n_5547;
wire n_4772;
wire n_3467;
wire n_6225;
wire n_4322;
wire n_8920;
wire n_8267;
wire n_12758;
wire n_10972;
wire n_7297;
wire n_6291;
wire n_2830;
wire n_5893;
wire n_4354;
wire n_4653;
wire n_12883;
wire n_9734;
wire n_9505;
wire n_9664;
wire n_12672;
wire n_7199;
wire n_5273;
wire n_10262;
wire n_10826;
wire n_8360;
wire n_4677;
wire n_3901;
wire n_8036;
wire n_9510;
wire n_5261;
wire n_11423;
wire n_6520;
wire n_7853;
wire n_7648;
wire n_9413;
wire n_9888;
wire n_3757;
wire n_8393;
wire n_11484;
wire n_8821;
wire n_11760;
wire n_9863;
wire n_12946;
wire n_10881;
wire n_8160;
wire n_9199;
wire n_3381;
wire n_11370;
wire n_5193;
wire n_10707;
wire n_9014;
wire n_10204;
wire n_9411;
wire n_12394;
wire n_12613;
wire n_12706;
wire n_4909;
wire n_11909;
wire n_9336;
wire n_9360;
wire n_10556;
wire n_9543;
wire n_2965;
wire n_3635;
wire n_6024;
wire n_7866;
wire n_5022;
wire n_5005;
wire n_2814;
wire n_3882;
wire n_3046;
wire n_7487;
wire n_10717;
wire n_6425;
wire n_5993;
wire n_3826;
wire n_3211;
wire n_12978;
wire n_12253;
wire n_3121;
wire n_7638;
wire n_8833;
wire n_5703;
wire n_8240;
wire n_12450;
wire n_4634;
wire n_3337;
wire n_7988;
wire n_9404;
wire n_8579;
wire n_6432;
wire n_5534;
wire n_9678;
wire n_3204;
wire n_12444;
wire n_8258;
wire n_9854;
wire n_7259;
wire n_11071;
wire n_11979;
wire n_8626;
wire n_12289;
wire n_6540;
wire n_6955;
wire n_9481;
wire n_5174;
wire n_10862;
wire n_4952;
wire n_12583;
wire n_5157;
wire n_3005;
wire n_4380;
wire n_9672;
wire n_3129;
wire n_9893;
wire n_4126;
wire n_7237;
wire n_8935;
wire n_11928;
wire n_5087;
wire n_3043;
wire n_12590;
wire n_3802;
wire n_4506;
wire n_6388;
wire n_12596;
wire n_10240;
wire n_5904;
wire n_9478;
wire n_4880;
wire n_11792;
wire n_9266;
wire n_9813;
wire n_12551;
wire n_6760;
wire n_8009;
wire n_11329;
wire n_3892;
wire n_4896;
wire n_5620;
wire n_5061;
wire n_5750;
wire n_7063;
wire n_5572;
wire n_10338;
wire n_10205;
wire n_12034;
wire n_3219;
wire n_11573;
wire n_11703;
wire n_9042;
wire n_2906;
wire n_4943;
wire n_11671;
wire n_8012;
wire n_11445;
wire n_7576;
wire n_9506;
wire n_8608;
wire n_8008;
wire n_12498;
wire n_10285;
wire n_3023;
wire n_6795;
wire n_5881;
wire n_8079;
wire n_6664;
wire n_12228;
wire n_5815;
wire n_12378;
wire n_11832;
wire n_6261;
wire n_4193;
wire n_5873;
wire n_4075;
wire n_9666;
wire n_3104;
wire n_10112;
wire n_6487;
wire n_9146;
wire n_4737;
wire n_7734;
wire n_6729;
wire n_3647;
wire n_10056;
wire n_9862;
wire n_5755;
wire n_10283;
wire n_9274;
wire n_2819;
wire n_8702;
wire n_5949;
wire n_10469;
wire n_5195;
wire n_7483;
wire n_3609;
wire n_4136;
wire n_6608;
wire n_7858;
wire n_9619;
wire n_12742;
wire n_4393;
wire n_7385;
wire n_11088;
wire n_12423;
wire n_10618;
wire n_3720;
wire n_8576;
wire n_9508;
wire n_4535;
wire n_10105;
wire n_7668;
wire n_13008;
wire n_8662;
wire n_4522;
wire n_6663;
wire n_4794;
wire n_5955;
wire n_7476;
wire n_3959;
wire n_7327;
wire n_5763;
wire n_6656;
wire n_8436;
wire n_11154;
wire n_9987;
wire n_8124;
wire n_8148;
wire n_12518;
wire n_8033;
wire n_6843;
wire n_12764;
wire n_3140;
wire n_7953;
wire n_8343;
wire n_5246;
wire n_5964;
wire n_11065;
wire n_12417;
wire n_3724;
wire n_8118;
wire n_12209;
wire n_12882;
wire n_3011;
wire n_7266;
wire n_5164;
wire n_11449;
wire n_4196;
wire n_6969;
wire n_11447;
wire n_8741;
wire n_12427;
wire n_4592;
wire n_4675;
wire n_5665;
wire n_5340;
wire n_6485;
wire n_3069;
wire n_5498;
wire n_7100;
wire n_4370;
wire n_5783;
wire n_11123;
wire n_8478;
wire n_5183;
wire n_11319;
wire n_11676;
wire n_6075;
wire n_7082;
wire n_9569;
wire n_3084;
wire n_6120;
wire n_6659;
wire n_6750;
wire n_3412;
wire n_11018;
wire n_5549;
wire n_9935;
wire n_9707;
wire n_8376;
wire n_3761;
wire n_9827;
wire n_7689;
wire n_4889;
wire n_7132;
wire n_11537;
wire n_8763;
wire n_2986;
wire n_5442;
wire n_5739;
wire n_7824;
wire n_8996;
wire n_12707;
wire n_3184;
wire n_9007;
wire n_4828;
wire n_9797;
wire n_6003;
wire n_5385;
wire n_8726;
wire n_8799;
wire n_4558;
wire n_7796;
wire n_10670;
wire n_9053;
wire n_6478;
wire n_6066;
wire n_9450;
wire n_12437;
wire n_7034;
wire n_6086;
wire n_9121;
wire n_4722;
wire n_6650;
wire n_6224;
wire n_10789;
wire n_10387;
wire n_8303;
wire n_8796;
wire n_4768;
wire n_3626;
wire n_12941;
wire n_10661;
wire n_11638;
wire n_4100;
wire n_10088;
wire n_12026;
wire n_10629;
wire n_7084;
wire n_5845;
wire n_9617;
wire n_9089;
wire n_8883;
wire n_7293;
wire n_10505;
wire n_8251;
wire n_10247;
wire n_9236;
wire n_4092;
wire n_5990;
wire n_6175;
wire n_3908;
wire n_10860;
wire n_6060;
wire n_7253;
wire n_3671;
wire n_6891;
wire n_5663;
wire n_12537;
wire n_9493;
wire n_8860;
wire n_8003;
wire n_6410;
wire n_12607;
wire n_3344;
wire n_4465;
wire n_5973;
wire n_12958;
wire n_12849;
wire n_3302;
wire n_5537;
wire n_5304;
wire n_8524;
wire n_6059;
wire n_5130;
wire n_12329;
wire n_8914;
wire n_10524;
wire n_7520;
wire n_12032;
wire n_12159;
wire n_3122;
wire n_5162;
wire n_4808;
wire n_8520;
wire n_9490;
wire n_3842;
wire n_6103;
wire n_6809;
wire n_10376;
wire n_3265;
wire n_12737;
wire n_4482;
wire n_11213;
wire n_10986;
wire n_12504;
wire n_12987;
wire n_6267;
wire n_8165;
wire n_11523;
wire n_9525;
wire n_2957;
wire n_9127;
wire n_9119;
wire n_12521;
wire n_5855;
wire n_11903;
wire n_9002;
wire n_10069;
wire n_10697;
wire n_11100;
wire n_12866;
wire n_8330;
wire n_12226;
wire n_8682;
wire n_5757;
wire n_6437;
wire n_3309;
wire n_7331;
wire n_6610;
wire n_7918;
wire n_12170;
wire n_11440;
wire n_10259;
wire n_8467;
wire n_8886;
wire n_8775;
wire n_10844;
wire n_3260;
wire n_12482;
wire n_4926;
wire n_3357;
wire n_11476;
wire n_8696;
wire n_4116;
wire n_6957;
wire n_5704;
wire n_7514;
wire n_11966;
wire n_10330;
wire n_7163;
wire n_7620;
wire n_11115;
wire n_9867;
wire n_2815;
wire n_5473;
wire n_11765;
wire n_4612;
wire n_3754;
wire n_5946;
wire n_10197;
wire n_6711;
wire n_8464;
wire n_12440;
wire n_4287;
wire n_7445;
wire n_10584;
wire n_6847;
wire n_9131;
wire n_3063;
wire n_9790;
wire n_5177;
wire n_3617;
wire n_10522;
wire n_11200;
wire n_10752;
wire n_11332;
wire n_7123;
wire n_6384;
wire n_10854;
wire n_4516;
wire n_11189;
wire n_12834;
wire n_3794;
wire n_10768;
wire n_8720;
wire n_4505;
wire n_7959;
wire n_10542;
wire n_9611;
wire n_7563;
wire n_6298;
wire n_11170;
wire n_11337;
wire n_9032;
wire n_9428;
wire n_3384;
wire n_9990;
wire n_7361;
wire n_12929;
wire n_11278;
wire n_4602;
wire n_5172;
wire n_8186;
wire n_4449;
wire n_9705;
wire n_8890;
wire n_7322;
wire n_8219;
wire n_5710;
wire n_7453;
wire n_6067;
wire n_9774;
wire n_5070;
wire n_12022;
wire n_6377;
wire n_12358;
wire n_12242;
wire n_4445;
wire n_5566;
wire n_10419;
wire n_5414;
wire n_8738;
wire n_4870;
wire n_10645;
wire n_11713;
wire n_2832;
wire n_12214;
wire n_6348;
wire n_3181;
wire n_7713;
wire n_10412;
wire n_4915;
wire n_5296;
wire n_6129;
wire n_5450;
wire n_3493;
wire n_11195;
wire n_6834;
wire n_10124;
wire n_11975;
wire n_5313;
wire n_12254;
wire n_3323;
wire n_12320;
wire n_9374;
wire n_4914;
wire n_10737;
wire n_9792;
wire n_6136;
wire n_7261;
wire n_6723;
wire n_5834;
wire n_2823;
wire n_8066;
wire n_5874;
wire n_7977;
wire n_10294;
wire n_10687;
wire n_12763;
wire n_11402;
wire n_8342;
wire n_7508;
wire n_9771;
wire n_10480;
wire n_9712;
wire n_7021;
wire n_12627;
wire n_5270;
wire n_11345;
wire n_5956;
wire n_7834;
wire n_4345;
wire n_5188;
wire n_9905;
wire n_3281;
wire n_6078;
wire n_3307;
wire n_7000;
wire n_8571;
wire n_9308;
wire n_9163;
wire n_4318;
wire n_10721;
wire n_10038;
wire n_7921;
wire n_8877;
wire n_4185;
wire n_8862;
wire n_10144;
wire n_8402;
wire n_10410;
wire n_4797;
wire n_7130;
wire n_10823;
wire n_10176;
wire n_11714;
wire n_5823;
wire n_3997;
wire n_5465;
wire n_4032;
wire n_3582;
wire n_9387;
wire n_7538;
wire n_11778;
wire n_12492;
wire n_7517;
wire n_5853;
wire n_2826;
wire n_3539;
wire n_10799;
wire n_10315;
wire n_7077;
wire n_11300;
wire n_12561;
wire n_4343;
wire n_11338;
wire n_4212;
wire n_12359;
wire n_6642;
wire n_4124;
wire n_11577;
wire n_5467;
wire n_5522;
wire n_4492;
wire n_7346;
wire n_10525;
wire n_5148;
wire n_11930;
wire n_4994;
wire n_7333;
wire n_4245;
wire n_4364;
wire n_4928;
wire n_11334;
wire n_4378;
wire n_3406;
wire n_3604;
wire n_7546;
wire n_3853;
wire n_4216;
wire n_9847;
wire n_12688;
wire n_5934;
wire n_6942;
wire n_8418;
wire n_10932;
wire n_10227;
wire n_11096;
wire n_9577;
wire n_10951;
wire n_2938;
wire n_4309;
wire n_3594;
wire n_8805;
wire n_9111;
wire n_10646;
wire n_6511;
wire n_3721;
wire n_12635;
wire n_6507;
wire n_12677;
wire n_9513;
wire n_12568;
wire n_11482;
wire n_9853;
wire n_11759;
wire n_10710;
wire n_7319;
wire n_7997;
wire n_2991;
wire n_12639;
wire n_6497;
wire n_12610;
wire n_6001;
wire n_6007;
wire n_9130;
wire n_10409;
wire n_9941;
wire n_2894;
wire n_9135;
wire n_6606;
wire n_4560;
wire n_3473;
wire n_10709;
wire n_10633;
wire n_5318;
wire n_11829;
wire n_2839;
wire n_5395;
wire n_7078;
wire n_3463;
wire n_7047;
wire n_8144;
wire n_5067;
wire n_3699;
wire n_7107;
wire n_10606;
wire n_3360;
wire n_3873;
wire n_11936;
wire n_3693;
wire n_10325;
wire n_7469;
wire n_3857;
wire n_8111;
wire n_11308;

BUFx2_ASAP7_75t_L g2814 ( 
.A(n_2158),
.Y(n_2814)
);

CKINVDCx5p33_ASAP7_75t_R g2815 ( 
.A(n_1048),
.Y(n_2815)
);

INVxp67_ASAP7_75t_SL g2816 ( 
.A(n_2249),
.Y(n_2816)
);

CKINVDCx5p33_ASAP7_75t_R g2817 ( 
.A(n_2498),
.Y(n_2817)
);

CKINVDCx20_ASAP7_75t_R g2818 ( 
.A(n_744),
.Y(n_2818)
);

CKINVDCx5p33_ASAP7_75t_R g2819 ( 
.A(n_2586),
.Y(n_2819)
);

CKINVDCx20_ASAP7_75t_R g2820 ( 
.A(n_505),
.Y(n_2820)
);

CKINVDCx5p33_ASAP7_75t_R g2821 ( 
.A(n_2628),
.Y(n_2821)
);

INVx1_ASAP7_75t_L g2822 ( 
.A(n_2719),
.Y(n_2822)
);

INVx1_ASAP7_75t_L g2823 ( 
.A(n_581),
.Y(n_2823)
);

INVx1_ASAP7_75t_L g2824 ( 
.A(n_1844),
.Y(n_2824)
);

INVx1_ASAP7_75t_L g2825 ( 
.A(n_2713),
.Y(n_2825)
);

INVx1_ASAP7_75t_L g2826 ( 
.A(n_1867),
.Y(n_2826)
);

CKINVDCx5p33_ASAP7_75t_R g2827 ( 
.A(n_390),
.Y(n_2827)
);

INVx1_ASAP7_75t_L g2828 ( 
.A(n_2681),
.Y(n_2828)
);

CKINVDCx5p33_ASAP7_75t_R g2829 ( 
.A(n_841),
.Y(n_2829)
);

CKINVDCx5p33_ASAP7_75t_R g2830 ( 
.A(n_2746),
.Y(n_2830)
);

INVx1_ASAP7_75t_L g2831 ( 
.A(n_68),
.Y(n_2831)
);

CKINVDCx5p33_ASAP7_75t_R g2832 ( 
.A(n_2169),
.Y(n_2832)
);

CKINVDCx5p33_ASAP7_75t_R g2833 ( 
.A(n_2580),
.Y(n_2833)
);

CKINVDCx5p33_ASAP7_75t_R g2834 ( 
.A(n_1726),
.Y(n_2834)
);

INVx1_ASAP7_75t_L g2835 ( 
.A(n_216),
.Y(n_2835)
);

CKINVDCx5p33_ASAP7_75t_R g2836 ( 
.A(n_1716),
.Y(n_2836)
);

CKINVDCx5p33_ASAP7_75t_R g2837 ( 
.A(n_2197),
.Y(n_2837)
);

CKINVDCx5p33_ASAP7_75t_R g2838 ( 
.A(n_425),
.Y(n_2838)
);

CKINVDCx5p33_ASAP7_75t_R g2839 ( 
.A(n_2526),
.Y(n_2839)
);

INVx1_ASAP7_75t_L g2840 ( 
.A(n_2092),
.Y(n_2840)
);

INVx1_ASAP7_75t_L g2841 ( 
.A(n_666),
.Y(n_2841)
);

INVx2_ASAP7_75t_SL g2842 ( 
.A(n_2777),
.Y(n_2842)
);

BUFx5_ASAP7_75t_L g2843 ( 
.A(n_598),
.Y(n_2843)
);

CKINVDCx5p33_ASAP7_75t_R g2844 ( 
.A(n_1583),
.Y(n_2844)
);

CKINVDCx5p33_ASAP7_75t_R g2845 ( 
.A(n_1854),
.Y(n_2845)
);

CKINVDCx5p33_ASAP7_75t_R g2846 ( 
.A(n_2689),
.Y(n_2846)
);

INVx1_ASAP7_75t_L g2847 ( 
.A(n_251),
.Y(n_2847)
);

INVx2_ASAP7_75t_L g2848 ( 
.A(n_2036),
.Y(n_2848)
);

CKINVDCx5p33_ASAP7_75t_R g2849 ( 
.A(n_2264),
.Y(n_2849)
);

CKINVDCx5p33_ASAP7_75t_R g2850 ( 
.A(n_731),
.Y(n_2850)
);

INVx1_ASAP7_75t_L g2851 ( 
.A(n_2177),
.Y(n_2851)
);

INVx1_ASAP7_75t_L g2852 ( 
.A(n_747),
.Y(n_2852)
);

INVx1_ASAP7_75t_L g2853 ( 
.A(n_1805),
.Y(n_2853)
);

INVx3_ASAP7_75t_L g2854 ( 
.A(n_2728),
.Y(n_2854)
);

CKINVDCx5p33_ASAP7_75t_R g2855 ( 
.A(n_2258),
.Y(n_2855)
);

CKINVDCx5p33_ASAP7_75t_R g2856 ( 
.A(n_2268),
.Y(n_2856)
);

CKINVDCx5p33_ASAP7_75t_R g2857 ( 
.A(n_1799),
.Y(n_2857)
);

INVx1_ASAP7_75t_L g2858 ( 
.A(n_2223),
.Y(n_2858)
);

INVx1_ASAP7_75t_L g2859 ( 
.A(n_546),
.Y(n_2859)
);

INVx2_ASAP7_75t_L g2860 ( 
.A(n_1667),
.Y(n_2860)
);

CKINVDCx20_ASAP7_75t_R g2861 ( 
.A(n_14),
.Y(n_2861)
);

CKINVDCx20_ASAP7_75t_R g2862 ( 
.A(n_1488),
.Y(n_2862)
);

CKINVDCx5p33_ASAP7_75t_R g2863 ( 
.A(n_1034),
.Y(n_2863)
);

INVx2_ASAP7_75t_L g2864 ( 
.A(n_675),
.Y(n_2864)
);

CKINVDCx5p33_ASAP7_75t_R g2865 ( 
.A(n_1926),
.Y(n_2865)
);

INVx2_ASAP7_75t_L g2866 ( 
.A(n_2366),
.Y(n_2866)
);

CKINVDCx5p33_ASAP7_75t_R g2867 ( 
.A(n_2112),
.Y(n_2867)
);

CKINVDCx5p33_ASAP7_75t_R g2868 ( 
.A(n_203),
.Y(n_2868)
);

INVx1_ASAP7_75t_L g2869 ( 
.A(n_1610),
.Y(n_2869)
);

CKINVDCx5p33_ASAP7_75t_R g2870 ( 
.A(n_1956),
.Y(n_2870)
);

CKINVDCx20_ASAP7_75t_R g2871 ( 
.A(n_1947),
.Y(n_2871)
);

INVx1_ASAP7_75t_L g2872 ( 
.A(n_1497),
.Y(n_2872)
);

CKINVDCx20_ASAP7_75t_R g2873 ( 
.A(n_1033),
.Y(n_2873)
);

CKINVDCx20_ASAP7_75t_R g2874 ( 
.A(n_1429),
.Y(n_2874)
);

CKINVDCx16_ASAP7_75t_R g2875 ( 
.A(n_2605),
.Y(n_2875)
);

INVx1_ASAP7_75t_L g2876 ( 
.A(n_583),
.Y(n_2876)
);

BUFx3_ASAP7_75t_L g2877 ( 
.A(n_2401),
.Y(n_2877)
);

CKINVDCx5p33_ASAP7_75t_R g2878 ( 
.A(n_1485),
.Y(n_2878)
);

CKINVDCx5p33_ASAP7_75t_R g2879 ( 
.A(n_830),
.Y(n_2879)
);

CKINVDCx20_ASAP7_75t_R g2880 ( 
.A(n_725),
.Y(n_2880)
);

INVx1_ASAP7_75t_L g2881 ( 
.A(n_2803),
.Y(n_2881)
);

INVx1_ASAP7_75t_SL g2882 ( 
.A(n_1063),
.Y(n_2882)
);

CKINVDCx5p33_ASAP7_75t_R g2883 ( 
.A(n_1385),
.Y(n_2883)
);

INVx1_ASAP7_75t_L g2884 ( 
.A(n_643),
.Y(n_2884)
);

CKINVDCx5p33_ASAP7_75t_R g2885 ( 
.A(n_2722),
.Y(n_2885)
);

CKINVDCx5p33_ASAP7_75t_R g2886 ( 
.A(n_2710),
.Y(n_2886)
);

INVx1_ASAP7_75t_L g2887 ( 
.A(n_2577),
.Y(n_2887)
);

CKINVDCx5p33_ASAP7_75t_R g2888 ( 
.A(n_359),
.Y(n_2888)
);

CKINVDCx5p33_ASAP7_75t_R g2889 ( 
.A(n_183),
.Y(n_2889)
);

BUFx2_ASAP7_75t_SL g2890 ( 
.A(n_2612),
.Y(n_2890)
);

CKINVDCx5p33_ASAP7_75t_R g2891 ( 
.A(n_2584),
.Y(n_2891)
);

INVx1_ASAP7_75t_L g2892 ( 
.A(n_2356),
.Y(n_2892)
);

INVx1_ASAP7_75t_L g2893 ( 
.A(n_1325),
.Y(n_2893)
);

CKINVDCx5p33_ASAP7_75t_R g2894 ( 
.A(n_250),
.Y(n_2894)
);

CKINVDCx5p33_ASAP7_75t_R g2895 ( 
.A(n_2596),
.Y(n_2895)
);

INVx1_ASAP7_75t_L g2896 ( 
.A(n_2592),
.Y(n_2896)
);

CKINVDCx5p33_ASAP7_75t_R g2897 ( 
.A(n_1809),
.Y(n_2897)
);

CKINVDCx5p33_ASAP7_75t_R g2898 ( 
.A(n_2194),
.Y(n_2898)
);

BUFx5_ASAP7_75t_L g2899 ( 
.A(n_2486),
.Y(n_2899)
);

CKINVDCx20_ASAP7_75t_R g2900 ( 
.A(n_2651),
.Y(n_2900)
);

CKINVDCx5p33_ASAP7_75t_R g2901 ( 
.A(n_102),
.Y(n_2901)
);

CKINVDCx5p33_ASAP7_75t_R g2902 ( 
.A(n_2280),
.Y(n_2902)
);

INVx1_ASAP7_75t_SL g2903 ( 
.A(n_2639),
.Y(n_2903)
);

INVx2_ASAP7_75t_L g2904 ( 
.A(n_535),
.Y(n_2904)
);

INVx1_ASAP7_75t_L g2905 ( 
.A(n_2714),
.Y(n_2905)
);

CKINVDCx5p33_ASAP7_75t_R g2906 ( 
.A(n_2554),
.Y(n_2906)
);

CKINVDCx5p33_ASAP7_75t_R g2907 ( 
.A(n_854),
.Y(n_2907)
);

CKINVDCx5p33_ASAP7_75t_R g2908 ( 
.A(n_2204),
.Y(n_2908)
);

CKINVDCx5p33_ASAP7_75t_R g2909 ( 
.A(n_1584),
.Y(n_2909)
);

CKINVDCx5p33_ASAP7_75t_R g2910 ( 
.A(n_2591),
.Y(n_2910)
);

CKINVDCx5p33_ASAP7_75t_R g2911 ( 
.A(n_2484),
.Y(n_2911)
);

CKINVDCx5p33_ASAP7_75t_R g2912 ( 
.A(n_1192),
.Y(n_2912)
);

INVx1_ASAP7_75t_L g2913 ( 
.A(n_2609),
.Y(n_2913)
);

INVx3_ASAP7_75t_L g2914 ( 
.A(n_1795),
.Y(n_2914)
);

CKINVDCx5p33_ASAP7_75t_R g2915 ( 
.A(n_1324),
.Y(n_2915)
);

CKINVDCx5p33_ASAP7_75t_R g2916 ( 
.A(n_1166),
.Y(n_2916)
);

INVx1_ASAP7_75t_L g2917 ( 
.A(n_2701),
.Y(n_2917)
);

CKINVDCx5p33_ASAP7_75t_R g2918 ( 
.A(n_2122),
.Y(n_2918)
);

INVx1_ASAP7_75t_L g2919 ( 
.A(n_2194),
.Y(n_2919)
);

INVx1_ASAP7_75t_SL g2920 ( 
.A(n_2687),
.Y(n_2920)
);

INVx1_ASAP7_75t_L g2921 ( 
.A(n_380),
.Y(n_2921)
);

CKINVDCx5p33_ASAP7_75t_R g2922 ( 
.A(n_2563),
.Y(n_2922)
);

CKINVDCx5p33_ASAP7_75t_R g2923 ( 
.A(n_39),
.Y(n_2923)
);

CKINVDCx5p33_ASAP7_75t_R g2924 ( 
.A(n_2394),
.Y(n_2924)
);

INVx2_ASAP7_75t_L g2925 ( 
.A(n_500),
.Y(n_2925)
);

INVx1_ASAP7_75t_L g2926 ( 
.A(n_2566),
.Y(n_2926)
);

CKINVDCx20_ASAP7_75t_R g2927 ( 
.A(n_1148),
.Y(n_2927)
);

CKINVDCx5p33_ASAP7_75t_R g2928 ( 
.A(n_2453),
.Y(n_2928)
);

INVx1_ASAP7_75t_L g2929 ( 
.A(n_1454),
.Y(n_2929)
);

CKINVDCx5p33_ASAP7_75t_R g2930 ( 
.A(n_2095),
.Y(n_2930)
);

INVx2_ASAP7_75t_L g2931 ( 
.A(n_1773),
.Y(n_2931)
);

INVx1_ASAP7_75t_L g2932 ( 
.A(n_2732),
.Y(n_2932)
);

INVx1_ASAP7_75t_L g2933 ( 
.A(n_2034),
.Y(n_2933)
);

CKINVDCx5p33_ASAP7_75t_R g2934 ( 
.A(n_2767),
.Y(n_2934)
);

CKINVDCx5p33_ASAP7_75t_R g2935 ( 
.A(n_904),
.Y(n_2935)
);

CKINVDCx5p33_ASAP7_75t_R g2936 ( 
.A(n_139),
.Y(n_2936)
);

INVx1_ASAP7_75t_L g2937 ( 
.A(n_864),
.Y(n_2937)
);

CKINVDCx5p33_ASAP7_75t_R g2938 ( 
.A(n_1362),
.Y(n_2938)
);

INVx1_ASAP7_75t_SL g2939 ( 
.A(n_1984),
.Y(n_2939)
);

CKINVDCx5p33_ASAP7_75t_R g2940 ( 
.A(n_1964),
.Y(n_2940)
);

CKINVDCx5p33_ASAP7_75t_R g2941 ( 
.A(n_2618),
.Y(n_2941)
);

CKINVDCx5p33_ASAP7_75t_R g2942 ( 
.A(n_1507),
.Y(n_2942)
);

INVxp67_ASAP7_75t_L g2943 ( 
.A(n_507),
.Y(n_2943)
);

CKINVDCx5p33_ASAP7_75t_R g2944 ( 
.A(n_2510),
.Y(n_2944)
);

INVx1_ASAP7_75t_L g2945 ( 
.A(n_2725),
.Y(n_2945)
);

INVx1_ASAP7_75t_L g2946 ( 
.A(n_1951),
.Y(n_2946)
);

INVx2_ASAP7_75t_SL g2947 ( 
.A(n_2271),
.Y(n_2947)
);

CKINVDCx5p33_ASAP7_75t_R g2948 ( 
.A(n_2095),
.Y(n_2948)
);

INVx1_ASAP7_75t_L g2949 ( 
.A(n_70),
.Y(n_2949)
);

CKINVDCx5p33_ASAP7_75t_R g2950 ( 
.A(n_154),
.Y(n_2950)
);

INVx1_ASAP7_75t_L g2951 ( 
.A(n_2746),
.Y(n_2951)
);

CKINVDCx5p33_ASAP7_75t_R g2952 ( 
.A(n_2353),
.Y(n_2952)
);

CKINVDCx5p33_ASAP7_75t_R g2953 ( 
.A(n_2526),
.Y(n_2953)
);

CKINVDCx20_ASAP7_75t_R g2954 ( 
.A(n_2754),
.Y(n_2954)
);

CKINVDCx5p33_ASAP7_75t_R g2955 ( 
.A(n_2405),
.Y(n_2955)
);

INVx2_ASAP7_75t_L g2956 ( 
.A(n_2569),
.Y(n_2956)
);

CKINVDCx5p33_ASAP7_75t_R g2957 ( 
.A(n_704),
.Y(n_2957)
);

CKINVDCx5p33_ASAP7_75t_R g2958 ( 
.A(n_80),
.Y(n_2958)
);

CKINVDCx5p33_ASAP7_75t_R g2959 ( 
.A(n_200),
.Y(n_2959)
);

CKINVDCx5p33_ASAP7_75t_R g2960 ( 
.A(n_2346),
.Y(n_2960)
);

CKINVDCx5p33_ASAP7_75t_R g2961 ( 
.A(n_2402),
.Y(n_2961)
);

CKINVDCx5p33_ASAP7_75t_R g2962 ( 
.A(n_2682),
.Y(n_2962)
);

CKINVDCx5p33_ASAP7_75t_R g2963 ( 
.A(n_2603),
.Y(n_2963)
);

CKINVDCx5p33_ASAP7_75t_R g2964 ( 
.A(n_2813),
.Y(n_2964)
);

BUFx3_ASAP7_75t_L g2965 ( 
.A(n_765),
.Y(n_2965)
);

INVx1_ASAP7_75t_L g2966 ( 
.A(n_2379),
.Y(n_2966)
);

CKINVDCx5p33_ASAP7_75t_R g2967 ( 
.A(n_1823),
.Y(n_2967)
);

BUFx3_ASAP7_75t_L g2968 ( 
.A(n_1217),
.Y(n_2968)
);

CKINVDCx5p33_ASAP7_75t_R g2969 ( 
.A(n_1708),
.Y(n_2969)
);

CKINVDCx5p33_ASAP7_75t_R g2970 ( 
.A(n_1214),
.Y(n_2970)
);

CKINVDCx5p33_ASAP7_75t_R g2971 ( 
.A(n_888),
.Y(n_2971)
);

INVx1_ASAP7_75t_L g2972 ( 
.A(n_629),
.Y(n_2972)
);

CKINVDCx20_ASAP7_75t_R g2973 ( 
.A(n_680),
.Y(n_2973)
);

INVx1_ASAP7_75t_L g2974 ( 
.A(n_65),
.Y(n_2974)
);

BUFx3_ASAP7_75t_L g2975 ( 
.A(n_1414),
.Y(n_2975)
);

CKINVDCx5p33_ASAP7_75t_R g2976 ( 
.A(n_2642),
.Y(n_2976)
);

CKINVDCx5p33_ASAP7_75t_R g2977 ( 
.A(n_932),
.Y(n_2977)
);

INVx1_ASAP7_75t_L g2978 ( 
.A(n_2549),
.Y(n_2978)
);

CKINVDCx5p33_ASAP7_75t_R g2979 ( 
.A(n_571),
.Y(n_2979)
);

INVx1_ASAP7_75t_L g2980 ( 
.A(n_2716),
.Y(n_2980)
);

INVx2_ASAP7_75t_L g2981 ( 
.A(n_2401),
.Y(n_2981)
);

INVx1_ASAP7_75t_L g2982 ( 
.A(n_1692),
.Y(n_2982)
);

INVx1_ASAP7_75t_L g2983 ( 
.A(n_981),
.Y(n_2983)
);

BUFx2_ASAP7_75t_L g2984 ( 
.A(n_941),
.Y(n_2984)
);

BUFx3_ASAP7_75t_L g2985 ( 
.A(n_2594),
.Y(n_2985)
);

INVx2_ASAP7_75t_L g2986 ( 
.A(n_2467),
.Y(n_2986)
);

CKINVDCx5p33_ASAP7_75t_R g2987 ( 
.A(n_360),
.Y(n_2987)
);

INVx2_ASAP7_75t_L g2988 ( 
.A(n_1936),
.Y(n_2988)
);

CKINVDCx5p33_ASAP7_75t_R g2989 ( 
.A(n_1473),
.Y(n_2989)
);

CKINVDCx5p33_ASAP7_75t_R g2990 ( 
.A(n_1729),
.Y(n_2990)
);

CKINVDCx5p33_ASAP7_75t_R g2991 ( 
.A(n_2570),
.Y(n_2991)
);

CKINVDCx5p33_ASAP7_75t_R g2992 ( 
.A(n_1060),
.Y(n_2992)
);

CKINVDCx20_ASAP7_75t_R g2993 ( 
.A(n_1001),
.Y(n_2993)
);

INVx1_ASAP7_75t_L g2994 ( 
.A(n_2657),
.Y(n_2994)
);

INVx1_ASAP7_75t_SL g2995 ( 
.A(n_2630),
.Y(n_2995)
);

BUFx2_ASAP7_75t_SL g2996 ( 
.A(n_1439),
.Y(n_2996)
);

CKINVDCx5p33_ASAP7_75t_R g2997 ( 
.A(n_1769),
.Y(n_2997)
);

CKINVDCx5p33_ASAP7_75t_R g2998 ( 
.A(n_625),
.Y(n_2998)
);

INVx1_ASAP7_75t_SL g2999 ( 
.A(n_1686),
.Y(n_2999)
);

INVx1_ASAP7_75t_L g3000 ( 
.A(n_1098),
.Y(n_3000)
);

CKINVDCx5p33_ASAP7_75t_R g3001 ( 
.A(n_625),
.Y(n_3001)
);

CKINVDCx16_ASAP7_75t_R g3002 ( 
.A(n_291),
.Y(n_3002)
);

CKINVDCx5p33_ASAP7_75t_R g3003 ( 
.A(n_2724),
.Y(n_3003)
);

CKINVDCx5p33_ASAP7_75t_R g3004 ( 
.A(n_1663),
.Y(n_3004)
);

BUFx3_ASAP7_75t_L g3005 ( 
.A(n_1694),
.Y(n_3005)
);

CKINVDCx5p33_ASAP7_75t_R g3006 ( 
.A(n_771),
.Y(n_3006)
);

INVx1_ASAP7_75t_L g3007 ( 
.A(n_145),
.Y(n_3007)
);

INVx1_ASAP7_75t_L g3008 ( 
.A(n_977),
.Y(n_3008)
);

INVx1_ASAP7_75t_L g3009 ( 
.A(n_1367),
.Y(n_3009)
);

INVx1_ASAP7_75t_L g3010 ( 
.A(n_1384),
.Y(n_3010)
);

BUFx3_ASAP7_75t_L g3011 ( 
.A(n_1606),
.Y(n_3011)
);

CKINVDCx20_ASAP7_75t_R g3012 ( 
.A(n_390),
.Y(n_3012)
);

INVx1_ASAP7_75t_L g3013 ( 
.A(n_381),
.Y(n_3013)
);

INVx1_ASAP7_75t_L g3014 ( 
.A(n_1827),
.Y(n_3014)
);

CKINVDCx5p33_ASAP7_75t_R g3015 ( 
.A(n_2553),
.Y(n_3015)
);

CKINVDCx5p33_ASAP7_75t_R g3016 ( 
.A(n_861),
.Y(n_3016)
);

CKINVDCx14_ASAP7_75t_R g3017 ( 
.A(n_1837),
.Y(n_3017)
);

INVx1_ASAP7_75t_L g3018 ( 
.A(n_709),
.Y(n_3018)
);

CKINVDCx5p33_ASAP7_75t_R g3019 ( 
.A(n_233),
.Y(n_3019)
);

INVx1_ASAP7_75t_L g3020 ( 
.A(n_1387),
.Y(n_3020)
);

CKINVDCx5p33_ASAP7_75t_R g3021 ( 
.A(n_1088),
.Y(n_3021)
);

INVx1_ASAP7_75t_SL g3022 ( 
.A(n_382),
.Y(n_3022)
);

CKINVDCx5p33_ASAP7_75t_R g3023 ( 
.A(n_2162),
.Y(n_3023)
);

CKINVDCx16_ASAP7_75t_R g3024 ( 
.A(n_1682),
.Y(n_3024)
);

CKINVDCx5p33_ASAP7_75t_R g3025 ( 
.A(n_2058),
.Y(n_3025)
);

INVx1_ASAP7_75t_L g3026 ( 
.A(n_739),
.Y(n_3026)
);

CKINVDCx5p33_ASAP7_75t_R g3027 ( 
.A(n_2779),
.Y(n_3027)
);

CKINVDCx5p33_ASAP7_75t_R g3028 ( 
.A(n_2800),
.Y(n_3028)
);

BUFx6f_ASAP7_75t_L g3029 ( 
.A(n_239),
.Y(n_3029)
);

CKINVDCx5p33_ASAP7_75t_R g3030 ( 
.A(n_2187),
.Y(n_3030)
);

CKINVDCx5p33_ASAP7_75t_R g3031 ( 
.A(n_1999),
.Y(n_3031)
);

INVx1_ASAP7_75t_L g3032 ( 
.A(n_34),
.Y(n_3032)
);

CKINVDCx20_ASAP7_75t_R g3033 ( 
.A(n_425),
.Y(n_3033)
);

INVx1_ASAP7_75t_L g3034 ( 
.A(n_468),
.Y(n_3034)
);

CKINVDCx16_ASAP7_75t_R g3035 ( 
.A(n_1165),
.Y(n_3035)
);

CKINVDCx5p33_ASAP7_75t_R g3036 ( 
.A(n_2418),
.Y(n_3036)
);

CKINVDCx5p33_ASAP7_75t_R g3037 ( 
.A(n_1746),
.Y(n_3037)
);

CKINVDCx5p33_ASAP7_75t_R g3038 ( 
.A(n_2733),
.Y(n_3038)
);

INVx1_ASAP7_75t_L g3039 ( 
.A(n_1995),
.Y(n_3039)
);

CKINVDCx5p33_ASAP7_75t_R g3040 ( 
.A(n_1289),
.Y(n_3040)
);

CKINVDCx5p33_ASAP7_75t_R g3041 ( 
.A(n_365),
.Y(n_3041)
);

INVx1_ASAP7_75t_L g3042 ( 
.A(n_81),
.Y(n_3042)
);

CKINVDCx14_ASAP7_75t_R g3043 ( 
.A(n_839),
.Y(n_3043)
);

INVx2_ASAP7_75t_SL g3044 ( 
.A(n_421),
.Y(n_3044)
);

CKINVDCx5p33_ASAP7_75t_R g3045 ( 
.A(n_156),
.Y(n_3045)
);

CKINVDCx5p33_ASAP7_75t_R g3046 ( 
.A(n_1849),
.Y(n_3046)
);

INVx1_ASAP7_75t_L g3047 ( 
.A(n_343),
.Y(n_3047)
);

CKINVDCx5p33_ASAP7_75t_R g3048 ( 
.A(n_2540),
.Y(n_3048)
);

CKINVDCx5p33_ASAP7_75t_R g3049 ( 
.A(n_1406),
.Y(n_3049)
);

INVx1_ASAP7_75t_L g3050 ( 
.A(n_1898),
.Y(n_3050)
);

INVx1_ASAP7_75t_L g3051 ( 
.A(n_1500),
.Y(n_3051)
);

BUFx3_ASAP7_75t_L g3052 ( 
.A(n_1226),
.Y(n_3052)
);

BUFx6f_ASAP7_75t_L g3053 ( 
.A(n_1981),
.Y(n_3053)
);

CKINVDCx5p33_ASAP7_75t_R g3054 ( 
.A(n_764),
.Y(n_3054)
);

INVx2_ASAP7_75t_SL g3055 ( 
.A(n_1),
.Y(n_3055)
);

CKINVDCx5p33_ASAP7_75t_R g3056 ( 
.A(n_134),
.Y(n_3056)
);

BUFx3_ASAP7_75t_L g3057 ( 
.A(n_555),
.Y(n_3057)
);

CKINVDCx20_ASAP7_75t_R g3058 ( 
.A(n_2137),
.Y(n_3058)
);

INVx1_ASAP7_75t_L g3059 ( 
.A(n_701),
.Y(n_3059)
);

BUFx5_ASAP7_75t_L g3060 ( 
.A(n_1655),
.Y(n_3060)
);

INVx1_ASAP7_75t_L g3061 ( 
.A(n_2780),
.Y(n_3061)
);

INVx2_ASAP7_75t_SL g3062 ( 
.A(n_2416),
.Y(n_3062)
);

INVx1_ASAP7_75t_L g3063 ( 
.A(n_2607),
.Y(n_3063)
);

CKINVDCx5p33_ASAP7_75t_R g3064 ( 
.A(n_1590),
.Y(n_3064)
);

INVx1_ASAP7_75t_L g3065 ( 
.A(n_997),
.Y(n_3065)
);

CKINVDCx5p33_ASAP7_75t_R g3066 ( 
.A(n_2153),
.Y(n_3066)
);

CKINVDCx5p33_ASAP7_75t_R g3067 ( 
.A(n_1959),
.Y(n_3067)
);

CKINVDCx5p33_ASAP7_75t_R g3068 ( 
.A(n_387),
.Y(n_3068)
);

CKINVDCx5p33_ASAP7_75t_R g3069 ( 
.A(n_131),
.Y(n_3069)
);

INVx1_ASAP7_75t_L g3070 ( 
.A(n_1928),
.Y(n_3070)
);

CKINVDCx5p33_ASAP7_75t_R g3071 ( 
.A(n_928),
.Y(n_3071)
);

INVx1_ASAP7_75t_L g3072 ( 
.A(n_2802),
.Y(n_3072)
);

CKINVDCx16_ASAP7_75t_R g3073 ( 
.A(n_2323),
.Y(n_3073)
);

INVx1_ASAP7_75t_L g3074 ( 
.A(n_2196),
.Y(n_3074)
);

INVx1_ASAP7_75t_L g3075 ( 
.A(n_2423),
.Y(n_3075)
);

CKINVDCx5p33_ASAP7_75t_R g3076 ( 
.A(n_76),
.Y(n_3076)
);

INVx1_ASAP7_75t_L g3077 ( 
.A(n_1937),
.Y(n_3077)
);

INVx3_ASAP7_75t_L g3078 ( 
.A(n_428),
.Y(n_3078)
);

CKINVDCx5p33_ASAP7_75t_R g3079 ( 
.A(n_1561),
.Y(n_3079)
);

CKINVDCx5p33_ASAP7_75t_R g3080 ( 
.A(n_2291),
.Y(n_3080)
);

CKINVDCx5p33_ASAP7_75t_R g3081 ( 
.A(n_1502),
.Y(n_3081)
);

INVx1_ASAP7_75t_SL g3082 ( 
.A(n_2038),
.Y(n_3082)
);

CKINVDCx5p33_ASAP7_75t_R g3083 ( 
.A(n_1056),
.Y(n_3083)
);

CKINVDCx5p33_ASAP7_75t_R g3084 ( 
.A(n_441),
.Y(n_3084)
);

INVx1_ASAP7_75t_L g3085 ( 
.A(n_2449),
.Y(n_3085)
);

CKINVDCx5p33_ASAP7_75t_R g3086 ( 
.A(n_1254),
.Y(n_3086)
);

CKINVDCx5p33_ASAP7_75t_R g3087 ( 
.A(n_2277),
.Y(n_3087)
);

CKINVDCx20_ASAP7_75t_R g3088 ( 
.A(n_1947),
.Y(n_3088)
);

CKINVDCx5p33_ASAP7_75t_R g3089 ( 
.A(n_2372),
.Y(n_3089)
);

INVx1_ASAP7_75t_L g3090 ( 
.A(n_936),
.Y(n_3090)
);

CKINVDCx5p33_ASAP7_75t_R g3091 ( 
.A(n_663),
.Y(n_3091)
);

CKINVDCx5p33_ASAP7_75t_R g3092 ( 
.A(n_2486),
.Y(n_3092)
);

CKINVDCx5p33_ASAP7_75t_R g3093 ( 
.A(n_142),
.Y(n_3093)
);

INVx2_ASAP7_75t_L g3094 ( 
.A(n_2610),
.Y(n_3094)
);

INVx1_ASAP7_75t_L g3095 ( 
.A(n_422),
.Y(n_3095)
);

CKINVDCx5p33_ASAP7_75t_R g3096 ( 
.A(n_414),
.Y(n_3096)
);

CKINVDCx5p33_ASAP7_75t_R g3097 ( 
.A(n_2686),
.Y(n_3097)
);

INVx1_ASAP7_75t_L g3098 ( 
.A(n_1192),
.Y(n_3098)
);

CKINVDCx5p33_ASAP7_75t_R g3099 ( 
.A(n_2793),
.Y(n_3099)
);

CKINVDCx5p33_ASAP7_75t_R g3100 ( 
.A(n_583),
.Y(n_3100)
);

INVx1_ASAP7_75t_L g3101 ( 
.A(n_2753),
.Y(n_3101)
);

CKINVDCx5p33_ASAP7_75t_R g3102 ( 
.A(n_2808),
.Y(n_3102)
);

INVx1_ASAP7_75t_L g3103 ( 
.A(n_2087),
.Y(n_3103)
);

CKINVDCx5p33_ASAP7_75t_R g3104 ( 
.A(n_1594),
.Y(n_3104)
);

CKINVDCx5p33_ASAP7_75t_R g3105 ( 
.A(n_734),
.Y(n_3105)
);

CKINVDCx5p33_ASAP7_75t_R g3106 ( 
.A(n_276),
.Y(n_3106)
);

CKINVDCx5p33_ASAP7_75t_R g3107 ( 
.A(n_671),
.Y(n_3107)
);

INVx2_ASAP7_75t_L g3108 ( 
.A(n_1677),
.Y(n_3108)
);

CKINVDCx5p33_ASAP7_75t_R g3109 ( 
.A(n_1567),
.Y(n_3109)
);

CKINVDCx5p33_ASAP7_75t_R g3110 ( 
.A(n_1695),
.Y(n_3110)
);

CKINVDCx20_ASAP7_75t_R g3111 ( 
.A(n_1550),
.Y(n_3111)
);

INVx1_ASAP7_75t_L g3112 ( 
.A(n_219),
.Y(n_3112)
);

INVx1_ASAP7_75t_L g3113 ( 
.A(n_1081),
.Y(n_3113)
);

CKINVDCx5p33_ASAP7_75t_R g3114 ( 
.A(n_968),
.Y(n_3114)
);

INVx2_ASAP7_75t_SL g3115 ( 
.A(n_1247),
.Y(n_3115)
);

CKINVDCx16_ASAP7_75t_R g3116 ( 
.A(n_147),
.Y(n_3116)
);

BUFx6f_ASAP7_75t_L g3117 ( 
.A(n_346),
.Y(n_3117)
);

BUFx5_ASAP7_75t_L g3118 ( 
.A(n_2330),
.Y(n_3118)
);

CKINVDCx5p33_ASAP7_75t_R g3119 ( 
.A(n_2109),
.Y(n_3119)
);

BUFx10_ASAP7_75t_L g3120 ( 
.A(n_2707),
.Y(n_3120)
);

INVx1_ASAP7_75t_L g3121 ( 
.A(n_2370),
.Y(n_3121)
);

CKINVDCx5p33_ASAP7_75t_R g3122 ( 
.A(n_623),
.Y(n_3122)
);

CKINVDCx5p33_ASAP7_75t_R g3123 ( 
.A(n_2106),
.Y(n_3123)
);

CKINVDCx5p33_ASAP7_75t_R g3124 ( 
.A(n_2208),
.Y(n_3124)
);

INVx1_ASAP7_75t_L g3125 ( 
.A(n_142),
.Y(n_3125)
);

INVx1_ASAP7_75t_L g3126 ( 
.A(n_459),
.Y(n_3126)
);

CKINVDCx5p33_ASAP7_75t_R g3127 ( 
.A(n_2115),
.Y(n_3127)
);

CKINVDCx5p33_ASAP7_75t_R g3128 ( 
.A(n_2461),
.Y(n_3128)
);

INVx1_ASAP7_75t_L g3129 ( 
.A(n_1524),
.Y(n_3129)
);

CKINVDCx5p33_ASAP7_75t_R g3130 ( 
.A(n_1297),
.Y(n_3130)
);

INVx1_ASAP7_75t_SL g3131 ( 
.A(n_879),
.Y(n_3131)
);

CKINVDCx5p33_ASAP7_75t_R g3132 ( 
.A(n_1911),
.Y(n_3132)
);

INVx1_ASAP7_75t_L g3133 ( 
.A(n_2152),
.Y(n_3133)
);

CKINVDCx5p33_ASAP7_75t_R g3134 ( 
.A(n_2078),
.Y(n_3134)
);

CKINVDCx20_ASAP7_75t_R g3135 ( 
.A(n_528),
.Y(n_3135)
);

CKINVDCx5p33_ASAP7_75t_R g3136 ( 
.A(n_505),
.Y(n_3136)
);

CKINVDCx5p33_ASAP7_75t_R g3137 ( 
.A(n_1533),
.Y(n_3137)
);

INVx1_ASAP7_75t_L g3138 ( 
.A(n_1177),
.Y(n_3138)
);

CKINVDCx5p33_ASAP7_75t_R g3139 ( 
.A(n_2328),
.Y(n_3139)
);

INVx1_ASAP7_75t_L g3140 ( 
.A(n_713),
.Y(n_3140)
);

CKINVDCx5p33_ASAP7_75t_R g3141 ( 
.A(n_2675),
.Y(n_3141)
);

INVx1_ASAP7_75t_L g3142 ( 
.A(n_2601),
.Y(n_3142)
);

INVx1_ASAP7_75t_L g3143 ( 
.A(n_1817),
.Y(n_3143)
);

INVx2_ASAP7_75t_L g3144 ( 
.A(n_486),
.Y(n_3144)
);

CKINVDCx5p33_ASAP7_75t_R g3145 ( 
.A(n_411),
.Y(n_3145)
);

BUFx10_ASAP7_75t_L g3146 ( 
.A(n_2201),
.Y(n_3146)
);

CKINVDCx20_ASAP7_75t_R g3147 ( 
.A(n_420),
.Y(n_3147)
);

BUFx6f_ASAP7_75t_L g3148 ( 
.A(n_563),
.Y(n_3148)
);

CKINVDCx5p33_ASAP7_75t_R g3149 ( 
.A(n_458),
.Y(n_3149)
);

CKINVDCx5p33_ASAP7_75t_R g3150 ( 
.A(n_70),
.Y(n_3150)
);

CKINVDCx5p33_ASAP7_75t_R g3151 ( 
.A(n_2058),
.Y(n_3151)
);

INVx1_ASAP7_75t_L g3152 ( 
.A(n_1353),
.Y(n_3152)
);

INVx1_ASAP7_75t_L g3153 ( 
.A(n_640),
.Y(n_3153)
);

CKINVDCx5p33_ASAP7_75t_R g3154 ( 
.A(n_2086),
.Y(n_3154)
);

CKINVDCx5p33_ASAP7_75t_R g3155 ( 
.A(n_2196),
.Y(n_3155)
);

INVx1_ASAP7_75t_L g3156 ( 
.A(n_230),
.Y(n_3156)
);

INVx1_ASAP7_75t_L g3157 ( 
.A(n_2281),
.Y(n_3157)
);

CKINVDCx5p33_ASAP7_75t_R g3158 ( 
.A(n_2752),
.Y(n_3158)
);

CKINVDCx5p33_ASAP7_75t_R g3159 ( 
.A(n_2734),
.Y(n_3159)
);

CKINVDCx5p33_ASAP7_75t_R g3160 ( 
.A(n_2669),
.Y(n_3160)
);

CKINVDCx5p33_ASAP7_75t_R g3161 ( 
.A(n_1946),
.Y(n_3161)
);

CKINVDCx5p33_ASAP7_75t_R g3162 ( 
.A(n_2717),
.Y(n_3162)
);

CKINVDCx5p33_ASAP7_75t_R g3163 ( 
.A(n_2106),
.Y(n_3163)
);

CKINVDCx5p33_ASAP7_75t_R g3164 ( 
.A(n_777),
.Y(n_3164)
);

CKINVDCx5p33_ASAP7_75t_R g3165 ( 
.A(n_358),
.Y(n_3165)
);

CKINVDCx5p33_ASAP7_75t_R g3166 ( 
.A(n_2149),
.Y(n_3166)
);

BUFx3_ASAP7_75t_L g3167 ( 
.A(n_1364),
.Y(n_3167)
);

CKINVDCx5p33_ASAP7_75t_R g3168 ( 
.A(n_377),
.Y(n_3168)
);

CKINVDCx5p33_ASAP7_75t_R g3169 ( 
.A(n_1938),
.Y(n_3169)
);

CKINVDCx5p33_ASAP7_75t_R g3170 ( 
.A(n_2667),
.Y(n_3170)
);

CKINVDCx5p33_ASAP7_75t_R g3171 ( 
.A(n_553),
.Y(n_3171)
);

CKINVDCx5p33_ASAP7_75t_R g3172 ( 
.A(n_2076),
.Y(n_3172)
);

CKINVDCx5p33_ASAP7_75t_R g3173 ( 
.A(n_2644),
.Y(n_3173)
);

CKINVDCx5p33_ASAP7_75t_R g3174 ( 
.A(n_604),
.Y(n_3174)
);

CKINVDCx5p33_ASAP7_75t_R g3175 ( 
.A(n_2626),
.Y(n_3175)
);

CKINVDCx5p33_ASAP7_75t_R g3176 ( 
.A(n_496),
.Y(n_3176)
);

CKINVDCx5p33_ASAP7_75t_R g3177 ( 
.A(n_2661),
.Y(n_3177)
);

CKINVDCx5p33_ASAP7_75t_R g3178 ( 
.A(n_1383),
.Y(n_3178)
);

CKINVDCx5p33_ASAP7_75t_R g3179 ( 
.A(n_385),
.Y(n_3179)
);

INVx1_ASAP7_75t_L g3180 ( 
.A(n_1168),
.Y(n_3180)
);

INVx1_ASAP7_75t_L g3181 ( 
.A(n_878),
.Y(n_3181)
);

CKINVDCx5p33_ASAP7_75t_R g3182 ( 
.A(n_2731),
.Y(n_3182)
);

BUFx5_ASAP7_75t_L g3183 ( 
.A(n_2748),
.Y(n_3183)
);

INVx1_ASAP7_75t_L g3184 ( 
.A(n_1244),
.Y(n_3184)
);

INVx1_ASAP7_75t_L g3185 ( 
.A(n_1496),
.Y(n_3185)
);

CKINVDCx5p33_ASAP7_75t_R g3186 ( 
.A(n_1217),
.Y(n_3186)
);

CKINVDCx5p33_ASAP7_75t_R g3187 ( 
.A(n_2605),
.Y(n_3187)
);

INVx1_ASAP7_75t_L g3188 ( 
.A(n_2442),
.Y(n_3188)
);

CKINVDCx5p33_ASAP7_75t_R g3189 ( 
.A(n_1784),
.Y(n_3189)
);

CKINVDCx5p33_ASAP7_75t_R g3190 ( 
.A(n_269),
.Y(n_3190)
);

CKINVDCx5p33_ASAP7_75t_R g3191 ( 
.A(n_2093),
.Y(n_3191)
);

INVx1_ASAP7_75t_SL g3192 ( 
.A(n_1401),
.Y(n_3192)
);

CKINVDCx5p33_ASAP7_75t_R g3193 ( 
.A(n_421),
.Y(n_3193)
);

CKINVDCx5p33_ASAP7_75t_R g3194 ( 
.A(n_2394),
.Y(n_3194)
);

CKINVDCx5p33_ASAP7_75t_R g3195 ( 
.A(n_2809),
.Y(n_3195)
);

INVx1_ASAP7_75t_L g3196 ( 
.A(n_89),
.Y(n_3196)
);

CKINVDCx5p33_ASAP7_75t_R g3197 ( 
.A(n_2311),
.Y(n_3197)
);

CKINVDCx5p33_ASAP7_75t_R g3198 ( 
.A(n_2304),
.Y(n_3198)
);

CKINVDCx5p33_ASAP7_75t_R g3199 ( 
.A(n_2678),
.Y(n_3199)
);

CKINVDCx5p33_ASAP7_75t_R g3200 ( 
.A(n_2357),
.Y(n_3200)
);

INVx1_ASAP7_75t_L g3201 ( 
.A(n_1316),
.Y(n_3201)
);

INVx2_ASAP7_75t_SL g3202 ( 
.A(n_627),
.Y(n_3202)
);

CKINVDCx5p33_ASAP7_75t_R g3203 ( 
.A(n_850),
.Y(n_3203)
);

INVx1_ASAP7_75t_L g3204 ( 
.A(n_1912),
.Y(n_3204)
);

CKINVDCx5p33_ASAP7_75t_R g3205 ( 
.A(n_994),
.Y(n_3205)
);

CKINVDCx5p33_ASAP7_75t_R g3206 ( 
.A(n_207),
.Y(n_3206)
);

HB1xp67_ASAP7_75t_L g3207 ( 
.A(n_2719),
.Y(n_3207)
);

CKINVDCx5p33_ASAP7_75t_R g3208 ( 
.A(n_448),
.Y(n_3208)
);

INVx2_ASAP7_75t_L g3209 ( 
.A(n_2671),
.Y(n_3209)
);

CKINVDCx5p33_ASAP7_75t_R g3210 ( 
.A(n_2805),
.Y(n_3210)
);

CKINVDCx5p33_ASAP7_75t_R g3211 ( 
.A(n_1436),
.Y(n_3211)
);

CKINVDCx5p33_ASAP7_75t_R g3212 ( 
.A(n_941),
.Y(n_3212)
);

INVx2_ASAP7_75t_L g3213 ( 
.A(n_1140),
.Y(n_3213)
);

CKINVDCx5p33_ASAP7_75t_R g3214 ( 
.A(n_989),
.Y(n_3214)
);

CKINVDCx5p33_ASAP7_75t_R g3215 ( 
.A(n_2625),
.Y(n_3215)
);

CKINVDCx5p33_ASAP7_75t_R g3216 ( 
.A(n_2726),
.Y(n_3216)
);

CKINVDCx20_ASAP7_75t_R g3217 ( 
.A(n_668),
.Y(n_3217)
);

INVx1_ASAP7_75t_SL g3218 ( 
.A(n_2280),
.Y(n_3218)
);

CKINVDCx5p33_ASAP7_75t_R g3219 ( 
.A(n_1995),
.Y(n_3219)
);

INVx1_ASAP7_75t_SL g3220 ( 
.A(n_1939),
.Y(n_3220)
);

CKINVDCx20_ASAP7_75t_R g3221 ( 
.A(n_2295),
.Y(n_3221)
);

CKINVDCx5p33_ASAP7_75t_R g3222 ( 
.A(n_1109),
.Y(n_3222)
);

CKINVDCx20_ASAP7_75t_R g3223 ( 
.A(n_834),
.Y(n_3223)
);

BUFx5_ASAP7_75t_L g3224 ( 
.A(n_1623),
.Y(n_3224)
);

CKINVDCx5p33_ASAP7_75t_R g3225 ( 
.A(n_1090),
.Y(n_3225)
);

INVx1_ASAP7_75t_L g3226 ( 
.A(n_2450),
.Y(n_3226)
);

INVx1_ASAP7_75t_SL g3227 ( 
.A(n_2739),
.Y(n_3227)
);

INVx2_ASAP7_75t_L g3228 ( 
.A(n_2625),
.Y(n_3228)
);

CKINVDCx5p33_ASAP7_75t_R g3229 ( 
.A(n_2427),
.Y(n_3229)
);

CKINVDCx20_ASAP7_75t_R g3230 ( 
.A(n_1025),
.Y(n_3230)
);

CKINVDCx5p33_ASAP7_75t_R g3231 ( 
.A(n_2549),
.Y(n_3231)
);

CKINVDCx5p33_ASAP7_75t_R g3232 ( 
.A(n_1809),
.Y(n_3232)
);

CKINVDCx5p33_ASAP7_75t_R g3233 ( 
.A(n_746),
.Y(n_3233)
);

CKINVDCx5p33_ASAP7_75t_R g3234 ( 
.A(n_2425),
.Y(n_3234)
);

CKINVDCx14_ASAP7_75t_R g3235 ( 
.A(n_688),
.Y(n_3235)
);

INVx1_ASAP7_75t_L g3236 ( 
.A(n_2495),
.Y(n_3236)
);

CKINVDCx20_ASAP7_75t_R g3237 ( 
.A(n_2624),
.Y(n_3237)
);

CKINVDCx5p33_ASAP7_75t_R g3238 ( 
.A(n_582),
.Y(n_3238)
);

INVx1_ASAP7_75t_L g3239 ( 
.A(n_2651),
.Y(n_3239)
);

CKINVDCx5p33_ASAP7_75t_R g3240 ( 
.A(n_660),
.Y(n_3240)
);

CKINVDCx5p33_ASAP7_75t_R g3241 ( 
.A(n_2645),
.Y(n_3241)
);

CKINVDCx5p33_ASAP7_75t_R g3242 ( 
.A(n_1455),
.Y(n_3242)
);

INVx1_ASAP7_75t_L g3243 ( 
.A(n_1388),
.Y(n_3243)
);

CKINVDCx5p33_ASAP7_75t_R g3244 ( 
.A(n_2314),
.Y(n_3244)
);

INVx1_ASAP7_75t_L g3245 ( 
.A(n_2117),
.Y(n_3245)
);

CKINVDCx5p33_ASAP7_75t_R g3246 ( 
.A(n_1597),
.Y(n_3246)
);

CKINVDCx20_ASAP7_75t_R g3247 ( 
.A(n_2759),
.Y(n_3247)
);

CKINVDCx5p33_ASAP7_75t_R g3248 ( 
.A(n_586),
.Y(n_3248)
);

INVx2_ASAP7_75t_SL g3249 ( 
.A(n_1545),
.Y(n_3249)
);

BUFx2_ASAP7_75t_L g3250 ( 
.A(n_1355),
.Y(n_3250)
);

CKINVDCx20_ASAP7_75t_R g3251 ( 
.A(n_1047),
.Y(n_3251)
);

CKINVDCx5p33_ASAP7_75t_R g3252 ( 
.A(n_1726),
.Y(n_3252)
);

CKINVDCx5p33_ASAP7_75t_R g3253 ( 
.A(n_1385),
.Y(n_3253)
);

CKINVDCx5p33_ASAP7_75t_R g3254 ( 
.A(n_1696),
.Y(n_3254)
);

BUFx2_ASAP7_75t_L g3255 ( 
.A(n_2421),
.Y(n_3255)
);

INVx1_ASAP7_75t_L g3256 ( 
.A(n_370),
.Y(n_3256)
);

CKINVDCx5p33_ASAP7_75t_R g3257 ( 
.A(n_2030),
.Y(n_3257)
);

CKINVDCx5p33_ASAP7_75t_R g3258 ( 
.A(n_2229),
.Y(n_3258)
);

CKINVDCx5p33_ASAP7_75t_R g3259 ( 
.A(n_62),
.Y(n_3259)
);

CKINVDCx5p33_ASAP7_75t_R g3260 ( 
.A(n_1814),
.Y(n_3260)
);

BUFx10_ASAP7_75t_L g3261 ( 
.A(n_2068),
.Y(n_3261)
);

INVx1_ASAP7_75t_SL g3262 ( 
.A(n_81),
.Y(n_3262)
);

CKINVDCx5p33_ASAP7_75t_R g3263 ( 
.A(n_2206),
.Y(n_3263)
);

CKINVDCx20_ASAP7_75t_R g3264 ( 
.A(n_1970),
.Y(n_3264)
);

BUFx10_ASAP7_75t_L g3265 ( 
.A(n_1620),
.Y(n_3265)
);

INVx2_ASAP7_75t_L g3266 ( 
.A(n_1500),
.Y(n_3266)
);

INVx1_ASAP7_75t_L g3267 ( 
.A(n_1616),
.Y(n_3267)
);

CKINVDCx5p33_ASAP7_75t_R g3268 ( 
.A(n_838),
.Y(n_3268)
);

BUFx5_ASAP7_75t_L g3269 ( 
.A(n_1399),
.Y(n_3269)
);

BUFx2_ASAP7_75t_L g3270 ( 
.A(n_1355),
.Y(n_3270)
);

CKINVDCx5p33_ASAP7_75t_R g3271 ( 
.A(n_1670),
.Y(n_3271)
);

BUFx10_ASAP7_75t_L g3272 ( 
.A(n_2372),
.Y(n_3272)
);

BUFx2_ASAP7_75t_L g3273 ( 
.A(n_459),
.Y(n_3273)
);

CKINVDCx5p33_ASAP7_75t_R g3274 ( 
.A(n_2707),
.Y(n_3274)
);

CKINVDCx5p33_ASAP7_75t_R g3275 ( 
.A(n_523),
.Y(n_3275)
);

CKINVDCx20_ASAP7_75t_R g3276 ( 
.A(n_1073),
.Y(n_3276)
);

INVx1_ASAP7_75t_L g3277 ( 
.A(n_1418),
.Y(n_3277)
);

CKINVDCx5p33_ASAP7_75t_R g3278 ( 
.A(n_425),
.Y(n_3278)
);

CKINVDCx5p33_ASAP7_75t_R g3279 ( 
.A(n_1183),
.Y(n_3279)
);

INVx1_ASAP7_75t_L g3280 ( 
.A(n_811),
.Y(n_3280)
);

CKINVDCx5p33_ASAP7_75t_R g3281 ( 
.A(n_378),
.Y(n_3281)
);

INVx1_ASAP7_75t_L g3282 ( 
.A(n_2432),
.Y(n_3282)
);

CKINVDCx20_ASAP7_75t_R g3283 ( 
.A(n_2629),
.Y(n_3283)
);

INVx2_ASAP7_75t_L g3284 ( 
.A(n_1483),
.Y(n_3284)
);

INVx1_ASAP7_75t_L g3285 ( 
.A(n_2477),
.Y(n_3285)
);

CKINVDCx5p33_ASAP7_75t_R g3286 ( 
.A(n_36),
.Y(n_3286)
);

INVx1_ASAP7_75t_L g3287 ( 
.A(n_341),
.Y(n_3287)
);

CKINVDCx5p33_ASAP7_75t_R g3288 ( 
.A(n_428),
.Y(n_3288)
);

CKINVDCx5p33_ASAP7_75t_R g3289 ( 
.A(n_2652),
.Y(n_3289)
);

INVx4_ASAP7_75t_R g3290 ( 
.A(n_241),
.Y(n_3290)
);

CKINVDCx5p33_ASAP7_75t_R g3291 ( 
.A(n_354),
.Y(n_3291)
);

CKINVDCx5p33_ASAP7_75t_R g3292 ( 
.A(n_2641),
.Y(n_3292)
);

CKINVDCx5p33_ASAP7_75t_R g3293 ( 
.A(n_1968),
.Y(n_3293)
);

CKINVDCx5p33_ASAP7_75t_R g3294 ( 
.A(n_2567),
.Y(n_3294)
);

BUFx3_ASAP7_75t_L g3295 ( 
.A(n_2016),
.Y(n_3295)
);

CKINVDCx5p33_ASAP7_75t_R g3296 ( 
.A(n_215),
.Y(n_3296)
);

CKINVDCx5p33_ASAP7_75t_R g3297 ( 
.A(n_2635),
.Y(n_3297)
);

INVx1_ASAP7_75t_L g3298 ( 
.A(n_2629),
.Y(n_3298)
);

BUFx3_ASAP7_75t_L g3299 ( 
.A(n_397),
.Y(n_3299)
);

CKINVDCx5p33_ASAP7_75t_R g3300 ( 
.A(n_2690),
.Y(n_3300)
);

INVx1_ASAP7_75t_L g3301 ( 
.A(n_1433),
.Y(n_3301)
);

INVx1_ASAP7_75t_L g3302 ( 
.A(n_468),
.Y(n_3302)
);

INVx2_ASAP7_75t_SL g3303 ( 
.A(n_181),
.Y(n_3303)
);

INVx1_ASAP7_75t_L g3304 ( 
.A(n_2048),
.Y(n_3304)
);

BUFx10_ASAP7_75t_L g3305 ( 
.A(n_1245),
.Y(n_3305)
);

CKINVDCx5p33_ASAP7_75t_R g3306 ( 
.A(n_996),
.Y(n_3306)
);

INVx1_ASAP7_75t_L g3307 ( 
.A(n_1027),
.Y(n_3307)
);

CKINVDCx5p33_ASAP7_75t_R g3308 ( 
.A(n_715),
.Y(n_3308)
);

CKINVDCx20_ASAP7_75t_R g3309 ( 
.A(n_2157),
.Y(n_3309)
);

CKINVDCx5p33_ASAP7_75t_R g3310 ( 
.A(n_1395),
.Y(n_3310)
);

CKINVDCx5p33_ASAP7_75t_R g3311 ( 
.A(n_1700),
.Y(n_3311)
);

BUFx10_ASAP7_75t_L g3312 ( 
.A(n_2623),
.Y(n_3312)
);

CKINVDCx20_ASAP7_75t_R g3313 ( 
.A(n_417),
.Y(n_3313)
);

CKINVDCx5p33_ASAP7_75t_R g3314 ( 
.A(n_2410),
.Y(n_3314)
);

HB1xp67_ASAP7_75t_L g3315 ( 
.A(n_2631),
.Y(n_3315)
);

INVx1_ASAP7_75t_L g3316 ( 
.A(n_1490),
.Y(n_3316)
);

INVx1_ASAP7_75t_L g3317 ( 
.A(n_2274),
.Y(n_3317)
);

CKINVDCx5p33_ASAP7_75t_R g3318 ( 
.A(n_834),
.Y(n_3318)
);

CKINVDCx5p33_ASAP7_75t_R g3319 ( 
.A(n_1480),
.Y(n_3319)
);

CKINVDCx5p33_ASAP7_75t_R g3320 ( 
.A(n_2654),
.Y(n_3320)
);

INVx1_ASAP7_75t_L g3321 ( 
.A(n_1534),
.Y(n_3321)
);

CKINVDCx5p33_ASAP7_75t_R g3322 ( 
.A(n_1233),
.Y(n_3322)
);

INVx1_ASAP7_75t_L g3323 ( 
.A(n_2),
.Y(n_3323)
);

CKINVDCx5p33_ASAP7_75t_R g3324 ( 
.A(n_1695),
.Y(n_3324)
);

INVx1_ASAP7_75t_L g3325 ( 
.A(n_2175),
.Y(n_3325)
);

CKINVDCx5p33_ASAP7_75t_R g3326 ( 
.A(n_578),
.Y(n_3326)
);

INVx2_ASAP7_75t_L g3327 ( 
.A(n_2539),
.Y(n_3327)
);

INVx2_ASAP7_75t_L g3328 ( 
.A(n_1872),
.Y(n_3328)
);

INVx2_ASAP7_75t_SL g3329 ( 
.A(n_713),
.Y(n_3329)
);

INVx1_ASAP7_75t_SL g3330 ( 
.A(n_2699),
.Y(n_3330)
);

BUFx5_ASAP7_75t_L g3331 ( 
.A(n_2744),
.Y(n_3331)
);

CKINVDCx5p33_ASAP7_75t_R g3332 ( 
.A(n_656),
.Y(n_3332)
);

CKINVDCx5p33_ASAP7_75t_R g3333 ( 
.A(n_2295),
.Y(n_3333)
);

CKINVDCx5p33_ASAP7_75t_R g3334 ( 
.A(n_1023),
.Y(n_3334)
);

CKINVDCx5p33_ASAP7_75t_R g3335 ( 
.A(n_2703),
.Y(n_3335)
);

INVx1_ASAP7_75t_L g3336 ( 
.A(n_2598),
.Y(n_3336)
);

INVx1_ASAP7_75t_SL g3337 ( 
.A(n_94),
.Y(n_3337)
);

CKINVDCx5p33_ASAP7_75t_R g3338 ( 
.A(n_2616),
.Y(n_3338)
);

INVx1_ASAP7_75t_L g3339 ( 
.A(n_1647),
.Y(n_3339)
);

CKINVDCx5p33_ASAP7_75t_R g3340 ( 
.A(n_2747),
.Y(n_3340)
);

CKINVDCx5p33_ASAP7_75t_R g3341 ( 
.A(n_603),
.Y(n_3341)
);

INVx1_ASAP7_75t_L g3342 ( 
.A(n_2461),
.Y(n_3342)
);

CKINVDCx5p33_ASAP7_75t_R g3343 ( 
.A(n_496),
.Y(n_3343)
);

BUFx10_ASAP7_75t_L g3344 ( 
.A(n_2311),
.Y(n_3344)
);

CKINVDCx5p33_ASAP7_75t_R g3345 ( 
.A(n_552),
.Y(n_3345)
);

CKINVDCx20_ASAP7_75t_R g3346 ( 
.A(n_149),
.Y(n_3346)
);

CKINVDCx5p33_ASAP7_75t_R g3347 ( 
.A(n_2273),
.Y(n_3347)
);

CKINVDCx5p33_ASAP7_75t_R g3348 ( 
.A(n_2051),
.Y(n_3348)
);

CKINVDCx14_ASAP7_75t_R g3349 ( 
.A(n_762),
.Y(n_3349)
);

INVx2_ASAP7_75t_SL g3350 ( 
.A(n_2428),
.Y(n_3350)
);

CKINVDCx16_ASAP7_75t_R g3351 ( 
.A(n_128),
.Y(n_3351)
);

INVx1_ASAP7_75t_L g3352 ( 
.A(n_2708),
.Y(n_3352)
);

INVx1_ASAP7_75t_L g3353 ( 
.A(n_55),
.Y(n_3353)
);

BUFx10_ASAP7_75t_L g3354 ( 
.A(n_1510),
.Y(n_3354)
);

INVx2_ASAP7_75t_SL g3355 ( 
.A(n_1274),
.Y(n_3355)
);

CKINVDCx5p33_ASAP7_75t_R g3356 ( 
.A(n_1900),
.Y(n_3356)
);

CKINVDCx20_ASAP7_75t_R g3357 ( 
.A(n_2030),
.Y(n_3357)
);

CKINVDCx5p33_ASAP7_75t_R g3358 ( 
.A(n_1944),
.Y(n_3358)
);

CKINVDCx5p33_ASAP7_75t_R g3359 ( 
.A(n_1003),
.Y(n_3359)
);

CKINVDCx20_ASAP7_75t_R g3360 ( 
.A(n_1601),
.Y(n_3360)
);

CKINVDCx5p33_ASAP7_75t_R g3361 ( 
.A(n_1597),
.Y(n_3361)
);

CKINVDCx5p33_ASAP7_75t_R g3362 ( 
.A(n_1331),
.Y(n_3362)
);

INVx1_ASAP7_75t_L g3363 ( 
.A(n_1228),
.Y(n_3363)
);

CKINVDCx5p33_ASAP7_75t_R g3364 ( 
.A(n_1530),
.Y(n_3364)
);

INVx1_ASAP7_75t_SL g3365 ( 
.A(n_557),
.Y(n_3365)
);

CKINVDCx5p33_ASAP7_75t_R g3366 ( 
.A(n_384),
.Y(n_3366)
);

CKINVDCx5p33_ASAP7_75t_R g3367 ( 
.A(n_1918),
.Y(n_3367)
);

CKINVDCx20_ASAP7_75t_R g3368 ( 
.A(n_23),
.Y(n_3368)
);

BUFx2_ASAP7_75t_L g3369 ( 
.A(n_2656),
.Y(n_3369)
);

CKINVDCx5p33_ASAP7_75t_R g3370 ( 
.A(n_2259),
.Y(n_3370)
);

CKINVDCx5p33_ASAP7_75t_R g3371 ( 
.A(n_2056),
.Y(n_3371)
);

CKINVDCx5p33_ASAP7_75t_R g3372 ( 
.A(n_2309),
.Y(n_3372)
);

INVx1_ASAP7_75t_L g3373 ( 
.A(n_356),
.Y(n_3373)
);

INVx1_ASAP7_75t_L g3374 ( 
.A(n_1043),
.Y(n_3374)
);

CKINVDCx5p33_ASAP7_75t_R g3375 ( 
.A(n_1347),
.Y(n_3375)
);

CKINVDCx5p33_ASAP7_75t_R g3376 ( 
.A(n_2570),
.Y(n_3376)
);

INVx1_ASAP7_75t_L g3377 ( 
.A(n_1494),
.Y(n_3377)
);

INVx1_ASAP7_75t_L g3378 ( 
.A(n_608),
.Y(n_3378)
);

CKINVDCx20_ASAP7_75t_R g3379 ( 
.A(n_1814),
.Y(n_3379)
);

INVx1_ASAP7_75t_L g3380 ( 
.A(n_2749),
.Y(n_3380)
);

INVx1_ASAP7_75t_SL g3381 ( 
.A(n_1241),
.Y(n_3381)
);

CKINVDCx5p33_ASAP7_75t_R g3382 ( 
.A(n_508),
.Y(n_3382)
);

INVx1_ASAP7_75t_L g3383 ( 
.A(n_2617),
.Y(n_3383)
);

CKINVDCx5p33_ASAP7_75t_R g3384 ( 
.A(n_2608),
.Y(n_3384)
);

BUFx2_ASAP7_75t_L g3385 ( 
.A(n_1561),
.Y(n_3385)
);

INVx1_ASAP7_75t_L g3386 ( 
.A(n_2615),
.Y(n_3386)
);

CKINVDCx5p33_ASAP7_75t_R g3387 ( 
.A(n_303),
.Y(n_3387)
);

CKINVDCx5p33_ASAP7_75t_R g3388 ( 
.A(n_2612),
.Y(n_3388)
);

CKINVDCx20_ASAP7_75t_R g3389 ( 
.A(n_1600),
.Y(n_3389)
);

INVx1_ASAP7_75t_L g3390 ( 
.A(n_1878),
.Y(n_3390)
);

INVx1_ASAP7_75t_L g3391 ( 
.A(n_339),
.Y(n_3391)
);

INVx2_ASAP7_75t_L g3392 ( 
.A(n_2417),
.Y(n_3392)
);

CKINVDCx20_ASAP7_75t_R g3393 ( 
.A(n_2278),
.Y(n_3393)
);

CKINVDCx5p33_ASAP7_75t_R g3394 ( 
.A(n_2662),
.Y(n_3394)
);

CKINVDCx5p33_ASAP7_75t_R g3395 ( 
.A(n_2052),
.Y(n_3395)
);

INVx1_ASAP7_75t_L g3396 ( 
.A(n_2633),
.Y(n_3396)
);

INVx2_ASAP7_75t_L g3397 ( 
.A(n_2716),
.Y(n_3397)
);

INVx1_ASAP7_75t_SL g3398 ( 
.A(n_2235),
.Y(n_3398)
);

CKINVDCx5p33_ASAP7_75t_R g3399 ( 
.A(n_2743),
.Y(n_3399)
);

INVx1_ASAP7_75t_L g3400 ( 
.A(n_1485),
.Y(n_3400)
);

BUFx6f_ASAP7_75t_L g3401 ( 
.A(n_1746),
.Y(n_3401)
);

CKINVDCx5p33_ASAP7_75t_R g3402 ( 
.A(n_2653),
.Y(n_3402)
);

CKINVDCx5p33_ASAP7_75t_R g3403 ( 
.A(n_501),
.Y(n_3403)
);

CKINVDCx20_ASAP7_75t_R g3404 ( 
.A(n_1993),
.Y(n_3404)
);

INVx1_ASAP7_75t_L g3405 ( 
.A(n_2575),
.Y(n_3405)
);

INVx1_ASAP7_75t_L g3406 ( 
.A(n_419),
.Y(n_3406)
);

CKINVDCx5p33_ASAP7_75t_R g3407 ( 
.A(n_1403),
.Y(n_3407)
);

INVx1_ASAP7_75t_L g3408 ( 
.A(n_2125),
.Y(n_3408)
);

INVx2_ASAP7_75t_SL g3409 ( 
.A(n_974),
.Y(n_3409)
);

CKINVDCx5p33_ASAP7_75t_R g3410 ( 
.A(n_1489),
.Y(n_3410)
);

INVx1_ASAP7_75t_L g3411 ( 
.A(n_1134),
.Y(n_3411)
);

CKINVDCx5p33_ASAP7_75t_R g3412 ( 
.A(n_744),
.Y(n_3412)
);

CKINVDCx16_ASAP7_75t_R g3413 ( 
.A(n_1235),
.Y(n_3413)
);

INVx1_ASAP7_75t_L g3414 ( 
.A(n_2754),
.Y(n_3414)
);

BUFx8_ASAP7_75t_SL g3415 ( 
.A(n_1496),
.Y(n_3415)
);

INVx2_ASAP7_75t_SL g3416 ( 
.A(n_1955),
.Y(n_3416)
);

INVx1_ASAP7_75t_L g3417 ( 
.A(n_325),
.Y(n_3417)
);

CKINVDCx5p33_ASAP7_75t_R g3418 ( 
.A(n_2435),
.Y(n_3418)
);

CKINVDCx5p33_ASAP7_75t_R g3419 ( 
.A(n_802),
.Y(n_3419)
);

CKINVDCx20_ASAP7_75t_R g3420 ( 
.A(n_1265),
.Y(n_3420)
);

INVx1_ASAP7_75t_SL g3421 ( 
.A(n_2381),
.Y(n_3421)
);

CKINVDCx5p33_ASAP7_75t_R g3422 ( 
.A(n_482),
.Y(n_3422)
);

INVx1_ASAP7_75t_SL g3423 ( 
.A(n_1403),
.Y(n_3423)
);

CKINVDCx5p33_ASAP7_75t_R g3424 ( 
.A(n_2714),
.Y(n_3424)
);

INVx1_ASAP7_75t_L g3425 ( 
.A(n_1607),
.Y(n_3425)
);

INVx1_ASAP7_75t_L g3426 ( 
.A(n_849),
.Y(n_3426)
);

CKINVDCx5p33_ASAP7_75t_R g3427 ( 
.A(n_2361),
.Y(n_3427)
);

INVx1_ASAP7_75t_L g3428 ( 
.A(n_2750),
.Y(n_3428)
);

CKINVDCx5p33_ASAP7_75t_R g3429 ( 
.A(n_517),
.Y(n_3429)
);

CKINVDCx5p33_ASAP7_75t_R g3430 ( 
.A(n_1789),
.Y(n_3430)
);

CKINVDCx5p33_ASAP7_75t_R g3431 ( 
.A(n_2269),
.Y(n_3431)
);

CKINVDCx5p33_ASAP7_75t_R g3432 ( 
.A(n_1858),
.Y(n_3432)
);

INVx2_ASAP7_75t_L g3433 ( 
.A(n_1862),
.Y(n_3433)
);

INVx2_ASAP7_75t_L g3434 ( 
.A(n_2671),
.Y(n_3434)
);

INVx1_ASAP7_75t_L g3435 ( 
.A(n_2504),
.Y(n_3435)
);

CKINVDCx5p33_ASAP7_75t_R g3436 ( 
.A(n_2737),
.Y(n_3436)
);

INVx1_ASAP7_75t_L g3437 ( 
.A(n_1330),
.Y(n_3437)
);

CKINVDCx20_ASAP7_75t_R g3438 ( 
.A(n_1194),
.Y(n_3438)
);

CKINVDCx5p33_ASAP7_75t_R g3439 ( 
.A(n_445),
.Y(n_3439)
);

INVx1_ASAP7_75t_L g3440 ( 
.A(n_1547),
.Y(n_3440)
);

INVxp67_ASAP7_75t_SL g3441 ( 
.A(n_934),
.Y(n_3441)
);

BUFx3_ASAP7_75t_L g3442 ( 
.A(n_1253),
.Y(n_3442)
);

CKINVDCx5p33_ASAP7_75t_R g3443 ( 
.A(n_2731),
.Y(n_3443)
);

CKINVDCx20_ASAP7_75t_R g3444 ( 
.A(n_2774),
.Y(n_3444)
);

CKINVDCx5p33_ASAP7_75t_R g3445 ( 
.A(n_1913),
.Y(n_3445)
);

CKINVDCx5p33_ASAP7_75t_R g3446 ( 
.A(n_1664),
.Y(n_3446)
);

INVx1_ASAP7_75t_L g3447 ( 
.A(n_2684),
.Y(n_3447)
);

HB1xp67_ASAP7_75t_L g3448 ( 
.A(n_1172),
.Y(n_3448)
);

CKINVDCx5p33_ASAP7_75t_R g3449 ( 
.A(n_1380),
.Y(n_3449)
);

CKINVDCx5p33_ASAP7_75t_R g3450 ( 
.A(n_2332),
.Y(n_3450)
);

CKINVDCx5p33_ASAP7_75t_R g3451 ( 
.A(n_2074),
.Y(n_3451)
);

INVx1_ASAP7_75t_L g3452 ( 
.A(n_2571),
.Y(n_3452)
);

CKINVDCx5p33_ASAP7_75t_R g3453 ( 
.A(n_256),
.Y(n_3453)
);

CKINVDCx5p33_ASAP7_75t_R g3454 ( 
.A(n_370),
.Y(n_3454)
);

CKINVDCx5p33_ASAP7_75t_R g3455 ( 
.A(n_1433),
.Y(n_3455)
);

CKINVDCx5p33_ASAP7_75t_R g3456 ( 
.A(n_1669),
.Y(n_3456)
);

INVx1_ASAP7_75t_L g3457 ( 
.A(n_1161),
.Y(n_3457)
);

BUFx2_ASAP7_75t_L g3458 ( 
.A(n_2514),
.Y(n_3458)
);

CKINVDCx5p33_ASAP7_75t_R g3459 ( 
.A(n_707),
.Y(n_3459)
);

CKINVDCx5p33_ASAP7_75t_R g3460 ( 
.A(n_1599),
.Y(n_3460)
);

CKINVDCx5p33_ASAP7_75t_R g3461 ( 
.A(n_697),
.Y(n_3461)
);

CKINVDCx5p33_ASAP7_75t_R g3462 ( 
.A(n_2742),
.Y(n_3462)
);

HB1xp67_ASAP7_75t_L g3463 ( 
.A(n_2532),
.Y(n_3463)
);

CKINVDCx5p33_ASAP7_75t_R g3464 ( 
.A(n_979),
.Y(n_3464)
);

CKINVDCx5p33_ASAP7_75t_R g3465 ( 
.A(n_676),
.Y(n_3465)
);

BUFx3_ASAP7_75t_L g3466 ( 
.A(n_758),
.Y(n_3466)
);

CKINVDCx16_ASAP7_75t_R g3467 ( 
.A(n_427),
.Y(n_3467)
);

INVx1_ASAP7_75t_L g3468 ( 
.A(n_1453),
.Y(n_3468)
);

CKINVDCx5p33_ASAP7_75t_R g3469 ( 
.A(n_74),
.Y(n_3469)
);

CKINVDCx5p33_ASAP7_75t_R g3470 ( 
.A(n_2660),
.Y(n_3470)
);

CKINVDCx5p33_ASAP7_75t_R g3471 ( 
.A(n_2588),
.Y(n_3471)
);

CKINVDCx5p33_ASAP7_75t_R g3472 ( 
.A(n_1646),
.Y(n_3472)
);

BUFx10_ASAP7_75t_L g3473 ( 
.A(n_993),
.Y(n_3473)
);

CKINVDCx5p33_ASAP7_75t_R g3474 ( 
.A(n_1307),
.Y(n_3474)
);

CKINVDCx5p33_ASAP7_75t_R g3475 ( 
.A(n_2753),
.Y(n_3475)
);

CKINVDCx5p33_ASAP7_75t_R g3476 ( 
.A(n_1456),
.Y(n_3476)
);

BUFx10_ASAP7_75t_L g3477 ( 
.A(n_338),
.Y(n_3477)
);

CKINVDCx20_ASAP7_75t_R g3478 ( 
.A(n_2382),
.Y(n_3478)
);

CKINVDCx5p33_ASAP7_75t_R g3479 ( 
.A(n_2801),
.Y(n_3479)
);

CKINVDCx20_ASAP7_75t_R g3480 ( 
.A(n_555),
.Y(n_3480)
);

CKINVDCx5p33_ASAP7_75t_R g3481 ( 
.A(n_2738),
.Y(n_3481)
);

BUFx6f_ASAP7_75t_L g3482 ( 
.A(n_849),
.Y(n_3482)
);

CKINVDCx5p33_ASAP7_75t_R g3483 ( 
.A(n_1923),
.Y(n_3483)
);

BUFx2_ASAP7_75t_L g3484 ( 
.A(n_1590),
.Y(n_3484)
);

INVx1_ASAP7_75t_L g3485 ( 
.A(n_1245),
.Y(n_3485)
);

INVx1_ASAP7_75t_L g3486 ( 
.A(n_1767),
.Y(n_3486)
);

INVx1_ASAP7_75t_L g3487 ( 
.A(n_1129),
.Y(n_3487)
);

BUFx3_ASAP7_75t_L g3488 ( 
.A(n_169),
.Y(n_3488)
);

BUFx3_ASAP7_75t_L g3489 ( 
.A(n_416),
.Y(n_3489)
);

INVxp33_ASAP7_75t_L g3490 ( 
.A(n_1653),
.Y(n_3490)
);

INVx1_ASAP7_75t_L g3491 ( 
.A(n_1890),
.Y(n_3491)
);

INVx1_ASAP7_75t_L g3492 ( 
.A(n_1294),
.Y(n_3492)
);

INVx1_ASAP7_75t_L g3493 ( 
.A(n_2741),
.Y(n_3493)
);

BUFx6f_ASAP7_75t_L g3494 ( 
.A(n_464),
.Y(n_3494)
);

INVx1_ASAP7_75t_L g3495 ( 
.A(n_2211),
.Y(n_3495)
);

CKINVDCx5p33_ASAP7_75t_R g3496 ( 
.A(n_234),
.Y(n_3496)
);

CKINVDCx16_ASAP7_75t_R g3497 ( 
.A(n_2698),
.Y(n_3497)
);

CKINVDCx5p33_ASAP7_75t_R g3498 ( 
.A(n_2509),
.Y(n_3498)
);

INVx1_ASAP7_75t_L g3499 ( 
.A(n_2562),
.Y(n_3499)
);

HB1xp67_ASAP7_75t_L g3500 ( 
.A(n_2079),
.Y(n_3500)
);

CKINVDCx20_ASAP7_75t_R g3501 ( 
.A(n_1359),
.Y(n_3501)
);

INVx1_ASAP7_75t_L g3502 ( 
.A(n_1284),
.Y(n_3502)
);

CKINVDCx5p33_ASAP7_75t_R g3503 ( 
.A(n_684),
.Y(n_3503)
);

BUFx6f_ASAP7_75t_L g3504 ( 
.A(n_1846),
.Y(n_3504)
);

CKINVDCx20_ASAP7_75t_R g3505 ( 
.A(n_794),
.Y(n_3505)
);

INVx1_ASAP7_75t_L g3506 ( 
.A(n_2406),
.Y(n_3506)
);

INVx1_ASAP7_75t_L g3507 ( 
.A(n_385),
.Y(n_3507)
);

CKINVDCx5p33_ASAP7_75t_R g3508 ( 
.A(n_1982),
.Y(n_3508)
);

INVx1_ASAP7_75t_L g3509 ( 
.A(n_402),
.Y(n_3509)
);

INVx1_ASAP7_75t_SL g3510 ( 
.A(n_2153),
.Y(n_3510)
);

CKINVDCx20_ASAP7_75t_R g3511 ( 
.A(n_1611),
.Y(n_3511)
);

INVx1_ASAP7_75t_SL g3512 ( 
.A(n_2715),
.Y(n_3512)
);

INVx1_ASAP7_75t_L g3513 ( 
.A(n_1281),
.Y(n_3513)
);

CKINVDCx5p33_ASAP7_75t_R g3514 ( 
.A(n_888),
.Y(n_3514)
);

CKINVDCx5p33_ASAP7_75t_R g3515 ( 
.A(n_2341),
.Y(n_3515)
);

CKINVDCx5p33_ASAP7_75t_R g3516 ( 
.A(n_2490),
.Y(n_3516)
);

INVx1_ASAP7_75t_L g3517 ( 
.A(n_918),
.Y(n_3517)
);

INVx1_ASAP7_75t_L g3518 ( 
.A(n_2016),
.Y(n_3518)
);

BUFx10_ASAP7_75t_L g3519 ( 
.A(n_2456),
.Y(n_3519)
);

CKINVDCx5p33_ASAP7_75t_R g3520 ( 
.A(n_333),
.Y(n_3520)
);

CKINVDCx5p33_ASAP7_75t_R g3521 ( 
.A(n_1232),
.Y(n_3521)
);

CKINVDCx5p33_ASAP7_75t_R g3522 ( 
.A(n_2634),
.Y(n_3522)
);

CKINVDCx5p33_ASAP7_75t_R g3523 ( 
.A(n_411),
.Y(n_3523)
);

CKINVDCx5p33_ASAP7_75t_R g3524 ( 
.A(n_2519),
.Y(n_3524)
);

CKINVDCx5p33_ASAP7_75t_R g3525 ( 
.A(n_1184),
.Y(n_3525)
);

INVx1_ASAP7_75t_L g3526 ( 
.A(n_2384),
.Y(n_3526)
);

CKINVDCx5p33_ASAP7_75t_R g3527 ( 
.A(n_259),
.Y(n_3527)
);

CKINVDCx5p33_ASAP7_75t_R g3528 ( 
.A(n_2582),
.Y(n_3528)
);

BUFx6f_ASAP7_75t_L g3529 ( 
.A(n_365),
.Y(n_3529)
);

INVx1_ASAP7_75t_L g3530 ( 
.A(n_1939),
.Y(n_3530)
);

INVx1_ASAP7_75t_L g3531 ( 
.A(n_2729),
.Y(n_3531)
);

CKINVDCx5p33_ASAP7_75t_R g3532 ( 
.A(n_570),
.Y(n_3532)
);

INVx1_ASAP7_75t_L g3533 ( 
.A(n_903),
.Y(n_3533)
);

INVx1_ASAP7_75t_L g3534 ( 
.A(n_1449),
.Y(n_3534)
);

CKINVDCx5p33_ASAP7_75t_R g3535 ( 
.A(n_706),
.Y(n_3535)
);

CKINVDCx5p33_ASAP7_75t_R g3536 ( 
.A(n_965),
.Y(n_3536)
);

CKINVDCx5p33_ASAP7_75t_R g3537 ( 
.A(n_2205),
.Y(n_3537)
);

CKINVDCx5p33_ASAP7_75t_R g3538 ( 
.A(n_247),
.Y(n_3538)
);

CKINVDCx5p33_ASAP7_75t_R g3539 ( 
.A(n_2125),
.Y(n_3539)
);

INVx1_ASAP7_75t_L g3540 ( 
.A(n_2460),
.Y(n_3540)
);

CKINVDCx5p33_ASAP7_75t_R g3541 ( 
.A(n_112),
.Y(n_3541)
);

CKINVDCx5p33_ASAP7_75t_R g3542 ( 
.A(n_628),
.Y(n_3542)
);

INVx1_ASAP7_75t_L g3543 ( 
.A(n_2659),
.Y(n_3543)
);

CKINVDCx5p33_ASAP7_75t_R g3544 ( 
.A(n_2474),
.Y(n_3544)
);

INVx2_ASAP7_75t_L g3545 ( 
.A(n_1582),
.Y(n_3545)
);

CKINVDCx5p33_ASAP7_75t_R g3546 ( 
.A(n_1891),
.Y(n_3546)
);

CKINVDCx5p33_ASAP7_75t_R g3547 ( 
.A(n_2677),
.Y(n_3547)
);

CKINVDCx14_ASAP7_75t_R g3548 ( 
.A(n_1646),
.Y(n_3548)
);

INVx1_ASAP7_75t_L g3549 ( 
.A(n_1341),
.Y(n_3549)
);

CKINVDCx20_ASAP7_75t_R g3550 ( 
.A(n_2668),
.Y(n_3550)
);

CKINVDCx5p33_ASAP7_75t_R g3551 ( 
.A(n_1636),
.Y(n_3551)
);

CKINVDCx5p33_ASAP7_75t_R g3552 ( 
.A(n_1909),
.Y(n_3552)
);

BUFx3_ASAP7_75t_L g3553 ( 
.A(n_2042),
.Y(n_3553)
);

CKINVDCx5p33_ASAP7_75t_R g3554 ( 
.A(n_586),
.Y(n_3554)
);

INVx1_ASAP7_75t_L g3555 ( 
.A(n_1211),
.Y(n_3555)
);

CKINVDCx5p33_ASAP7_75t_R g3556 ( 
.A(n_2711),
.Y(n_3556)
);

CKINVDCx5p33_ASAP7_75t_R g3557 ( 
.A(n_143),
.Y(n_3557)
);

CKINVDCx20_ASAP7_75t_R g3558 ( 
.A(n_31),
.Y(n_3558)
);

CKINVDCx5p33_ASAP7_75t_R g3559 ( 
.A(n_1429),
.Y(n_3559)
);

CKINVDCx5p33_ASAP7_75t_R g3560 ( 
.A(n_2613),
.Y(n_3560)
);

CKINVDCx5p33_ASAP7_75t_R g3561 ( 
.A(n_2155),
.Y(n_3561)
);

CKINVDCx20_ASAP7_75t_R g3562 ( 
.A(n_2720),
.Y(n_3562)
);

CKINVDCx20_ASAP7_75t_R g3563 ( 
.A(n_335),
.Y(n_3563)
);

CKINVDCx5p33_ASAP7_75t_R g3564 ( 
.A(n_1146),
.Y(n_3564)
);

INVx1_ASAP7_75t_L g3565 ( 
.A(n_1937),
.Y(n_3565)
);

CKINVDCx5p33_ASAP7_75t_R g3566 ( 
.A(n_958),
.Y(n_3566)
);

CKINVDCx5p33_ASAP7_75t_R g3567 ( 
.A(n_2700),
.Y(n_3567)
);

INVx2_ASAP7_75t_L g3568 ( 
.A(n_1554),
.Y(n_3568)
);

INVx1_ASAP7_75t_L g3569 ( 
.A(n_1662),
.Y(n_3569)
);

CKINVDCx5p33_ASAP7_75t_R g3570 ( 
.A(n_631),
.Y(n_3570)
);

CKINVDCx5p33_ASAP7_75t_R g3571 ( 
.A(n_2692),
.Y(n_3571)
);

CKINVDCx5p33_ASAP7_75t_R g3572 ( 
.A(n_1019),
.Y(n_3572)
);

CKINVDCx5p33_ASAP7_75t_R g3573 ( 
.A(n_288),
.Y(n_3573)
);

CKINVDCx5p33_ASAP7_75t_R g3574 ( 
.A(n_2744),
.Y(n_3574)
);

CKINVDCx5p33_ASAP7_75t_R g3575 ( 
.A(n_905),
.Y(n_3575)
);

CKINVDCx5p33_ASAP7_75t_R g3576 ( 
.A(n_1909),
.Y(n_3576)
);

INVxp67_ASAP7_75t_L g3577 ( 
.A(n_109),
.Y(n_3577)
);

INVx1_ASAP7_75t_SL g3578 ( 
.A(n_1077),
.Y(n_3578)
);

BUFx3_ASAP7_75t_L g3579 ( 
.A(n_2186),
.Y(n_3579)
);

INVx1_ASAP7_75t_SL g3580 ( 
.A(n_1147),
.Y(n_3580)
);

BUFx2_ASAP7_75t_L g3581 ( 
.A(n_592),
.Y(n_3581)
);

CKINVDCx20_ASAP7_75t_R g3582 ( 
.A(n_1397),
.Y(n_3582)
);

CKINVDCx5p33_ASAP7_75t_R g3583 ( 
.A(n_244),
.Y(n_3583)
);

INVx1_ASAP7_75t_L g3584 ( 
.A(n_646),
.Y(n_3584)
);

INVx1_ASAP7_75t_L g3585 ( 
.A(n_2256),
.Y(n_3585)
);

INVxp67_ASAP7_75t_L g3586 ( 
.A(n_2521),
.Y(n_3586)
);

INVx2_ASAP7_75t_SL g3587 ( 
.A(n_106),
.Y(n_3587)
);

CKINVDCx5p33_ASAP7_75t_R g3588 ( 
.A(n_998),
.Y(n_3588)
);

CKINVDCx5p33_ASAP7_75t_R g3589 ( 
.A(n_1828),
.Y(n_3589)
);

CKINVDCx20_ASAP7_75t_R g3590 ( 
.A(n_2503),
.Y(n_3590)
);

CKINVDCx5p33_ASAP7_75t_R g3591 ( 
.A(n_1244),
.Y(n_3591)
);

INVx1_ASAP7_75t_SL g3592 ( 
.A(n_2249),
.Y(n_3592)
);

INVx2_ASAP7_75t_L g3593 ( 
.A(n_526),
.Y(n_3593)
);

CKINVDCx5p33_ASAP7_75t_R g3594 ( 
.A(n_2286),
.Y(n_3594)
);

CKINVDCx5p33_ASAP7_75t_R g3595 ( 
.A(n_347),
.Y(n_3595)
);

CKINVDCx5p33_ASAP7_75t_R g3596 ( 
.A(n_1412),
.Y(n_3596)
);

CKINVDCx14_ASAP7_75t_R g3597 ( 
.A(n_1095),
.Y(n_3597)
);

INVx2_ASAP7_75t_SL g3598 ( 
.A(n_1083),
.Y(n_3598)
);

CKINVDCx5p33_ASAP7_75t_R g3599 ( 
.A(n_2021),
.Y(n_3599)
);

CKINVDCx20_ASAP7_75t_R g3600 ( 
.A(n_1375),
.Y(n_3600)
);

INVx1_ASAP7_75t_L g3601 ( 
.A(n_1124),
.Y(n_3601)
);

CKINVDCx5p33_ASAP7_75t_R g3602 ( 
.A(n_171),
.Y(n_3602)
);

INVx1_ASAP7_75t_L g3603 ( 
.A(n_2593),
.Y(n_3603)
);

INVx2_ASAP7_75t_SL g3604 ( 
.A(n_55),
.Y(n_3604)
);

INVx1_ASAP7_75t_L g3605 ( 
.A(n_145),
.Y(n_3605)
);

INVxp33_ASAP7_75t_R g3606 ( 
.A(n_986),
.Y(n_3606)
);

INVx1_ASAP7_75t_L g3607 ( 
.A(n_2564),
.Y(n_3607)
);

CKINVDCx5p33_ASAP7_75t_R g3608 ( 
.A(n_1841),
.Y(n_3608)
);

CKINVDCx5p33_ASAP7_75t_R g3609 ( 
.A(n_1530),
.Y(n_3609)
);

CKINVDCx5p33_ASAP7_75t_R g3610 ( 
.A(n_565),
.Y(n_3610)
);

CKINVDCx5p33_ASAP7_75t_R g3611 ( 
.A(n_647),
.Y(n_3611)
);

CKINVDCx5p33_ASAP7_75t_R g3612 ( 
.A(n_2037),
.Y(n_3612)
);

CKINVDCx5p33_ASAP7_75t_R g3613 ( 
.A(n_2206),
.Y(n_3613)
);

BUFx10_ASAP7_75t_L g3614 ( 
.A(n_2301),
.Y(n_3614)
);

CKINVDCx5p33_ASAP7_75t_R g3615 ( 
.A(n_1458),
.Y(n_3615)
);

CKINVDCx5p33_ASAP7_75t_R g3616 ( 
.A(n_2364),
.Y(n_3616)
);

CKINVDCx20_ASAP7_75t_R g3617 ( 
.A(n_2088),
.Y(n_3617)
);

CKINVDCx20_ASAP7_75t_R g3618 ( 
.A(n_1659),
.Y(n_3618)
);

CKINVDCx5p33_ASAP7_75t_R g3619 ( 
.A(n_365),
.Y(n_3619)
);

CKINVDCx5p33_ASAP7_75t_R g3620 ( 
.A(n_479),
.Y(n_3620)
);

INVx1_ASAP7_75t_SL g3621 ( 
.A(n_2371),
.Y(n_3621)
);

INVx1_ASAP7_75t_L g3622 ( 
.A(n_2565),
.Y(n_3622)
);

INVx1_ASAP7_75t_L g3623 ( 
.A(n_2774),
.Y(n_3623)
);

CKINVDCx5p33_ASAP7_75t_R g3624 ( 
.A(n_2298),
.Y(n_3624)
);

INVx1_ASAP7_75t_L g3625 ( 
.A(n_2636),
.Y(n_3625)
);

CKINVDCx5p33_ASAP7_75t_R g3626 ( 
.A(n_2721),
.Y(n_3626)
);

INVx2_ASAP7_75t_L g3627 ( 
.A(n_2253),
.Y(n_3627)
);

INVx1_ASAP7_75t_L g3628 ( 
.A(n_865),
.Y(n_3628)
);

BUFx10_ASAP7_75t_L g3629 ( 
.A(n_1201),
.Y(n_3629)
);

CKINVDCx5p33_ASAP7_75t_R g3630 ( 
.A(n_1643),
.Y(n_3630)
);

BUFx3_ASAP7_75t_L g3631 ( 
.A(n_571),
.Y(n_3631)
);

CKINVDCx20_ASAP7_75t_R g3632 ( 
.A(n_1507),
.Y(n_3632)
);

INVx2_ASAP7_75t_L g3633 ( 
.A(n_826),
.Y(n_3633)
);

CKINVDCx5p33_ASAP7_75t_R g3634 ( 
.A(n_1708),
.Y(n_3634)
);

CKINVDCx5p33_ASAP7_75t_R g3635 ( 
.A(n_2059),
.Y(n_3635)
);

INVx2_ASAP7_75t_L g3636 ( 
.A(n_667),
.Y(n_3636)
);

CKINVDCx5p33_ASAP7_75t_R g3637 ( 
.A(n_2000),
.Y(n_3637)
);

CKINVDCx5p33_ASAP7_75t_R g3638 ( 
.A(n_2694),
.Y(n_3638)
);

CKINVDCx5p33_ASAP7_75t_R g3639 ( 
.A(n_2395),
.Y(n_3639)
);

INVx2_ASAP7_75t_L g3640 ( 
.A(n_2695),
.Y(n_3640)
);

CKINVDCx5p33_ASAP7_75t_R g3641 ( 
.A(n_731),
.Y(n_3641)
);

CKINVDCx5p33_ASAP7_75t_R g3642 ( 
.A(n_638),
.Y(n_3642)
);

CKINVDCx5p33_ASAP7_75t_R g3643 ( 
.A(n_2632),
.Y(n_3643)
);

CKINVDCx20_ASAP7_75t_R g3644 ( 
.A(n_2164),
.Y(n_3644)
);

CKINVDCx20_ASAP7_75t_R g3645 ( 
.A(n_2644),
.Y(n_3645)
);

INVx1_ASAP7_75t_L g3646 ( 
.A(n_1128),
.Y(n_3646)
);

CKINVDCx5p33_ASAP7_75t_R g3647 ( 
.A(n_2561),
.Y(n_3647)
);

CKINVDCx5p33_ASAP7_75t_R g3648 ( 
.A(n_2376),
.Y(n_3648)
);

CKINVDCx5p33_ASAP7_75t_R g3649 ( 
.A(n_2585),
.Y(n_3649)
);

CKINVDCx5p33_ASAP7_75t_R g3650 ( 
.A(n_1476),
.Y(n_3650)
);

CKINVDCx5p33_ASAP7_75t_R g3651 ( 
.A(n_2492),
.Y(n_3651)
);

INVx1_ASAP7_75t_SL g3652 ( 
.A(n_2159),
.Y(n_3652)
);

CKINVDCx20_ASAP7_75t_R g3653 ( 
.A(n_1512),
.Y(n_3653)
);

CKINVDCx5p33_ASAP7_75t_R g3654 ( 
.A(n_2648),
.Y(n_3654)
);

BUFx5_ASAP7_75t_L g3655 ( 
.A(n_2459),
.Y(n_3655)
);

INVx1_ASAP7_75t_L g3656 ( 
.A(n_978),
.Y(n_3656)
);

INVx1_ASAP7_75t_L g3657 ( 
.A(n_1777),
.Y(n_3657)
);

BUFx5_ASAP7_75t_L g3658 ( 
.A(n_184),
.Y(n_3658)
);

INVx1_ASAP7_75t_L g3659 ( 
.A(n_1979),
.Y(n_3659)
);

CKINVDCx5p33_ASAP7_75t_R g3660 ( 
.A(n_1264),
.Y(n_3660)
);

INVx2_ASAP7_75t_L g3661 ( 
.A(n_214),
.Y(n_3661)
);

CKINVDCx5p33_ASAP7_75t_R g3662 ( 
.A(n_1987),
.Y(n_3662)
);

CKINVDCx5p33_ASAP7_75t_R g3663 ( 
.A(n_2428),
.Y(n_3663)
);

CKINVDCx5p33_ASAP7_75t_R g3664 ( 
.A(n_2530),
.Y(n_3664)
);

CKINVDCx20_ASAP7_75t_R g3665 ( 
.A(n_1334),
.Y(n_3665)
);

CKINVDCx5p33_ASAP7_75t_R g3666 ( 
.A(n_742),
.Y(n_3666)
);

CKINVDCx5p33_ASAP7_75t_R g3667 ( 
.A(n_574),
.Y(n_3667)
);

CKINVDCx5p33_ASAP7_75t_R g3668 ( 
.A(n_222),
.Y(n_3668)
);

INVx1_ASAP7_75t_L g3669 ( 
.A(n_1416),
.Y(n_3669)
);

INVx1_ASAP7_75t_L g3670 ( 
.A(n_1827),
.Y(n_3670)
);

INVx1_ASAP7_75t_L g3671 ( 
.A(n_939),
.Y(n_3671)
);

CKINVDCx5p33_ASAP7_75t_R g3672 ( 
.A(n_2313),
.Y(n_3672)
);

CKINVDCx5p33_ASAP7_75t_R g3673 ( 
.A(n_1020),
.Y(n_3673)
);

INVx1_ASAP7_75t_L g3674 ( 
.A(n_1732),
.Y(n_3674)
);

CKINVDCx5p33_ASAP7_75t_R g3675 ( 
.A(n_1891),
.Y(n_3675)
);

CKINVDCx5p33_ASAP7_75t_R g3676 ( 
.A(n_116),
.Y(n_3676)
);

INVx1_ASAP7_75t_L g3677 ( 
.A(n_2578),
.Y(n_3677)
);

CKINVDCx5p33_ASAP7_75t_R g3678 ( 
.A(n_2208),
.Y(n_3678)
);

INVx1_ASAP7_75t_L g3679 ( 
.A(n_2694),
.Y(n_3679)
);

CKINVDCx20_ASAP7_75t_R g3680 ( 
.A(n_2673),
.Y(n_3680)
);

CKINVDCx5p33_ASAP7_75t_R g3681 ( 
.A(n_281),
.Y(n_3681)
);

CKINVDCx5p33_ASAP7_75t_R g3682 ( 
.A(n_2168),
.Y(n_3682)
);

CKINVDCx5p33_ASAP7_75t_R g3683 ( 
.A(n_984),
.Y(n_3683)
);

INVx1_ASAP7_75t_L g3684 ( 
.A(n_2611),
.Y(n_3684)
);

CKINVDCx5p33_ASAP7_75t_R g3685 ( 
.A(n_2429),
.Y(n_3685)
);

INVx1_ASAP7_75t_L g3686 ( 
.A(n_2556),
.Y(n_3686)
);

CKINVDCx20_ASAP7_75t_R g3687 ( 
.A(n_860),
.Y(n_3687)
);

INVxp33_ASAP7_75t_SL g3688 ( 
.A(n_1479),
.Y(n_3688)
);

INVx1_ASAP7_75t_L g3689 ( 
.A(n_2730),
.Y(n_3689)
);

CKINVDCx5p33_ASAP7_75t_R g3690 ( 
.A(n_95),
.Y(n_3690)
);

INVx1_ASAP7_75t_L g3691 ( 
.A(n_1021),
.Y(n_3691)
);

INVx1_ASAP7_75t_L g3692 ( 
.A(n_916),
.Y(n_3692)
);

CKINVDCx5p33_ASAP7_75t_R g3693 ( 
.A(n_400),
.Y(n_3693)
);

CKINVDCx5p33_ASAP7_75t_R g3694 ( 
.A(n_2736),
.Y(n_3694)
);

CKINVDCx5p33_ASAP7_75t_R g3695 ( 
.A(n_1320),
.Y(n_3695)
);

INVx1_ASAP7_75t_SL g3696 ( 
.A(n_815),
.Y(n_3696)
);

CKINVDCx5p33_ASAP7_75t_R g3697 ( 
.A(n_1324),
.Y(n_3697)
);

BUFx2_ASAP7_75t_SL g3698 ( 
.A(n_1308),
.Y(n_3698)
);

CKINVDCx5p33_ASAP7_75t_R g3699 ( 
.A(n_1211),
.Y(n_3699)
);

CKINVDCx5p33_ASAP7_75t_R g3700 ( 
.A(n_2321),
.Y(n_3700)
);

CKINVDCx20_ASAP7_75t_R g3701 ( 
.A(n_2471),
.Y(n_3701)
);

BUFx3_ASAP7_75t_L g3702 ( 
.A(n_1209),
.Y(n_3702)
);

CKINVDCx5p33_ASAP7_75t_R g3703 ( 
.A(n_208),
.Y(n_3703)
);

INVx1_ASAP7_75t_L g3704 ( 
.A(n_2643),
.Y(n_3704)
);

BUFx6f_ASAP7_75t_L g3705 ( 
.A(n_1232),
.Y(n_3705)
);

CKINVDCx16_ASAP7_75t_R g3706 ( 
.A(n_289),
.Y(n_3706)
);

CKINVDCx14_ASAP7_75t_R g3707 ( 
.A(n_376),
.Y(n_3707)
);

CKINVDCx16_ASAP7_75t_R g3708 ( 
.A(n_2484),
.Y(n_3708)
);

CKINVDCx5p33_ASAP7_75t_R g3709 ( 
.A(n_2018),
.Y(n_3709)
);

CKINVDCx5p33_ASAP7_75t_R g3710 ( 
.A(n_1113),
.Y(n_3710)
);

INVx2_ASAP7_75t_L g3711 ( 
.A(n_1862),
.Y(n_3711)
);

BUFx3_ASAP7_75t_L g3712 ( 
.A(n_1384),
.Y(n_3712)
);

CKINVDCx5p33_ASAP7_75t_R g3713 ( 
.A(n_2665),
.Y(n_3713)
);

CKINVDCx5p33_ASAP7_75t_R g3714 ( 
.A(n_1682),
.Y(n_3714)
);

CKINVDCx5p33_ASAP7_75t_R g3715 ( 
.A(n_671),
.Y(n_3715)
);

CKINVDCx5p33_ASAP7_75t_R g3716 ( 
.A(n_2202),
.Y(n_3716)
);

INVx1_ASAP7_75t_L g3717 ( 
.A(n_2663),
.Y(n_3717)
);

CKINVDCx5p33_ASAP7_75t_R g3718 ( 
.A(n_2622),
.Y(n_3718)
);

CKINVDCx5p33_ASAP7_75t_R g3719 ( 
.A(n_603),
.Y(n_3719)
);

CKINVDCx5p33_ASAP7_75t_R g3720 ( 
.A(n_2611),
.Y(n_3720)
);

INVx1_ASAP7_75t_L g3721 ( 
.A(n_1150),
.Y(n_3721)
);

INVx1_ASAP7_75t_L g3722 ( 
.A(n_1443),
.Y(n_3722)
);

CKINVDCx5p33_ASAP7_75t_R g3723 ( 
.A(n_1389),
.Y(n_3723)
);

INVx1_ASAP7_75t_SL g3724 ( 
.A(n_62),
.Y(n_3724)
);

CKINVDCx5p33_ASAP7_75t_R g3725 ( 
.A(n_2562),
.Y(n_3725)
);

CKINVDCx5p33_ASAP7_75t_R g3726 ( 
.A(n_651),
.Y(n_3726)
);

CKINVDCx16_ASAP7_75t_R g3727 ( 
.A(n_1396),
.Y(n_3727)
);

CKINVDCx20_ASAP7_75t_R g3728 ( 
.A(n_901),
.Y(n_3728)
);

INVx4_ASAP7_75t_R g3729 ( 
.A(n_97),
.Y(n_3729)
);

INVx1_ASAP7_75t_L g3730 ( 
.A(n_526),
.Y(n_3730)
);

BUFx3_ASAP7_75t_L g3731 ( 
.A(n_346),
.Y(n_3731)
);

CKINVDCx5p33_ASAP7_75t_R g3732 ( 
.A(n_2260),
.Y(n_3732)
);

CKINVDCx5p33_ASAP7_75t_R g3733 ( 
.A(n_1714),
.Y(n_3733)
);

BUFx10_ASAP7_75t_L g3734 ( 
.A(n_1710),
.Y(n_3734)
);

INVx1_ASAP7_75t_L g3735 ( 
.A(n_2344),
.Y(n_3735)
);

CKINVDCx5p33_ASAP7_75t_R g3736 ( 
.A(n_2039),
.Y(n_3736)
);

BUFx5_ASAP7_75t_L g3737 ( 
.A(n_1103),
.Y(n_3737)
);

CKINVDCx5p33_ASAP7_75t_R g3738 ( 
.A(n_2752),
.Y(n_3738)
);

CKINVDCx5p33_ASAP7_75t_R g3739 ( 
.A(n_2649),
.Y(n_3739)
);

CKINVDCx5p33_ASAP7_75t_R g3740 ( 
.A(n_1304),
.Y(n_3740)
);

INVx1_ASAP7_75t_L g3741 ( 
.A(n_1535),
.Y(n_3741)
);

CKINVDCx5p33_ASAP7_75t_R g3742 ( 
.A(n_277),
.Y(n_3742)
);

INVx2_ASAP7_75t_SL g3743 ( 
.A(n_1523),
.Y(n_3743)
);

INVx1_ASAP7_75t_L g3744 ( 
.A(n_2356),
.Y(n_3744)
);

CKINVDCx5p33_ASAP7_75t_R g3745 ( 
.A(n_424),
.Y(n_3745)
);

CKINVDCx5p33_ASAP7_75t_R g3746 ( 
.A(n_2706),
.Y(n_3746)
);

CKINVDCx5p33_ASAP7_75t_R g3747 ( 
.A(n_1195),
.Y(n_3747)
);

CKINVDCx5p33_ASAP7_75t_R g3748 ( 
.A(n_1610),
.Y(n_3748)
);

INVx1_ASAP7_75t_L g3749 ( 
.A(n_2014),
.Y(n_3749)
);

CKINVDCx5p33_ASAP7_75t_R g3750 ( 
.A(n_2124),
.Y(n_3750)
);

CKINVDCx5p33_ASAP7_75t_R g3751 ( 
.A(n_2574),
.Y(n_3751)
);

INVx1_ASAP7_75t_SL g3752 ( 
.A(n_637),
.Y(n_3752)
);

BUFx10_ASAP7_75t_L g3753 ( 
.A(n_445),
.Y(n_3753)
);

BUFx10_ASAP7_75t_L g3754 ( 
.A(n_1113),
.Y(n_3754)
);

INVx1_ASAP7_75t_L g3755 ( 
.A(n_372),
.Y(n_3755)
);

INVx1_ASAP7_75t_SL g3756 ( 
.A(n_1674),
.Y(n_3756)
);

CKINVDCx5p33_ASAP7_75t_R g3757 ( 
.A(n_1752),
.Y(n_3757)
);

CKINVDCx5p33_ASAP7_75t_R g3758 ( 
.A(n_2780),
.Y(n_3758)
);

CKINVDCx5p33_ASAP7_75t_R g3759 ( 
.A(n_818),
.Y(n_3759)
);

INVx1_ASAP7_75t_L g3760 ( 
.A(n_2029),
.Y(n_3760)
);

CKINVDCx5p33_ASAP7_75t_R g3761 ( 
.A(n_2643),
.Y(n_3761)
);

INVx1_ASAP7_75t_L g3762 ( 
.A(n_2591),
.Y(n_3762)
);

INVx1_ASAP7_75t_L g3763 ( 
.A(n_660),
.Y(n_3763)
);

INVx1_ASAP7_75t_L g3764 ( 
.A(n_307),
.Y(n_3764)
);

INVx1_ASAP7_75t_L g3765 ( 
.A(n_374),
.Y(n_3765)
);

CKINVDCx5p33_ASAP7_75t_R g3766 ( 
.A(n_269),
.Y(n_3766)
);

CKINVDCx5p33_ASAP7_75t_R g3767 ( 
.A(n_2655),
.Y(n_3767)
);

CKINVDCx5p33_ASAP7_75t_R g3768 ( 
.A(n_1978),
.Y(n_3768)
);

INVx1_ASAP7_75t_L g3769 ( 
.A(n_196),
.Y(n_3769)
);

HB1xp67_ASAP7_75t_L g3770 ( 
.A(n_2772),
.Y(n_3770)
);

INVx1_ASAP7_75t_L g3771 ( 
.A(n_1576),
.Y(n_3771)
);

CKINVDCx5p33_ASAP7_75t_R g3772 ( 
.A(n_653),
.Y(n_3772)
);

INVx1_ASAP7_75t_L g3773 ( 
.A(n_1843),
.Y(n_3773)
);

INVx2_ASAP7_75t_L g3774 ( 
.A(n_2502),
.Y(n_3774)
);

CKINVDCx5p33_ASAP7_75t_R g3775 ( 
.A(n_1123),
.Y(n_3775)
);

INVx1_ASAP7_75t_SL g3776 ( 
.A(n_228),
.Y(n_3776)
);

CKINVDCx5p33_ASAP7_75t_R g3777 ( 
.A(n_1223),
.Y(n_3777)
);

CKINVDCx5p33_ASAP7_75t_R g3778 ( 
.A(n_2602),
.Y(n_3778)
);

CKINVDCx5p33_ASAP7_75t_R g3779 ( 
.A(n_749),
.Y(n_3779)
);

CKINVDCx5p33_ASAP7_75t_R g3780 ( 
.A(n_2465),
.Y(n_3780)
);

CKINVDCx5p33_ASAP7_75t_R g3781 ( 
.A(n_1076),
.Y(n_3781)
);

BUFx3_ASAP7_75t_L g3782 ( 
.A(n_2056),
.Y(n_3782)
);

CKINVDCx5p33_ASAP7_75t_R g3783 ( 
.A(n_1105),
.Y(n_3783)
);

CKINVDCx5p33_ASAP7_75t_R g3784 ( 
.A(n_971),
.Y(n_3784)
);

CKINVDCx20_ASAP7_75t_R g3785 ( 
.A(n_697),
.Y(n_3785)
);

CKINVDCx5p33_ASAP7_75t_R g3786 ( 
.A(n_1153),
.Y(n_3786)
);

CKINVDCx20_ASAP7_75t_R g3787 ( 
.A(n_2771),
.Y(n_3787)
);

CKINVDCx16_ASAP7_75t_R g3788 ( 
.A(n_2747),
.Y(n_3788)
);

CKINVDCx5p33_ASAP7_75t_R g3789 ( 
.A(n_1717),
.Y(n_3789)
);

INVx1_ASAP7_75t_L g3790 ( 
.A(n_2437),
.Y(n_3790)
);

CKINVDCx5p33_ASAP7_75t_R g3791 ( 
.A(n_2476),
.Y(n_3791)
);

CKINVDCx5p33_ASAP7_75t_R g3792 ( 
.A(n_2144),
.Y(n_3792)
);

INVx1_ASAP7_75t_L g3793 ( 
.A(n_2658),
.Y(n_3793)
);

CKINVDCx5p33_ASAP7_75t_R g3794 ( 
.A(n_675),
.Y(n_3794)
);

CKINVDCx5p33_ASAP7_75t_R g3795 ( 
.A(n_2735),
.Y(n_3795)
);

CKINVDCx5p33_ASAP7_75t_R g3796 ( 
.A(n_1138),
.Y(n_3796)
);

INVx1_ASAP7_75t_L g3797 ( 
.A(n_1285),
.Y(n_3797)
);

BUFx3_ASAP7_75t_L g3798 ( 
.A(n_1851),
.Y(n_3798)
);

INVx2_ASAP7_75t_L g3799 ( 
.A(n_2320),
.Y(n_3799)
);

CKINVDCx5p33_ASAP7_75t_R g3800 ( 
.A(n_1571),
.Y(n_3800)
);

CKINVDCx5p33_ASAP7_75t_R g3801 ( 
.A(n_2197),
.Y(n_3801)
);

INVx1_ASAP7_75t_L g3802 ( 
.A(n_869),
.Y(n_3802)
);

CKINVDCx5p33_ASAP7_75t_R g3803 ( 
.A(n_1185),
.Y(n_3803)
);

INVx1_ASAP7_75t_L g3804 ( 
.A(n_1),
.Y(n_3804)
);

INVx1_ASAP7_75t_SL g3805 ( 
.A(n_2450),
.Y(n_3805)
);

INVx1_ASAP7_75t_SL g3806 ( 
.A(n_408),
.Y(n_3806)
);

CKINVDCx5p33_ASAP7_75t_R g3807 ( 
.A(n_786),
.Y(n_3807)
);

CKINVDCx5p33_ASAP7_75t_R g3808 ( 
.A(n_238),
.Y(n_3808)
);

INVx1_ASAP7_75t_L g3809 ( 
.A(n_2478),
.Y(n_3809)
);

INVx1_ASAP7_75t_L g3810 ( 
.A(n_2763),
.Y(n_3810)
);

INVx1_ASAP7_75t_L g3811 ( 
.A(n_2462),
.Y(n_3811)
);

CKINVDCx5p33_ASAP7_75t_R g3812 ( 
.A(n_830),
.Y(n_3812)
);

CKINVDCx5p33_ASAP7_75t_R g3813 ( 
.A(n_1034),
.Y(n_3813)
);

INVx1_ASAP7_75t_L g3814 ( 
.A(n_178),
.Y(n_3814)
);

INVx1_ASAP7_75t_SL g3815 ( 
.A(n_1386),
.Y(n_3815)
);

CKINVDCx5p33_ASAP7_75t_R g3816 ( 
.A(n_2670),
.Y(n_3816)
);

INVx1_ASAP7_75t_L g3817 ( 
.A(n_661),
.Y(n_3817)
);

BUFx2_ASAP7_75t_L g3818 ( 
.A(n_1803),
.Y(n_3818)
);

INVx1_ASAP7_75t_L g3819 ( 
.A(n_1944),
.Y(n_3819)
);

CKINVDCx5p33_ASAP7_75t_R g3820 ( 
.A(n_580),
.Y(n_3820)
);

INVx1_ASAP7_75t_L g3821 ( 
.A(n_67),
.Y(n_3821)
);

INVx1_ASAP7_75t_L g3822 ( 
.A(n_58),
.Y(n_3822)
);

INVx1_ASAP7_75t_L g3823 ( 
.A(n_807),
.Y(n_3823)
);

BUFx3_ASAP7_75t_L g3824 ( 
.A(n_2412),
.Y(n_3824)
);

INVx1_ASAP7_75t_L g3825 ( 
.A(n_2666),
.Y(n_3825)
);

CKINVDCx20_ASAP7_75t_R g3826 ( 
.A(n_750),
.Y(n_3826)
);

CKINVDCx5p33_ASAP7_75t_R g3827 ( 
.A(n_2001),
.Y(n_3827)
);

INVx1_ASAP7_75t_L g3828 ( 
.A(n_505),
.Y(n_3828)
);

INVx1_ASAP7_75t_L g3829 ( 
.A(n_2650),
.Y(n_3829)
);

INVx1_ASAP7_75t_L g3830 ( 
.A(n_2568),
.Y(n_3830)
);

BUFx6f_ASAP7_75t_L g3831 ( 
.A(n_832),
.Y(n_3831)
);

INVx1_ASAP7_75t_L g3832 ( 
.A(n_1977),
.Y(n_3832)
);

INVx2_ASAP7_75t_L g3833 ( 
.A(n_1716),
.Y(n_3833)
);

INVx1_ASAP7_75t_SL g3834 ( 
.A(n_1881),
.Y(n_3834)
);

CKINVDCx5p33_ASAP7_75t_R g3835 ( 
.A(n_1168),
.Y(n_3835)
);

CKINVDCx20_ASAP7_75t_R g3836 ( 
.A(n_2034),
.Y(n_3836)
);

INVx1_ASAP7_75t_L g3837 ( 
.A(n_70),
.Y(n_3837)
);

CKINVDCx5p33_ASAP7_75t_R g3838 ( 
.A(n_2536),
.Y(n_3838)
);

INVx2_ASAP7_75t_SL g3839 ( 
.A(n_1455),
.Y(n_3839)
);

INVx1_ASAP7_75t_L g3840 ( 
.A(n_820),
.Y(n_3840)
);

CKINVDCx5p33_ASAP7_75t_R g3841 ( 
.A(n_2015),
.Y(n_3841)
);

INVx1_ASAP7_75t_L g3842 ( 
.A(n_914),
.Y(n_3842)
);

CKINVDCx5p33_ASAP7_75t_R g3843 ( 
.A(n_2462),
.Y(n_3843)
);

CKINVDCx5p33_ASAP7_75t_R g3844 ( 
.A(n_2606),
.Y(n_3844)
);

CKINVDCx5p33_ASAP7_75t_R g3845 ( 
.A(n_345),
.Y(n_3845)
);

CKINVDCx5p33_ASAP7_75t_R g3846 ( 
.A(n_2004),
.Y(n_3846)
);

CKINVDCx5p33_ASAP7_75t_R g3847 ( 
.A(n_768),
.Y(n_3847)
);

CKINVDCx5p33_ASAP7_75t_R g3848 ( 
.A(n_2599),
.Y(n_3848)
);

CKINVDCx5p33_ASAP7_75t_R g3849 ( 
.A(n_1159),
.Y(n_3849)
);

CKINVDCx5p33_ASAP7_75t_R g3850 ( 
.A(n_1931),
.Y(n_3850)
);

CKINVDCx20_ASAP7_75t_R g3851 ( 
.A(n_1333),
.Y(n_3851)
);

CKINVDCx5p33_ASAP7_75t_R g3852 ( 
.A(n_1467),
.Y(n_3852)
);

CKINVDCx5p33_ASAP7_75t_R g3853 ( 
.A(n_983),
.Y(n_3853)
);

INVx1_ASAP7_75t_L g3854 ( 
.A(n_2734),
.Y(n_3854)
);

CKINVDCx5p33_ASAP7_75t_R g3855 ( 
.A(n_2185),
.Y(n_3855)
);

INVx1_ASAP7_75t_L g3856 ( 
.A(n_1043),
.Y(n_3856)
);

CKINVDCx5p33_ASAP7_75t_R g3857 ( 
.A(n_61),
.Y(n_3857)
);

BUFx3_ASAP7_75t_L g3858 ( 
.A(n_1364),
.Y(n_3858)
);

CKINVDCx5p33_ASAP7_75t_R g3859 ( 
.A(n_2013),
.Y(n_3859)
);

CKINVDCx5p33_ASAP7_75t_R g3860 ( 
.A(n_1643),
.Y(n_3860)
);

CKINVDCx5p33_ASAP7_75t_R g3861 ( 
.A(n_1022),
.Y(n_3861)
);

CKINVDCx5p33_ASAP7_75t_R g3862 ( 
.A(n_1768),
.Y(n_3862)
);

CKINVDCx5p33_ASAP7_75t_R g3863 ( 
.A(n_2662),
.Y(n_3863)
);

CKINVDCx5p33_ASAP7_75t_R g3864 ( 
.A(n_415),
.Y(n_3864)
);

CKINVDCx5p33_ASAP7_75t_R g3865 ( 
.A(n_516),
.Y(n_3865)
);

HB1xp67_ASAP7_75t_L g3866 ( 
.A(n_424),
.Y(n_3866)
);

INVx1_ASAP7_75t_L g3867 ( 
.A(n_1473),
.Y(n_3867)
);

CKINVDCx5p33_ASAP7_75t_R g3868 ( 
.A(n_1477),
.Y(n_3868)
);

CKINVDCx5p33_ASAP7_75t_R g3869 ( 
.A(n_581),
.Y(n_3869)
);

BUFx5_ASAP7_75t_L g3870 ( 
.A(n_539),
.Y(n_3870)
);

CKINVDCx5p33_ASAP7_75t_R g3871 ( 
.A(n_596),
.Y(n_3871)
);

BUFx5_ASAP7_75t_L g3872 ( 
.A(n_2672),
.Y(n_3872)
);

BUFx2_ASAP7_75t_L g3873 ( 
.A(n_1025),
.Y(n_3873)
);

INVx1_ASAP7_75t_L g3874 ( 
.A(n_1187),
.Y(n_3874)
);

BUFx10_ASAP7_75t_L g3875 ( 
.A(n_268),
.Y(n_3875)
);

CKINVDCx16_ASAP7_75t_R g3876 ( 
.A(n_2314),
.Y(n_3876)
);

BUFx3_ASAP7_75t_L g3877 ( 
.A(n_1340),
.Y(n_3877)
);

CKINVDCx5p33_ASAP7_75t_R g3878 ( 
.A(n_115),
.Y(n_3878)
);

BUFx2_ASAP7_75t_L g3879 ( 
.A(n_1265),
.Y(n_3879)
);

CKINVDCx5p33_ASAP7_75t_R g3880 ( 
.A(n_1222),
.Y(n_3880)
);

CKINVDCx5p33_ASAP7_75t_R g3881 ( 
.A(n_82),
.Y(n_3881)
);

INVx1_ASAP7_75t_L g3882 ( 
.A(n_1552),
.Y(n_3882)
);

HB1xp67_ASAP7_75t_L g3883 ( 
.A(n_2384),
.Y(n_3883)
);

INVx1_ASAP7_75t_L g3884 ( 
.A(n_304),
.Y(n_3884)
);

CKINVDCx5p33_ASAP7_75t_R g3885 ( 
.A(n_533),
.Y(n_3885)
);

CKINVDCx5p33_ASAP7_75t_R g3886 ( 
.A(n_2524),
.Y(n_3886)
);

CKINVDCx5p33_ASAP7_75t_R g3887 ( 
.A(n_1115),
.Y(n_3887)
);

CKINVDCx5p33_ASAP7_75t_R g3888 ( 
.A(n_2619),
.Y(n_3888)
);

CKINVDCx5p33_ASAP7_75t_R g3889 ( 
.A(n_1109),
.Y(n_3889)
);

CKINVDCx5p33_ASAP7_75t_R g3890 ( 
.A(n_1468),
.Y(n_3890)
);

CKINVDCx5p33_ASAP7_75t_R g3891 ( 
.A(n_237),
.Y(n_3891)
);

INVx1_ASAP7_75t_L g3892 ( 
.A(n_2614),
.Y(n_3892)
);

INVx2_ASAP7_75t_L g3893 ( 
.A(n_466),
.Y(n_3893)
);

CKINVDCx5p33_ASAP7_75t_R g3894 ( 
.A(n_1831),
.Y(n_3894)
);

CKINVDCx5p33_ASAP7_75t_R g3895 ( 
.A(n_2572),
.Y(n_3895)
);

CKINVDCx5p33_ASAP7_75t_R g3896 ( 
.A(n_803),
.Y(n_3896)
);

CKINVDCx5p33_ASAP7_75t_R g3897 ( 
.A(n_2698),
.Y(n_3897)
);

CKINVDCx5p33_ASAP7_75t_R g3898 ( 
.A(n_1951),
.Y(n_3898)
);

INVx2_ASAP7_75t_SL g3899 ( 
.A(n_2723),
.Y(n_3899)
);

INVx1_ASAP7_75t_L g3900 ( 
.A(n_1194),
.Y(n_3900)
);

CKINVDCx5p33_ASAP7_75t_R g3901 ( 
.A(n_1158),
.Y(n_3901)
);

INVx2_ASAP7_75t_L g3902 ( 
.A(n_1839),
.Y(n_3902)
);

INVx1_ASAP7_75t_L g3903 ( 
.A(n_2760),
.Y(n_3903)
);

CKINVDCx5p33_ASAP7_75t_R g3904 ( 
.A(n_20),
.Y(n_3904)
);

CKINVDCx5p33_ASAP7_75t_R g3905 ( 
.A(n_305),
.Y(n_3905)
);

INVx1_ASAP7_75t_L g3906 ( 
.A(n_2085),
.Y(n_3906)
);

CKINVDCx5p33_ASAP7_75t_R g3907 ( 
.A(n_2096),
.Y(n_3907)
);

CKINVDCx5p33_ASAP7_75t_R g3908 ( 
.A(n_1436),
.Y(n_3908)
);

INVxp33_ASAP7_75t_R g3909 ( 
.A(n_1805),
.Y(n_3909)
);

BUFx6f_ASAP7_75t_L g3910 ( 
.A(n_1804),
.Y(n_3910)
);

CKINVDCx20_ASAP7_75t_R g3911 ( 
.A(n_2236),
.Y(n_3911)
);

CKINVDCx5p33_ASAP7_75t_R g3912 ( 
.A(n_4),
.Y(n_3912)
);

INVx1_ASAP7_75t_L g3913 ( 
.A(n_1711),
.Y(n_3913)
);

CKINVDCx5p33_ASAP7_75t_R g3914 ( 
.A(n_2778),
.Y(n_3914)
);

CKINVDCx5p33_ASAP7_75t_R g3915 ( 
.A(n_2676),
.Y(n_3915)
);

INVx2_ASAP7_75t_L g3916 ( 
.A(n_135),
.Y(n_3916)
);

CKINVDCx5p33_ASAP7_75t_R g3917 ( 
.A(n_2325),
.Y(n_3917)
);

CKINVDCx5p33_ASAP7_75t_R g3918 ( 
.A(n_288),
.Y(n_3918)
);

BUFx2_ASAP7_75t_L g3919 ( 
.A(n_2391),
.Y(n_3919)
);

CKINVDCx5p33_ASAP7_75t_R g3920 ( 
.A(n_34),
.Y(n_3920)
);

INVx2_ASAP7_75t_SL g3921 ( 
.A(n_1584),
.Y(n_3921)
);

CKINVDCx5p33_ASAP7_75t_R g3922 ( 
.A(n_1721),
.Y(n_3922)
);

INVx1_ASAP7_75t_L g3923 ( 
.A(n_1567),
.Y(n_3923)
);

INVx1_ASAP7_75t_L g3924 ( 
.A(n_1122),
.Y(n_3924)
);

BUFx2_ASAP7_75t_SL g3925 ( 
.A(n_767),
.Y(n_3925)
);

HB1xp67_ASAP7_75t_L g3926 ( 
.A(n_610),
.Y(n_3926)
);

INVx1_ASAP7_75t_L g3927 ( 
.A(n_1456),
.Y(n_3927)
);

CKINVDCx5p33_ASAP7_75t_R g3928 ( 
.A(n_1525),
.Y(n_3928)
);

BUFx5_ASAP7_75t_L g3929 ( 
.A(n_2417),
.Y(n_3929)
);

CKINVDCx5p33_ASAP7_75t_R g3930 ( 
.A(n_1225),
.Y(n_3930)
);

CKINVDCx5p33_ASAP7_75t_R g3931 ( 
.A(n_1058),
.Y(n_3931)
);

INVx1_ASAP7_75t_L g3932 ( 
.A(n_2362),
.Y(n_3932)
);

CKINVDCx5p33_ASAP7_75t_R g3933 ( 
.A(n_2569),
.Y(n_3933)
);

CKINVDCx20_ASAP7_75t_R g3934 ( 
.A(n_2433),
.Y(n_3934)
);

CKINVDCx5p33_ASAP7_75t_R g3935 ( 
.A(n_2718),
.Y(n_3935)
);

CKINVDCx5p33_ASAP7_75t_R g3936 ( 
.A(n_712),
.Y(n_3936)
);

CKINVDCx5p33_ASAP7_75t_R g3937 ( 
.A(n_1050),
.Y(n_3937)
);

CKINVDCx5p33_ASAP7_75t_R g3938 ( 
.A(n_2518),
.Y(n_3938)
);

BUFx10_ASAP7_75t_L g3939 ( 
.A(n_937),
.Y(n_3939)
);

CKINVDCx20_ASAP7_75t_R g3940 ( 
.A(n_211),
.Y(n_3940)
);

INVx2_ASAP7_75t_L g3941 ( 
.A(n_569),
.Y(n_3941)
);

CKINVDCx5p33_ASAP7_75t_R g3942 ( 
.A(n_349),
.Y(n_3942)
);

CKINVDCx14_ASAP7_75t_R g3943 ( 
.A(n_2108),
.Y(n_3943)
);

CKINVDCx5p33_ASAP7_75t_R g3944 ( 
.A(n_1857),
.Y(n_3944)
);

CKINVDCx5p33_ASAP7_75t_R g3945 ( 
.A(n_2110),
.Y(n_3945)
);

CKINVDCx5p33_ASAP7_75t_R g3946 ( 
.A(n_592),
.Y(n_3946)
);

INVx1_ASAP7_75t_L g3947 ( 
.A(n_463),
.Y(n_3947)
);

CKINVDCx20_ASAP7_75t_R g3948 ( 
.A(n_2261),
.Y(n_3948)
);

INVx1_ASAP7_75t_SL g3949 ( 
.A(n_749),
.Y(n_3949)
);

INVx1_ASAP7_75t_L g3950 ( 
.A(n_1296),
.Y(n_3950)
);

INVx2_ASAP7_75t_L g3951 ( 
.A(n_1451),
.Y(n_3951)
);

BUFx6f_ASAP7_75t_L g3952 ( 
.A(n_2583),
.Y(n_3952)
);

INVx1_ASAP7_75t_L g3953 ( 
.A(n_345),
.Y(n_3953)
);

CKINVDCx5p33_ASAP7_75t_R g3954 ( 
.A(n_2581),
.Y(n_3954)
);

CKINVDCx5p33_ASAP7_75t_R g3955 ( 
.A(n_2033),
.Y(n_3955)
);

CKINVDCx5p33_ASAP7_75t_R g3956 ( 
.A(n_2709),
.Y(n_3956)
);

INVx1_ASAP7_75t_L g3957 ( 
.A(n_947),
.Y(n_3957)
);

CKINVDCx5p33_ASAP7_75t_R g3958 ( 
.A(n_2158),
.Y(n_3958)
);

CKINVDCx5p33_ASAP7_75t_R g3959 ( 
.A(n_2334),
.Y(n_3959)
);

INVx1_ASAP7_75t_L g3960 ( 
.A(n_2627),
.Y(n_3960)
);

CKINVDCx5p33_ASAP7_75t_R g3961 ( 
.A(n_1753),
.Y(n_3961)
);

CKINVDCx5p33_ASAP7_75t_R g3962 ( 
.A(n_677),
.Y(n_3962)
);

INVx1_ASAP7_75t_L g3963 ( 
.A(n_653),
.Y(n_3963)
);

CKINVDCx5p33_ASAP7_75t_R g3964 ( 
.A(n_2365),
.Y(n_3964)
);

INVx1_ASAP7_75t_SL g3965 ( 
.A(n_2540),
.Y(n_3965)
);

INVx1_ASAP7_75t_L g3966 ( 
.A(n_514),
.Y(n_3966)
);

CKINVDCx5p33_ASAP7_75t_R g3967 ( 
.A(n_1425),
.Y(n_3967)
);

CKINVDCx5p33_ASAP7_75t_R g3968 ( 
.A(n_1800),
.Y(n_3968)
);

INVx1_ASAP7_75t_L g3969 ( 
.A(n_156),
.Y(n_3969)
);

INVx1_ASAP7_75t_L g3970 ( 
.A(n_1930),
.Y(n_3970)
);

CKINVDCx5p33_ASAP7_75t_R g3971 ( 
.A(n_372),
.Y(n_3971)
);

INVx1_ASAP7_75t_SL g3972 ( 
.A(n_2517),
.Y(n_3972)
);

CKINVDCx5p33_ASAP7_75t_R g3973 ( 
.A(n_1645),
.Y(n_3973)
);

INVx1_ASAP7_75t_L g3974 ( 
.A(n_2595),
.Y(n_3974)
);

INVx1_ASAP7_75t_L g3975 ( 
.A(n_2202),
.Y(n_3975)
);

INVx1_ASAP7_75t_L g3976 ( 
.A(n_1273),
.Y(n_3976)
);

INVx2_ASAP7_75t_SL g3977 ( 
.A(n_2751),
.Y(n_3977)
);

INVx2_ASAP7_75t_L g3978 ( 
.A(n_2576),
.Y(n_3978)
);

CKINVDCx5p33_ASAP7_75t_R g3979 ( 
.A(n_206),
.Y(n_3979)
);

CKINVDCx20_ASAP7_75t_R g3980 ( 
.A(n_91),
.Y(n_3980)
);

INVx1_ASAP7_75t_L g3981 ( 
.A(n_39),
.Y(n_3981)
);

CKINVDCx5p33_ASAP7_75t_R g3982 ( 
.A(n_1578),
.Y(n_3982)
);

CKINVDCx5p33_ASAP7_75t_R g3983 ( 
.A(n_2634),
.Y(n_3983)
);

CKINVDCx5p33_ASAP7_75t_R g3984 ( 
.A(n_2164),
.Y(n_3984)
);

CKINVDCx5p33_ASAP7_75t_R g3985 ( 
.A(n_638),
.Y(n_3985)
);

HB1xp67_ASAP7_75t_L g3986 ( 
.A(n_636),
.Y(n_3986)
);

CKINVDCx5p33_ASAP7_75t_R g3987 ( 
.A(n_1544),
.Y(n_3987)
);

INVx1_ASAP7_75t_L g3988 ( 
.A(n_1488),
.Y(n_3988)
);

INVx2_ASAP7_75t_L g3989 ( 
.A(n_2712),
.Y(n_3989)
);

BUFx6f_ASAP7_75t_L g3990 ( 
.A(n_2307),
.Y(n_3990)
);

CKINVDCx5p33_ASAP7_75t_R g3991 ( 
.A(n_2496),
.Y(n_3991)
);

CKINVDCx5p33_ASAP7_75t_R g3992 ( 
.A(n_2781),
.Y(n_3992)
);

BUFx2_ASAP7_75t_L g3993 ( 
.A(n_1857),
.Y(n_3993)
);

CKINVDCx5p33_ASAP7_75t_R g3994 ( 
.A(n_2705),
.Y(n_3994)
);

BUFx10_ASAP7_75t_L g3995 ( 
.A(n_1293),
.Y(n_3995)
);

CKINVDCx5p33_ASAP7_75t_R g3996 ( 
.A(n_2664),
.Y(n_3996)
);

BUFx8_ASAP7_75t_SL g3997 ( 
.A(n_1969),
.Y(n_3997)
);

CKINVDCx5p33_ASAP7_75t_R g3998 ( 
.A(n_1365),
.Y(n_3998)
);

CKINVDCx5p33_ASAP7_75t_R g3999 ( 
.A(n_68),
.Y(n_3999)
);

INVx1_ASAP7_75t_L g4000 ( 
.A(n_2702),
.Y(n_4000)
);

INVx1_ASAP7_75t_L g4001 ( 
.A(n_1772),
.Y(n_4001)
);

CKINVDCx5p33_ASAP7_75t_R g4002 ( 
.A(n_2727),
.Y(n_4002)
);

INVx1_ASAP7_75t_L g4003 ( 
.A(n_677),
.Y(n_4003)
);

BUFx5_ASAP7_75t_L g4004 ( 
.A(n_2273),
.Y(n_4004)
);

BUFx3_ASAP7_75t_L g4005 ( 
.A(n_1425),
.Y(n_4005)
);

CKINVDCx5p33_ASAP7_75t_R g4006 ( 
.A(n_1861),
.Y(n_4006)
);

INVx1_ASAP7_75t_L g4007 ( 
.A(n_1470),
.Y(n_4007)
);

CKINVDCx5p33_ASAP7_75t_R g4008 ( 
.A(n_2554),
.Y(n_4008)
);

INVx1_ASAP7_75t_L g4009 ( 
.A(n_2499),
.Y(n_4009)
);

CKINVDCx5p33_ASAP7_75t_R g4010 ( 
.A(n_324),
.Y(n_4010)
);

CKINVDCx16_ASAP7_75t_R g4011 ( 
.A(n_1688),
.Y(n_4011)
);

HB1xp67_ASAP7_75t_L g4012 ( 
.A(n_994),
.Y(n_4012)
);

CKINVDCx5p33_ASAP7_75t_R g4013 ( 
.A(n_1628),
.Y(n_4013)
);

CKINVDCx5p33_ASAP7_75t_R g4014 ( 
.A(n_2563),
.Y(n_4014)
);

CKINVDCx5p33_ASAP7_75t_R g4015 ( 
.A(n_1864),
.Y(n_4015)
);

INVx1_ASAP7_75t_L g4016 ( 
.A(n_171),
.Y(n_4016)
);

CKINVDCx5p33_ASAP7_75t_R g4017 ( 
.A(n_2545),
.Y(n_4017)
);

INVx2_ASAP7_75t_L g4018 ( 
.A(n_271),
.Y(n_4018)
);

CKINVDCx20_ASAP7_75t_R g4019 ( 
.A(n_1310),
.Y(n_4019)
);

BUFx3_ASAP7_75t_L g4020 ( 
.A(n_1529),
.Y(n_4020)
);

INVx1_ASAP7_75t_L g4021 ( 
.A(n_579),
.Y(n_4021)
);

CKINVDCx5p33_ASAP7_75t_R g4022 ( 
.A(n_58),
.Y(n_4022)
);

INVx1_ASAP7_75t_L g4023 ( 
.A(n_2573),
.Y(n_4023)
);

INVx1_ASAP7_75t_L g4024 ( 
.A(n_2326),
.Y(n_4024)
);

INVx2_ASAP7_75t_L g4025 ( 
.A(n_1305),
.Y(n_4025)
);

INVx1_ASAP7_75t_L g4026 ( 
.A(n_2495),
.Y(n_4026)
);

CKINVDCx5p33_ASAP7_75t_R g4027 ( 
.A(n_2763),
.Y(n_4027)
);

CKINVDCx5p33_ASAP7_75t_R g4028 ( 
.A(n_2688),
.Y(n_4028)
);

CKINVDCx5p33_ASAP7_75t_R g4029 ( 
.A(n_2697),
.Y(n_4029)
);

BUFx6f_ASAP7_75t_L g4030 ( 
.A(n_2008),
.Y(n_4030)
);

CKINVDCx5p33_ASAP7_75t_R g4031 ( 
.A(n_2458),
.Y(n_4031)
);

CKINVDCx20_ASAP7_75t_R g4032 ( 
.A(n_2680),
.Y(n_4032)
);

CKINVDCx20_ASAP7_75t_R g4033 ( 
.A(n_2483),
.Y(n_4033)
);

CKINVDCx5p33_ASAP7_75t_R g4034 ( 
.A(n_399),
.Y(n_4034)
);

CKINVDCx20_ASAP7_75t_R g4035 ( 
.A(n_1967),
.Y(n_4035)
);

CKINVDCx5p33_ASAP7_75t_R g4036 ( 
.A(n_2718),
.Y(n_4036)
);

CKINVDCx5p33_ASAP7_75t_R g4037 ( 
.A(n_2638),
.Y(n_4037)
);

CKINVDCx16_ASAP7_75t_R g4038 ( 
.A(n_2290),
.Y(n_4038)
);

INVx1_ASAP7_75t_SL g4039 ( 
.A(n_1967),
.Y(n_4039)
);

CKINVDCx20_ASAP7_75t_R g4040 ( 
.A(n_1119),
.Y(n_4040)
);

INVx1_ASAP7_75t_L g4041 ( 
.A(n_2668),
.Y(n_4041)
);

INVx1_ASAP7_75t_L g4042 ( 
.A(n_1627),
.Y(n_4042)
);

CKINVDCx5p33_ASAP7_75t_R g4043 ( 
.A(n_901),
.Y(n_4043)
);

CKINVDCx20_ASAP7_75t_R g4044 ( 
.A(n_205),
.Y(n_4044)
);

CKINVDCx5p33_ASAP7_75t_R g4045 ( 
.A(n_1560),
.Y(n_4045)
);

BUFx2_ASAP7_75t_L g4046 ( 
.A(n_1638),
.Y(n_4046)
);

INVx1_ASAP7_75t_L g4047 ( 
.A(n_214),
.Y(n_4047)
);

CKINVDCx5p33_ASAP7_75t_R g4048 ( 
.A(n_311),
.Y(n_4048)
);

CKINVDCx5p33_ASAP7_75t_R g4049 ( 
.A(n_565),
.Y(n_4049)
);

CKINVDCx5p33_ASAP7_75t_R g4050 ( 
.A(n_270),
.Y(n_4050)
);

BUFx3_ASAP7_75t_L g4051 ( 
.A(n_2033),
.Y(n_4051)
);

CKINVDCx20_ASAP7_75t_R g4052 ( 
.A(n_2588),
.Y(n_4052)
);

BUFx10_ASAP7_75t_L g4053 ( 
.A(n_1269),
.Y(n_4053)
);

CKINVDCx5p33_ASAP7_75t_R g4054 ( 
.A(n_2640),
.Y(n_4054)
);

INVx1_ASAP7_75t_L g4055 ( 
.A(n_991),
.Y(n_4055)
);

CKINVDCx14_ASAP7_75t_R g4056 ( 
.A(n_2646),
.Y(n_4056)
);

CKINVDCx5p33_ASAP7_75t_R g4057 ( 
.A(n_787),
.Y(n_4057)
);

CKINVDCx5p33_ASAP7_75t_R g4058 ( 
.A(n_2679),
.Y(n_4058)
);

INVx2_ASAP7_75t_L g4059 ( 
.A(n_2579),
.Y(n_4059)
);

CKINVDCx5p33_ASAP7_75t_R g4060 ( 
.A(n_2169),
.Y(n_4060)
);

CKINVDCx16_ASAP7_75t_R g4061 ( 
.A(n_1129),
.Y(n_4061)
);

CKINVDCx20_ASAP7_75t_R g4062 ( 
.A(n_151),
.Y(n_4062)
);

CKINVDCx20_ASAP7_75t_R g4063 ( 
.A(n_882),
.Y(n_4063)
);

INVx2_ASAP7_75t_SL g4064 ( 
.A(n_1803),
.Y(n_4064)
);

INVx2_ASAP7_75t_L g4065 ( 
.A(n_1896),
.Y(n_4065)
);

CKINVDCx5p33_ASAP7_75t_R g4066 ( 
.A(n_142),
.Y(n_4066)
);

CKINVDCx5p33_ASAP7_75t_R g4067 ( 
.A(n_1189),
.Y(n_4067)
);

CKINVDCx5p33_ASAP7_75t_R g4068 ( 
.A(n_1832),
.Y(n_4068)
);

INVx1_ASAP7_75t_L g4069 ( 
.A(n_1114),
.Y(n_4069)
);

CKINVDCx11_ASAP7_75t_R g4070 ( 
.A(n_921),
.Y(n_4070)
);

CKINVDCx5p33_ASAP7_75t_R g4071 ( 
.A(n_2704),
.Y(n_4071)
);

CKINVDCx5p33_ASAP7_75t_R g4072 ( 
.A(n_1578),
.Y(n_4072)
);

CKINVDCx5p33_ASAP7_75t_R g4073 ( 
.A(n_2685),
.Y(n_4073)
);

CKINVDCx5p33_ASAP7_75t_R g4074 ( 
.A(n_2795),
.Y(n_4074)
);

CKINVDCx5p33_ASAP7_75t_R g4075 ( 
.A(n_1685),
.Y(n_4075)
);

BUFx5_ASAP7_75t_L g4076 ( 
.A(n_2143),
.Y(n_4076)
);

INVx1_ASAP7_75t_SL g4077 ( 
.A(n_2696),
.Y(n_4077)
);

CKINVDCx5p33_ASAP7_75t_R g4078 ( 
.A(n_1784),
.Y(n_4078)
);

BUFx3_ASAP7_75t_L g4079 ( 
.A(n_1861),
.Y(n_4079)
);

BUFx10_ASAP7_75t_L g4080 ( 
.A(n_1539),
.Y(n_4080)
);

CKINVDCx5p33_ASAP7_75t_R g4081 ( 
.A(n_1054),
.Y(n_4081)
);

INVx1_ASAP7_75t_L g4082 ( 
.A(n_2693),
.Y(n_4082)
);

CKINVDCx5p33_ASAP7_75t_R g4083 ( 
.A(n_2779),
.Y(n_4083)
);

CKINVDCx5p33_ASAP7_75t_R g4084 ( 
.A(n_2620),
.Y(n_4084)
);

CKINVDCx20_ASAP7_75t_R g4085 ( 
.A(n_591),
.Y(n_4085)
);

CKINVDCx16_ASAP7_75t_R g4086 ( 
.A(n_135),
.Y(n_4086)
);

INVx2_ASAP7_75t_L g4087 ( 
.A(n_12),
.Y(n_4087)
);

CKINVDCx16_ASAP7_75t_R g4088 ( 
.A(n_674),
.Y(n_4088)
);

CKINVDCx5p33_ASAP7_75t_R g4089 ( 
.A(n_474),
.Y(n_4089)
);

CKINVDCx5p33_ASAP7_75t_R g4090 ( 
.A(n_2682),
.Y(n_4090)
);

CKINVDCx5p33_ASAP7_75t_R g4091 ( 
.A(n_2114),
.Y(n_4091)
);

INVx1_ASAP7_75t_SL g4092 ( 
.A(n_980),
.Y(n_4092)
);

INVx2_ASAP7_75t_L g4093 ( 
.A(n_1957),
.Y(n_4093)
);

BUFx5_ASAP7_75t_L g4094 ( 
.A(n_2254),
.Y(n_4094)
);

CKINVDCx5p33_ASAP7_75t_R g4095 ( 
.A(n_1322),
.Y(n_4095)
);

CKINVDCx5p33_ASAP7_75t_R g4096 ( 
.A(n_1832),
.Y(n_4096)
);

CKINVDCx5p33_ASAP7_75t_R g4097 ( 
.A(n_2621),
.Y(n_4097)
);

INVx1_ASAP7_75t_L g4098 ( 
.A(n_806),
.Y(n_4098)
);

CKINVDCx5p33_ASAP7_75t_R g4099 ( 
.A(n_1250),
.Y(n_4099)
);

CKINVDCx5p33_ASAP7_75t_R g4100 ( 
.A(n_1760),
.Y(n_4100)
);

CKINVDCx5p33_ASAP7_75t_R g4101 ( 
.A(n_1430),
.Y(n_4101)
);

CKINVDCx5p33_ASAP7_75t_R g4102 ( 
.A(n_2448),
.Y(n_4102)
);

CKINVDCx5p33_ASAP7_75t_R g4103 ( 
.A(n_2597),
.Y(n_4103)
);

INVx1_ASAP7_75t_L g4104 ( 
.A(n_453),
.Y(n_4104)
);

INVx1_ASAP7_75t_L g4105 ( 
.A(n_852),
.Y(n_4105)
);

INVx2_ASAP7_75t_L g4106 ( 
.A(n_434),
.Y(n_4106)
);

CKINVDCx5p33_ASAP7_75t_R g4107 ( 
.A(n_2173),
.Y(n_4107)
);

CKINVDCx5p33_ASAP7_75t_R g4108 ( 
.A(n_2749),
.Y(n_4108)
);

INVx1_ASAP7_75t_L g4109 ( 
.A(n_2604),
.Y(n_4109)
);

CKINVDCx5p33_ASAP7_75t_R g4110 ( 
.A(n_2600),
.Y(n_4110)
);

CKINVDCx20_ASAP7_75t_R g4111 ( 
.A(n_389),
.Y(n_4111)
);

INVx2_ASAP7_75t_L g4112 ( 
.A(n_1894),
.Y(n_4112)
);

CKINVDCx5p33_ASAP7_75t_R g4113 ( 
.A(n_938),
.Y(n_4113)
);

CKINVDCx20_ASAP7_75t_R g4114 ( 
.A(n_1062),
.Y(n_4114)
);

CKINVDCx5p33_ASAP7_75t_R g4115 ( 
.A(n_214),
.Y(n_4115)
);

INVx1_ASAP7_75t_L g4116 ( 
.A(n_1528),
.Y(n_4116)
);

CKINVDCx5p33_ASAP7_75t_R g4117 ( 
.A(n_876),
.Y(n_4117)
);

CKINVDCx5p33_ASAP7_75t_R g4118 ( 
.A(n_2587),
.Y(n_4118)
);

CKINVDCx5p33_ASAP7_75t_R g4119 ( 
.A(n_1349),
.Y(n_4119)
);

INVx2_ASAP7_75t_L g4120 ( 
.A(n_113),
.Y(n_4120)
);

CKINVDCx20_ASAP7_75t_R g4121 ( 
.A(n_2026),
.Y(n_4121)
);

CKINVDCx5p33_ASAP7_75t_R g4122 ( 
.A(n_2637),
.Y(n_4122)
);

CKINVDCx16_ASAP7_75t_R g4123 ( 
.A(n_2590),
.Y(n_4123)
);

CKINVDCx5p33_ASAP7_75t_R g4124 ( 
.A(n_641),
.Y(n_4124)
);

INVx1_ASAP7_75t_L g4125 ( 
.A(n_2291),
.Y(n_4125)
);

CKINVDCx5p33_ASAP7_75t_R g4126 ( 
.A(n_699),
.Y(n_4126)
);

CKINVDCx16_ASAP7_75t_R g4127 ( 
.A(n_2509),
.Y(n_4127)
);

CKINVDCx5p33_ASAP7_75t_R g4128 ( 
.A(n_2492),
.Y(n_4128)
);

CKINVDCx5p33_ASAP7_75t_R g4129 ( 
.A(n_1863),
.Y(n_4129)
);

CKINVDCx5p33_ASAP7_75t_R g4130 ( 
.A(n_2114),
.Y(n_4130)
);

INVx1_ASAP7_75t_L g4131 ( 
.A(n_1302),
.Y(n_4131)
);

CKINVDCx5p33_ASAP7_75t_R g4132 ( 
.A(n_1841),
.Y(n_4132)
);

INVx1_ASAP7_75t_SL g4133 ( 
.A(n_887),
.Y(n_4133)
);

CKINVDCx5p33_ASAP7_75t_R g4134 ( 
.A(n_108),
.Y(n_4134)
);

CKINVDCx5p33_ASAP7_75t_R g4135 ( 
.A(n_2432),
.Y(n_4135)
);

CKINVDCx20_ASAP7_75t_R g4136 ( 
.A(n_1842),
.Y(n_4136)
);

CKINVDCx5p33_ASAP7_75t_R g4137 ( 
.A(n_1107),
.Y(n_4137)
);

INVx2_ASAP7_75t_SL g4138 ( 
.A(n_1851),
.Y(n_4138)
);

INVx1_ASAP7_75t_L g4139 ( 
.A(n_2242),
.Y(n_4139)
);

CKINVDCx5p33_ASAP7_75t_R g4140 ( 
.A(n_2435),
.Y(n_4140)
);

INVx1_ASAP7_75t_L g4141 ( 
.A(n_988),
.Y(n_4141)
);

CKINVDCx5p33_ASAP7_75t_R g4142 ( 
.A(n_2804),
.Y(n_4142)
);

CKINVDCx5p33_ASAP7_75t_R g4143 ( 
.A(n_1703),
.Y(n_4143)
);

CKINVDCx5p33_ASAP7_75t_R g4144 ( 
.A(n_2647),
.Y(n_4144)
);

CKINVDCx5p33_ASAP7_75t_R g4145 ( 
.A(n_307),
.Y(n_4145)
);

INVx1_ASAP7_75t_L g4146 ( 
.A(n_824),
.Y(n_4146)
);

CKINVDCx5p33_ASAP7_75t_R g4147 ( 
.A(n_2087),
.Y(n_4147)
);

INVx1_ASAP7_75t_L g4148 ( 
.A(n_1587),
.Y(n_4148)
);

INVx1_ASAP7_75t_SL g4149 ( 
.A(n_135),
.Y(n_4149)
);

CKINVDCx5p33_ASAP7_75t_R g4150 ( 
.A(n_1281),
.Y(n_4150)
);

INVx1_ASAP7_75t_L g4151 ( 
.A(n_706),
.Y(n_4151)
);

INVx1_ASAP7_75t_L g4152 ( 
.A(n_2353),
.Y(n_4152)
);

CKINVDCx5p33_ASAP7_75t_R g4153 ( 
.A(n_2691),
.Y(n_4153)
);

INVx1_ASAP7_75t_L g4154 ( 
.A(n_1164),
.Y(n_4154)
);

BUFx3_ASAP7_75t_L g4155 ( 
.A(n_1926),
.Y(n_4155)
);

CKINVDCx5p33_ASAP7_75t_R g4156 ( 
.A(n_2340),
.Y(n_4156)
);

CKINVDCx5p33_ASAP7_75t_R g4157 ( 
.A(n_1421),
.Y(n_4157)
);

INVx1_ASAP7_75t_L g4158 ( 
.A(n_2674),
.Y(n_4158)
);

CKINVDCx5p33_ASAP7_75t_R g4159 ( 
.A(n_2589),
.Y(n_4159)
);

CKINVDCx5p33_ASAP7_75t_R g4160 ( 
.A(n_1012),
.Y(n_4160)
);

BUFx8_ASAP7_75t_SL g4161 ( 
.A(n_977),
.Y(n_4161)
);

INVx1_ASAP7_75t_L g4162 ( 
.A(n_2740),
.Y(n_4162)
);

INVx1_ASAP7_75t_L g4163 ( 
.A(n_2382),
.Y(n_4163)
);

INVx1_ASAP7_75t_L g4164 ( 
.A(n_2398),
.Y(n_4164)
);

CKINVDCx5p33_ASAP7_75t_R g4165 ( 
.A(n_878),
.Y(n_4165)
);

INVx1_ASAP7_75t_L g4166 ( 
.A(n_2630),
.Y(n_4166)
);

INVx1_ASAP7_75t_L g4167 ( 
.A(n_2423),
.Y(n_4167)
);

BUFx3_ASAP7_75t_L g4168 ( 
.A(n_69),
.Y(n_4168)
);

CKINVDCx5p33_ASAP7_75t_R g4169 ( 
.A(n_2017),
.Y(n_4169)
);

CKINVDCx5p33_ASAP7_75t_R g4170 ( 
.A(n_1775),
.Y(n_4170)
);

CKINVDCx5p33_ASAP7_75t_R g4171 ( 
.A(n_313),
.Y(n_4171)
);

INVx1_ASAP7_75t_L g4172 ( 
.A(n_1333),
.Y(n_4172)
);

CKINVDCx5p33_ASAP7_75t_R g4173 ( 
.A(n_2360),
.Y(n_4173)
);

INVx1_ASAP7_75t_L g4174 ( 
.A(n_893),
.Y(n_4174)
);

CKINVDCx5p33_ASAP7_75t_R g4175 ( 
.A(n_2066),
.Y(n_4175)
);

CKINVDCx5p33_ASAP7_75t_R g4176 ( 
.A(n_2581),
.Y(n_4176)
);

CKINVDCx5p33_ASAP7_75t_R g4177 ( 
.A(n_719),
.Y(n_4177)
);

INVx1_ASAP7_75t_L g4178 ( 
.A(n_144),
.Y(n_4178)
);

INVx1_ASAP7_75t_L g4179 ( 
.A(n_2334),
.Y(n_4179)
);

BUFx10_ASAP7_75t_L g4180 ( 
.A(n_2359),
.Y(n_4180)
);

CKINVDCx5p33_ASAP7_75t_R g4181 ( 
.A(n_974),
.Y(n_4181)
);

CKINVDCx5p33_ASAP7_75t_R g4182 ( 
.A(n_2268),
.Y(n_4182)
);

INVx2_ASAP7_75t_L g4183 ( 
.A(n_1654),
.Y(n_4183)
);

CKINVDCx5p33_ASAP7_75t_R g4184 ( 
.A(n_1348),
.Y(n_4184)
);

CKINVDCx16_ASAP7_75t_R g4185 ( 
.A(n_2761),
.Y(n_4185)
);

CKINVDCx5p33_ASAP7_75t_R g4186 ( 
.A(n_1854),
.Y(n_4186)
);

CKINVDCx5p33_ASAP7_75t_R g4187 ( 
.A(n_150),
.Y(n_4187)
);

INVx2_ASAP7_75t_L g4188 ( 
.A(n_1306),
.Y(n_4188)
);

CKINVDCx5p33_ASAP7_75t_R g4189 ( 
.A(n_2683),
.Y(n_4189)
);

INVx1_ASAP7_75t_L g4190 ( 
.A(n_551),
.Y(n_4190)
);

INVx2_ASAP7_75t_L g4191 ( 
.A(n_1815),
.Y(n_4191)
);

CKINVDCx16_ASAP7_75t_R g4192 ( 
.A(n_2745),
.Y(n_4192)
);

CKINVDCx5p33_ASAP7_75t_R g4193 ( 
.A(n_529),
.Y(n_4193)
);

CKINVDCx5p33_ASAP7_75t_R g4194 ( 
.A(n_1085),
.Y(n_4194)
);

BUFx6f_ASAP7_75t_L g4195 ( 
.A(n_119),
.Y(n_4195)
);

INVx1_ASAP7_75t_L g4196 ( 
.A(n_2151),
.Y(n_4196)
);

CKINVDCx20_ASAP7_75t_R g4197 ( 
.A(n_2004),
.Y(n_4197)
);

INVx1_ASAP7_75t_L g4198 ( 
.A(n_3658),
.Y(n_4198)
);

CKINVDCx5p33_ASAP7_75t_R g4199 ( 
.A(n_4070),
.Y(n_4199)
);

INVx1_ASAP7_75t_L g4200 ( 
.A(n_3658),
.Y(n_4200)
);

BUFx5_ASAP7_75t_L g4201 ( 
.A(n_2822),
.Y(n_4201)
);

CKINVDCx5p33_ASAP7_75t_R g4202 ( 
.A(n_3415),
.Y(n_4202)
);

INVxp33_ASAP7_75t_SL g4203 ( 
.A(n_3866),
.Y(n_4203)
);

INVx1_ASAP7_75t_L g4204 ( 
.A(n_3658),
.Y(n_4204)
);

INVx1_ASAP7_75t_L g4205 ( 
.A(n_3658),
.Y(n_4205)
);

INVx1_ASAP7_75t_L g4206 ( 
.A(n_3658),
.Y(n_4206)
);

CKINVDCx5p33_ASAP7_75t_R g4207 ( 
.A(n_3997),
.Y(n_4207)
);

NOR2xp67_ASAP7_75t_L g4208 ( 
.A(n_2854),
.B(n_0),
.Y(n_4208)
);

CKINVDCx5p33_ASAP7_75t_R g4209 ( 
.A(n_4161),
.Y(n_4209)
);

INVx1_ASAP7_75t_L g4210 ( 
.A(n_3870),
.Y(n_4210)
);

INVx1_ASAP7_75t_L g4211 ( 
.A(n_3870),
.Y(n_4211)
);

INVx1_ASAP7_75t_L g4212 ( 
.A(n_3870),
.Y(n_4212)
);

INVxp67_ASAP7_75t_L g4213 ( 
.A(n_3273),
.Y(n_4213)
);

NOR2xp33_ASAP7_75t_L g4214 ( 
.A(n_3707),
.B(n_0),
.Y(n_4214)
);

INVx1_ASAP7_75t_L g4215 ( 
.A(n_3870),
.Y(n_4215)
);

INVx1_ASAP7_75t_L g4216 ( 
.A(n_3870),
.Y(n_4216)
);

BUFx3_ASAP7_75t_L g4217 ( 
.A(n_3057),
.Y(n_4217)
);

INVx1_ASAP7_75t_L g4218 ( 
.A(n_2843),
.Y(n_4218)
);

INVx1_ASAP7_75t_L g4219 ( 
.A(n_2843),
.Y(n_4219)
);

CKINVDCx5p33_ASAP7_75t_R g4220 ( 
.A(n_3002),
.Y(n_4220)
);

CKINVDCx16_ASAP7_75t_R g4221 ( 
.A(n_3116),
.Y(n_4221)
);

CKINVDCx5p33_ASAP7_75t_R g4222 ( 
.A(n_3351),
.Y(n_4222)
);

NAND2xp5_ASAP7_75t_L g4223 ( 
.A(n_3017),
.B(n_0),
.Y(n_4223)
);

INVx1_ASAP7_75t_L g4224 ( 
.A(n_2843),
.Y(n_4224)
);

INVx1_ASAP7_75t_L g4225 ( 
.A(n_2843),
.Y(n_4225)
);

INVxp67_ASAP7_75t_SL g4226 ( 
.A(n_3078),
.Y(n_4226)
);

INVx1_ASAP7_75t_L g4227 ( 
.A(n_2843),
.Y(n_4227)
);

INVx1_ASAP7_75t_L g4228 ( 
.A(n_2899),
.Y(n_4228)
);

INVx1_ASAP7_75t_SL g4229 ( 
.A(n_2814),
.Y(n_4229)
);

INVxp67_ASAP7_75t_L g4230 ( 
.A(n_2984),
.Y(n_4230)
);

INVx1_ASAP7_75t_L g4231 ( 
.A(n_2899),
.Y(n_4231)
);

INVx1_ASAP7_75t_L g4232 ( 
.A(n_2899),
.Y(n_4232)
);

INVx1_ASAP7_75t_L g4233 ( 
.A(n_2899),
.Y(n_4233)
);

CKINVDCx5p33_ASAP7_75t_R g4234 ( 
.A(n_3467),
.Y(n_4234)
);

CKINVDCx5p33_ASAP7_75t_R g4235 ( 
.A(n_3706),
.Y(n_4235)
);

INVx1_ASAP7_75t_L g4236 ( 
.A(n_2899),
.Y(n_4236)
);

INVx1_ASAP7_75t_L g4237 ( 
.A(n_3060),
.Y(n_4237)
);

INVx1_ASAP7_75t_L g4238 ( 
.A(n_3060),
.Y(n_4238)
);

INVx1_ASAP7_75t_L g4239 ( 
.A(n_3060),
.Y(n_4239)
);

CKINVDCx16_ASAP7_75t_R g4240 ( 
.A(n_4086),
.Y(n_4240)
);

INVx1_ASAP7_75t_L g4241 ( 
.A(n_3060),
.Y(n_4241)
);

CKINVDCx5p33_ASAP7_75t_R g4242 ( 
.A(n_3043),
.Y(n_4242)
);

INVx1_ASAP7_75t_L g4243 ( 
.A(n_3060),
.Y(n_4243)
);

CKINVDCx5p33_ASAP7_75t_R g4244 ( 
.A(n_3235),
.Y(n_4244)
);

INVx1_ASAP7_75t_L g4245 ( 
.A(n_3118),
.Y(n_4245)
);

CKINVDCx5p33_ASAP7_75t_R g4246 ( 
.A(n_3349),
.Y(n_4246)
);

CKINVDCx16_ASAP7_75t_R g4247 ( 
.A(n_2875),
.Y(n_4247)
);

CKINVDCx5p33_ASAP7_75t_R g4248 ( 
.A(n_3548),
.Y(n_4248)
);

INVx1_ASAP7_75t_L g4249 ( 
.A(n_3118),
.Y(n_4249)
);

INVx1_ASAP7_75t_L g4250 ( 
.A(n_3118),
.Y(n_4250)
);

INVx1_ASAP7_75t_L g4251 ( 
.A(n_3118),
.Y(n_4251)
);

INVxp67_ASAP7_75t_SL g4252 ( 
.A(n_3078),
.Y(n_4252)
);

CKINVDCx5p33_ASAP7_75t_R g4253 ( 
.A(n_3597),
.Y(n_4253)
);

INVx2_ASAP7_75t_L g4254 ( 
.A(n_3118),
.Y(n_4254)
);

INVx1_ASAP7_75t_L g4255 ( 
.A(n_3183),
.Y(n_4255)
);

CKINVDCx5p33_ASAP7_75t_R g4256 ( 
.A(n_3943),
.Y(n_4256)
);

INVx1_ASAP7_75t_L g4257 ( 
.A(n_3183),
.Y(n_4257)
);

INVx1_ASAP7_75t_L g4258 ( 
.A(n_3183),
.Y(n_4258)
);

CKINVDCx20_ASAP7_75t_R g4259 ( 
.A(n_4056),
.Y(n_4259)
);

INVx1_ASAP7_75t_L g4260 ( 
.A(n_3183),
.Y(n_4260)
);

BUFx6f_ASAP7_75t_L g4261 ( 
.A(n_3029),
.Y(n_4261)
);

INVx1_ASAP7_75t_L g4262 ( 
.A(n_3183),
.Y(n_4262)
);

CKINVDCx5p33_ASAP7_75t_R g4263 ( 
.A(n_3024),
.Y(n_4263)
);

INVx1_ASAP7_75t_L g4264 ( 
.A(n_3224),
.Y(n_4264)
);

INVx1_ASAP7_75t_L g4265 ( 
.A(n_3224),
.Y(n_4265)
);

CKINVDCx5p33_ASAP7_75t_R g4266 ( 
.A(n_3035),
.Y(n_4266)
);

INVx1_ASAP7_75t_L g4267 ( 
.A(n_3224),
.Y(n_4267)
);

CKINVDCx5p33_ASAP7_75t_R g4268 ( 
.A(n_3073),
.Y(n_4268)
);

CKINVDCx5p33_ASAP7_75t_R g4269 ( 
.A(n_3413),
.Y(n_4269)
);

HB1xp67_ASAP7_75t_L g4270 ( 
.A(n_3497),
.Y(n_4270)
);

BUFx3_ASAP7_75t_L g4271 ( 
.A(n_3299),
.Y(n_4271)
);

INVx1_ASAP7_75t_L g4272 ( 
.A(n_3224),
.Y(n_4272)
);

CKINVDCx20_ASAP7_75t_R g4273 ( 
.A(n_3708),
.Y(n_4273)
);

CKINVDCx5p33_ASAP7_75t_R g4274 ( 
.A(n_3727),
.Y(n_4274)
);

INVx1_ASAP7_75t_L g4275 ( 
.A(n_3224),
.Y(n_4275)
);

INVx1_ASAP7_75t_L g4276 ( 
.A(n_3269),
.Y(n_4276)
);

CKINVDCx20_ASAP7_75t_R g4277 ( 
.A(n_3788),
.Y(n_4277)
);

INVx1_ASAP7_75t_L g4278 ( 
.A(n_3269),
.Y(n_4278)
);

CKINVDCx5p33_ASAP7_75t_R g4279 ( 
.A(n_3876),
.Y(n_4279)
);

INVxp67_ASAP7_75t_L g4280 ( 
.A(n_3250),
.Y(n_4280)
);

INVx2_ASAP7_75t_L g4281 ( 
.A(n_3269),
.Y(n_4281)
);

CKINVDCx5p33_ASAP7_75t_R g4282 ( 
.A(n_4011),
.Y(n_4282)
);

CKINVDCx5p33_ASAP7_75t_R g4283 ( 
.A(n_4038),
.Y(n_4283)
);

INVx1_ASAP7_75t_L g4284 ( 
.A(n_3269),
.Y(n_4284)
);

INVx1_ASAP7_75t_L g4285 ( 
.A(n_3269),
.Y(n_4285)
);

CKINVDCx20_ASAP7_75t_R g4286 ( 
.A(n_4061),
.Y(n_4286)
);

INVx1_ASAP7_75t_L g4287 ( 
.A(n_3331),
.Y(n_4287)
);

INVx1_ASAP7_75t_L g4288 ( 
.A(n_3331),
.Y(n_4288)
);

CKINVDCx5p33_ASAP7_75t_R g4289 ( 
.A(n_4088),
.Y(n_4289)
);

CKINVDCx16_ASAP7_75t_R g4290 ( 
.A(n_4123),
.Y(n_4290)
);

INVx2_ASAP7_75t_L g4291 ( 
.A(n_3331),
.Y(n_4291)
);

CKINVDCx5p33_ASAP7_75t_R g4292 ( 
.A(n_4127),
.Y(n_4292)
);

INVx2_ASAP7_75t_L g4293 ( 
.A(n_3331),
.Y(n_4293)
);

INVx1_ASAP7_75t_L g4294 ( 
.A(n_3331),
.Y(n_4294)
);

INVx1_ASAP7_75t_L g4295 ( 
.A(n_3655),
.Y(n_4295)
);

INVx1_ASAP7_75t_L g4296 ( 
.A(n_3655),
.Y(n_4296)
);

INVx1_ASAP7_75t_L g4297 ( 
.A(n_3655),
.Y(n_4297)
);

CKINVDCx5p33_ASAP7_75t_R g4298 ( 
.A(n_4185),
.Y(n_4298)
);

CKINVDCx5p33_ASAP7_75t_R g4299 ( 
.A(n_4192),
.Y(n_4299)
);

INVx1_ASAP7_75t_L g4300 ( 
.A(n_3655),
.Y(n_4300)
);

INVx1_ASAP7_75t_L g4301 ( 
.A(n_3655),
.Y(n_4301)
);

INVxp67_ASAP7_75t_L g4302 ( 
.A(n_3255),
.Y(n_4302)
);

INVxp33_ASAP7_75t_SL g4303 ( 
.A(n_3207),
.Y(n_4303)
);

INVx1_ASAP7_75t_L g4304 ( 
.A(n_3737),
.Y(n_4304)
);

BUFx3_ASAP7_75t_L g4305 ( 
.A(n_3488),
.Y(n_4305)
);

NOR2xp67_ASAP7_75t_L g4306 ( 
.A(n_2854),
.B(n_1),
.Y(n_4306)
);

INVx1_ASAP7_75t_L g4307 ( 
.A(n_3737),
.Y(n_4307)
);

INVx1_ASAP7_75t_L g4308 ( 
.A(n_3737),
.Y(n_4308)
);

INVx1_ASAP7_75t_SL g4309 ( 
.A(n_3270),
.Y(n_4309)
);

INVx1_ASAP7_75t_L g4310 ( 
.A(n_3737),
.Y(n_4310)
);

CKINVDCx5p33_ASAP7_75t_R g4311 ( 
.A(n_2827),
.Y(n_4311)
);

INVx1_ASAP7_75t_L g4312 ( 
.A(n_3737),
.Y(n_4312)
);

INVx1_ASAP7_75t_L g4313 ( 
.A(n_3872),
.Y(n_4313)
);

INVx1_ASAP7_75t_L g4314 ( 
.A(n_3872),
.Y(n_4314)
);

BUFx3_ASAP7_75t_L g4315 ( 
.A(n_3489),
.Y(n_4315)
);

INVx1_ASAP7_75t_L g4316 ( 
.A(n_3872),
.Y(n_4316)
);

INVx1_ASAP7_75t_L g4317 ( 
.A(n_3872),
.Y(n_4317)
);

CKINVDCx16_ASAP7_75t_R g4318 ( 
.A(n_3477),
.Y(n_4318)
);

INVx1_ASAP7_75t_L g4319 ( 
.A(n_3872),
.Y(n_4319)
);

CKINVDCx5p33_ASAP7_75t_R g4320 ( 
.A(n_2838),
.Y(n_4320)
);

INVx1_ASAP7_75t_L g4321 ( 
.A(n_3929),
.Y(n_4321)
);

BUFx2_ASAP7_75t_L g4322 ( 
.A(n_3369),
.Y(n_4322)
);

INVx1_ASAP7_75t_L g4323 ( 
.A(n_3929),
.Y(n_4323)
);

INVx2_ASAP7_75t_L g4324 ( 
.A(n_3929),
.Y(n_4324)
);

INVx1_ASAP7_75t_L g4325 ( 
.A(n_3929),
.Y(n_4325)
);

NOR2xp67_ASAP7_75t_L g4326 ( 
.A(n_2914),
.B(n_2),
.Y(n_4326)
);

INVx1_ASAP7_75t_L g4327 ( 
.A(n_3929),
.Y(n_4327)
);

INVxp33_ASAP7_75t_L g4328 ( 
.A(n_3315),
.Y(n_4328)
);

INVx1_ASAP7_75t_L g4329 ( 
.A(n_4004),
.Y(n_4329)
);

INVxp33_ASAP7_75t_SL g4330 ( 
.A(n_3448),
.Y(n_4330)
);

CKINVDCx20_ASAP7_75t_R g4331 ( 
.A(n_2818),
.Y(n_4331)
);

INVxp67_ASAP7_75t_SL g4332 ( 
.A(n_2914),
.Y(n_4332)
);

CKINVDCx5p33_ASAP7_75t_R g4333 ( 
.A(n_2868),
.Y(n_4333)
);

INVx2_ASAP7_75t_L g4334 ( 
.A(n_4004),
.Y(n_4334)
);

BUFx3_ASAP7_75t_L g4335 ( 
.A(n_3731),
.Y(n_4335)
);

BUFx2_ASAP7_75t_L g4336 ( 
.A(n_3385),
.Y(n_4336)
);

INVxp67_ASAP7_75t_L g4337 ( 
.A(n_3458),
.Y(n_4337)
);

INVx1_ASAP7_75t_L g4338 ( 
.A(n_4004),
.Y(n_4338)
);

CKINVDCx5p33_ASAP7_75t_R g4339 ( 
.A(n_2888),
.Y(n_4339)
);

CKINVDCx5p33_ASAP7_75t_R g4340 ( 
.A(n_2889),
.Y(n_4340)
);

INVxp67_ASAP7_75t_SL g4341 ( 
.A(n_3029),
.Y(n_4341)
);

INVx1_ASAP7_75t_L g4342 ( 
.A(n_4004),
.Y(n_4342)
);

BUFx10_ASAP7_75t_L g4343 ( 
.A(n_2894),
.Y(n_4343)
);

HB1xp67_ASAP7_75t_L g4344 ( 
.A(n_3463),
.Y(n_4344)
);

NOR2xp67_ASAP7_75t_L g4345 ( 
.A(n_3586),
.B(n_2),
.Y(n_4345)
);

INVx1_ASAP7_75t_L g4346 ( 
.A(n_4004),
.Y(n_4346)
);

INVx1_ASAP7_75t_L g4347 ( 
.A(n_4076),
.Y(n_4347)
);

INVx1_ASAP7_75t_L g4348 ( 
.A(n_4076),
.Y(n_4348)
);

INVx1_ASAP7_75t_L g4349 ( 
.A(n_4076),
.Y(n_4349)
);

INVxp33_ASAP7_75t_SL g4350 ( 
.A(n_3500),
.Y(n_4350)
);

CKINVDCx5p33_ASAP7_75t_R g4351 ( 
.A(n_2901),
.Y(n_4351)
);

CKINVDCx5p33_ASAP7_75t_R g4352 ( 
.A(n_2923),
.Y(n_4352)
);

INVx1_ASAP7_75t_L g4353 ( 
.A(n_4076),
.Y(n_4353)
);

INVx2_ASAP7_75t_L g4354 ( 
.A(n_4076),
.Y(n_4354)
);

INVx2_ASAP7_75t_L g4355 ( 
.A(n_4094),
.Y(n_4355)
);

CKINVDCx16_ASAP7_75t_R g4356 ( 
.A(n_3477),
.Y(n_4356)
);

INVx2_ASAP7_75t_L g4357 ( 
.A(n_4094),
.Y(n_4357)
);

INVx1_ASAP7_75t_SL g4358 ( 
.A(n_3484),
.Y(n_4358)
);

BUFx6f_ASAP7_75t_L g4359 ( 
.A(n_3029),
.Y(n_4359)
);

INVx1_ASAP7_75t_L g4360 ( 
.A(n_4094),
.Y(n_4360)
);

INVx1_ASAP7_75t_L g4361 ( 
.A(n_4094),
.Y(n_4361)
);

INVx2_ASAP7_75t_L g4362 ( 
.A(n_4094),
.Y(n_4362)
);

INVx1_ASAP7_75t_L g4363 ( 
.A(n_4190),
.Y(n_4363)
);

INVx1_ASAP7_75t_L g4364 ( 
.A(n_2831),
.Y(n_4364)
);

CKINVDCx20_ASAP7_75t_R g4365 ( 
.A(n_2862),
.Y(n_4365)
);

INVx1_ASAP7_75t_L g4366 ( 
.A(n_2835),
.Y(n_4366)
);

INVx2_ASAP7_75t_L g4367 ( 
.A(n_2847),
.Y(n_4367)
);

CKINVDCx20_ASAP7_75t_R g4368 ( 
.A(n_2871),
.Y(n_4368)
);

INVx1_ASAP7_75t_L g4369 ( 
.A(n_2859),
.Y(n_4369)
);

INVx1_ASAP7_75t_L g4370 ( 
.A(n_2921),
.Y(n_4370)
);

CKINVDCx16_ASAP7_75t_R g4371 ( 
.A(n_3753),
.Y(n_4371)
);

INVx1_ASAP7_75t_L g4372 ( 
.A(n_2949),
.Y(n_4372)
);

CKINVDCx5p33_ASAP7_75t_R g4373 ( 
.A(n_2936),
.Y(n_4373)
);

CKINVDCx5p33_ASAP7_75t_R g4374 ( 
.A(n_2950),
.Y(n_4374)
);

HB1xp67_ASAP7_75t_L g4375 ( 
.A(n_3770),
.Y(n_4375)
);

CKINVDCx5p33_ASAP7_75t_R g4376 ( 
.A(n_2958),
.Y(n_4376)
);

INVx1_ASAP7_75t_L g4377 ( 
.A(n_2974),
.Y(n_4377)
);

BUFx3_ASAP7_75t_L g4378 ( 
.A(n_4168),
.Y(n_4378)
);

INVx1_ASAP7_75t_L g4379 ( 
.A(n_3007),
.Y(n_4379)
);

INVx1_ASAP7_75t_L g4380 ( 
.A(n_3013),
.Y(n_4380)
);

INVx2_ASAP7_75t_L g4381 ( 
.A(n_3032),
.Y(n_4381)
);

INVxp33_ASAP7_75t_L g4382 ( 
.A(n_3883),
.Y(n_4382)
);

CKINVDCx5p33_ASAP7_75t_R g4383 ( 
.A(n_2959),
.Y(n_4383)
);

INVx1_ASAP7_75t_L g4384 ( 
.A(n_3034),
.Y(n_4384)
);

INVx1_ASAP7_75t_L g4385 ( 
.A(n_3042),
.Y(n_4385)
);

INVx1_ASAP7_75t_L g4386 ( 
.A(n_3047),
.Y(n_4386)
);

CKINVDCx20_ASAP7_75t_R g4387 ( 
.A(n_2873),
.Y(n_4387)
);

CKINVDCx5p33_ASAP7_75t_R g4388 ( 
.A(n_2987),
.Y(n_4388)
);

CKINVDCx5p33_ASAP7_75t_R g4389 ( 
.A(n_3019),
.Y(n_4389)
);

INVx1_ASAP7_75t_L g4390 ( 
.A(n_3095),
.Y(n_4390)
);

INVx1_ASAP7_75t_L g4391 ( 
.A(n_3112),
.Y(n_4391)
);

CKINVDCx5p33_ASAP7_75t_R g4392 ( 
.A(n_3041),
.Y(n_4392)
);

INVx1_ASAP7_75t_L g4393 ( 
.A(n_3125),
.Y(n_4393)
);

INVx1_ASAP7_75t_L g4394 ( 
.A(n_3126),
.Y(n_4394)
);

CKINVDCx5p33_ASAP7_75t_R g4395 ( 
.A(n_3045),
.Y(n_4395)
);

CKINVDCx16_ASAP7_75t_R g4396 ( 
.A(n_3753),
.Y(n_4396)
);

INVx2_ASAP7_75t_L g4397 ( 
.A(n_3156),
.Y(n_4397)
);

INVx1_ASAP7_75t_L g4398 ( 
.A(n_3196),
.Y(n_4398)
);

BUFx3_ASAP7_75t_L g4399 ( 
.A(n_2877),
.Y(n_4399)
);

CKINVDCx5p33_ASAP7_75t_R g4400 ( 
.A(n_3056),
.Y(n_4400)
);

INVx1_ASAP7_75t_L g4401 ( 
.A(n_3256),
.Y(n_4401)
);

INVx1_ASAP7_75t_L g4402 ( 
.A(n_3287),
.Y(n_4402)
);

INVx1_ASAP7_75t_L g4403 ( 
.A(n_3302),
.Y(n_4403)
);

CKINVDCx5p33_ASAP7_75t_R g4404 ( 
.A(n_3068),
.Y(n_4404)
);

INVx1_ASAP7_75t_L g4405 ( 
.A(n_3323),
.Y(n_4405)
);

CKINVDCx16_ASAP7_75t_R g4406 ( 
.A(n_3875),
.Y(n_4406)
);

CKINVDCx20_ASAP7_75t_R g4407 ( 
.A(n_2874),
.Y(n_4407)
);

INVx1_ASAP7_75t_L g4408 ( 
.A(n_3353),
.Y(n_4408)
);

CKINVDCx5p33_ASAP7_75t_R g4409 ( 
.A(n_3069),
.Y(n_4409)
);

CKINVDCx5p33_ASAP7_75t_R g4410 ( 
.A(n_3076),
.Y(n_4410)
);

CKINVDCx5p33_ASAP7_75t_R g4411 ( 
.A(n_3084),
.Y(n_4411)
);

INVx1_ASAP7_75t_L g4412 ( 
.A(n_3373),
.Y(n_4412)
);

INVx1_ASAP7_75t_L g4413 ( 
.A(n_3391),
.Y(n_4413)
);

INVx1_ASAP7_75t_L g4414 ( 
.A(n_3406),
.Y(n_4414)
);

INVx1_ASAP7_75t_L g4415 ( 
.A(n_3417),
.Y(n_4415)
);

INVxp33_ASAP7_75t_L g4416 ( 
.A(n_3926),
.Y(n_4416)
);

CKINVDCx20_ASAP7_75t_R g4417 ( 
.A(n_2880),
.Y(n_4417)
);

CKINVDCx16_ASAP7_75t_R g4418 ( 
.A(n_3875),
.Y(n_4418)
);

INVx2_ASAP7_75t_L g4419 ( 
.A(n_3507),
.Y(n_4419)
);

INVx1_ASAP7_75t_L g4420 ( 
.A(n_3509),
.Y(n_4420)
);

INVx1_ASAP7_75t_L g4421 ( 
.A(n_3605),
.Y(n_4421)
);

INVx1_ASAP7_75t_L g4422 ( 
.A(n_3730),
.Y(n_4422)
);

INVx1_ASAP7_75t_L g4423 ( 
.A(n_3755),
.Y(n_4423)
);

HB1xp67_ASAP7_75t_L g4424 ( 
.A(n_3986),
.Y(n_4424)
);

INVx2_ASAP7_75t_L g4425 ( 
.A(n_3764),
.Y(n_4425)
);

INVx1_ASAP7_75t_L g4426 ( 
.A(n_3765),
.Y(n_4426)
);

INVx1_ASAP7_75t_L g4427 ( 
.A(n_3769),
.Y(n_4427)
);

INVx1_ASAP7_75t_L g4428 ( 
.A(n_3804),
.Y(n_4428)
);

CKINVDCx5p33_ASAP7_75t_R g4429 ( 
.A(n_3093),
.Y(n_4429)
);

CKINVDCx5p33_ASAP7_75t_R g4430 ( 
.A(n_3096),
.Y(n_4430)
);

INVx1_ASAP7_75t_L g4431 ( 
.A(n_3814),
.Y(n_4431)
);

INVx1_ASAP7_75t_L g4432 ( 
.A(n_3821),
.Y(n_4432)
);

INVx2_ASAP7_75t_L g4433 ( 
.A(n_3822),
.Y(n_4433)
);

CKINVDCx5p33_ASAP7_75t_R g4434 ( 
.A(n_3106),
.Y(n_4434)
);

INVxp33_ASAP7_75t_L g4435 ( 
.A(n_4012),
.Y(n_4435)
);

INVx1_ASAP7_75t_L g4436 ( 
.A(n_3828),
.Y(n_4436)
);

INVx1_ASAP7_75t_SL g4437 ( 
.A(n_3581),
.Y(n_4437)
);

CKINVDCx5p33_ASAP7_75t_R g4438 ( 
.A(n_3136),
.Y(n_4438)
);

CKINVDCx14_ASAP7_75t_R g4439 ( 
.A(n_3818),
.Y(n_4439)
);

INVx1_ASAP7_75t_L g4440 ( 
.A(n_3837),
.Y(n_4440)
);

INVx1_ASAP7_75t_L g4441 ( 
.A(n_3884),
.Y(n_4441)
);

INVxp67_ASAP7_75t_L g4442 ( 
.A(n_3873),
.Y(n_4442)
);

INVx3_ASAP7_75t_L g4443 ( 
.A(n_3053),
.Y(n_4443)
);

CKINVDCx5p33_ASAP7_75t_R g4444 ( 
.A(n_3145),
.Y(n_4444)
);

BUFx3_ASAP7_75t_L g4445 ( 
.A(n_2965),
.Y(n_4445)
);

INVxp67_ASAP7_75t_SL g4446 ( 
.A(n_3117),
.Y(n_4446)
);

INVx2_ASAP7_75t_L g4447 ( 
.A(n_3947),
.Y(n_4447)
);

INVx2_ASAP7_75t_L g4448 ( 
.A(n_3953),
.Y(n_4448)
);

INVx1_ASAP7_75t_L g4449 ( 
.A(n_3966),
.Y(n_4449)
);

INVx1_ASAP7_75t_L g4450 ( 
.A(n_3969),
.Y(n_4450)
);

INVx1_ASAP7_75t_L g4451 ( 
.A(n_3981),
.Y(n_4451)
);

INVx2_ASAP7_75t_L g4452 ( 
.A(n_4016),
.Y(n_4452)
);

CKINVDCx5p33_ASAP7_75t_R g4453 ( 
.A(n_3149),
.Y(n_4453)
);

INVx1_ASAP7_75t_L g4454 ( 
.A(n_4047),
.Y(n_4454)
);

INVxp67_ASAP7_75t_L g4455 ( 
.A(n_3879),
.Y(n_4455)
);

CKINVDCx5p33_ASAP7_75t_R g4456 ( 
.A(n_3150),
.Y(n_4456)
);

INVx1_ASAP7_75t_L g4457 ( 
.A(n_4104),
.Y(n_4457)
);

HB1xp67_ASAP7_75t_L g4458 ( 
.A(n_3165),
.Y(n_4458)
);

INVx1_ASAP7_75t_L g4459 ( 
.A(n_4178),
.Y(n_4459)
);

INVx1_ASAP7_75t_L g4460 ( 
.A(n_3117),
.Y(n_4460)
);

INVx1_ASAP7_75t_L g4461 ( 
.A(n_3117),
.Y(n_4461)
);

CKINVDCx5p33_ASAP7_75t_R g4462 ( 
.A(n_3168),
.Y(n_4462)
);

NOR2xp33_ASAP7_75t_L g4463 ( 
.A(n_3688),
.B(n_3490),
.Y(n_4463)
);

INVx2_ASAP7_75t_L g4464 ( 
.A(n_2904),
.Y(n_4464)
);

INVx1_ASAP7_75t_L g4465 ( 
.A(n_4195),
.Y(n_4465)
);

CKINVDCx5p33_ASAP7_75t_R g4466 ( 
.A(n_3171),
.Y(n_4466)
);

NOR2xp67_ASAP7_75t_L g4467 ( 
.A(n_2842),
.B(n_3),
.Y(n_4467)
);

INVx1_ASAP7_75t_L g4468 ( 
.A(n_4195),
.Y(n_4468)
);

CKINVDCx5p33_ASAP7_75t_R g4469 ( 
.A(n_3176),
.Y(n_4469)
);

INVxp67_ASAP7_75t_SL g4470 ( 
.A(n_3148),
.Y(n_4470)
);

INVx1_ASAP7_75t_L g4471 ( 
.A(n_4195),
.Y(n_4471)
);

CKINVDCx5p33_ASAP7_75t_R g4472 ( 
.A(n_3179),
.Y(n_4472)
);

INVxp67_ASAP7_75t_SL g4473 ( 
.A(n_3148),
.Y(n_4473)
);

HB1xp67_ASAP7_75t_L g4474 ( 
.A(n_4193),
.Y(n_4474)
);

BUFx2_ASAP7_75t_L g4475 ( 
.A(n_3919),
.Y(n_4475)
);

BUFx6f_ASAP7_75t_L g4476 ( 
.A(n_3148),
.Y(n_4476)
);

INVx1_ASAP7_75t_L g4477 ( 
.A(n_3494),
.Y(n_4477)
);

INVx1_ASAP7_75t_L g4478 ( 
.A(n_3494),
.Y(n_4478)
);

CKINVDCx5p33_ASAP7_75t_R g4479 ( 
.A(n_3190),
.Y(n_4479)
);

INVx1_ASAP7_75t_L g4480 ( 
.A(n_3494),
.Y(n_4480)
);

BUFx2_ASAP7_75t_L g4481 ( 
.A(n_3993),
.Y(n_4481)
);

INVx1_ASAP7_75t_L g4482 ( 
.A(n_3529),
.Y(n_4482)
);

INVx1_ASAP7_75t_L g4483 ( 
.A(n_3529),
.Y(n_4483)
);

NOR2xp33_ASAP7_75t_L g4484 ( 
.A(n_4046),
.B(n_3),
.Y(n_4484)
);

INVx1_ASAP7_75t_L g4485 ( 
.A(n_3529),
.Y(n_4485)
);

CKINVDCx5p33_ASAP7_75t_R g4486 ( 
.A(n_3193),
.Y(n_4486)
);

INVx1_ASAP7_75t_L g4487 ( 
.A(n_2925),
.Y(n_4487)
);

INVx1_ASAP7_75t_L g4488 ( 
.A(n_3144),
.Y(n_4488)
);

INVx1_ASAP7_75t_L g4489 ( 
.A(n_3593),
.Y(n_4489)
);

INVx1_ASAP7_75t_SL g4490 ( 
.A(n_3135),
.Y(n_4490)
);

INVx1_ASAP7_75t_L g4491 ( 
.A(n_3661),
.Y(n_4491)
);

CKINVDCx5p33_ASAP7_75t_R g4492 ( 
.A(n_3206),
.Y(n_4492)
);

BUFx6f_ASAP7_75t_L g4493 ( 
.A(n_3053),
.Y(n_4493)
);

INVx1_ASAP7_75t_L g4494 ( 
.A(n_3893),
.Y(n_4494)
);

INVx1_ASAP7_75t_L g4495 ( 
.A(n_3916),
.Y(n_4495)
);

INVxp67_ASAP7_75t_SL g4496 ( 
.A(n_3053),
.Y(n_4496)
);

INVx1_ASAP7_75t_L g4497 ( 
.A(n_4018),
.Y(n_4497)
);

CKINVDCx5p33_ASAP7_75t_R g4498 ( 
.A(n_3208),
.Y(n_4498)
);

INVx1_ASAP7_75t_L g4499 ( 
.A(n_4087),
.Y(n_4499)
);

CKINVDCx5p33_ASAP7_75t_R g4500 ( 
.A(n_3259),
.Y(n_4500)
);

INVx1_ASAP7_75t_L g4501 ( 
.A(n_4106),
.Y(n_4501)
);

INVx1_ASAP7_75t_L g4502 ( 
.A(n_4120),
.Y(n_4502)
);

INVx2_ASAP7_75t_L g4503 ( 
.A(n_3401),
.Y(n_4503)
);

CKINVDCx5p33_ASAP7_75t_R g4504 ( 
.A(n_3275),
.Y(n_4504)
);

INVx1_ASAP7_75t_L g4505 ( 
.A(n_3401),
.Y(n_4505)
);

BUFx2_ASAP7_75t_SL g4506 ( 
.A(n_2947),
.Y(n_4506)
);

BUFx3_ASAP7_75t_L g4507 ( 
.A(n_2968),
.Y(n_4507)
);

BUFx3_ASAP7_75t_L g4508 ( 
.A(n_2975),
.Y(n_4508)
);

INVx1_ASAP7_75t_L g4509 ( 
.A(n_3401),
.Y(n_4509)
);

INVx1_ASAP7_75t_L g4510 ( 
.A(n_3482),
.Y(n_4510)
);

CKINVDCx16_ASAP7_75t_R g4511 ( 
.A(n_3120),
.Y(n_4511)
);

INVx2_ASAP7_75t_L g4512 ( 
.A(n_3482),
.Y(n_4512)
);

BUFx3_ASAP7_75t_L g4513 ( 
.A(n_2985),
.Y(n_4513)
);

INVx1_ASAP7_75t_L g4514 ( 
.A(n_3482),
.Y(n_4514)
);

INVx1_ASAP7_75t_L g4515 ( 
.A(n_3504),
.Y(n_4515)
);

INVx1_ASAP7_75t_L g4516 ( 
.A(n_3504),
.Y(n_4516)
);

BUFx3_ASAP7_75t_L g4517 ( 
.A(n_3005),
.Y(n_4517)
);

CKINVDCx5p33_ASAP7_75t_R g4518 ( 
.A(n_3278),
.Y(n_4518)
);

INVx1_ASAP7_75t_L g4519 ( 
.A(n_3504),
.Y(n_4519)
);

BUFx2_ASAP7_75t_L g4520 ( 
.A(n_3281),
.Y(n_4520)
);

CKINVDCx20_ASAP7_75t_R g4521 ( 
.A(n_2900),
.Y(n_4521)
);

BUFx2_ASAP7_75t_L g4522 ( 
.A(n_3286),
.Y(n_4522)
);

INVx2_ASAP7_75t_L g4523 ( 
.A(n_3705),
.Y(n_4523)
);

INVxp33_ASAP7_75t_SL g4524 ( 
.A(n_3288),
.Y(n_4524)
);

INVx1_ASAP7_75t_L g4525 ( 
.A(n_3705),
.Y(n_4525)
);

INVx1_ASAP7_75t_L g4526 ( 
.A(n_3705),
.Y(n_4526)
);

BUFx2_ASAP7_75t_SL g4527 ( 
.A(n_3062),
.Y(n_4527)
);

INVx1_ASAP7_75t_L g4528 ( 
.A(n_3831),
.Y(n_4528)
);

HB1xp67_ASAP7_75t_L g4529 ( 
.A(n_4187),
.Y(n_4529)
);

INVx2_ASAP7_75t_L g4530 ( 
.A(n_3831),
.Y(n_4530)
);

CKINVDCx14_ASAP7_75t_R g4531 ( 
.A(n_3120),
.Y(n_4531)
);

BUFx2_ASAP7_75t_L g4532 ( 
.A(n_3291),
.Y(n_4532)
);

INVx1_ASAP7_75t_L g4533 ( 
.A(n_3831),
.Y(n_4533)
);

INVx1_ASAP7_75t_L g4534 ( 
.A(n_3910),
.Y(n_4534)
);

INVx1_ASAP7_75t_L g4535 ( 
.A(n_3910),
.Y(n_4535)
);

NOR2xp33_ASAP7_75t_L g4536 ( 
.A(n_3044),
.B(n_3),
.Y(n_4536)
);

INVx1_ASAP7_75t_L g4537 ( 
.A(n_3910),
.Y(n_4537)
);

CKINVDCx5p33_ASAP7_75t_R g4538 ( 
.A(n_3296),
.Y(n_4538)
);

CKINVDCx5p33_ASAP7_75t_R g4539 ( 
.A(n_3343),
.Y(n_4539)
);

INVx1_ASAP7_75t_L g4540 ( 
.A(n_3952),
.Y(n_4540)
);

INVx1_ASAP7_75t_L g4541 ( 
.A(n_3952),
.Y(n_4541)
);

INVx1_ASAP7_75t_L g4542 ( 
.A(n_3952),
.Y(n_4542)
);

INVx1_ASAP7_75t_L g4543 ( 
.A(n_3990),
.Y(n_4543)
);

INVx1_ASAP7_75t_L g4544 ( 
.A(n_3990),
.Y(n_4544)
);

CKINVDCx5p33_ASAP7_75t_R g4545 ( 
.A(n_3345),
.Y(n_4545)
);

INVxp67_ASAP7_75t_SL g4546 ( 
.A(n_3990),
.Y(n_4546)
);

CKINVDCx16_ASAP7_75t_R g4547 ( 
.A(n_3146),
.Y(n_4547)
);

INVx1_ASAP7_75t_L g4548 ( 
.A(n_4030),
.Y(n_4548)
);

INVx1_ASAP7_75t_L g4549 ( 
.A(n_4030),
.Y(n_4549)
);

CKINVDCx5p33_ASAP7_75t_R g4550 ( 
.A(n_3366),
.Y(n_4550)
);

NOR2xp67_ASAP7_75t_L g4551 ( 
.A(n_3115),
.B(n_4),
.Y(n_4551)
);

INVx1_ASAP7_75t_L g4552 ( 
.A(n_4030),
.Y(n_4552)
);

BUFx3_ASAP7_75t_L g4553 ( 
.A(n_3011),
.Y(n_4553)
);

INVx1_ASAP7_75t_L g4554 ( 
.A(n_3052),
.Y(n_4554)
);

INVx1_ASAP7_75t_L g4555 ( 
.A(n_3167),
.Y(n_4555)
);

INVx1_ASAP7_75t_L g4556 ( 
.A(n_3295),
.Y(n_4556)
);

INVx1_ASAP7_75t_L g4557 ( 
.A(n_3442),
.Y(n_4557)
);

BUFx6f_ASAP7_75t_L g4558 ( 
.A(n_3466),
.Y(n_4558)
);

HB1xp67_ASAP7_75t_L g4559 ( 
.A(n_3382),
.Y(n_4559)
);

INVx1_ASAP7_75t_L g4560 ( 
.A(n_3553),
.Y(n_4560)
);

CKINVDCx16_ASAP7_75t_R g4561 ( 
.A(n_3146),
.Y(n_4561)
);

INVx1_ASAP7_75t_L g4562 ( 
.A(n_3579),
.Y(n_4562)
);

INVxp67_ASAP7_75t_L g4563 ( 
.A(n_3261),
.Y(n_4563)
);

INVx1_ASAP7_75t_L g4564 ( 
.A(n_3631),
.Y(n_4564)
);

INVxp67_ASAP7_75t_L g4565 ( 
.A(n_3261),
.Y(n_4565)
);

INVx1_ASAP7_75t_L g4566 ( 
.A(n_3702),
.Y(n_4566)
);

NOR2xp33_ASAP7_75t_L g4567 ( 
.A(n_3055),
.B(n_4),
.Y(n_4567)
);

INVx1_ASAP7_75t_L g4568 ( 
.A(n_3712),
.Y(n_4568)
);

INVx1_ASAP7_75t_L g4569 ( 
.A(n_3782),
.Y(n_4569)
);

INVx1_ASAP7_75t_L g4570 ( 
.A(n_3798),
.Y(n_4570)
);

CKINVDCx5p33_ASAP7_75t_R g4571 ( 
.A(n_3387),
.Y(n_4571)
);

HB1xp67_ASAP7_75t_L g4572 ( 
.A(n_3403),
.Y(n_4572)
);

INVx1_ASAP7_75t_L g4573 ( 
.A(n_3824),
.Y(n_4573)
);

INVxp67_ASAP7_75t_L g4574 ( 
.A(n_3265),
.Y(n_4574)
);

CKINVDCx16_ASAP7_75t_R g4575 ( 
.A(n_4180),
.Y(n_4575)
);

INVxp67_ASAP7_75t_L g4576 ( 
.A(n_3265),
.Y(n_4576)
);

INVx1_ASAP7_75t_L g4577 ( 
.A(n_3858),
.Y(n_4577)
);

INVx1_ASAP7_75t_L g4578 ( 
.A(n_3877),
.Y(n_4578)
);

CKINVDCx5p33_ASAP7_75t_R g4579 ( 
.A(n_3422),
.Y(n_4579)
);

INVx1_ASAP7_75t_L g4580 ( 
.A(n_4005),
.Y(n_4580)
);

INVxp33_ASAP7_75t_SL g4581 ( 
.A(n_3429),
.Y(n_4581)
);

INVx1_ASAP7_75t_L g4582 ( 
.A(n_4020),
.Y(n_4582)
);

INVxp33_ASAP7_75t_L g4583 ( 
.A(n_2823),
.Y(n_4583)
);

CKINVDCx5p33_ASAP7_75t_R g4584 ( 
.A(n_3439),
.Y(n_4584)
);

INVx1_ASAP7_75t_L g4585 ( 
.A(n_4051),
.Y(n_4585)
);

INVx1_ASAP7_75t_L g4586 ( 
.A(n_4079),
.Y(n_4586)
);

INVx1_ASAP7_75t_L g4587 ( 
.A(n_4155),
.Y(n_4587)
);

CKINVDCx5p33_ASAP7_75t_R g4588 ( 
.A(n_3453),
.Y(n_4588)
);

INVx1_ASAP7_75t_L g4589 ( 
.A(n_4179),
.Y(n_4589)
);

INVx2_ASAP7_75t_L g4590 ( 
.A(n_2824),
.Y(n_4590)
);

CKINVDCx20_ASAP7_75t_R g4591 ( 
.A(n_2927),
.Y(n_4591)
);

INVx1_ASAP7_75t_SL g4592 ( 
.A(n_2820),
.Y(n_4592)
);

INVx1_ASAP7_75t_L g4593 ( 
.A(n_4196),
.Y(n_4593)
);

INVx1_ASAP7_75t_L g4594 ( 
.A(n_2825),
.Y(n_4594)
);

INVx1_ASAP7_75t_L g4595 ( 
.A(n_2826),
.Y(n_4595)
);

INVx1_ASAP7_75t_L g4596 ( 
.A(n_2828),
.Y(n_4596)
);

INVx1_ASAP7_75t_L g4597 ( 
.A(n_2840),
.Y(n_4597)
);

INVx1_ASAP7_75t_L g4598 ( 
.A(n_2841),
.Y(n_4598)
);

INVx1_ASAP7_75t_L g4599 ( 
.A(n_2851),
.Y(n_4599)
);

INVx1_ASAP7_75t_L g4600 ( 
.A(n_2852),
.Y(n_4600)
);

INVx1_ASAP7_75t_L g4601 ( 
.A(n_2853),
.Y(n_4601)
);

INVx2_ASAP7_75t_L g4602 ( 
.A(n_2858),
.Y(n_4602)
);

INVx1_ASAP7_75t_SL g4603 ( 
.A(n_3033),
.Y(n_4603)
);

CKINVDCx16_ASAP7_75t_R g4604 ( 
.A(n_3272),
.Y(n_4604)
);

CKINVDCx5p33_ASAP7_75t_R g4605 ( 
.A(n_3454),
.Y(n_4605)
);

INVx1_ASAP7_75t_L g4606 ( 
.A(n_4174),
.Y(n_4606)
);

INVx1_ASAP7_75t_L g4607 ( 
.A(n_2869),
.Y(n_4607)
);

NAND2xp5_ASAP7_75t_L g4608 ( 
.A(n_3303),
.B(n_5),
.Y(n_4608)
);

INVx1_ASAP7_75t_L g4609 ( 
.A(n_2872),
.Y(n_4609)
);

INVx1_ASAP7_75t_L g4610 ( 
.A(n_2876),
.Y(n_4610)
);

BUFx6f_ASAP7_75t_L g4611 ( 
.A(n_2848),
.Y(n_4611)
);

INVx1_ASAP7_75t_SL g4612 ( 
.A(n_3563),
.Y(n_4612)
);

OR2x2_ASAP7_75t_L g4613 ( 
.A(n_3022),
.B(n_5),
.Y(n_4613)
);

INVx1_ASAP7_75t_L g4614 ( 
.A(n_2881),
.Y(n_4614)
);

INVx1_ASAP7_75t_L g4615 ( 
.A(n_2884),
.Y(n_4615)
);

CKINVDCx5p33_ASAP7_75t_R g4616 ( 
.A(n_3469),
.Y(n_4616)
);

CKINVDCx16_ASAP7_75t_R g4617 ( 
.A(n_3272),
.Y(n_4617)
);

CKINVDCx5p33_ASAP7_75t_R g4618 ( 
.A(n_3496),
.Y(n_4618)
);

CKINVDCx5p33_ASAP7_75t_R g4619 ( 
.A(n_3520),
.Y(n_4619)
);

INVx1_ASAP7_75t_L g4620 ( 
.A(n_2887),
.Y(n_4620)
);

CKINVDCx20_ASAP7_75t_R g4621 ( 
.A(n_4331),
.Y(n_4621)
);

HB1xp67_ASAP7_75t_L g4622 ( 
.A(n_4263),
.Y(n_4622)
);

CKINVDCx20_ASAP7_75t_R g4623 ( 
.A(n_4365),
.Y(n_4623)
);

INVx1_ASAP7_75t_L g4624 ( 
.A(n_4496),
.Y(n_4624)
);

CKINVDCx5p33_ASAP7_75t_R g4625 ( 
.A(n_4202),
.Y(n_4625)
);

CKINVDCx5p33_ASAP7_75t_R g4626 ( 
.A(n_4207),
.Y(n_4626)
);

CKINVDCx5p33_ASAP7_75t_R g4627 ( 
.A(n_4209),
.Y(n_4627)
);

CKINVDCx20_ASAP7_75t_R g4628 ( 
.A(n_4368),
.Y(n_4628)
);

INVx1_ASAP7_75t_L g4629 ( 
.A(n_4546),
.Y(n_4629)
);

CKINVDCx20_ASAP7_75t_R g4630 ( 
.A(n_4387),
.Y(n_4630)
);

CKINVDCx20_ASAP7_75t_R g4631 ( 
.A(n_4407),
.Y(n_4631)
);

INVx1_ASAP7_75t_L g4632 ( 
.A(n_4341),
.Y(n_4632)
);

CKINVDCx20_ASAP7_75t_R g4633 ( 
.A(n_4417),
.Y(n_4633)
);

CKINVDCx5p33_ASAP7_75t_R g4634 ( 
.A(n_4311),
.Y(n_4634)
);

CKINVDCx5p33_ASAP7_75t_R g4635 ( 
.A(n_4320),
.Y(n_4635)
);

INVx1_ASAP7_75t_L g4636 ( 
.A(n_4446),
.Y(n_4636)
);

CKINVDCx20_ASAP7_75t_R g4637 ( 
.A(n_4521),
.Y(n_4637)
);

INVx1_ASAP7_75t_L g4638 ( 
.A(n_4470),
.Y(n_4638)
);

INVx1_ASAP7_75t_L g4639 ( 
.A(n_4473),
.Y(n_4639)
);

CKINVDCx5p33_ASAP7_75t_R g4640 ( 
.A(n_4333),
.Y(n_4640)
);

NOR2xp67_ASAP7_75t_L g4641 ( 
.A(n_4339),
.B(n_3202),
.Y(n_4641)
);

INVx1_ASAP7_75t_L g4642 ( 
.A(n_4198),
.Y(n_4642)
);

INVx1_ASAP7_75t_L g4643 ( 
.A(n_4200),
.Y(n_4643)
);

INVxp33_ASAP7_75t_SL g4644 ( 
.A(n_4199),
.Y(n_4644)
);

NOR2xp33_ASAP7_75t_L g4645 ( 
.A(n_4463),
.B(n_3587),
.Y(n_4645)
);

CKINVDCx20_ASAP7_75t_R g4646 ( 
.A(n_4591),
.Y(n_4646)
);

CKINVDCx5p33_ASAP7_75t_R g4647 ( 
.A(n_4340),
.Y(n_4647)
);

INVx1_ASAP7_75t_L g4648 ( 
.A(n_4204),
.Y(n_4648)
);

INVx1_ASAP7_75t_L g4649 ( 
.A(n_4205),
.Y(n_4649)
);

INVx1_ASAP7_75t_L g4650 ( 
.A(n_4206),
.Y(n_4650)
);

INVxp67_ASAP7_75t_SL g4651 ( 
.A(n_4399),
.Y(n_4651)
);

NOR2xp33_ASAP7_75t_L g4652 ( 
.A(n_4524),
.B(n_3604),
.Y(n_4652)
);

CKINVDCx20_ASAP7_75t_R g4653 ( 
.A(n_4259),
.Y(n_4653)
);

CKINVDCx5p33_ASAP7_75t_R g4654 ( 
.A(n_4351),
.Y(n_4654)
);

INVx1_ASAP7_75t_L g4655 ( 
.A(n_4210),
.Y(n_4655)
);

INVx1_ASAP7_75t_L g4656 ( 
.A(n_4211),
.Y(n_4656)
);

HB1xp67_ASAP7_75t_L g4657 ( 
.A(n_4266),
.Y(n_4657)
);

INVx1_ASAP7_75t_L g4658 ( 
.A(n_4212),
.Y(n_4658)
);

INVx1_ASAP7_75t_L g4659 ( 
.A(n_4215),
.Y(n_4659)
);

CKINVDCx5p33_ASAP7_75t_R g4660 ( 
.A(n_4352),
.Y(n_4660)
);

CKINVDCx5p33_ASAP7_75t_R g4661 ( 
.A(n_4373),
.Y(n_4661)
);

CKINVDCx20_ASAP7_75t_R g4662 ( 
.A(n_4273),
.Y(n_4662)
);

INVx1_ASAP7_75t_L g4663 ( 
.A(n_4216),
.Y(n_4663)
);

INVx1_ASAP7_75t_L g4664 ( 
.A(n_4493),
.Y(n_4664)
);

INVx1_ASAP7_75t_L g4665 ( 
.A(n_4493),
.Y(n_4665)
);

CKINVDCx5p33_ASAP7_75t_R g4666 ( 
.A(n_4374),
.Y(n_4666)
);

INVx1_ASAP7_75t_L g4667 ( 
.A(n_4493),
.Y(n_4667)
);

INVx1_ASAP7_75t_L g4668 ( 
.A(n_4460),
.Y(n_4668)
);

CKINVDCx5p33_ASAP7_75t_R g4669 ( 
.A(n_4376),
.Y(n_4669)
);

NOR2xp67_ASAP7_75t_L g4670 ( 
.A(n_4383),
.B(n_3249),
.Y(n_4670)
);

CKINVDCx20_ASAP7_75t_R g4671 ( 
.A(n_4277),
.Y(n_4671)
);

INVxp67_ASAP7_75t_L g4672 ( 
.A(n_4270),
.Y(n_4672)
);

INVx1_ASAP7_75t_L g4673 ( 
.A(n_4461),
.Y(n_4673)
);

INVx1_ASAP7_75t_L g4674 ( 
.A(n_4465),
.Y(n_4674)
);

CKINVDCx5p33_ASAP7_75t_R g4675 ( 
.A(n_4388),
.Y(n_4675)
);

INVx1_ASAP7_75t_L g4676 ( 
.A(n_4468),
.Y(n_4676)
);

INVx1_ASAP7_75t_SL g4677 ( 
.A(n_4490),
.Y(n_4677)
);

CKINVDCx5p33_ASAP7_75t_R g4678 ( 
.A(n_4389),
.Y(n_4678)
);

INVxp33_ASAP7_75t_SL g4679 ( 
.A(n_4268),
.Y(n_4679)
);

INVx1_ASAP7_75t_L g4680 ( 
.A(n_4471),
.Y(n_4680)
);

INVx1_ASAP7_75t_L g4681 ( 
.A(n_4477),
.Y(n_4681)
);

INVx1_ASAP7_75t_L g4682 ( 
.A(n_4478),
.Y(n_4682)
);

INVx1_ASAP7_75t_L g4683 ( 
.A(n_4480),
.Y(n_4683)
);

CKINVDCx20_ASAP7_75t_R g4684 ( 
.A(n_4286),
.Y(n_4684)
);

INVxp33_ASAP7_75t_SL g4685 ( 
.A(n_4269),
.Y(n_4685)
);

CKINVDCx20_ASAP7_75t_R g4686 ( 
.A(n_4247),
.Y(n_4686)
);

INVx1_ASAP7_75t_L g4687 ( 
.A(n_4482),
.Y(n_4687)
);

CKINVDCx20_ASAP7_75t_R g4688 ( 
.A(n_4290),
.Y(n_4688)
);

INVx1_ASAP7_75t_L g4689 ( 
.A(n_4483),
.Y(n_4689)
);

BUFx3_ASAP7_75t_L g4690 ( 
.A(n_4217),
.Y(n_4690)
);

CKINVDCx5p33_ASAP7_75t_R g4691 ( 
.A(n_4392),
.Y(n_4691)
);

INVx1_ASAP7_75t_L g4692 ( 
.A(n_4485),
.Y(n_4692)
);

INVx1_ASAP7_75t_L g4693 ( 
.A(n_4261),
.Y(n_4693)
);

HB1xp67_ASAP7_75t_L g4694 ( 
.A(n_4274),
.Y(n_4694)
);

CKINVDCx5p33_ASAP7_75t_R g4695 ( 
.A(n_4395),
.Y(n_4695)
);

INVx1_ASAP7_75t_L g4696 ( 
.A(n_4261),
.Y(n_4696)
);

INVxp67_ASAP7_75t_SL g4697 ( 
.A(n_4445),
.Y(n_4697)
);

CKINVDCx5p33_ASAP7_75t_R g4698 ( 
.A(n_4400),
.Y(n_4698)
);

INVx1_ASAP7_75t_L g4699 ( 
.A(n_4261),
.Y(n_4699)
);

INVx1_ASAP7_75t_L g4700 ( 
.A(n_4359),
.Y(n_4700)
);

CKINVDCx5p33_ASAP7_75t_R g4701 ( 
.A(n_4404),
.Y(n_4701)
);

NOR2xp33_ASAP7_75t_L g4702 ( 
.A(n_4581),
.B(n_4242),
.Y(n_4702)
);

CKINVDCx20_ASAP7_75t_R g4703 ( 
.A(n_4221),
.Y(n_4703)
);

INVx1_ASAP7_75t_L g4704 ( 
.A(n_4359),
.Y(n_4704)
);

HB1xp67_ASAP7_75t_L g4705 ( 
.A(n_4279),
.Y(n_4705)
);

CKINVDCx5p33_ASAP7_75t_R g4706 ( 
.A(n_4409),
.Y(n_4706)
);

INVx1_ASAP7_75t_L g4707 ( 
.A(n_4359),
.Y(n_4707)
);

INVx1_ASAP7_75t_L g4708 ( 
.A(n_4476),
.Y(n_4708)
);

INVx1_ASAP7_75t_L g4709 ( 
.A(n_4476),
.Y(n_4709)
);

CKINVDCx20_ASAP7_75t_R g4710 ( 
.A(n_4240),
.Y(n_4710)
);

INVxp33_ASAP7_75t_L g4711 ( 
.A(n_4458),
.Y(n_4711)
);

INVx1_ASAP7_75t_L g4712 ( 
.A(n_4476),
.Y(n_4712)
);

CKINVDCx5p33_ASAP7_75t_R g4713 ( 
.A(n_4410),
.Y(n_4713)
);

INVx1_ASAP7_75t_L g4714 ( 
.A(n_4503),
.Y(n_4714)
);

INVx1_ASAP7_75t_L g4715 ( 
.A(n_4512),
.Y(n_4715)
);

INVxp67_ASAP7_75t_L g4716 ( 
.A(n_4474),
.Y(n_4716)
);

INVx1_ASAP7_75t_L g4717 ( 
.A(n_4523),
.Y(n_4717)
);

CKINVDCx5p33_ASAP7_75t_R g4718 ( 
.A(n_4411),
.Y(n_4718)
);

CKINVDCx5p33_ASAP7_75t_R g4719 ( 
.A(n_4429),
.Y(n_4719)
);

INVx1_ASAP7_75t_L g4720 ( 
.A(n_4530),
.Y(n_4720)
);

CKINVDCx20_ASAP7_75t_R g4721 ( 
.A(n_4282),
.Y(n_4721)
);

INVx1_ASAP7_75t_L g4722 ( 
.A(n_4226),
.Y(n_4722)
);

BUFx6f_ASAP7_75t_SL g4723 ( 
.A(n_4343),
.Y(n_4723)
);

INVx1_ASAP7_75t_L g4724 ( 
.A(n_4252),
.Y(n_4724)
);

INVx1_ASAP7_75t_L g4725 ( 
.A(n_4505),
.Y(n_4725)
);

CKINVDCx5p33_ASAP7_75t_R g4726 ( 
.A(n_4430),
.Y(n_4726)
);

CKINVDCx5p33_ASAP7_75t_R g4727 ( 
.A(n_4434),
.Y(n_4727)
);

CKINVDCx5p33_ASAP7_75t_R g4728 ( 
.A(n_4438),
.Y(n_4728)
);

INVx1_ASAP7_75t_L g4729 ( 
.A(n_4509),
.Y(n_4729)
);

CKINVDCx20_ASAP7_75t_R g4730 ( 
.A(n_4283),
.Y(n_4730)
);

INVx2_ASAP7_75t_L g4731 ( 
.A(n_4443),
.Y(n_4731)
);

CKINVDCx5p33_ASAP7_75t_R g4732 ( 
.A(n_4444),
.Y(n_4732)
);

CKINVDCx20_ASAP7_75t_R g4733 ( 
.A(n_4289),
.Y(n_4733)
);

CKINVDCx5p33_ASAP7_75t_R g4734 ( 
.A(n_4453),
.Y(n_4734)
);

NOR2xp33_ASAP7_75t_L g4735 ( 
.A(n_4244),
.B(n_3523),
.Y(n_4735)
);

CKINVDCx14_ASAP7_75t_R g4736 ( 
.A(n_4531),
.Y(n_4736)
);

NOR2xp33_ASAP7_75t_L g4737 ( 
.A(n_4246),
.B(n_3527),
.Y(n_4737)
);

INVx1_ASAP7_75t_L g4738 ( 
.A(n_4510),
.Y(n_4738)
);

INVx1_ASAP7_75t_L g4739 ( 
.A(n_4514),
.Y(n_4739)
);

INVx1_ASAP7_75t_L g4740 ( 
.A(n_4515),
.Y(n_4740)
);

NAND2xp5_ASAP7_75t_L g4741 ( 
.A(n_4332),
.B(n_3329),
.Y(n_4741)
);

INVxp67_ASAP7_75t_SL g4742 ( 
.A(n_4507),
.Y(n_4742)
);

CKINVDCx20_ASAP7_75t_R g4743 ( 
.A(n_4292),
.Y(n_4743)
);

INVx1_ASAP7_75t_L g4744 ( 
.A(n_4516),
.Y(n_4744)
);

CKINVDCx5p33_ASAP7_75t_R g4745 ( 
.A(n_4456),
.Y(n_4745)
);

INVx1_ASAP7_75t_L g4746 ( 
.A(n_4519),
.Y(n_4746)
);

CKINVDCx20_ASAP7_75t_R g4747 ( 
.A(n_4298),
.Y(n_4747)
);

INVx1_ASAP7_75t_L g4748 ( 
.A(n_4525),
.Y(n_4748)
);

CKINVDCx20_ASAP7_75t_R g4749 ( 
.A(n_4299),
.Y(n_4749)
);

INVxp67_ASAP7_75t_SL g4750 ( 
.A(n_4508),
.Y(n_4750)
);

INVxp33_ASAP7_75t_SL g4751 ( 
.A(n_4220),
.Y(n_4751)
);

INVx1_ASAP7_75t_L g4752 ( 
.A(n_4526),
.Y(n_4752)
);

CKINVDCx20_ASAP7_75t_R g4753 ( 
.A(n_4222),
.Y(n_4753)
);

INVx1_ASAP7_75t_L g4754 ( 
.A(n_4528),
.Y(n_4754)
);

BUFx3_ASAP7_75t_L g4755 ( 
.A(n_4271),
.Y(n_4755)
);

INVxp67_ASAP7_75t_L g4756 ( 
.A(n_4529),
.Y(n_4756)
);

INVx1_ASAP7_75t_L g4757 ( 
.A(n_4533),
.Y(n_4757)
);

INVx1_ASAP7_75t_L g4758 ( 
.A(n_4534),
.Y(n_4758)
);

INVx1_ASAP7_75t_L g4759 ( 
.A(n_4535),
.Y(n_4759)
);

INVx1_ASAP7_75t_L g4760 ( 
.A(n_4537),
.Y(n_4760)
);

CKINVDCx5p33_ASAP7_75t_R g4761 ( 
.A(n_4462),
.Y(n_4761)
);

CKINVDCx20_ASAP7_75t_R g4762 ( 
.A(n_4234),
.Y(n_4762)
);

INVx1_ASAP7_75t_L g4763 ( 
.A(n_4540),
.Y(n_4763)
);

INVx1_ASAP7_75t_L g4764 ( 
.A(n_4541),
.Y(n_4764)
);

CKINVDCx20_ASAP7_75t_R g4765 ( 
.A(n_4235),
.Y(n_4765)
);

CKINVDCx5p33_ASAP7_75t_R g4766 ( 
.A(n_4466),
.Y(n_4766)
);

INVx1_ASAP7_75t_L g4767 ( 
.A(n_4542),
.Y(n_4767)
);

INVx1_ASAP7_75t_L g4768 ( 
.A(n_4543),
.Y(n_4768)
);

INVx1_ASAP7_75t_L g4769 ( 
.A(n_4544),
.Y(n_4769)
);

NOR2xp67_ASAP7_75t_L g4770 ( 
.A(n_4469),
.B(n_3350),
.Y(n_4770)
);

NOR2xp67_ASAP7_75t_L g4771 ( 
.A(n_4472),
.B(n_3355),
.Y(n_4771)
);

INVx1_ASAP7_75t_L g4772 ( 
.A(n_4548),
.Y(n_4772)
);

CKINVDCx5p33_ASAP7_75t_R g4773 ( 
.A(n_4479),
.Y(n_4773)
);

XOR2xp5_ASAP7_75t_L g4774 ( 
.A(n_4511),
.B(n_4547),
.Y(n_4774)
);

CKINVDCx16_ASAP7_75t_R g4775 ( 
.A(n_4318),
.Y(n_4775)
);

CKINVDCx20_ASAP7_75t_R g4776 ( 
.A(n_4439),
.Y(n_4776)
);

BUFx3_ASAP7_75t_L g4777 ( 
.A(n_4305),
.Y(n_4777)
);

CKINVDCx5p33_ASAP7_75t_R g4778 ( 
.A(n_4486),
.Y(n_4778)
);

CKINVDCx20_ASAP7_75t_R g4779 ( 
.A(n_4248),
.Y(n_4779)
);

INVxp33_ASAP7_75t_L g4780 ( 
.A(n_4559),
.Y(n_4780)
);

CKINVDCx20_ASAP7_75t_R g4781 ( 
.A(n_4253),
.Y(n_4781)
);

INVx3_ASAP7_75t_L g4782 ( 
.A(n_4443),
.Y(n_4782)
);

INVx1_ASAP7_75t_L g4783 ( 
.A(n_4549),
.Y(n_4783)
);

INVx1_ASAP7_75t_L g4784 ( 
.A(n_4552),
.Y(n_4784)
);

CKINVDCx5p33_ASAP7_75t_R g4785 ( 
.A(n_4492),
.Y(n_4785)
);

CKINVDCx20_ASAP7_75t_R g4786 ( 
.A(n_4256),
.Y(n_4786)
);

INVxp67_ASAP7_75t_SL g4787 ( 
.A(n_4513),
.Y(n_4787)
);

INVx1_ASAP7_75t_L g4788 ( 
.A(n_4558),
.Y(n_4788)
);

INVx1_ASAP7_75t_L g4789 ( 
.A(n_4558),
.Y(n_4789)
);

CKINVDCx5p33_ASAP7_75t_R g4790 ( 
.A(n_4498),
.Y(n_4790)
);

CKINVDCx5p33_ASAP7_75t_R g4791 ( 
.A(n_4500),
.Y(n_4791)
);

CKINVDCx5p33_ASAP7_75t_R g4792 ( 
.A(n_4504),
.Y(n_4792)
);

CKINVDCx5p33_ASAP7_75t_R g4793 ( 
.A(n_4518),
.Y(n_4793)
);

INVx1_ASAP7_75t_L g4794 ( 
.A(n_4558),
.Y(n_4794)
);

CKINVDCx5p33_ASAP7_75t_R g4795 ( 
.A(n_4538),
.Y(n_4795)
);

CKINVDCx20_ASAP7_75t_R g4796 ( 
.A(n_4592),
.Y(n_4796)
);

INVxp67_ASAP7_75t_L g4797 ( 
.A(n_4572),
.Y(n_4797)
);

BUFx3_ASAP7_75t_L g4798 ( 
.A(n_4315),
.Y(n_4798)
);

INVx1_ASAP7_75t_L g4799 ( 
.A(n_4218),
.Y(n_4799)
);

INVx1_ASAP7_75t_L g4800 ( 
.A(n_4219),
.Y(n_4800)
);

CKINVDCx5p33_ASAP7_75t_R g4801 ( 
.A(n_4539),
.Y(n_4801)
);

CKINVDCx20_ASAP7_75t_R g4802 ( 
.A(n_4603),
.Y(n_4802)
);

HB1xp67_ASAP7_75t_L g4803 ( 
.A(n_4545),
.Y(n_4803)
);

CKINVDCx20_ASAP7_75t_R g4804 ( 
.A(n_4612),
.Y(n_4804)
);

INVx1_ASAP7_75t_L g4805 ( 
.A(n_4224),
.Y(n_4805)
);

CKINVDCx5p33_ASAP7_75t_R g4806 ( 
.A(n_4550),
.Y(n_4806)
);

CKINVDCx20_ASAP7_75t_R g4807 ( 
.A(n_4571),
.Y(n_4807)
);

INVx1_ASAP7_75t_L g4808 ( 
.A(n_4225),
.Y(n_4808)
);

CKINVDCx5p33_ASAP7_75t_R g4809 ( 
.A(n_4579),
.Y(n_4809)
);

CKINVDCx5p33_ASAP7_75t_R g4810 ( 
.A(n_4584),
.Y(n_4810)
);

HB1xp67_ASAP7_75t_L g4811 ( 
.A(n_4588),
.Y(n_4811)
);

INVx1_ASAP7_75t_L g4812 ( 
.A(n_4227),
.Y(n_4812)
);

CKINVDCx5p33_ASAP7_75t_R g4813 ( 
.A(n_4605),
.Y(n_4813)
);

INVx1_ASAP7_75t_L g4814 ( 
.A(n_4228),
.Y(n_4814)
);

CKINVDCx5p33_ASAP7_75t_R g4815 ( 
.A(n_4616),
.Y(n_4815)
);

CKINVDCx5p33_ASAP7_75t_R g4816 ( 
.A(n_4618),
.Y(n_4816)
);

BUFx6f_ASAP7_75t_SL g4817 ( 
.A(n_4343),
.Y(n_4817)
);

CKINVDCx5p33_ASAP7_75t_R g4818 ( 
.A(n_4619),
.Y(n_4818)
);

NOR2xp33_ASAP7_75t_L g4819 ( 
.A(n_4223),
.B(n_3538),
.Y(n_4819)
);

INVx1_ASAP7_75t_L g4820 ( 
.A(n_4231),
.Y(n_4820)
);

CKINVDCx5p33_ASAP7_75t_R g4821 ( 
.A(n_4561),
.Y(n_4821)
);

INVx1_ASAP7_75t_L g4822 ( 
.A(n_4232),
.Y(n_4822)
);

CKINVDCx5p33_ASAP7_75t_R g4823 ( 
.A(n_4575),
.Y(n_4823)
);

CKINVDCx5p33_ASAP7_75t_R g4824 ( 
.A(n_4604),
.Y(n_4824)
);

CKINVDCx20_ASAP7_75t_R g4825 ( 
.A(n_4356),
.Y(n_4825)
);

CKINVDCx20_ASAP7_75t_R g4826 ( 
.A(n_4371),
.Y(n_4826)
);

INVx1_ASAP7_75t_L g4827 ( 
.A(n_4233),
.Y(n_4827)
);

INVx1_ASAP7_75t_L g4828 ( 
.A(n_4236),
.Y(n_4828)
);

CKINVDCx5p33_ASAP7_75t_R g4829 ( 
.A(n_4617),
.Y(n_4829)
);

INVx1_ASAP7_75t_L g4830 ( 
.A(n_4237),
.Y(n_4830)
);

CKINVDCx20_ASAP7_75t_R g4831 ( 
.A(n_4396),
.Y(n_4831)
);

CKINVDCx5p33_ASAP7_75t_R g4832 ( 
.A(n_4406),
.Y(n_4832)
);

BUFx3_ASAP7_75t_L g4833 ( 
.A(n_4335),
.Y(n_4833)
);

INVx1_ASAP7_75t_L g4834 ( 
.A(n_4238),
.Y(n_4834)
);

INVxp67_ASAP7_75t_L g4835 ( 
.A(n_4520),
.Y(n_4835)
);

NOR2xp33_ASAP7_75t_L g4836 ( 
.A(n_4303),
.B(n_3541),
.Y(n_4836)
);

CKINVDCx5p33_ASAP7_75t_R g4837 ( 
.A(n_4418),
.Y(n_4837)
);

CKINVDCx20_ASAP7_75t_R g4838 ( 
.A(n_4522),
.Y(n_4838)
);

INVx1_ASAP7_75t_L g4839 ( 
.A(n_4239),
.Y(n_4839)
);

INVx1_ASAP7_75t_L g4840 ( 
.A(n_4241),
.Y(n_4840)
);

CKINVDCx20_ASAP7_75t_R g4841 ( 
.A(n_4532),
.Y(n_4841)
);

XOR2xp5_ASAP7_75t_L g4842 ( 
.A(n_4330),
.B(n_2861),
.Y(n_4842)
);

CKINVDCx5p33_ASAP7_75t_R g4843 ( 
.A(n_4229),
.Y(n_4843)
);

CKINVDCx20_ASAP7_75t_R g4844 ( 
.A(n_4322),
.Y(n_4844)
);

CKINVDCx5p33_ASAP7_75t_R g4845 ( 
.A(n_4309),
.Y(n_4845)
);

CKINVDCx5p33_ASAP7_75t_R g4846 ( 
.A(n_4358),
.Y(n_4846)
);

CKINVDCx20_ASAP7_75t_R g4847 ( 
.A(n_4336),
.Y(n_4847)
);

INVx1_ASAP7_75t_L g4848 ( 
.A(n_4243),
.Y(n_4848)
);

CKINVDCx20_ASAP7_75t_R g4849 ( 
.A(n_4475),
.Y(n_4849)
);

CKINVDCx16_ASAP7_75t_R g4850 ( 
.A(n_4437),
.Y(n_4850)
);

INVx1_ASAP7_75t_L g4851 ( 
.A(n_4245),
.Y(n_4851)
);

CKINVDCx20_ASAP7_75t_R g4852 ( 
.A(n_4481),
.Y(n_4852)
);

CKINVDCx5p33_ASAP7_75t_R g4853 ( 
.A(n_4350),
.Y(n_4853)
);

CKINVDCx20_ASAP7_75t_R g4854 ( 
.A(n_4344),
.Y(n_4854)
);

CKINVDCx20_ASAP7_75t_R g4855 ( 
.A(n_4375),
.Y(n_4855)
);

INVx1_ASAP7_75t_L g4856 ( 
.A(n_4249),
.Y(n_4856)
);

INVx1_ASAP7_75t_L g4857 ( 
.A(n_4250),
.Y(n_4857)
);

CKINVDCx5p33_ASAP7_75t_R g4858 ( 
.A(n_4203),
.Y(n_4858)
);

INVx1_ASAP7_75t_L g4859 ( 
.A(n_4251),
.Y(n_4859)
);

NOR2xp67_ASAP7_75t_L g4860 ( 
.A(n_4563),
.B(n_3409),
.Y(n_4860)
);

CKINVDCx20_ASAP7_75t_R g4861 ( 
.A(n_4424),
.Y(n_4861)
);

NOR2xp33_ASAP7_75t_L g4862 ( 
.A(n_4214),
.B(n_3557),
.Y(n_4862)
);

BUFx3_ASAP7_75t_L g4863 ( 
.A(n_4378),
.Y(n_4863)
);

CKINVDCx5p33_ASAP7_75t_R g4864 ( 
.A(n_4506),
.Y(n_4864)
);

HB1xp67_ASAP7_75t_L g4865 ( 
.A(n_4565),
.Y(n_4865)
);

CKINVDCx5p33_ASAP7_75t_R g4866 ( 
.A(n_4527),
.Y(n_4866)
);

INVx1_ASAP7_75t_L g4867 ( 
.A(n_4255),
.Y(n_4867)
);

INVxp67_ASAP7_75t_L g4868 ( 
.A(n_4517),
.Y(n_4868)
);

CKINVDCx5p33_ASAP7_75t_R g4869 ( 
.A(n_4553),
.Y(n_4869)
);

CKINVDCx20_ASAP7_75t_R g4870 ( 
.A(n_4230),
.Y(n_4870)
);

CKINVDCx20_ASAP7_75t_R g4871 ( 
.A(n_4280),
.Y(n_4871)
);

CKINVDCx5p33_ASAP7_75t_R g4872 ( 
.A(n_4302),
.Y(n_4872)
);

INVx1_ASAP7_75t_L g4873 ( 
.A(n_4257),
.Y(n_4873)
);

CKINVDCx5p33_ASAP7_75t_R g4874 ( 
.A(n_4337),
.Y(n_4874)
);

CKINVDCx20_ASAP7_75t_R g4875 ( 
.A(n_4442),
.Y(n_4875)
);

CKINVDCx5p33_ASAP7_75t_R g4876 ( 
.A(n_4455),
.Y(n_4876)
);

INVx1_ASAP7_75t_L g4877 ( 
.A(n_4258),
.Y(n_4877)
);

CKINVDCx5p33_ASAP7_75t_R g4878 ( 
.A(n_4213),
.Y(n_4878)
);

CKINVDCx14_ASAP7_75t_R g4879 ( 
.A(n_4613),
.Y(n_4879)
);

NOR2xp33_ASAP7_75t_L g4880 ( 
.A(n_4328),
.B(n_3573),
.Y(n_4880)
);

INVx1_ASAP7_75t_L g4881 ( 
.A(n_4260),
.Y(n_4881)
);

CKINVDCx20_ASAP7_75t_R g4882 ( 
.A(n_4574),
.Y(n_4882)
);

CKINVDCx5p33_ASAP7_75t_R g4883 ( 
.A(n_4576),
.Y(n_4883)
);

NOR2xp33_ASAP7_75t_L g4884 ( 
.A(n_4382),
.B(n_3583),
.Y(n_4884)
);

INVx1_ASAP7_75t_L g4885 ( 
.A(n_4262),
.Y(n_4885)
);

NOR2xp67_ASAP7_75t_L g4886 ( 
.A(n_4264),
.B(n_3416),
.Y(n_4886)
);

INVx1_ASAP7_75t_SL g4887 ( 
.A(n_4416),
.Y(n_4887)
);

CKINVDCx5p33_ASAP7_75t_R g4888 ( 
.A(n_4554),
.Y(n_4888)
);

CKINVDCx20_ASAP7_75t_R g4889 ( 
.A(n_4555),
.Y(n_4889)
);

CKINVDCx5p33_ASAP7_75t_R g4890 ( 
.A(n_4556),
.Y(n_4890)
);

CKINVDCx20_ASAP7_75t_R g4891 ( 
.A(n_4557),
.Y(n_4891)
);

NOR2xp33_ASAP7_75t_L g4892 ( 
.A(n_4435),
.B(n_3595),
.Y(n_4892)
);

CKINVDCx20_ASAP7_75t_R g4893 ( 
.A(n_4560),
.Y(n_4893)
);

INVx1_ASAP7_75t_L g4894 ( 
.A(n_4265),
.Y(n_4894)
);

CKINVDCx20_ASAP7_75t_R g4895 ( 
.A(n_4562),
.Y(n_4895)
);

INVx1_ASAP7_75t_L g4896 ( 
.A(n_4267),
.Y(n_4896)
);

INVx1_ASAP7_75t_L g4897 ( 
.A(n_4272),
.Y(n_4897)
);

INVx1_ASAP7_75t_L g4898 ( 
.A(n_4275),
.Y(n_4898)
);

CKINVDCx5p33_ASAP7_75t_R g4899 ( 
.A(n_4564),
.Y(n_4899)
);

CKINVDCx20_ASAP7_75t_R g4900 ( 
.A(n_4566),
.Y(n_4900)
);

CKINVDCx16_ASAP7_75t_R g4901 ( 
.A(n_4568),
.Y(n_4901)
);

CKINVDCx5p33_ASAP7_75t_R g4902 ( 
.A(n_4569),
.Y(n_4902)
);

CKINVDCx20_ASAP7_75t_R g4903 ( 
.A(n_4570),
.Y(n_4903)
);

CKINVDCx20_ASAP7_75t_R g4904 ( 
.A(n_4573),
.Y(n_4904)
);

HB1xp67_ASAP7_75t_L g4905 ( 
.A(n_4577),
.Y(n_4905)
);

CKINVDCx14_ASAP7_75t_R g4906 ( 
.A(n_4484),
.Y(n_4906)
);

INVx1_ASAP7_75t_L g4907 ( 
.A(n_4276),
.Y(n_4907)
);

CKINVDCx16_ASAP7_75t_R g4908 ( 
.A(n_4578),
.Y(n_4908)
);

CKINVDCx20_ASAP7_75t_R g4909 ( 
.A(n_4580),
.Y(n_4909)
);

INVxp33_ASAP7_75t_L g4910 ( 
.A(n_4583),
.Y(n_4910)
);

INVx1_ASAP7_75t_L g4911 ( 
.A(n_4278),
.Y(n_4911)
);

INVxp67_ASAP7_75t_SL g4912 ( 
.A(n_4582),
.Y(n_4912)
);

CKINVDCx5p33_ASAP7_75t_R g4913 ( 
.A(n_4585),
.Y(n_4913)
);

CKINVDCx20_ASAP7_75t_R g4914 ( 
.A(n_4586),
.Y(n_4914)
);

CKINVDCx20_ASAP7_75t_R g4915 ( 
.A(n_4587),
.Y(n_4915)
);

CKINVDCx5p33_ASAP7_75t_R g4916 ( 
.A(n_4201),
.Y(n_4916)
);

BUFx6f_ASAP7_75t_L g4917 ( 
.A(n_4611),
.Y(n_4917)
);

BUFx6f_ASAP7_75t_L g4918 ( 
.A(n_4611),
.Y(n_4918)
);

CKINVDCx20_ASAP7_75t_R g4919 ( 
.A(n_4608),
.Y(n_4919)
);

INVx1_ASAP7_75t_L g4920 ( 
.A(n_4284),
.Y(n_4920)
);

CKINVDCx20_ASAP7_75t_R g4921 ( 
.A(n_4201),
.Y(n_4921)
);

NOR2xp33_ASAP7_75t_L g4922 ( 
.A(n_4536),
.B(n_3602),
.Y(n_4922)
);

INVx1_ASAP7_75t_L g4923 ( 
.A(n_4285),
.Y(n_4923)
);

INVxp67_ASAP7_75t_L g4924 ( 
.A(n_4567),
.Y(n_4924)
);

INVx1_ASAP7_75t_L g4925 ( 
.A(n_4287),
.Y(n_4925)
);

INVx1_ASAP7_75t_L g4926 ( 
.A(n_4288),
.Y(n_4926)
);

INVx1_ASAP7_75t_L g4927 ( 
.A(n_4294),
.Y(n_4927)
);

INVx1_ASAP7_75t_L g4928 ( 
.A(n_4295),
.Y(n_4928)
);

INVx3_ASAP7_75t_L g4929 ( 
.A(n_4611),
.Y(n_4929)
);

INVx1_ASAP7_75t_L g4930 ( 
.A(n_4296),
.Y(n_4930)
);

INVx1_ASAP7_75t_L g4931 ( 
.A(n_4297),
.Y(n_4931)
);

NAND2xp5_ASAP7_75t_L g4932 ( 
.A(n_4201),
.B(n_3598),
.Y(n_4932)
);

XNOR2xp5_ASAP7_75t_L g4933 ( 
.A(n_4345),
.B(n_3012),
.Y(n_4933)
);

INVxp33_ASAP7_75t_SL g4934 ( 
.A(n_4467),
.Y(n_4934)
);

CKINVDCx20_ASAP7_75t_R g4935 ( 
.A(n_4201),
.Y(n_4935)
);

INVx1_ASAP7_75t_L g4936 ( 
.A(n_4300),
.Y(n_4936)
);

NAND2xp5_ASAP7_75t_L g4937 ( 
.A(n_4201),
.B(n_4301),
.Y(n_4937)
);

INVx1_ASAP7_75t_L g4938 ( 
.A(n_4304),
.Y(n_4938)
);

INVx1_ASAP7_75t_L g4939 ( 
.A(n_4307),
.Y(n_4939)
);

HB1xp67_ASAP7_75t_L g4940 ( 
.A(n_4363),
.Y(n_4940)
);

INVx1_ASAP7_75t_L g4941 ( 
.A(n_4308),
.Y(n_4941)
);

INVx1_ASAP7_75t_L g4942 ( 
.A(n_4310),
.Y(n_4942)
);

INVx2_ASAP7_75t_L g4943 ( 
.A(n_4254),
.Y(n_4943)
);

INVx1_ASAP7_75t_L g4944 ( 
.A(n_4312),
.Y(n_4944)
);

INVx1_ASAP7_75t_SL g4945 ( 
.A(n_4464),
.Y(n_4945)
);

CKINVDCx16_ASAP7_75t_R g4946 ( 
.A(n_4364),
.Y(n_4946)
);

NOR2xp67_ASAP7_75t_L g4947 ( 
.A(n_4313),
.B(n_3743),
.Y(n_4947)
);

CKINVDCx20_ASAP7_75t_R g4948 ( 
.A(n_4589),
.Y(n_4948)
);

CKINVDCx5p33_ASAP7_75t_R g4949 ( 
.A(n_4281),
.Y(n_4949)
);

CKINVDCx20_ASAP7_75t_R g4950 ( 
.A(n_4593),
.Y(n_4950)
);

INVx1_ASAP7_75t_L g4951 ( 
.A(n_4314),
.Y(n_4951)
);

CKINVDCx5p33_ASAP7_75t_R g4952 ( 
.A(n_4291),
.Y(n_4952)
);

CKINVDCx20_ASAP7_75t_R g4953 ( 
.A(n_4594),
.Y(n_4953)
);

INVxp33_ASAP7_75t_SL g4954 ( 
.A(n_4551),
.Y(n_4954)
);

INVxp67_ASAP7_75t_L g4955 ( 
.A(n_4366),
.Y(n_4955)
);

BUFx3_ASAP7_75t_L g4956 ( 
.A(n_4316),
.Y(n_4956)
);

INVx1_ASAP7_75t_L g4957 ( 
.A(n_4317),
.Y(n_4957)
);

CKINVDCx5p33_ASAP7_75t_R g4958 ( 
.A(n_4293),
.Y(n_4958)
);

CKINVDCx5p33_ASAP7_75t_R g4959 ( 
.A(n_4324),
.Y(n_4959)
);

CKINVDCx5p33_ASAP7_75t_R g4960 ( 
.A(n_4334),
.Y(n_4960)
);

INVx1_ASAP7_75t_L g4961 ( 
.A(n_4319),
.Y(n_4961)
);

INVx1_ASAP7_75t_L g4962 ( 
.A(n_4321),
.Y(n_4962)
);

INVx1_ASAP7_75t_L g4963 ( 
.A(n_4323),
.Y(n_4963)
);

CKINVDCx5p33_ASAP7_75t_R g4964 ( 
.A(n_4354),
.Y(n_4964)
);

INVx1_ASAP7_75t_SL g4965 ( 
.A(n_4595),
.Y(n_4965)
);

CKINVDCx5p33_ASAP7_75t_R g4966 ( 
.A(n_4355),
.Y(n_4966)
);

CKINVDCx5p33_ASAP7_75t_R g4967 ( 
.A(n_4357),
.Y(n_4967)
);

NOR2xp33_ASAP7_75t_L g4968 ( 
.A(n_4208),
.B(n_3610),
.Y(n_4968)
);

INVx1_ASAP7_75t_L g4969 ( 
.A(n_4325),
.Y(n_4969)
);

NOR2xp33_ASAP7_75t_R g4970 ( 
.A(n_4327),
.B(n_2815),
.Y(n_4970)
);

CKINVDCx5p33_ASAP7_75t_R g4971 ( 
.A(n_4362),
.Y(n_4971)
);

CKINVDCx20_ASAP7_75t_R g4972 ( 
.A(n_4596),
.Y(n_4972)
);

INVx1_ASAP7_75t_L g4973 ( 
.A(n_4329),
.Y(n_4973)
);

INVx1_ASAP7_75t_L g4974 ( 
.A(n_4338),
.Y(n_4974)
);

INVxp33_ASAP7_75t_SL g4975 ( 
.A(n_4306),
.Y(n_4975)
);

INVxp67_ASAP7_75t_SL g4976 ( 
.A(n_4326),
.Y(n_4976)
);

INVx1_ASAP7_75t_L g4977 ( 
.A(n_4342),
.Y(n_4977)
);

NAND2xp5_ASAP7_75t_L g4978 ( 
.A(n_4346),
.B(n_3839),
.Y(n_4978)
);

INVx2_ASAP7_75t_L g4979 ( 
.A(n_4367),
.Y(n_4979)
);

INVx1_ASAP7_75t_L g4980 ( 
.A(n_4347),
.Y(n_4980)
);

CKINVDCx5p33_ASAP7_75t_R g4981 ( 
.A(n_4348),
.Y(n_4981)
);

BUFx10_ASAP7_75t_L g4982 ( 
.A(n_4369),
.Y(n_4982)
);

INVx1_ASAP7_75t_L g4983 ( 
.A(n_4349),
.Y(n_4983)
);

AND2x2_ASAP7_75t_L g4984 ( 
.A(n_4381),
.B(n_2816),
.Y(n_4984)
);

HB1xp67_ASAP7_75t_L g4985 ( 
.A(n_4370),
.Y(n_4985)
);

NOR2xp67_ASAP7_75t_L g4986 ( 
.A(n_4353),
.B(n_3899),
.Y(n_4986)
);

INVx1_ASAP7_75t_L g4987 ( 
.A(n_4360),
.Y(n_4987)
);

CKINVDCx20_ASAP7_75t_R g4988 ( 
.A(n_4597),
.Y(n_4988)
);

CKINVDCx20_ASAP7_75t_R g4989 ( 
.A(n_4598),
.Y(n_4989)
);

CKINVDCx5p33_ASAP7_75t_R g4990 ( 
.A(n_4361),
.Y(n_4990)
);

CKINVDCx20_ASAP7_75t_R g4991 ( 
.A(n_4599),
.Y(n_4991)
);

INVx1_ASAP7_75t_L g4992 ( 
.A(n_4600),
.Y(n_4992)
);

INVx1_ASAP7_75t_L g4993 ( 
.A(n_4601),
.Y(n_4993)
);

CKINVDCx5p33_ASAP7_75t_R g4994 ( 
.A(n_4590),
.Y(n_4994)
);

INVx1_ASAP7_75t_L g4995 ( 
.A(n_4606),
.Y(n_4995)
);

INVx1_ASAP7_75t_L g4996 ( 
.A(n_4607),
.Y(n_4996)
);

INVx1_ASAP7_75t_L g4997 ( 
.A(n_4609),
.Y(n_4997)
);

INVxp67_ASAP7_75t_L g4998 ( 
.A(n_4372),
.Y(n_4998)
);

NOR2xp33_ASAP7_75t_L g4999 ( 
.A(n_4610),
.B(n_3619),
.Y(n_4999)
);

CKINVDCx5p33_ASAP7_75t_R g5000 ( 
.A(n_4602),
.Y(n_5000)
);

CKINVDCx20_ASAP7_75t_R g5001 ( 
.A(n_4614),
.Y(n_5001)
);

INVx1_ASAP7_75t_L g5002 ( 
.A(n_4615),
.Y(n_5002)
);

CKINVDCx5p33_ASAP7_75t_R g5003 ( 
.A(n_4397),
.Y(n_5003)
);

INVxp67_ASAP7_75t_SL g5004 ( 
.A(n_4620),
.Y(n_5004)
);

CKINVDCx20_ASAP7_75t_R g5005 ( 
.A(n_4377),
.Y(n_5005)
);

CKINVDCx20_ASAP7_75t_R g5006 ( 
.A(n_4379),
.Y(n_5006)
);

INVx1_ASAP7_75t_L g5007 ( 
.A(n_4380),
.Y(n_5007)
);

INVx1_ASAP7_75t_L g5008 ( 
.A(n_4384),
.Y(n_5008)
);

INVx1_ASAP7_75t_L g5009 ( 
.A(n_4385),
.Y(n_5009)
);

CKINVDCx5p33_ASAP7_75t_R g5010 ( 
.A(n_4419),
.Y(n_5010)
);

CKINVDCx5p33_ASAP7_75t_R g5011 ( 
.A(n_4425),
.Y(n_5011)
);

INVx2_ASAP7_75t_L g5012 ( 
.A(n_4433),
.Y(n_5012)
);

INVx1_ASAP7_75t_L g5013 ( 
.A(n_4386),
.Y(n_5013)
);

INVxp67_ASAP7_75t_SL g5014 ( 
.A(n_4447),
.Y(n_5014)
);

CKINVDCx5p33_ASAP7_75t_R g5015 ( 
.A(n_4448),
.Y(n_5015)
);

INVx1_ASAP7_75t_L g5016 ( 
.A(n_4390),
.Y(n_5016)
);

CKINVDCx20_ASAP7_75t_R g5017 ( 
.A(n_4391),
.Y(n_5017)
);

INVx1_ASAP7_75t_L g5018 ( 
.A(n_4393),
.Y(n_5018)
);

INVx1_ASAP7_75t_SL g5019 ( 
.A(n_4394),
.Y(n_5019)
);

NOR2xp67_ASAP7_75t_L g5020 ( 
.A(n_4487),
.B(n_3921),
.Y(n_5020)
);

CKINVDCx20_ASAP7_75t_R g5021 ( 
.A(n_4398),
.Y(n_5021)
);

INVxp67_ASAP7_75t_SL g5022 ( 
.A(n_4452),
.Y(n_5022)
);

NOR2xp67_ASAP7_75t_L g5023 ( 
.A(n_4488),
.B(n_3977),
.Y(n_5023)
);

NOR2xp67_ASAP7_75t_L g5024 ( 
.A(n_4489),
.B(n_4064),
.Y(n_5024)
);

NOR2xp33_ASAP7_75t_L g5025 ( 
.A(n_4401),
.B(n_3620),
.Y(n_5025)
);

INVxp67_ASAP7_75t_L g5026 ( 
.A(n_4402),
.Y(n_5026)
);

INVx1_ASAP7_75t_L g5027 ( 
.A(n_4403),
.Y(n_5027)
);

CKINVDCx20_ASAP7_75t_R g5028 ( 
.A(n_4405),
.Y(n_5028)
);

NOR2xp33_ASAP7_75t_L g5029 ( 
.A(n_4408),
.B(n_3668),
.Y(n_5029)
);

CKINVDCx5p33_ASAP7_75t_R g5030 ( 
.A(n_4412),
.Y(n_5030)
);

INVxp67_ASAP7_75t_SL g5031 ( 
.A(n_4413),
.Y(n_5031)
);

INVxp67_ASAP7_75t_SL g5032 ( 
.A(n_4414),
.Y(n_5032)
);

INVx1_ASAP7_75t_L g5033 ( 
.A(n_4415),
.Y(n_5033)
);

CKINVDCx5p33_ASAP7_75t_R g5034 ( 
.A(n_4420),
.Y(n_5034)
);

INVxp67_ASAP7_75t_SL g5035 ( 
.A(n_4421),
.Y(n_5035)
);

INVx1_ASAP7_75t_L g5036 ( 
.A(n_4422),
.Y(n_5036)
);

INVxp67_ASAP7_75t_SL g5037 ( 
.A(n_4423),
.Y(n_5037)
);

CKINVDCx14_ASAP7_75t_R g5038 ( 
.A(n_4426),
.Y(n_5038)
);

INVx1_ASAP7_75t_L g5039 ( 
.A(n_4427),
.Y(n_5039)
);

INVxp67_ASAP7_75t_L g5040 ( 
.A(n_4428),
.Y(n_5040)
);

INVx1_ASAP7_75t_L g5041 ( 
.A(n_4431),
.Y(n_5041)
);

NAND2xp33_ASAP7_75t_R g5042 ( 
.A(n_4432),
.B(n_3676),
.Y(n_5042)
);

NOR2xp33_ASAP7_75t_L g5043 ( 
.A(n_4436),
.B(n_3681),
.Y(n_5043)
);

INVx1_ASAP7_75t_L g5044 ( 
.A(n_4440),
.Y(n_5044)
);

INVx1_ASAP7_75t_L g5045 ( 
.A(n_4441),
.Y(n_5045)
);

INVx1_ASAP7_75t_L g5046 ( 
.A(n_4449),
.Y(n_5046)
);

INVx1_ASAP7_75t_L g5047 ( 
.A(n_4450),
.Y(n_5047)
);

CKINVDCx5p33_ASAP7_75t_R g5048 ( 
.A(n_4451),
.Y(n_5048)
);

CKINVDCx5p33_ASAP7_75t_R g5049 ( 
.A(n_4454),
.Y(n_5049)
);

CKINVDCx5p33_ASAP7_75t_R g5050 ( 
.A(n_4457),
.Y(n_5050)
);

HB1xp67_ASAP7_75t_L g5051 ( 
.A(n_4459),
.Y(n_5051)
);

NOR2xp33_ASAP7_75t_L g5052 ( 
.A(n_4491),
.B(n_3690),
.Y(n_5052)
);

INVxp33_ASAP7_75t_L g5053 ( 
.A(n_4494),
.Y(n_5053)
);

CKINVDCx20_ASAP7_75t_R g5054 ( 
.A(n_4495),
.Y(n_5054)
);

BUFx6f_ASAP7_75t_L g5055 ( 
.A(n_4497),
.Y(n_5055)
);

CKINVDCx5p33_ASAP7_75t_R g5056 ( 
.A(n_4499),
.Y(n_5056)
);

INVx1_ASAP7_75t_L g5057 ( 
.A(n_4501),
.Y(n_5057)
);

INVx1_ASAP7_75t_L g5058 ( 
.A(n_4502),
.Y(n_5058)
);

CKINVDCx5p33_ASAP7_75t_R g5059 ( 
.A(n_4202),
.Y(n_5059)
);

INVxp67_ASAP7_75t_SL g5060 ( 
.A(n_4496),
.Y(n_5060)
);

CKINVDCx5p33_ASAP7_75t_R g5061 ( 
.A(n_4202),
.Y(n_5061)
);

CKINVDCx5p33_ASAP7_75t_R g5062 ( 
.A(n_4202),
.Y(n_5062)
);

CKINVDCx5p33_ASAP7_75t_R g5063 ( 
.A(n_4202),
.Y(n_5063)
);

CKINVDCx20_ASAP7_75t_R g5064 ( 
.A(n_4331),
.Y(n_5064)
);

INVx1_ASAP7_75t_L g5065 ( 
.A(n_4496),
.Y(n_5065)
);

CKINVDCx5p33_ASAP7_75t_R g5066 ( 
.A(n_4202),
.Y(n_5066)
);

INVx1_ASAP7_75t_L g5067 ( 
.A(n_4496),
.Y(n_5067)
);

BUFx3_ASAP7_75t_L g5068 ( 
.A(n_4217),
.Y(n_5068)
);

INVx1_ASAP7_75t_L g5069 ( 
.A(n_4496),
.Y(n_5069)
);

CKINVDCx5p33_ASAP7_75t_R g5070 ( 
.A(n_4202),
.Y(n_5070)
);

INVxp33_ASAP7_75t_SL g5071 ( 
.A(n_4202),
.Y(n_5071)
);

INVxp67_ASAP7_75t_L g5072 ( 
.A(n_4270),
.Y(n_5072)
);

INVx2_ASAP7_75t_L g5073 ( 
.A(n_4503),
.Y(n_5073)
);

CKINVDCx5p33_ASAP7_75t_R g5074 ( 
.A(n_4202),
.Y(n_5074)
);

NOR2xp33_ASAP7_75t_R g5075 ( 
.A(n_4311),
.B(n_2817),
.Y(n_5075)
);

INVx1_ASAP7_75t_L g5076 ( 
.A(n_4496),
.Y(n_5076)
);

CKINVDCx5p33_ASAP7_75t_R g5077 ( 
.A(n_4202),
.Y(n_5077)
);

BUFx6f_ASAP7_75t_L g5078 ( 
.A(n_4261),
.Y(n_5078)
);

CKINVDCx5p33_ASAP7_75t_R g5079 ( 
.A(n_4202),
.Y(n_5079)
);

INVx1_ASAP7_75t_L g5080 ( 
.A(n_4496),
.Y(n_5080)
);

CKINVDCx20_ASAP7_75t_R g5081 ( 
.A(n_4331),
.Y(n_5081)
);

INVx1_ASAP7_75t_L g5082 ( 
.A(n_4496),
.Y(n_5082)
);

CKINVDCx5p33_ASAP7_75t_R g5083 ( 
.A(n_4202),
.Y(n_5083)
);

INVx1_ASAP7_75t_L g5084 ( 
.A(n_4496),
.Y(n_5084)
);

CKINVDCx5p33_ASAP7_75t_R g5085 ( 
.A(n_4202),
.Y(n_5085)
);

INVx1_ASAP7_75t_L g5086 ( 
.A(n_4496),
.Y(n_5086)
);

INVx1_ASAP7_75t_L g5087 ( 
.A(n_4496),
.Y(n_5087)
);

INVx1_ASAP7_75t_L g5088 ( 
.A(n_4496),
.Y(n_5088)
);

CKINVDCx20_ASAP7_75t_R g5089 ( 
.A(n_4331),
.Y(n_5089)
);

INVx1_ASAP7_75t_L g5090 ( 
.A(n_4496),
.Y(n_5090)
);

CKINVDCx5p33_ASAP7_75t_R g5091 ( 
.A(n_4202),
.Y(n_5091)
);

INVx2_ASAP7_75t_L g5092 ( 
.A(n_4503),
.Y(n_5092)
);

INVx1_ASAP7_75t_L g5093 ( 
.A(n_4496),
.Y(n_5093)
);

INVx1_ASAP7_75t_L g5094 ( 
.A(n_4496),
.Y(n_5094)
);

CKINVDCx5p33_ASAP7_75t_R g5095 ( 
.A(n_4202),
.Y(n_5095)
);

CKINVDCx20_ASAP7_75t_R g5096 ( 
.A(n_4331),
.Y(n_5096)
);

INVx1_ASAP7_75t_L g5097 ( 
.A(n_4496),
.Y(n_5097)
);

INVx1_ASAP7_75t_L g5098 ( 
.A(n_4496),
.Y(n_5098)
);

NOR2xp33_ASAP7_75t_L g5099 ( 
.A(n_4463),
.B(n_3693),
.Y(n_5099)
);

CKINVDCx5p33_ASAP7_75t_R g5100 ( 
.A(n_4202),
.Y(n_5100)
);

INVx1_ASAP7_75t_L g5101 ( 
.A(n_4496),
.Y(n_5101)
);

HB1xp67_ASAP7_75t_L g5102 ( 
.A(n_4263),
.Y(n_5102)
);

CKINVDCx5p33_ASAP7_75t_R g5103 ( 
.A(n_4202),
.Y(n_5103)
);

INVx1_ASAP7_75t_L g5104 ( 
.A(n_4496),
.Y(n_5104)
);

HB1xp67_ASAP7_75t_L g5105 ( 
.A(n_4263),
.Y(n_5105)
);

CKINVDCx5p33_ASAP7_75t_R g5106 ( 
.A(n_4202),
.Y(n_5106)
);

CKINVDCx20_ASAP7_75t_R g5107 ( 
.A(n_4331),
.Y(n_5107)
);

INVx1_ASAP7_75t_L g5108 ( 
.A(n_4496),
.Y(n_5108)
);

INVx1_ASAP7_75t_L g5109 ( 
.A(n_4496),
.Y(n_5109)
);

INVx1_ASAP7_75t_L g5110 ( 
.A(n_4496),
.Y(n_5110)
);

INVx2_ASAP7_75t_L g5111 ( 
.A(n_4503),
.Y(n_5111)
);

INVx1_ASAP7_75t_L g5112 ( 
.A(n_4496),
.Y(n_5112)
);

CKINVDCx5p33_ASAP7_75t_R g5113 ( 
.A(n_4202),
.Y(n_5113)
);

CKINVDCx5p33_ASAP7_75t_R g5114 ( 
.A(n_4202),
.Y(n_5114)
);

INVx1_ASAP7_75t_L g5115 ( 
.A(n_4496),
.Y(n_5115)
);

HB1xp67_ASAP7_75t_L g5116 ( 
.A(n_4263),
.Y(n_5116)
);

CKINVDCx20_ASAP7_75t_R g5117 ( 
.A(n_4331),
.Y(n_5117)
);

HB1xp67_ASAP7_75t_L g5118 ( 
.A(n_4263),
.Y(n_5118)
);

CKINVDCx5p33_ASAP7_75t_R g5119 ( 
.A(n_4202),
.Y(n_5119)
);

INVx1_ASAP7_75t_L g5120 ( 
.A(n_4496),
.Y(n_5120)
);

CKINVDCx20_ASAP7_75t_R g5121 ( 
.A(n_4331),
.Y(n_5121)
);

INVx2_ASAP7_75t_L g5122 ( 
.A(n_4929),
.Y(n_5122)
);

AND2x2_ASAP7_75t_L g5123 ( 
.A(n_4910),
.B(n_3305),
.Y(n_5123)
);

BUFx6f_ASAP7_75t_L g5124 ( 
.A(n_4917),
.Y(n_5124)
);

INVx1_ASAP7_75t_L g5125 ( 
.A(n_4992),
.Y(n_5125)
);

INVx2_ASAP7_75t_L g5126 ( 
.A(n_4929),
.Y(n_5126)
);

NOR2xp33_ASAP7_75t_L g5127 ( 
.A(n_4975),
.B(n_3703),
.Y(n_5127)
);

BUFx6f_ASAP7_75t_L g5128 ( 
.A(n_4917),
.Y(n_5128)
);

NAND2x1p5_ASAP7_75t_L g5129 ( 
.A(n_5019),
.B(n_2882),
.Y(n_5129)
);

INVx2_ASAP7_75t_L g5130 ( 
.A(n_4917),
.Y(n_5130)
);

INVx2_ASAP7_75t_L g5131 ( 
.A(n_4918),
.Y(n_5131)
);

NAND2xp5_ASAP7_75t_L g5132 ( 
.A(n_4916),
.B(n_4138),
.Y(n_5132)
);

BUFx3_ASAP7_75t_L g5133 ( 
.A(n_4690),
.Y(n_5133)
);

AND2x2_ASAP7_75t_L g5134 ( 
.A(n_4887),
.B(n_3305),
.Y(n_5134)
);

BUFx2_ASAP7_75t_L g5135 ( 
.A(n_4843),
.Y(n_5135)
);

NOR2x1_ASAP7_75t_L g5136 ( 
.A(n_4921),
.B(n_2890),
.Y(n_5136)
);

INVx2_ASAP7_75t_L g5137 ( 
.A(n_4918),
.Y(n_5137)
);

OA21x2_ASAP7_75t_L g5138 ( 
.A1(n_4937),
.A2(n_4932),
.B(n_4643),
.Y(n_5138)
);

BUFx8_ASAP7_75t_L g5139 ( 
.A(n_4723),
.Y(n_5139)
);

INVx1_ASAP7_75t_L g5140 ( 
.A(n_4993),
.Y(n_5140)
);

OAI22xp5_ASAP7_75t_SL g5141 ( 
.A1(n_4842),
.A2(n_3313),
.B1(n_3346),
.B2(n_3147),
.Y(n_5141)
);

INVx1_ASAP7_75t_L g5142 ( 
.A(n_4995),
.Y(n_5142)
);

INVx1_ASAP7_75t_L g5143 ( 
.A(n_4996),
.Y(n_5143)
);

AND2x2_ASAP7_75t_L g5144 ( 
.A(n_4946),
.B(n_3312),
.Y(n_5144)
);

INVxp67_ASAP7_75t_L g5145 ( 
.A(n_4677),
.Y(n_5145)
);

HB1xp67_ASAP7_75t_L g5146 ( 
.A(n_4845),
.Y(n_5146)
);

INVx2_ASAP7_75t_L g5147 ( 
.A(n_4918),
.Y(n_5147)
);

BUFx6f_ASAP7_75t_L g5148 ( 
.A(n_5078),
.Y(n_5148)
);

AND2x4_ASAP7_75t_L g5149 ( 
.A(n_4755),
.B(n_3441),
.Y(n_5149)
);

NAND2xp5_ASAP7_75t_L g5150 ( 
.A(n_4976),
.B(n_2860),
.Y(n_5150)
);

NAND2xp5_ASAP7_75t_L g5151 ( 
.A(n_5060),
.B(n_2864),
.Y(n_5151)
);

CKINVDCx5p33_ASAP7_75t_R g5152 ( 
.A(n_4634),
.Y(n_5152)
);

CKINVDCx6p67_ASAP7_75t_R g5153 ( 
.A(n_4723),
.Y(n_5153)
);

BUFx6f_ASAP7_75t_L g5154 ( 
.A(n_5078),
.Y(n_5154)
);

INVx3_ASAP7_75t_L g5155 ( 
.A(n_4777),
.Y(n_5155)
);

INVx1_ASAP7_75t_L g5156 ( 
.A(n_4997),
.Y(n_5156)
);

INVx2_ASAP7_75t_L g5157 ( 
.A(n_5073),
.Y(n_5157)
);

OAI22xp5_ASAP7_75t_SL g5158 ( 
.A1(n_4850),
.A2(n_3480),
.B1(n_3558),
.B2(n_3368),
.Y(n_5158)
);

INVx2_ASAP7_75t_L g5159 ( 
.A(n_5092),
.Y(n_5159)
);

INVx2_ASAP7_75t_L g5160 ( 
.A(n_5111),
.Y(n_5160)
);

NAND2xp5_ASAP7_75t_SL g5161 ( 
.A(n_4864),
.B(n_4866),
.Y(n_5161)
);

AND2x2_ASAP7_75t_SL g5162 ( 
.A(n_5099),
.B(n_2866),
.Y(n_5162)
);

INVx1_ASAP7_75t_L g5163 ( 
.A(n_5002),
.Y(n_5163)
);

CKINVDCx6p67_ASAP7_75t_R g5164 ( 
.A(n_4817),
.Y(n_5164)
);

INVx1_ASAP7_75t_L g5165 ( 
.A(n_5007),
.Y(n_5165)
);

AND2x2_ASAP7_75t_L g5166 ( 
.A(n_4965),
.B(n_3312),
.Y(n_5166)
);

INVx1_ASAP7_75t_L g5167 ( 
.A(n_5008),
.Y(n_5167)
);

HB1xp67_ASAP7_75t_L g5168 ( 
.A(n_4846),
.Y(n_5168)
);

AND2x4_ASAP7_75t_L g5169 ( 
.A(n_4798),
.B(n_2943),
.Y(n_5169)
);

INVx1_ASAP7_75t_L g5170 ( 
.A(n_5009),
.Y(n_5170)
);

AND2x6_ASAP7_75t_L g5171 ( 
.A(n_4735),
.B(n_3262),
.Y(n_5171)
);

OAI22xp5_ASAP7_75t_L g5172 ( 
.A1(n_4924),
.A2(n_4819),
.B1(n_4935),
.B2(n_4645),
.Y(n_5172)
);

INVx2_ASAP7_75t_L g5173 ( 
.A(n_4943),
.Y(n_5173)
);

AND2x4_ASAP7_75t_L g5174 ( 
.A(n_4833),
.B(n_4863),
.Y(n_5174)
);

AOI22xp5_ASAP7_75t_L g5175 ( 
.A1(n_4919),
.A2(n_2920),
.B1(n_2939),
.B2(n_2903),
.Y(n_5175)
);

INVx3_ASAP7_75t_L g5176 ( 
.A(n_5068),
.Y(n_5176)
);

HB1xp67_ASAP7_75t_L g5177 ( 
.A(n_4796),
.Y(n_5177)
);

HB1xp67_ASAP7_75t_L g5178 ( 
.A(n_4802),
.Y(n_5178)
);

AND2x6_ASAP7_75t_L g5179 ( 
.A(n_4737),
.B(n_4702),
.Y(n_5179)
);

INVx1_ASAP7_75t_L g5180 ( 
.A(n_5013),
.Y(n_5180)
);

INVx1_ASAP7_75t_L g5181 ( 
.A(n_5016),
.Y(n_5181)
);

INVx2_ASAP7_75t_L g5182 ( 
.A(n_5078),
.Y(n_5182)
);

NOR2x1_ASAP7_75t_L g5183 ( 
.A(n_4641),
.B(n_2996),
.Y(n_5183)
);

OAI21x1_ASAP7_75t_L g5184 ( 
.A1(n_4741),
.A2(n_2956),
.B(n_2931),
.Y(n_5184)
);

INVx2_ASAP7_75t_L g5185 ( 
.A(n_4979),
.Y(n_5185)
);

BUFx6f_ASAP7_75t_L g5186 ( 
.A(n_5055),
.Y(n_5186)
);

INVx1_ASAP7_75t_L g5187 ( 
.A(n_5018),
.Y(n_5187)
);

INVx2_ASAP7_75t_L g5188 ( 
.A(n_5012),
.Y(n_5188)
);

AOI22xp5_ASAP7_75t_SL g5189 ( 
.A1(n_4933),
.A2(n_3980),
.B1(n_4044),
.B2(n_3940),
.Y(n_5189)
);

INVx1_ASAP7_75t_L g5190 ( 
.A(n_5027),
.Y(n_5190)
);

BUFx8_ASAP7_75t_L g5191 ( 
.A(n_4817),
.Y(n_5191)
);

INVx6_ASAP7_75t_L g5192 ( 
.A(n_4982),
.Y(n_5192)
);

INVx1_ASAP7_75t_L g5193 ( 
.A(n_5033),
.Y(n_5193)
);

BUFx6f_ASAP7_75t_L g5194 ( 
.A(n_5055),
.Y(n_5194)
);

AND2x2_ASAP7_75t_SL g5195 ( 
.A(n_4836),
.B(n_4862),
.Y(n_5195)
);

AOI22xp5_ASAP7_75t_L g5196 ( 
.A1(n_4906),
.A2(n_2999),
.B1(n_3082),
.B2(n_2995),
.Y(n_5196)
);

INVx1_ASAP7_75t_L g5197 ( 
.A(n_5036),
.Y(n_5197)
);

INVx3_ASAP7_75t_L g5198 ( 
.A(n_4782),
.Y(n_5198)
);

BUFx8_ASAP7_75t_L g5199 ( 
.A(n_5039),
.Y(n_5199)
);

INVx3_ASAP7_75t_L g5200 ( 
.A(n_4782),
.Y(n_5200)
);

AND2x2_ASAP7_75t_SL g5201 ( 
.A(n_4901),
.B(n_2981),
.Y(n_5201)
);

NAND2xp5_ASAP7_75t_L g5202 ( 
.A(n_4949),
.B(n_2986),
.Y(n_5202)
);

INVx4_ASAP7_75t_L g5203 ( 
.A(n_4869),
.Y(n_5203)
);

NAND2xp5_ASAP7_75t_SL g5204 ( 
.A(n_4934),
.B(n_3742),
.Y(n_5204)
);

OAI21x1_ASAP7_75t_L g5205 ( 
.A1(n_4642),
.A2(n_3094),
.B(n_2988),
.Y(n_5205)
);

AND2x2_ASAP7_75t_L g5206 ( 
.A(n_4945),
.B(n_3344),
.Y(n_5206)
);

AND2x4_ASAP7_75t_L g5207 ( 
.A(n_4651),
.B(n_3577),
.Y(n_5207)
);

AND2x6_ASAP7_75t_L g5208 ( 
.A(n_4652),
.B(n_4922),
.Y(n_5208)
);

AND2x2_ASAP7_75t_L g5209 ( 
.A(n_4880),
.B(n_3344),
.Y(n_5209)
);

BUFx6f_ASAP7_75t_L g5210 ( 
.A(n_5055),
.Y(n_5210)
);

INVx1_ASAP7_75t_L g5211 ( 
.A(n_5041),
.Y(n_5211)
);

AND2x4_ASAP7_75t_L g5212 ( 
.A(n_4697),
.B(n_2892),
.Y(n_5212)
);

INVx2_ASAP7_75t_SL g5213 ( 
.A(n_4908),
.Y(n_5213)
);

AND2x2_ASAP7_75t_L g5214 ( 
.A(n_4884),
.B(n_3354),
.Y(n_5214)
);

BUFx2_ASAP7_75t_L g5215 ( 
.A(n_4804),
.Y(n_5215)
);

INVx6_ASAP7_75t_L g5216 ( 
.A(n_4982),
.Y(n_5216)
);

NOR2xp33_ASAP7_75t_L g5217 ( 
.A(n_4954),
.B(n_3745),
.Y(n_5217)
);

BUFx6f_ASAP7_75t_L g5218 ( 
.A(n_4731),
.Y(n_5218)
);

INVx1_ASAP7_75t_L g5219 ( 
.A(n_5044),
.Y(n_5219)
);

AND2x4_ASAP7_75t_L g5220 ( 
.A(n_4742),
.B(n_2893),
.Y(n_5220)
);

INVx2_ASAP7_75t_L g5221 ( 
.A(n_4668),
.Y(n_5221)
);

AND2x2_ASAP7_75t_L g5222 ( 
.A(n_4892),
.B(n_3354),
.Y(n_5222)
);

AND2x2_ASAP7_75t_L g5223 ( 
.A(n_4711),
.B(n_3473),
.Y(n_5223)
);

INVx4_ASAP7_75t_L g5224 ( 
.A(n_4981),
.Y(n_5224)
);

NAND2xp5_ASAP7_75t_L g5225 ( 
.A(n_4952),
.B(n_4958),
.Y(n_5225)
);

NAND2xp5_ASAP7_75t_L g5226 ( 
.A(n_4959),
.B(n_4960),
.Y(n_5226)
);

BUFx6f_ASAP7_75t_L g5227 ( 
.A(n_4788),
.Y(n_5227)
);

BUFx6f_ASAP7_75t_L g5228 ( 
.A(n_4789),
.Y(n_5228)
);

OAI22xp5_ASAP7_75t_L g5229 ( 
.A1(n_4879),
.A2(n_4724),
.B1(n_4722),
.B2(n_4716),
.Y(n_5229)
);

INVx1_ASAP7_75t_L g5230 ( 
.A(n_5045),
.Y(n_5230)
);

INVx2_ASAP7_75t_L g5231 ( 
.A(n_4673),
.Y(n_5231)
);

AND2x6_ASAP7_75t_L g5232 ( 
.A(n_4968),
.B(n_3337),
.Y(n_5232)
);

INVx2_ASAP7_75t_L g5233 ( 
.A(n_4674),
.Y(n_5233)
);

NAND2xp5_ASAP7_75t_L g5234 ( 
.A(n_4964),
.B(n_3108),
.Y(n_5234)
);

INVx2_ASAP7_75t_L g5235 ( 
.A(n_4676),
.Y(n_5235)
);

OR2x6_ASAP7_75t_L g5236 ( 
.A(n_4868),
.B(n_3698),
.Y(n_5236)
);

INVx1_ASAP7_75t_L g5237 ( 
.A(n_5046),
.Y(n_5237)
);

INVx2_ASAP7_75t_L g5238 ( 
.A(n_4680),
.Y(n_5238)
);

BUFx6f_ASAP7_75t_L g5239 ( 
.A(n_4794),
.Y(n_5239)
);

INVx2_ASAP7_75t_L g5240 ( 
.A(n_4681),
.Y(n_5240)
);

AND2x4_ASAP7_75t_L g5241 ( 
.A(n_4750),
.B(n_4787),
.Y(n_5241)
);

INVx3_ASAP7_75t_L g5242 ( 
.A(n_4956),
.Y(n_5242)
);

AND2x2_ASAP7_75t_L g5243 ( 
.A(n_4780),
.B(n_3473),
.Y(n_5243)
);

INVx2_ASAP7_75t_L g5244 ( 
.A(n_4682),
.Y(n_5244)
);

INVxp67_ASAP7_75t_SL g5245 ( 
.A(n_4648),
.Y(n_5245)
);

AND2x6_ASAP7_75t_L g5246 ( 
.A(n_4984),
.B(n_3365),
.Y(n_5246)
);

BUFx6f_ASAP7_75t_L g5247 ( 
.A(n_4664),
.Y(n_5247)
);

XNOR2xp5_ASAP7_75t_L g5248 ( 
.A(n_4774),
.B(n_4062),
.Y(n_5248)
);

INVx1_ASAP7_75t_L g5249 ( 
.A(n_5047),
.Y(n_5249)
);

AND2x4_ASAP7_75t_L g5250 ( 
.A(n_4670),
.B(n_2896),
.Y(n_5250)
);

INVx2_ASAP7_75t_L g5251 ( 
.A(n_4683),
.Y(n_5251)
);

OAI22xp5_ASAP7_75t_L g5252 ( 
.A1(n_4756),
.A2(n_4797),
.B1(n_5038),
.B2(n_4835),
.Y(n_5252)
);

INVx2_ASAP7_75t_L g5253 ( 
.A(n_4687),
.Y(n_5253)
);

INVxp67_ASAP7_75t_L g5254 ( 
.A(n_4865),
.Y(n_5254)
);

INVx1_ASAP7_75t_L g5255 ( 
.A(n_5014),
.Y(n_5255)
);

INVx2_ASAP7_75t_L g5256 ( 
.A(n_4689),
.Y(n_5256)
);

INVx3_ASAP7_75t_L g5257 ( 
.A(n_4665),
.Y(n_5257)
);

BUFx6f_ASAP7_75t_L g5258 ( 
.A(n_4667),
.Y(n_5258)
);

AOI22xp5_ASAP7_75t_L g5259 ( 
.A1(n_4889),
.A2(n_3192),
.B1(n_3218),
.B2(n_3131),
.Y(n_5259)
);

AND2x2_ASAP7_75t_SL g5260 ( 
.A(n_4775),
.B(n_3209),
.Y(n_5260)
);

XNOR2x2_ASAP7_75t_L g5261 ( 
.A(n_5025),
.B(n_3724),
.Y(n_5261)
);

NOR2x1_ASAP7_75t_L g5262 ( 
.A(n_4770),
.B(n_4771),
.Y(n_5262)
);

AND2x2_ASAP7_75t_SL g5263 ( 
.A(n_4622),
.B(n_3213),
.Y(n_5263)
);

OAI22x1_ASAP7_75t_L g5264 ( 
.A1(n_4858),
.A2(n_3909),
.B1(n_3606),
.B2(n_3806),
.Y(n_5264)
);

INVx6_ASAP7_75t_L g5265 ( 
.A(n_4870),
.Y(n_5265)
);

INVx2_ASAP7_75t_L g5266 ( 
.A(n_4692),
.Y(n_5266)
);

AND2x2_ASAP7_75t_L g5267 ( 
.A(n_4736),
.B(n_3519),
.Y(n_5267)
);

INVx4_ASAP7_75t_L g5268 ( 
.A(n_4990),
.Y(n_5268)
);

AND2x2_ASAP7_75t_L g5269 ( 
.A(n_5053),
.B(n_3519),
.Y(n_5269)
);

INVx2_ASAP7_75t_L g5270 ( 
.A(n_4725),
.Y(n_5270)
);

INVx2_ASAP7_75t_L g5271 ( 
.A(n_4729),
.Y(n_5271)
);

BUFx6f_ASAP7_75t_L g5272 ( 
.A(n_4693),
.Y(n_5272)
);

HB1xp67_ASAP7_75t_L g5273 ( 
.A(n_4878),
.Y(n_5273)
);

AND2x2_ASAP7_75t_L g5274 ( 
.A(n_4632),
.B(n_3614),
.Y(n_5274)
);

INVx2_ASAP7_75t_L g5275 ( 
.A(n_4738),
.Y(n_5275)
);

HB1xp67_ASAP7_75t_L g5276 ( 
.A(n_4872),
.Y(n_5276)
);

AND2x2_ASAP7_75t_L g5277 ( 
.A(n_4636),
.B(n_3614),
.Y(n_5277)
);

INVx3_ASAP7_75t_L g5278 ( 
.A(n_4696),
.Y(n_5278)
);

INVx1_ASAP7_75t_L g5279 ( 
.A(n_5022),
.Y(n_5279)
);

OAI22x1_ASAP7_75t_R g5280 ( 
.A1(n_4662),
.A2(n_4111),
.B1(n_2973),
.B2(n_2993),
.Y(n_5280)
);

NOR2x1_ASAP7_75t_L g5281 ( 
.A(n_4649),
.B(n_3925),
.Y(n_5281)
);

INVx2_ASAP7_75t_L g5282 ( 
.A(n_4739),
.Y(n_5282)
);

INVx2_ASAP7_75t_L g5283 ( 
.A(n_4740),
.Y(n_5283)
);

AND2x4_ASAP7_75t_L g5284 ( 
.A(n_5031),
.B(n_2905),
.Y(n_5284)
);

OAI22xp5_ASAP7_75t_L g5285 ( 
.A1(n_5030),
.A2(n_3808),
.B1(n_3845),
.B2(n_3766),
.Y(n_5285)
);

AND2x6_ASAP7_75t_L g5286 ( 
.A(n_5052),
.B(n_3776),
.Y(n_5286)
);

BUFx6f_ASAP7_75t_L g5287 ( 
.A(n_4699),
.Y(n_5287)
);

OAI22xp5_ASAP7_75t_SL g5288 ( 
.A1(n_4844),
.A2(n_3058),
.B1(n_3088),
.B2(n_2954),
.Y(n_5288)
);

INVx1_ASAP7_75t_L g5289 ( 
.A(n_4650),
.Y(n_5289)
);

INVx1_ASAP7_75t_L g5290 ( 
.A(n_4655),
.Y(n_5290)
);

AND2x2_ASAP7_75t_L g5291 ( 
.A(n_4638),
.B(n_3629),
.Y(n_5291)
);

CKINVDCx5p33_ASAP7_75t_R g5292 ( 
.A(n_4635),
.Y(n_5292)
);

NAND2xp5_ASAP7_75t_L g5293 ( 
.A(n_4966),
.B(n_3228),
.Y(n_5293)
);

INVx1_ASAP7_75t_L g5294 ( 
.A(n_4656),
.Y(n_5294)
);

AND2x6_ASAP7_75t_L g5295 ( 
.A(n_5029),
.B(n_4149),
.Y(n_5295)
);

OA21x2_ASAP7_75t_L g5296 ( 
.A1(n_4658),
.A2(n_4663),
.B(n_4659),
.Y(n_5296)
);

NAND2xp5_ASAP7_75t_L g5297 ( 
.A(n_4967),
.B(n_3266),
.Y(n_5297)
);

BUFx6f_ASAP7_75t_L g5298 ( 
.A(n_4700),
.Y(n_5298)
);

HB1xp67_ASAP7_75t_L g5299 ( 
.A(n_4874),
.Y(n_5299)
);

OA21x2_ASAP7_75t_L g5300 ( 
.A1(n_4799),
.A2(n_4805),
.B(n_4800),
.Y(n_5300)
);

INVx1_ASAP7_75t_L g5301 ( 
.A(n_4808),
.Y(n_5301)
);

AOI22xp5_ASAP7_75t_L g5302 ( 
.A1(n_4891),
.A2(n_3227),
.B1(n_3330),
.B2(n_3220),
.Y(n_5302)
);

AND2x2_ASAP7_75t_L g5303 ( 
.A(n_4639),
.B(n_3629),
.Y(n_5303)
);

INVx3_ASAP7_75t_L g5304 ( 
.A(n_4704),
.Y(n_5304)
);

OA21x2_ASAP7_75t_L g5305 ( 
.A1(n_4812),
.A2(n_2917),
.B(n_2913),
.Y(n_5305)
);

AND2x4_ASAP7_75t_L g5306 ( 
.A(n_5032),
.B(n_2919),
.Y(n_5306)
);

INVx2_ASAP7_75t_L g5307 ( 
.A(n_4744),
.Y(n_5307)
);

INVx2_ASAP7_75t_L g5308 ( 
.A(n_4746),
.Y(n_5308)
);

AND2x4_ASAP7_75t_L g5309 ( 
.A(n_5035),
.B(n_2926),
.Y(n_5309)
);

INVx2_ASAP7_75t_L g5310 ( 
.A(n_4748),
.Y(n_5310)
);

INVx1_ASAP7_75t_L g5311 ( 
.A(n_4814),
.Y(n_5311)
);

OAI21x1_ASAP7_75t_L g5312 ( 
.A1(n_4820),
.A2(n_4827),
.B(n_4822),
.Y(n_5312)
);

INVx2_ASAP7_75t_L g5313 ( 
.A(n_4752),
.Y(n_5313)
);

INVx2_ASAP7_75t_L g5314 ( 
.A(n_4754),
.Y(n_5314)
);

XOR2xp5_ASAP7_75t_L g5315 ( 
.A(n_4621),
.B(n_4623),
.Y(n_5315)
);

AND2x4_ASAP7_75t_L g5316 ( 
.A(n_5037),
.B(n_2929),
.Y(n_5316)
);

INVx2_ASAP7_75t_L g5317 ( 
.A(n_4757),
.Y(n_5317)
);

AND2x2_ASAP7_75t_L g5318 ( 
.A(n_5034),
.B(n_3734),
.Y(n_5318)
);

CKINVDCx11_ASAP7_75t_R g5319 ( 
.A(n_4776),
.Y(n_5319)
);

INVx3_ASAP7_75t_L g5320 ( 
.A(n_4707),
.Y(n_5320)
);

INVx2_ASAP7_75t_L g5321 ( 
.A(n_4758),
.Y(n_5321)
);

INVx2_ASAP7_75t_L g5322 ( 
.A(n_4759),
.Y(n_5322)
);

NAND2xp5_ASAP7_75t_L g5323 ( 
.A(n_4971),
.B(n_3284),
.Y(n_5323)
);

BUFx6f_ASAP7_75t_L g5324 ( 
.A(n_4708),
.Y(n_5324)
);

NAND2xp5_ASAP7_75t_L g5325 ( 
.A(n_4828),
.B(n_3327),
.Y(n_5325)
);

INVx1_ASAP7_75t_L g5326 ( 
.A(n_4830),
.Y(n_5326)
);

AND2x6_ASAP7_75t_L g5327 ( 
.A(n_5043),
.B(n_3381),
.Y(n_5327)
);

CKINVDCx6p67_ASAP7_75t_R g5328 ( 
.A(n_4825),
.Y(n_5328)
);

OA21x2_ASAP7_75t_L g5329 ( 
.A1(n_4834),
.A2(n_2933),
.B(n_2932),
.Y(n_5329)
);

OAI22xp5_ASAP7_75t_L g5330 ( 
.A1(n_5048),
.A2(n_3864),
.B1(n_3865),
.B2(n_3857),
.Y(n_5330)
);

NAND2xp5_ASAP7_75t_L g5331 ( 
.A(n_4839),
.B(n_3328),
.Y(n_5331)
);

INVx3_ASAP7_75t_L g5332 ( 
.A(n_4709),
.Y(n_5332)
);

AND2x4_ASAP7_75t_L g5333 ( 
.A(n_5004),
.B(n_2937),
.Y(n_5333)
);

NAND3xp33_ASAP7_75t_L g5334 ( 
.A(n_4999),
.B(n_3881),
.C(n_3878),
.Y(n_5334)
);

AND2x4_ASAP7_75t_L g5335 ( 
.A(n_5054),
.B(n_2945),
.Y(n_5335)
);

AND2x4_ASAP7_75t_L g5336 ( 
.A(n_4912),
.B(n_4624),
.Y(n_5336)
);

INVx2_ASAP7_75t_L g5337 ( 
.A(n_4760),
.Y(n_5337)
);

INVx2_ASAP7_75t_L g5338 ( 
.A(n_4763),
.Y(n_5338)
);

BUFx3_ASAP7_75t_L g5339 ( 
.A(n_4629),
.Y(n_5339)
);

NAND2xp5_ASAP7_75t_L g5340 ( 
.A(n_4840),
.B(n_4848),
.Y(n_5340)
);

BUFx6f_ASAP7_75t_L g5341 ( 
.A(n_4712),
.Y(n_5341)
);

INVx2_ASAP7_75t_L g5342 ( 
.A(n_4764),
.Y(n_5342)
);

INVx2_ASAP7_75t_L g5343 ( 
.A(n_4767),
.Y(n_5343)
);

INVx3_ASAP7_75t_L g5344 ( 
.A(n_4851),
.Y(n_5344)
);

HB1xp67_ASAP7_75t_L g5345 ( 
.A(n_4876),
.Y(n_5345)
);

INVx3_ASAP7_75t_L g5346 ( 
.A(n_4856),
.Y(n_5346)
);

AND2x6_ASAP7_75t_L g5347 ( 
.A(n_5057),
.B(n_3398),
.Y(n_5347)
);

INVx3_ASAP7_75t_L g5348 ( 
.A(n_4857),
.Y(n_5348)
);

INVx1_ASAP7_75t_L g5349 ( 
.A(n_4859),
.Y(n_5349)
);

INVx1_ASAP7_75t_L g5350 ( 
.A(n_4867),
.Y(n_5350)
);

HB1xp67_ASAP7_75t_L g5351 ( 
.A(n_4970),
.Y(n_5351)
);

INVx1_ASAP7_75t_L g5352 ( 
.A(n_4873),
.Y(n_5352)
);

INVx3_ASAP7_75t_L g5353 ( 
.A(n_4877),
.Y(n_5353)
);

INVx1_ASAP7_75t_L g5354 ( 
.A(n_4881),
.Y(n_5354)
);

INVx2_ASAP7_75t_L g5355 ( 
.A(n_4768),
.Y(n_5355)
);

INVx2_ASAP7_75t_L g5356 ( 
.A(n_4769),
.Y(n_5356)
);

OA21x2_ASAP7_75t_L g5357 ( 
.A1(n_4885),
.A2(n_2951),
.B(n_2946),
.Y(n_5357)
);

INVx2_ASAP7_75t_L g5358 ( 
.A(n_4772),
.Y(n_5358)
);

INVx1_ASAP7_75t_L g5359 ( 
.A(n_4894),
.Y(n_5359)
);

INVx1_ASAP7_75t_SL g5360 ( 
.A(n_4847),
.Y(n_5360)
);

INVx3_ASAP7_75t_L g5361 ( 
.A(n_4896),
.Y(n_5361)
);

NOR2x1_ASAP7_75t_L g5362 ( 
.A(n_4897),
.B(n_2966),
.Y(n_5362)
);

INVx3_ASAP7_75t_L g5363 ( 
.A(n_4898),
.Y(n_5363)
);

INVx1_ASAP7_75t_L g5364 ( 
.A(n_4907),
.Y(n_5364)
);

INVx2_ASAP7_75t_L g5365 ( 
.A(n_4783),
.Y(n_5365)
);

INVx3_ASAP7_75t_L g5366 ( 
.A(n_4911),
.Y(n_5366)
);

NOR2xp33_ASAP7_75t_L g5367 ( 
.A(n_5065),
.B(n_3885),
.Y(n_5367)
);

BUFx6f_ASAP7_75t_L g5368 ( 
.A(n_5058),
.Y(n_5368)
);

AND2x2_ASAP7_75t_SL g5369 ( 
.A(n_4657),
.B(n_3392),
.Y(n_5369)
);

NOR2xp33_ASAP7_75t_L g5370 ( 
.A(n_5067),
.B(n_3891),
.Y(n_5370)
);

NAND2xp5_ASAP7_75t_L g5371 ( 
.A(n_4920),
.B(n_3397),
.Y(n_5371)
);

INVx1_ASAP7_75t_L g5372 ( 
.A(n_4923),
.Y(n_5372)
);

AND2x2_ASAP7_75t_L g5373 ( 
.A(n_5049),
.B(n_3734),
.Y(n_5373)
);

AND2x6_ASAP7_75t_L g5374 ( 
.A(n_4925),
.B(n_3421),
.Y(n_5374)
);

AND2x4_ASAP7_75t_L g5375 ( 
.A(n_5069),
.B(n_2972),
.Y(n_5375)
);

OAI21x1_ASAP7_75t_L g5376 ( 
.A1(n_4926),
.A2(n_3434),
.B(n_3433),
.Y(n_5376)
);

INVx2_ASAP7_75t_L g5377 ( 
.A(n_4784),
.Y(n_5377)
);

AND2x4_ASAP7_75t_L g5378 ( 
.A(n_5076),
.B(n_2978),
.Y(n_5378)
);

INVx2_ASAP7_75t_L g5379 ( 
.A(n_4714),
.Y(n_5379)
);

INVx2_ASAP7_75t_L g5380 ( 
.A(n_4715),
.Y(n_5380)
);

BUFx6f_ASAP7_75t_L g5381 ( 
.A(n_4927),
.Y(n_5381)
);

NOR2xp33_ASAP7_75t_L g5382 ( 
.A(n_5080),
.B(n_3904),
.Y(n_5382)
);

OAI22x1_ASAP7_75t_R g5383 ( 
.A1(n_4671),
.A2(n_3217),
.B1(n_3221),
.B2(n_3111),
.Y(n_5383)
);

INVx3_ASAP7_75t_L g5384 ( 
.A(n_4928),
.Y(n_5384)
);

INVx1_ASAP7_75t_L g5385 ( 
.A(n_4930),
.Y(n_5385)
);

INVx1_ASAP7_75t_L g5386 ( 
.A(n_4931),
.Y(n_5386)
);

INVx1_ASAP7_75t_L g5387 ( 
.A(n_4936),
.Y(n_5387)
);

OAI22xp5_ASAP7_75t_SL g5388 ( 
.A1(n_4849),
.A2(n_3230),
.B1(n_3237),
.B2(n_3223),
.Y(n_5388)
);

INVx1_ASAP7_75t_L g5389 ( 
.A(n_4938),
.Y(n_5389)
);

NAND2xp5_ASAP7_75t_L g5390 ( 
.A(n_4939),
.B(n_3545),
.Y(n_5390)
);

AND2x2_ASAP7_75t_L g5391 ( 
.A(n_5050),
.B(n_5082),
.Y(n_5391)
);

INVx6_ASAP7_75t_L g5392 ( 
.A(n_4871),
.Y(n_5392)
);

INVx1_ASAP7_75t_L g5393 ( 
.A(n_4941),
.Y(n_5393)
);

AOI22xp5_ASAP7_75t_L g5394 ( 
.A1(n_4893),
.A2(n_3510),
.B1(n_3512),
.B2(n_3423),
.Y(n_5394)
);

BUFx6f_ASAP7_75t_L g5395 ( 
.A(n_4942),
.Y(n_5395)
);

NAND2xp5_ASAP7_75t_L g5396 ( 
.A(n_4944),
.B(n_3568),
.Y(n_5396)
);

HB1xp67_ASAP7_75t_L g5397 ( 
.A(n_4672),
.Y(n_5397)
);

INVx1_ASAP7_75t_L g5398 ( 
.A(n_4951),
.Y(n_5398)
);

BUFx6f_ASAP7_75t_L g5399 ( 
.A(n_4957),
.Y(n_5399)
);

AND2x2_ASAP7_75t_L g5400 ( 
.A(n_5084),
.B(n_3754),
.Y(n_5400)
);

INVx1_ASAP7_75t_L g5401 ( 
.A(n_4961),
.Y(n_5401)
);

INVx1_ASAP7_75t_L g5402 ( 
.A(n_4962),
.Y(n_5402)
);

INVx1_ASAP7_75t_L g5403 ( 
.A(n_4963),
.Y(n_5403)
);

AND2x4_ASAP7_75t_L g5404 ( 
.A(n_5086),
.B(n_5087),
.Y(n_5404)
);

INVx6_ASAP7_75t_L g5405 ( 
.A(n_4875),
.Y(n_5405)
);

INVx2_ASAP7_75t_L g5406 ( 
.A(n_4717),
.Y(n_5406)
);

INVx2_ASAP7_75t_L g5407 ( 
.A(n_4720),
.Y(n_5407)
);

AND2x2_ASAP7_75t_L g5408 ( 
.A(n_5088),
.B(n_3754),
.Y(n_5408)
);

BUFx3_ASAP7_75t_L g5409 ( 
.A(n_5090),
.Y(n_5409)
);

INVx2_ASAP7_75t_L g5410 ( 
.A(n_4969),
.Y(n_5410)
);

AND2x4_ASAP7_75t_L g5411 ( 
.A(n_5093),
.B(n_2980),
.Y(n_5411)
);

OAI21x1_ASAP7_75t_L g5412 ( 
.A1(n_4973),
.A2(n_3633),
.B(n_3627),
.Y(n_5412)
);

INVx1_ASAP7_75t_L g5413 ( 
.A(n_4974),
.Y(n_5413)
);

INVx1_ASAP7_75t_L g5414 ( 
.A(n_4977),
.Y(n_5414)
);

BUFx2_ASAP7_75t_L g5415 ( 
.A(n_4852),
.Y(n_5415)
);

OAI22xp33_ASAP7_75t_L g5416 ( 
.A1(n_5042),
.A2(n_3580),
.B1(n_3592),
.B2(n_3578),
.Y(n_5416)
);

NAND2xp5_ASAP7_75t_L g5417 ( 
.A(n_4980),
.B(n_3636),
.Y(n_5417)
);

BUFx6f_ASAP7_75t_L g5418 ( 
.A(n_4983),
.Y(n_5418)
);

INVx2_ASAP7_75t_L g5419 ( 
.A(n_4987),
.Y(n_5419)
);

AND2x2_ASAP7_75t_L g5420 ( 
.A(n_5094),
.B(n_3939),
.Y(n_5420)
);

NOR2xp33_ASAP7_75t_L g5421 ( 
.A(n_5097),
.B(n_5098),
.Y(n_5421)
);

AND2x2_ASAP7_75t_L g5422 ( 
.A(n_5101),
.B(n_3939),
.Y(n_5422)
);

INVx1_ASAP7_75t_L g5423 ( 
.A(n_4940),
.Y(n_5423)
);

CKINVDCx6p67_ASAP7_75t_R g5424 ( 
.A(n_4826),
.Y(n_5424)
);

INVx1_ASAP7_75t_L g5425 ( 
.A(n_4985),
.Y(n_5425)
);

INVx3_ASAP7_75t_L g5426 ( 
.A(n_5104),
.Y(n_5426)
);

INVx2_ASAP7_75t_L g5427 ( 
.A(n_5108),
.Y(n_5427)
);

AND2x2_ASAP7_75t_SL g5428 ( 
.A(n_4694),
.B(n_3640),
.Y(n_5428)
);

NAND2xp33_ASAP7_75t_L g5429 ( 
.A(n_4888),
.B(n_3905),
.Y(n_5429)
);

BUFx6f_ASAP7_75t_L g5430 ( 
.A(n_5109),
.Y(n_5430)
);

AND2x2_ASAP7_75t_L g5431 ( 
.A(n_5110),
.B(n_3995),
.Y(n_5431)
);

OAI22xp5_ASAP7_75t_L g5432 ( 
.A1(n_5072),
.A2(n_3918),
.B1(n_3920),
.B2(n_3912),
.Y(n_5432)
);

INVxp67_ASAP7_75t_L g5433 ( 
.A(n_4860),
.Y(n_5433)
);

HB1xp67_ASAP7_75t_L g5434 ( 
.A(n_4890),
.Y(n_5434)
);

INVx1_ASAP7_75t_L g5435 ( 
.A(n_5051),
.Y(n_5435)
);

INVx2_ASAP7_75t_L g5436 ( 
.A(n_5112),
.Y(n_5436)
);

BUFx6f_ASAP7_75t_L g5437 ( 
.A(n_5115),
.Y(n_5437)
);

AND2x2_ASAP7_75t_L g5438 ( 
.A(n_5120),
.B(n_3995),
.Y(n_5438)
);

CKINVDCx11_ASAP7_75t_R g5439 ( 
.A(n_4831),
.Y(n_5439)
);

INVx1_ASAP7_75t_L g5440 ( 
.A(n_4905),
.Y(n_5440)
);

INVx1_ASAP7_75t_L g5441 ( 
.A(n_5003),
.Y(n_5441)
);

BUFx6f_ASAP7_75t_L g5442 ( 
.A(n_5010),
.Y(n_5442)
);

INVx3_ASAP7_75t_L g5443 ( 
.A(n_5011),
.Y(n_5443)
);

OAI21x1_ASAP7_75t_L g5444 ( 
.A1(n_4978),
.A2(n_3774),
.B(n_3711),
.Y(n_5444)
);

AND2x2_ASAP7_75t_L g5445 ( 
.A(n_5015),
.B(n_4053),
.Y(n_5445)
);

AND2x6_ASAP7_75t_L g5446 ( 
.A(n_4679),
.B(n_3621),
.Y(n_5446)
);

INVx1_ASAP7_75t_L g5447 ( 
.A(n_4994),
.Y(n_5447)
);

INVx1_ASAP7_75t_L g5448 ( 
.A(n_5000),
.Y(n_5448)
);

NOR2xp33_ASAP7_75t_L g5449 ( 
.A(n_4899),
.B(n_3942),
.Y(n_5449)
);

INVx1_ASAP7_75t_L g5450 ( 
.A(n_5056),
.Y(n_5450)
);

INVx2_ASAP7_75t_L g5451 ( 
.A(n_4955),
.Y(n_5451)
);

INVxp33_ASAP7_75t_SL g5452 ( 
.A(n_5075),
.Y(n_5452)
);

OA21x2_ASAP7_75t_L g5453 ( 
.A1(n_4998),
.A2(n_2983),
.B(n_2982),
.Y(n_5453)
);

NAND2xp5_ASAP7_75t_L g5454 ( 
.A(n_4902),
.B(n_3799),
.Y(n_5454)
);

OA21x2_ASAP7_75t_L g5455 ( 
.A1(n_5026),
.A2(n_3000),
.B(n_2994),
.Y(n_5455)
);

OAI22xp5_ASAP7_75t_SL g5456 ( 
.A1(n_4854),
.A2(n_3251),
.B1(n_3264),
.B2(n_3247),
.Y(n_5456)
);

HB1xp67_ASAP7_75t_L g5457 ( 
.A(n_4913),
.Y(n_5457)
);

AND2x2_ASAP7_75t_L g5458 ( 
.A(n_4803),
.B(n_4811),
.Y(n_5458)
);

CKINVDCx5p33_ASAP7_75t_R g5459 ( 
.A(n_4640),
.Y(n_5459)
);

INVx2_ASAP7_75t_L g5460 ( 
.A(n_5040),
.Y(n_5460)
);

NAND2xp5_ASAP7_75t_L g5461 ( 
.A(n_4886),
.B(n_4947),
.Y(n_5461)
);

INVx1_ASAP7_75t_L g5462 ( 
.A(n_4986),
.Y(n_5462)
);

INVx1_ASAP7_75t_L g5463 ( 
.A(n_4948),
.Y(n_5463)
);

INVx3_ASAP7_75t_L g5464 ( 
.A(n_4883),
.Y(n_5464)
);

INVx1_ASAP7_75t_L g5465 ( 
.A(n_4950),
.Y(n_5465)
);

NOR2xp33_ASAP7_75t_L g5466 ( 
.A(n_4647),
.B(n_3971),
.Y(n_5466)
);

HB1xp67_ASAP7_75t_L g5467 ( 
.A(n_4855),
.Y(n_5467)
);

NAND2xp5_ASAP7_75t_L g5468 ( 
.A(n_5020),
.B(n_3833),
.Y(n_5468)
);

INVx1_ASAP7_75t_L g5469 ( 
.A(n_4953),
.Y(n_5469)
);

INVx2_ASAP7_75t_L g5470 ( 
.A(n_4972),
.Y(n_5470)
);

INVx1_ASAP7_75t_L g5471 ( 
.A(n_4988),
.Y(n_5471)
);

INVx1_ASAP7_75t_L g5472 ( 
.A(n_4989),
.Y(n_5472)
);

BUFx2_ASAP7_75t_L g5473 ( 
.A(n_4861),
.Y(n_5473)
);

NAND2xp33_ASAP7_75t_L g5474 ( 
.A(n_4654),
.B(n_4660),
.Y(n_5474)
);

INVx1_ASAP7_75t_L g5475 ( 
.A(n_4991),
.Y(n_5475)
);

INVx1_ASAP7_75t_L g5476 ( 
.A(n_5001),
.Y(n_5476)
);

NAND2xp5_ASAP7_75t_L g5477 ( 
.A(n_5023),
.B(n_3902),
.Y(n_5477)
);

AOI22xp5_ASAP7_75t_L g5478 ( 
.A1(n_4895),
.A2(n_3696),
.B1(n_3752),
.B2(n_3652),
.Y(n_5478)
);

INVx1_ASAP7_75t_L g5479 ( 
.A(n_5005),
.Y(n_5479)
);

BUFx6f_ASAP7_75t_L g5480 ( 
.A(n_4661),
.Y(n_5480)
);

INVx2_ASAP7_75t_L g5481 ( 
.A(n_5006),
.Y(n_5481)
);

INVx1_ASAP7_75t_L g5482 ( 
.A(n_5017),
.Y(n_5482)
);

INVx2_ASAP7_75t_L g5483 ( 
.A(n_5021),
.Y(n_5483)
);

INVx3_ASAP7_75t_L g5484 ( 
.A(n_4853),
.Y(n_5484)
);

INVx1_ASAP7_75t_L g5485 ( 
.A(n_5028),
.Y(n_5485)
);

BUFx2_ASAP7_75t_L g5486 ( 
.A(n_4838),
.Y(n_5486)
);

AOI22xp5_ASAP7_75t_L g5487 ( 
.A1(n_4900),
.A2(n_3805),
.B1(n_3815),
.B2(n_3756),
.Y(n_5487)
);

OAI22xp5_ASAP7_75t_SL g5488 ( 
.A1(n_4841),
.A2(n_3283),
.B1(n_3309),
.B2(n_3276),
.Y(n_5488)
);

NAND2xp5_ASAP7_75t_SL g5489 ( 
.A(n_4666),
.B(n_3979),
.Y(n_5489)
);

NAND2xp5_ASAP7_75t_L g5490 ( 
.A(n_5024),
.B(n_3941),
.Y(n_5490)
);

OAI22xp5_ASAP7_75t_SL g5491 ( 
.A1(n_4703),
.A2(n_3360),
.B1(n_3379),
.B2(n_3357),
.Y(n_5491)
);

OA21x2_ASAP7_75t_L g5492 ( 
.A1(n_4669),
.A2(n_3009),
.B(n_3008),
.Y(n_5492)
);

INVx1_ASAP7_75t_L g5493 ( 
.A(n_4903),
.Y(n_5493)
);

INVx2_ASAP7_75t_L g5494 ( 
.A(n_4904),
.Y(n_5494)
);

AOI22xp5_ASAP7_75t_L g5495 ( 
.A1(n_4909),
.A2(n_3949),
.B1(n_3965),
.B2(n_3834),
.Y(n_5495)
);

INVx1_ASAP7_75t_L g5496 ( 
.A(n_4914),
.Y(n_5496)
);

OAI21x1_ASAP7_75t_L g5497 ( 
.A1(n_4705),
.A2(n_3978),
.B(n_3951),
.Y(n_5497)
);

OA21x2_ASAP7_75t_L g5498 ( 
.A1(n_4675),
.A2(n_3014),
.B(n_3010),
.Y(n_5498)
);

NOR2xp33_ASAP7_75t_L g5499 ( 
.A(n_4678),
.B(n_3999),
.Y(n_5499)
);

INVx1_ASAP7_75t_L g5500 ( 
.A(n_4915),
.Y(n_5500)
);

BUFx6f_ASAP7_75t_L g5501 ( 
.A(n_4691),
.Y(n_5501)
);

NOR2xp33_ASAP7_75t_R g5502 ( 
.A(n_4625),
.B(n_3389),
.Y(n_5502)
);

INVxp67_ASAP7_75t_L g5503 ( 
.A(n_5102),
.Y(n_5503)
);

INVx3_ASAP7_75t_L g5504 ( 
.A(n_4695),
.Y(n_5504)
);

INVx1_ASAP7_75t_L g5505 ( 
.A(n_5105),
.Y(n_5505)
);

NAND2xp5_ASAP7_75t_L g5506 ( 
.A(n_4698),
.B(n_3989),
.Y(n_5506)
);

INVx3_ASAP7_75t_L g5507 ( 
.A(n_4701),
.Y(n_5507)
);

INVx1_ASAP7_75t_L g5508 ( 
.A(n_5116),
.Y(n_5508)
);

BUFx6f_ASAP7_75t_L g5509 ( 
.A(n_4706),
.Y(n_5509)
);

INVx2_ASAP7_75t_L g5510 ( 
.A(n_4713),
.Y(n_5510)
);

INVx1_ASAP7_75t_L g5511 ( 
.A(n_5118),
.Y(n_5511)
);

INVx3_ASAP7_75t_L g5512 ( 
.A(n_4718),
.Y(n_5512)
);

CKINVDCx16_ASAP7_75t_R g5513 ( 
.A(n_4710),
.Y(n_5513)
);

INVx1_ASAP7_75t_L g5514 ( 
.A(n_4719),
.Y(n_5514)
);

OAI22xp5_ASAP7_75t_SL g5515 ( 
.A1(n_4686),
.A2(n_3404),
.B1(n_3420),
.B2(n_3393),
.Y(n_5515)
);

BUFx2_ASAP7_75t_L g5516 ( 
.A(n_4688),
.Y(n_5516)
);

NAND2xp5_ASAP7_75t_L g5517 ( 
.A(n_4726),
.B(n_4025),
.Y(n_5517)
);

INVx1_ASAP7_75t_L g5518 ( 
.A(n_4727),
.Y(n_5518)
);

INVx2_ASAP7_75t_L g5519 ( 
.A(n_4728),
.Y(n_5519)
);

OAI22xp5_ASAP7_75t_SL g5520 ( 
.A1(n_4684),
.A2(n_3444),
.B1(n_3478),
.B2(n_3438),
.Y(n_5520)
);

INVx1_ASAP7_75t_L g5521 ( 
.A(n_4732),
.Y(n_5521)
);

INVx1_ASAP7_75t_L g5522 ( 
.A(n_4734),
.Y(n_5522)
);

INVx1_ASAP7_75t_L g5523 ( 
.A(n_4745),
.Y(n_5523)
);

INVx1_ASAP7_75t_L g5524 ( 
.A(n_4761),
.Y(n_5524)
);

INVx3_ASAP7_75t_L g5525 ( 
.A(n_4766),
.Y(n_5525)
);

OAI22xp5_ASAP7_75t_SL g5526 ( 
.A1(n_4882),
.A2(n_3505),
.B1(n_3511),
.B2(n_3501),
.Y(n_5526)
);

AND2x2_ASAP7_75t_L g5527 ( 
.A(n_4773),
.B(n_4053),
.Y(n_5527)
);

AOI22xp5_ASAP7_75t_L g5528 ( 
.A1(n_4778),
.A2(n_4039),
.B1(n_4077),
.B2(n_3972),
.Y(n_5528)
);

BUFx2_ASAP7_75t_L g5529 ( 
.A(n_4753),
.Y(n_5529)
);

BUFx6f_ASAP7_75t_L g5530 ( 
.A(n_4785),
.Y(n_5530)
);

OAI21x1_ASAP7_75t_L g5531 ( 
.A1(n_4685),
.A2(n_4065),
.B(n_4059),
.Y(n_5531)
);

NOR2x1_ASAP7_75t_L g5532 ( 
.A(n_4807),
.B(n_3018),
.Y(n_5532)
);

BUFx8_ASAP7_75t_SL g5533 ( 
.A(n_4628),
.Y(n_5533)
);

AND2x4_ASAP7_75t_L g5534 ( 
.A(n_4790),
.B(n_3020),
.Y(n_5534)
);

OAI22xp5_ASAP7_75t_L g5535 ( 
.A1(n_4791),
.A2(n_4022),
.B1(n_4034),
.B2(n_4010),
.Y(n_5535)
);

INVx4_ASAP7_75t_L g5536 ( 
.A(n_4792),
.Y(n_5536)
);

INVx3_ASAP7_75t_L g5537 ( 
.A(n_4793),
.Y(n_5537)
);

AND2x2_ASAP7_75t_L g5538 ( 
.A(n_4795),
.B(n_4080),
.Y(n_5538)
);

INVx3_ASAP7_75t_L g5539 ( 
.A(n_4801),
.Y(n_5539)
);

INVx2_ASAP7_75t_L g5540 ( 
.A(n_4806),
.Y(n_5540)
);

BUFx6f_ASAP7_75t_L g5541 ( 
.A(n_4809),
.Y(n_5541)
);

NAND2xp5_ASAP7_75t_L g5542 ( 
.A(n_4810),
.B(n_4093),
.Y(n_5542)
);

INVx1_ASAP7_75t_L g5543 ( 
.A(n_4813),
.Y(n_5543)
);

OAI22xp5_ASAP7_75t_L g5544 ( 
.A1(n_4815),
.A2(n_4049),
.B1(n_4050),
.B2(n_4048),
.Y(n_5544)
);

INVx2_ASAP7_75t_L g5545 ( 
.A(n_4816),
.Y(n_5545)
);

CKINVDCx8_ASAP7_75t_R g5546 ( 
.A(n_4832),
.Y(n_5546)
);

XNOR2xp5_ASAP7_75t_L g5547 ( 
.A(n_4630),
.B(n_4631),
.Y(n_5547)
);

INVx3_ASAP7_75t_L g5548 ( 
.A(n_4818),
.Y(n_5548)
);

INVx1_ASAP7_75t_L g5549 ( 
.A(n_4751),
.Y(n_5549)
);

BUFx6f_ASAP7_75t_L g5550 ( 
.A(n_4837),
.Y(n_5550)
);

INVx4_ASAP7_75t_L g5551 ( 
.A(n_4626),
.Y(n_5551)
);

INVx3_ASAP7_75t_L g5552 ( 
.A(n_4821),
.Y(n_5552)
);

INVx2_ASAP7_75t_L g5553 ( 
.A(n_4627),
.Y(n_5553)
);

AOI22xp5_ASAP7_75t_L g5554 ( 
.A1(n_4779),
.A2(n_4133),
.B1(n_4092),
.B2(n_4089),
.Y(n_5554)
);

AND2x2_ASAP7_75t_L g5555 ( 
.A(n_4823),
.B(n_4080),
.Y(n_5555)
);

AND2x6_ASAP7_75t_L g5556 ( 
.A(n_5071),
.B(n_3026),
.Y(n_5556)
);

AND2x4_ASAP7_75t_L g5557 ( 
.A(n_4762),
.B(n_3039),
.Y(n_5557)
);

INVx2_ASAP7_75t_L g5558 ( 
.A(n_5059),
.Y(n_5558)
);

NOR2xp33_ASAP7_75t_L g5559 ( 
.A(n_4644),
.B(n_4066),
.Y(n_5559)
);

INVx1_ASAP7_75t_L g5560 ( 
.A(n_5061),
.Y(n_5560)
);

INVx3_ASAP7_75t_L g5561 ( 
.A(n_4824),
.Y(n_5561)
);

INVx1_ASAP7_75t_L g5562 ( 
.A(n_5062),
.Y(n_5562)
);

AND2x2_ASAP7_75t_L g5563 ( 
.A(n_4829),
.B(n_4180),
.Y(n_5563)
);

AND2x2_ASAP7_75t_L g5564 ( 
.A(n_5063),
.B(n_2819),
.Y(n_5564)
);

INVx6_ASAP7_75t_L g5565 ( 
.A(n_4633),
.Y(n_5565)
);

NAND2xp5_ASAP7_75t_L g5566 ( 
.A(n_5066),
.B(n_4112),
.Y(n_5566)
);

INVx1_ASAP7_75t_L g5567 ( 
.A(n_5070),
.Y(n_5567)
);

INVx1_ASAP7_75t_L g5568 ( 
.A(n_5074),
.Y(n_5568)
);

NOR2xp33_ASAP7_75t_L g5569 ( 
.A(n_5077),
.B(n_4115),
.Y(n_5569)
);

INVx6_ASAP7_75t_L g5570 ( 
.A(n_4637),
.Y(n_5570)
);

INVx1_ASAP7_75t_L g5571 ( 
.A(n_5079),
.Y(n_5571)
);

NAND2xp5_ASAP7_75t_L g5572 ( 
.A(n_5083),
.B(n_4183),
.Y(n_5572)
);

CKINVDCx6p67_ASAP7_75t_R g5573 ( 
.A(n_4653),
.Y(n_5573)
);

INVx1_ASAP7_75t_L g5574 ( 
.A(n_5085),
.Y(n_5574)
);

NAND2xp5_ASAP7_75t_L g5575 ( 
.A(n_5091),
.B(n_4188),
.Y(n_5575)
);

INVx2_ASAP7_75t_L g5576 ( 
.A(n_5095),
.Y(n_5576)
);

INVx1_ASAP7_75t_L g5577 ( 
.A(n_5100),
.Y(n_5577)
);

NAND2x1p5_ASAP7_75t_L g5578 ( 
.A(n_5103),
.B(n_3050),
.Y(n_5578)
);

INVx1_ASAP7_75t_L g5579 ( 
.A(n_5106),
.Y(n_5579)
);

NAND2xp5_ASAP7_75t_L g5580 ( 
.A(n_5113),
.B(n_4191),
.Y(n_5580)
);

AND2x4_ASAP7_75t_L g5581 ( 
.A(n_4765),
.B(n_3051),
.Y(n_5581)
);

BUFx6f_ASAP7_75t_L g5582 ( 
.A(n_5114),
.Y(n_5582)
);

OA21x2_ASAP7_75t_L g5583 ( 
.A1(n_5119),
.A2(n_3061),
.B(n_3059),
.Y(n_5583)
);

INVx1_ASAP7_75t_L g5584 ( 
.A(n_4781),
.Y(n_5584)
);

BUFx6f_ASAP7_75t_L g5585 ( 
.A(n_4721),
.Y(n_5585)
);

INVx1_ASAP7_75t_L g5586 ( 
.A(n_4786),
.Y(n_5586)
);

INVx2_ASAP7_75t_L g5587 ( 
.A(n_4730),
.Y(n_5587)
);

INVx3_ASAP7_75t_L g5588 ( 
.A(n_4733),
.Y(n_5588)
);

INVxp33_ASAP7_75t_SL g5589 ( 
.A(n_4646),
.Y(n_5589)
);

CKINVDCx11_ASAP7_75t_R g5590 ( 
.A(n_5064),
.Y(n_5590)
);

INVx1_ASAP7_75t_L g5591 ( 
.A(n_4743),
.Y(n_5591)
);

OAI22xp5_ASAP7_75t_SL g5592 ( 
.A1(n_4747),
.A2(n_3562),
.B1(n_3582),
.B2(n_3550),
.Y(n_5592)
);

BUFx3_ASAP7_75t_L g5593 ( 
.A(n_4749),
.Y(n_5593)
);

OAI22xp5_ASAP7_75t_L g5594 ( 
.A1(n_5081),
.A2(n_4145),
.B1(n_4171),
.B2(n_4134),
.Y(n_5594)
);

INVx1_ASAP7_75t_L g5595 ( 
.A(n_5121),
.Y(n_5595)
);

INVxp67_ASAP7_75t_L g5596 ( 
.A(n_5089),
.Y(n_5596)
);

NAND2xp5_ASAP7_75t_SL g5597 ( 
.A(n_5117),
.B(n_2821),
.Y(n_5597)
);

INVx2_ASAP7_75t_L g5598 ( 
.A(n_5096),
.Y(n_5598)
);

INVx2_ASAP7_75t_L g5599 ( 
.A(n_5107),
.Y(n_5599)
);

NAND2xp5_ASAP7_75t_L g5600 ( 
.A(n_4916),
.B(n_3063),
.Y(n_5600)
);

HB1xp67_ASAP7_75t_L g5601 ( 
.A(n_4887),
.Y(n_5601)
);

BUFx3_ASAP7_75t_L g5602 ( 
.A(n_4690),
.Y(n_5602)
);

AOI22xp5_ASAP7_75t_L g5603 ( 
.A1(n_5099),
.A2(n_2830),
.B1(n_2832),
.B2(n_2829),
.Y(n_5603)
);

BUFx6f_ASAP7_75t_L g5604 ( 
.A(n_4917),
.Y(n_5604)
);

AND2x2_ASAP7_75t_L g5605 ( 
.A(n_4910),
.B(n_2833),
.Y(n_5605)
);

AND2x4_ASAP7_75t_L g5606 ( 
.A(n_4690),
.B(n_3065),
.Y(n_5606)
);

OAI22xp5_ASAP7_75t_SL g5607 ( 
.A1(n_4842),
.A2(n_3600),
.B1(n_3617),
.B2(n_3590),
.Y(n_5607)
);

INVx1_ASAP7_75t_L g5608 ( 
.A(n_4992),
.Y(n_5608)
);

INVx2_ASAP7_75t_L g5609 ( 
.A(n_4929),
.Y(n_5609)
);

INVx1_ASAP7_75t_L g5610 ( 
.A(n_4992),
.Y(n_5610)
);

NAND2xp5_ASAP7_75t_L g5611 ( 
.A(n_4916),
.B(n_3070),
.Y(n_5611)
);

XOR2xp5_ASAP7_75t_L g5612 ( 
.A(n_4621),
.B(n_3618),
.Y(n_5612)
);

INVx1_ASAP7_75t_L g5613 ( 
.A(n_4992),
.Y(n_5613)
);

INVx2_ASAP7_75t_L g5614 ( 
.A(n_4929),
.Y(n_5614)
);

AOI22xp5_ASAP7_75t_L g5615 ( 
.A1(n_5099),
.A2(n_2836),
.B1(n_2837),
.B2(n_2834),
.Y(n_5615)
);

INVx1_ASAP7_75t_L g5616 ( 
.A(n_4992),
.Y(n_5616)
);

OAI22xp5_ASAP7_75t_SL g5617 ( 
.A1(n_4842),
.A2(n_3644),
.B1(n_3645),
.B2(n_3632),
.Y(n_5617)
);

AOI22xp5_ASAP7_75t_L g5618 ( 
.A1(n_5099),
.A2(n_2844),
.B1(n_2845),
.B2(n_2839),
.Y(n_5618)
);

INVx2_ASAP7_75t_L g5619 ( 
.A(n_4929),
.Y(n_5619)
);

INVx1_ASAP7_75t_L g5620 ( 
.A(n_4992),
.Y(n_5620)
);

OAI22xp5_ASAP7_75t_L g5621 ( 
.A1(n_4924),
.A2(n_2849),
.B1(n_2850),
.B2(n_2846),
.Y(n_5621)
);

INVx1_ASAP7_75t_L g5622 ( 
.A(n_4992),
.Y(n_5622)
);

BUFx6f_ASAP7_75t_L g5623 ( 
.A(n_4917),
.Y(n_5623)
);

INVx5_ASAP7_75t_L g5624 ( 
.A(n_4850),
.Y(n_5624)
);

INVx1_ASAP7_75t_L g5625 ( 
.A(n_4992),
.Y(n_5625)
);

INVx1_ASAP7_75t_L g5626 ( 
.A(n_4992),
.Y(n_5626)
);

INVx4_ASAP7_75t_L g5627 ( 
.A(n_4869),
.Y(n_5627)
);

AND2x6_ASAP7_75t_L g5628 ( 
.A(n_4735),
.B(n_3072),
.Y(n_5628)
);

INVx2_ASAP7_75t_L g5629 ( 
.A(n_4929),
.Y(n_5629)
);

BUFx2_ASAP7_75t_L g5630 ( 
.A(n_4843),
.Y(n_5630)
);

NAND2xp5_ASAP7_75t_L g5631 ( 
.A(n_4916),
.B(n_3074),
.Y(n_5631)
);

INVx2_ASAP7_75t_L g5632 ( 
.A(n_4929),
.Y(n_5632)
);

NAND2xp5_ASAP7_75t_L g5633 ( 
.A(n_4916),
.B(n_3075),
.Y(n_5633)
);

INVx2_ASAP7_75t_L g5634 ( 
.A(n_4929),
.Y(n_5634)
);

INVx1_ASAP7_75t_L g5635 ( 
.A(n_4992),
.Y(n_5635)
);

INVx1_ASAP7_75t_L g5636 ( 
.A(n_4992),
.Y(n_5636)
);

NAND2xp5_ASAP7_75t_L g5637 ( 
.A(n_4916),
.B(n_3077),
.Y(n_5637)
);

NAND2xp5_ASAP7_75t_L g5638 ( 
.A(n_4916),
.B(n_3085),
.Y(n_5638)
);

BUFx8_ASAP7_75t_L g5639 ( 
.A(n_4723),
.Y(n_5639)
);

AND2x4_ASAP7_75t_L g5640 ( 
.A(n_4690),
.B(n_3090),
.Y(n_5640)
);

BUFx3_ASAP7_75t_L g5641 ( 
.A(n_4690),
.Y(n_5641)
);

AND2x2_ASAP7_75t_SL g5642 ( 
.A(n_4850),
.B(n_3098),
.Y(n_5642)
);

INVx1_ASAP7_75t_L g5643 ( 
.A(n_4992),
.Y(n_5643)
);

NAND2xp33_ASAP7_75t_L g5644 ( 
.A(n_4981),
.B(n_2855),
.Y(n_5644)
);

NAND2xp5_ASAP7_75t_L g5645 ( 
.A(n_4916),
.B(n_3101),
.Y(n_5645)
);

INVx6_ASAP7_75t_L g5646 ( 
.A(n_4982),
.Y(n_5646)
);

HB1xp67_ASAP7_75t_L g5647 ( 
.A(n_4887),
.Y(n_5647)
);

BUFx6f_ASAP7_75t_L g5648 ( 
.A(n_4917),
.Y(n_5648)
);

INVx2_ASAP7_75t_L g5649 ( 
.A(n_4929),
.Y(n_5649)
);

OAI22xp5_ASAP7_75t_SL g5650 ( 
.A1(n_4842),
.A2(n_3665),
.B1(n_3680),
.B2(n_3653),
.Y(n_5650)
);

NOR2x1_ASAP7_75t_L g5651 ( 
.A(n_4921),
.B(n_3103),
.Y(n_5651)
);

NAND2xp5_ASAP7_75t_L g5652 ( 
.A(n_4916),
.B(n_3113),
.Y(n_5652)
);

OAI22xp5_ASAP7_75t_SL g5653 ( 
.A1(n_4842),
.A2(n_3701),
.B1(n_3728),
.B2(n_3687),
.Y(n_5653)
);

BUFx6f_ASAP7_75t_L g5654 ( 
.A(n_4917),
.Y(n_5654)
);

INVx3_ASAP7_75t_L g5655 ( 
.A(n_4917),
.Y(n_5655)
);

BUFx6f_ASAP7_75t_L g5656 ( 
.A(n_4917),
.Y(n_5656)
);

OAI21x1_ASAP7_75t_L g5657 ( 
.A1(n_4937),
.A2(n_3129),
.B(n_3121),
.Y(n_5657)
);

INVx1_ASAP7_75t_L g5658 ( 
.A(n_4992),
.Y(n_5658)
);

INVx1_ASAP7_75t_L g5659 ( 
.A(n_4992),
.Y(n_5659)
);

INVx2_ASAP7_75t_SL g5660 ( 
.A(n_4887),
.Y(n_5660)
);

INVx1_ASAP7_75t_L g5661 ( 
.A(n_4992),
.Y(n_5661)
);

INVx1_ASAP7_75t_L g5662 ( 
.A(n_4992),
.Y(n_5662)
);

INVx2_ASAP7_75t_L g5663 ( 
.A(n_4929),
.Y(n_5663)
);

NAND2xp5_ASAP7_75t_L g5664 ( 
.A(n_4916),
.B(n_3133),
.Y(n_5664)
);

INVx1_ASAP7_75t_L g5665 ( 
.A(n_4992),
.Y(n_5665)
);

INVx1_ASAP7_75t_L g5666 ( 
.A(n_4992),
.Y(n_5666)
);

AOI22xp5_ASAP7_75t_L g5667 ( 
.A1(n_5099),
.A2(n_2857),
.B1(n_2863),
.B2(n_2856),
.Y(n_5667)
);

AND2x4_ASAP7_75t_L g5668 ( 
.A(n_4690),
.B(n_3138),
.Y(n_5668)
);

INVx1_ASAP7_75t_L g5669 ( 
.A(n_4992),
.Y(n_5669)
);

BUFx6f_ASAP7_75t_L g5670 ( 
.A(n_4917),
.Y(n_5670)
);

INVx2_ASAP7_75t_L g5671 ( 
.A(n_4929),
.Y(n_5671)
);

AND2x2_ASAP7_75t_L g5672 ( 
.A(n_4910),
.B(n_2865),
.Y(n_5672)
);

INVx1_ASAP7_75t_L g5673 ( 
.A(n_4992),
.Y(n_5673)
);

AOI22xp5_ASAP7_75t_L g5674 ( 
.A1(n_5099),
.A2(n_2870),
.B1(n_2878),
.B2(n_2867),
.Y(n_5674)
);

INVx1_ASAP7_75t_L g5675 ( 
.A(n_4992),
.Y(n_5675)
);

INVxp67_ASAP7_75t_L g5676 ( 
.A(n_4887),
.Y(n_5676)
);

AOI22xp5_ASAP7_75t_L g5677 ( 
.A1(n_5099),
.A2(n_2883),
.B1(n_2885),
.B2(n_2879),
.Y(n_5677)
);

INVx2_ASAP7_75t_SL g5678 ( 
.A(n_4887),
.Y(n_5678)
);

INVx1_ASAP7_75t_L g5679 ( 
.A(n_4992),
.Y(n_5679)
);

NAND2xp5_ASAP7_75t_L g5680 ( 
.A(n_4916),
.B(n_3140),
.Y(n_5680)
);

INVx3_ASAP7_75t_L g5681 ( 
.A(n_4917),
.Y(n_5681)
);

OA21x2_ASAP7_75t_L g5682 ( 
.A1(n_4937),
.A2(n_3143),
.B(n_3142),
.Y(n_5682)
);

CKINVDCx5p33_ASAP7_75t_R g5683 ( 
.A(n_4634),
.Y(n_5683)
);

INVx2_ASAP7_75t_L g5684 ( 
.A(n_4929),
.Y(n_5684)
);

INVx1_ASAP7_75t_L g5685 ( 
.A(n_4992),
.Y(n_5685)
);

BUFx6f_ASAP7_75t_L g5686 ( 
.A(n_4917),
.Y(n_5686)
);

HB1xp67_ASAP7_75t_L g5687 ( 
.A(n_4887),
.Y(n_5687)
);

AND2x4_ASAP7_75t_L g5688 ( 
.A(n_4690),
.B(n_3152),
.Y(n_5688)
);

AND2x2_ASAP7_75t_L g5689 ( 
.A(n_4910),
.B(n_2886),
.Y(n_5689)
);

INVx1_ASAP7_75t_L g5690 ( 
.A(n_4992),
.Y(n_5690)
);

INVx1_ASAP7_75t_L g5691 ( 
.A(n_4992),
.Y(n_5691)
);

INVx1_ASAP7_75t_L g5692 ( 
.A(n_4992),
.Y(n_5692)
);

BUFx8_ASAP7_75t_L g5693 ( 
.A(n_4723),
.Y(n_5693)
);

AND2x2_ASAP7_75t_SL g5694 ( 
.A(n_4850),
.B(n_3153),
.Y(n_5694)
);

AND2x4_ASAP7_75t_L g5695 ( 
.A(n_4690),
.B(n_3157),
.Y(n_5695)
);

INVx1_ASAP7_75t_L g5696 ( 
.A(n_4992),
.Y(n_5696)
);

AND2x4_ASAP7_75t_L g5697 ( 
.A(n_4690),
.B(n_3180),
.Y(n_5697)
);

NAND2xp5_ASAP7_75t_L g5698 ( 
.A(n_4916),
.B(n_3181),
.Y(n_5698)
);

NOR2xp33_ASAP7_75t_R g5699 ( 
.A(n_5152),
.B(n_3785),
.Y(n_5699)
);

INVx1_ASAP7_75t_L g5700 ( 
.A(n_5125),
.Y(n_5700)
);

CKINVDCx20_ASAP7_75t_R g5701 ( 
.A(n_5533),
.Y(n_5701)
);

INVx3_ASAP7_75t_L g5702 ( 
.A(n_5198),
.Y(n_5702)
);

NAND2xp33_ASAP7_75t_R g5703 ( 
.A(n_5502),
.B(n_2891),
.Y(n_5703)
);

BUFx2_ASAP7_75t_L g5704 ( 
.A(n_5676),
.Y(n_5704)
);

INVx1_ASAP7_75t_L g5705 ( 
.A(n_5690),
.Y(n_5705)
);

INVx1_ASAP7_75t_L g5706 ( 
.A(n_5691),
.Y(n_5706)
);

INVx3_ASAP7_75t_L g5707 ( 
.A(n_5200),
.Y(n_5707)
);

INVx2_ASAP7_75t_L g5708 ( 
.A(n_5173),
.Y(n_5708)
);

NAND2xp33_ASAP7_75t_R g5709 ( 
.A(n_5215),
.B(n_2895),
.Y(n_5709)
);

CKINVDCx5p33_ASAP7_75t_R g5710 ( 
.A(n_5292),
.Y(n_5710)
);

INVx2_ASAP7_75t_L g5711 ( 
.A(n_5185),
.Y(n_5711)
);

CKINVDCx20_ASAP7_75t_R g5712 ( 
.A(n_5590),
.Y(n_5712)
);

CKINVDCx5p33_ASAP7_75t_R g5713 ( 
.A(n_5459),
.Y(n_5713)
);

INVx3_ASAP7_75t_L g5714 ( 
.A(n_5188),
.Y(n_5714)
);

INVx2_ASAP7_75t_L g5715 ( 
.A(n_5157),
.Y(n_5715)
);

BUFx6f_ASAP7_75t_L g5716 ( 
.A(n_5148),
.Y(n_5716)
);

CKINVDCx16_ASAP7_75t_R g5717 ( 
.A(n_5513),
.Y(n_5717)
);

CKINVDCx5p33_ASAP7_75t_R g5718 ( 
.A(n_5683),
.Y(n_5718)
);

INVx1_ASAP7_75t_L g5719 ( 
.A(n_5685),
.Y(n_5719)
);

INVx2_ASAP7_75t_L g5720 ( 
.A(n_5159),
.Y(n_5720)
);

INVx1_ASAP7_75t_L g5721 ( 
.A(n_5692),
.Y(n_5721)
);

CKINVDCx20_ASAP7_75t_R g5722 ( 
.A(n_5573),
.Y(n_5722)
);

HB1xp67_ASAP7_75t_L g5723 ( 
.A(n_5660),
.Y(n_5723)
);

CKINVDCx5p33_ASAP7_75t_R g5724 ( 
.A(n_5452),
.Y(n_5724)
);

CKINVDCx5p33_ASAP7_75t_R g5725 ( 
.A(n_5589),
.Y(n_5725)
);

CKINVDCx5p33_ASAP7_75t_R g5726 ( 
.A(n_5439),
.Y(n_5726)
);

NAND2xp5_ASAP7_75t_SL g5727 ( 
.A(n_5195),
.B(n_2897),
.Y(n_5727)
);

NAND2xp33_ASAP7_75t_R g5728 ( 
.A(n_5135),
.B(n_2898),
.Y(n_5728)
);

CKINVDCx5p33_ASAP7_75t_R g5729 ( 
.A(n_5319),
.Y(n_5729)
);

INVx2_ASAP7_75t_SL g5730 ( 
.A(n_5678),
.Y(n_5730)
);

INVx1_ASAP7_75t_L g5731 ( 
.A(n_5140),
.Y(n_5731)
);

CKINVDCx5p33_ASAP7_75t_R g5732 ( 
.A(n_5547),
.Y(n_5732)
);

INVx2_ASAP7_75t_L g5733 ( 
.A(n_5160),
.Y(n_5733)
);

CKINVDCx5p33_ASAP7_75t_R g5734 ( 
.A(n_5480),
.Y(n_5734)
);

CKINVDCx20_ASAP7_75t_R g5735 ( 
.A(n_5315),
.Y(n_5735)
);

CKINVDCx5p33_ASAP7_75t_R g5736 ( 
.A(n_5501),
.Y(n_5736)
);

CKINVDCx5p33_ASAP7_75t_R g5737 ( 
.A(n_5509),
.Y(n_5737)
);

NOR2x1p5_ASAP7_75t_L g5738 ( 
.A(n_5153),
.B(n_2902),
.Y(n_5738)
);

CKINVDCx5p33_ASAP7_75t_R g5739 ( 
.A(n_5530),
.Y(n_5739)
);

CKINVDCx5p33_ASAP7_75t_R g5740 ( 
.A(n_5541),
.Y(n_5740)
);

CKINVDCx5p33_ASAP7_75t_R g5741 ( 
.A(n_5630),
.Y(n_5741)
);

CKINVDCx5p33_ASAP7_75t_R g5742 ( 
.A(n_5582),
.Y(n_5742)
);

INVx2_ASAP7_75t_L g5743 ( 
.A(n_5410),
.Y(n_5743)
);

CKINVDCx5p33_ASAP7_75t_R g5744 ( 
.A(n_5565),
.Y(n_5744)
);

CKINVDCx20_ASAP7_75t_R g5745 ( 
.A(n_5328),
.Y(n_5745)
);

CKINVDCx5p33_ASAP7_75t_R g5746 ( 
.A(n_5570),
.Y(n_5746)
);

INVx1_ASAP7_75t_L g5747 ( 
.A(n_5142),
.Y(n_5747)
);

AND2x2_ASAP7_75t_L g5748 ( 
.A(n_5145),
.B(n_3787),
.Y(n_5748)
);

INVx2_ASAP7_75t_L g5749 ( 
.A(n_5419),
.Y(n_5749)
);

INVxp67_ASAP7_75t_L g5750 ( 
.A(n_5601),
.Y(n_5750)
);

CKINVDCx5p33_ASAP7_75t_R g5751 ( 
.A(n_5536),
.Y(n_5751)
);

CKINVDCx6p67_ASAP7_75t_R g5752 ( 
.A(n_5624),
.Y(n_5752)
);

NOR2xp33_ASAP7_75t_R g5753 ( 
.A(n_5546),
.B(n_3826),
.Y(n_5753)
);

NOR2xp33_ASAP7_75t_R g5754 ( 
.A(n_5552),
.B(n_5561),
.Y(n_5754)
);

CKINVDCx5p33_ASAP7_75t_R g5755 ( 
.A(n_5647),
.Y(n_5755)
);

INVx2_ASAP7_75t_L g5756 ( 
.A(n_5379),
.Y(n_5756)
);

INVx2_ASAP7_75t_SL g5757 ( 
.A(n_5687),
.Y(n_5757)
);

HB1xp67_ASAP7_75t_L g5758 ( 
.A(n_5134),
.Y(n_5758)
);

CKINVDCx5p33_ASAP7_75t_R g5759 ( 
.A(n_5424),
.Y(n_5759)
);

INVx1_ASAP7_75t_L g5760 ( 
.A(n_5696),
.Y(n_5760)
);

CKINVDCx5p33_ASAP7_75t_R g5761 ( 
.A(n_5593),
.Y(n_5761)
);

INVx1_ASAP7_75t_L g5762 ( 
.A(n_5143),
.Y(n_5762)
);

INVx2_ASAP7_75t_L g5763 ( 
.A(n_5380),
.Y(n_5763)
);

BUFx6f_ASAP7_75t_L g5764 ( 
.A(n_5154),
.Y(n_5764)
);

INVx1_ASAP7_75t_L g5765 ( 
.A(n_5156),
.Y(n_5765)
);

CKINVDCx5p33_ASAP7_75t_R g5766 ( 
.A(n_5504),
.Y(n_5766)
);

BUFx6f_ASAP7_75t_L g5767 ( 
.A(n_5124),
.Y(n_5767)
);

CKINVDCx5p33_ASAP7_75t_R g5768 ( 
.A(n_5507),
.Y(n_5768)
);

CKINVDCx5p33_ASAP7_75t_R g5769 ( 
.A(n_5512),
.Y(n_5769)
);

INVx2_ASAP7_75t_L g5770 ( 
.A(n_5406),
.Y(n_5770)
);

CKINVDCx5p33_ASAP7_75t_R g5771 ( 
.A(n_5525),
.Y(n_5771)
);

INVx2_ASAP7_75t_L g5772 ( 
.A(n_5407),
.Y(n_5772)
);

CKINVDCx5p33_ASAP7_75t_R g5773 ( 
.A(n_5537),
.Y(n_5773)
);

INVx1_ASAP7_75t_L g5774 ( 
.A(n_5163),
.Y(n_5774)
);

CKINVDCx5p33_ASAP7_75t_R g5775 ( 
.A(n_5539),
.Y(n_5775)
);

AOI22xp5_ASAP7_75t_L g5776 ( 
.A1(n_5208),
.A2(n_5172),
.B1(n_5162),
.B2(n_5179),
.Y(n_5776)
);

CKINVDCx5p33_ASAP7_75t_R g5777 ( 
.A(n_5548),
.Y(n_5777)
);

INVx2_ASAP7_75t_L g5778 ( 
.A(n_5221),
.Y(n_5778)
);

INVx1_ASAP7_75t_L g5779 ( 
.A(n_5165),
.Y(n_5779)
);

CKINVDCx5p33_ASAP7_75t_R g5780 ( 
.A(n_5551),
.Y(n_5780)
);

INVx1_ASAP7_75t_SL g5781 ( 
.A(n_5360),
.Y(n_5781)
);

BUFx6f_ASAP7_75t_L g5782 ( 
.A(n_5128),
.Y(n_5782)
);

BUFx10_ASAP7_75t_L g5783 ( 
.A(n_5569),
.Y(n_5783)
);

CKINVDCx5p33_ASAP7_75t_R g5784 ( 
.A(n_5585),
.Y(n_5784)
);

CKINVDCx5p33_ASAP7_75t_R g5785 ( 
.A(n_5164),
.Y(n_5785)
);

CKINVDCx5p33_ASAP7_75t_R g5786 ( 
.A(n_5529),
.Y(n_5786)
);

INVx3_ASAP7_75t_L g5787 ( 
.A(n_5682),
.Y(n_5787)
);

CKINVDCx5p33_ASAP7_75t_R g5788 ( 
.A(n_5146),
.Y(n_5788)
);

INVx2_ASAP7_75t_L g5789 ( 
.A(n_5231),
.Y(n_5789)
);

INVx1_ASAP7_75t_L g5790 ( 
.A(n_5167),
.Y(n_5790)
);

CKINVDCx5p33_ASAP7_75t_R g5791 ( 
.A(n_5168),
.Y(n_5791)
);

CKINVDCx5p33_ASAP7_75t_R g5792 ( 
.A(n_5203),
.Y(n_5792)
);

INVx3_ASAP7_75t_L g5793 ( 
.A(n_5130),
.Y(n_5793)
);

BUFx2_ASAP7_75t_L g5794 ( 
.A(n_5473),
.Y(n_5794)
);

CKINVDCx20_ASAP7_75t_R g5795 ( 
.A(n_5516),
.Y(n_5795)
);

INVx2_ASAP7_75t_L g5796 ( 
.A(n_5233),
.Y(n_5796)
);

CKINVDCx5p33_ASAP7_75t_R g5797 ( 
.A(n_5627),
.Y(n_5797)
);

INVx1_ASAP7_75t_L g5798 ( 
.A(n_5170),
.Y(n_5798)
);

INVx1_ASAP7_75t_L g5799 ( 
.A(n_5180),
.Y(n_5799)
);

CKINVDCx5p33_ASAP7_75t_R g5800 ( 
.A(n_5550),
.Y(n_5800)
);

INVx2_ASAP7_75t_L g5801 ( 
.A(n_5235),
.Y(n_5801)
);

NAND2xp33_ASAP7_75t_R g5802 ( 
.A(n_5415),
.B(n_2906),
.Y(n_5802)
);

CKINVDCx5p33_ASAP7_75t_R g5803 ( 
.A(n_5179),
.Y(n_5803)
);

BUFx10_ASAP7_75t_L g5804 ( 
.A(n_5559),
.Y(n_5804)
);

INVx1_ASAP7_75t_L g5805 ( 
.A(n_5181),
.Y(n_5805)
);

INVx2_ASAP7_75t_L g5806 ( 
.A(n_5238),
.Y(n_5806)
);

CKINVDCx5p33_ASAP7_75t_R g5807 ( 
.A(n_5442),
.Y(n_5807)
);

NOR2xp33_ASAP7_75t_R g5808 ( 
.A(n_5588),
.B(n_3836),
.Y(n_5808)
);

CKINVDCx5p33_ASAP7_75t_R g5809 ( 
.A(n_5139),
.Y(n_5809)
);

BUFx6f_ASAP7_75t_L g5810 ( 
.A(n_5604),
.Y(n_5810)
);

INVxp33_ASAP7_75t_SL g5811 ( 
.A(n_5612),
.Y(n_5811)
);

CKINVDCx5p33_ASAP7_75t_R g5812 ( 
.A(n_5191),
.Y(n_5812)
);

CKINVDCx5p33_ASAP7_75t_R g5813 ( 
.A(n_5639),
.Y(n_5813)
);

INVx1_ASAP7_75t_L g5814 ( 
.A(n_5187),
.Y(n_5814)
);

CKINVDCx5p33_ASAP7_75t_R g5815 ( 
.A(n_5693),
.Y(n_5815)
);

INVx2_ASAP7_75t_L g5816 ( 
.A(n_5240),
.Y(n_5816)
);

INVx2_ASAP7_75t_L g5817 ( 
.A(n_5244),
.Y(n_5817)
);

NOR2xp33_ASAP7_75t_L g5818 ( 
.A(n_5127),
.B(n_2907),
.Y(n_5818)
);

CKINVDCx5p33_ASAP7_75t_R g5819 ( 
.A(n_5351),
.Y(n_5819)
);

INVx1_ASAP7_75t_L g5820 ( 
.A(n_5190),
.Y(n_5820)
);

NOR2xp33_ASAP7_75t_R g5821 ( 
.A(n_5474),
.B(n_3851),
.Y(n_5821)
);

BUFx2_ASAP7_75t_L g5822 ( 
.A(n_5177),
.Y(n_5822)
);

BUFx3_ASAP7_75t_L g5823 ( 
.A(n_5133),
.Y(n_5823)
);

CKINVDCx20_ASAP7_75t_R g5824 ( 
.A(n_5178),
.Y(n_5824)
);

CKINVDCx20_ASAP7_75t_R g5825 ( 
.A(n_5486),
.Y(n_5825)
);

INVx3_ASAP7_75t_L g5826 ( 
.A(n_5131),
.Y(n_5826)
);

CKINVDCx5p33_ASAP7_75t_R g5827 ( 
.A(n_5265),
.Y(n_5827)
);

CKINVDCx5p33_ASAP7_75t_R g5828 ( 
.A(n_5392),
.Y(n_5828)
);

CKINVDCx5p33_ASAP7_75t_R g5829 ( 
.A(n_5405),
.Y(n_5829)
);

INVx1_ASAP7_75t_L g5830 ( 
.A(n_5193),
.Y(n_5830)
);

CKINVDCx20_ASAP7_75t_R g5831 ( 
.A(n_5273),
.Y(n_5831)
);

CKINVDCx20_ASAP7_75t_R g5832 ( 
.A(n_5276),
.Y(n_5832)
);

INVx2_ASAP7_75t_L g5833 ( 
.A(n_5251),
.Y(n_5833)
);

NAND2xp5_ASAP7_75t_L g5834 ( 
.A(n_5426),
.B(n_2908),
.Y(n_5834)
);

INVx1_ASAP7_75t_L g5835 ( 
.A(n_5197),
.Y(n_5835)
);

INVx1_ASAP7_75t_L g5836 ( 
.A(n_5211),
.Y(n_5836)
);

INVx2_ASAP7_75t_L g5837 ( 
.A(n_5253),
.Y(n_5837)
);

CKINVDCx5p33_ASAP7_75t_R g5838 ( 
.A(n_5510),
.Y(n_5838)
);

CKINVDCx5p33_ASAP7_75t_R g5839 ( 
.A(n_5519),
.Y(n_5839)
);

CKINVDCx5p33_ASAP7_75t_R g5840 ( 
.A(n_5540),
.Y(n_5840)
);

NOR2xp33_ASAP7_75t_R g5841 ( 
.A(n_5484),
.B(n_5464),
.Y(n_5841)
);

NAND2xp33_ASAP7_75t_R g5842 ( 
.A(n_5557),
.B(n_5581),
.Y(n_5842)
);

XOR2xp5_ASAP7_75t_L g5843 ( 
.A(n_5248),
.B(n_3911),
.Y(n_5843)
);

CKINVDCx20_ASAP7_75t_R g5844 ( 
.A(n_5299),
.Y(n_5844)
);

NAND2xp33_ASAP7_75t_R g5845 ( 
.A(n_5583),
.B(n_2909),
.Y(n_5845)
);

CKINVDCx5p33_ASAP7_75t_R g5846 ( 
.A(n_5545),
.Y(n_5846)
);

INVx1_ASAP7_75t_L g5847 ( 
.A(n_5219),
.Y(n_5847)
);

CKINVDCx5p33_ASAP7_75t_R g5848 ( 
.A(n_5192),
.Y(n_5848)
);

INVx3_ASAP7_75t_L g5849 ( 
.A(n_5137),
.Y(n_5849)
);

NOR2xp67_ASAP7_75t_L g5850 ( 
.A(n_5224),
.B(n_2910),
.Y(n_5850)
);

CKINVDCx5p33_ASAP7_75t_R g5851 ( 
.A(n_5216),
.Y(n_5851)
);

CKINVDCx20_ASAP7_75t_R g5852 ( 
.A(n_5345),
.Y(n_5852)
);

CKINVDCx5p33_ASAP7_75t_R g5853 ( 
.A(n_5646),
.Y(n_5853)
);

CKINVDCx5p33_ASAP7_75t_R g5854 ( 
.A(n_5602),
.Y(n_5854)
);

CKINVDCx5p33_ASAP7_75t_R g5855 ( 
.A(n_5641),
.Y(n_5855)
);

INVx1_ASAP7_75t_L g5856 ( 
.A(n_5230),
.Y(n_5856)
);

AND3x2_ASAP7_75t_L g5857 ( 
.A(n_5467),
.B(n_3185),
.C(n_3184),
.Y(n_5857)
);

CKINVDCx5p33_ASAP7_75t_R g5858 ( 
.A(n_5553),
.Y(n_5858)
);

CKINVDCx5p33_ASAP7_75t_R g5859 ( 
.A(n_5558),
.Y(n_5859)
);

CKINVDCx5p33_ASAP7_75t_R g5860 ( 
.A(n_5576),
.Y(n_5860)
);

INVx1_ASAP7_75t_L g5861 ( 
.A(n_5237),
.Y(n_5861)
);

INVx2_ASAP7_75t_L g5862 ( 
.A(n_5256),
.Y(n_5862)
);

CKINVDCx5p33_ASAP7_75t_R g5863 ( 
.A(n_5466),
.Y(n_5863)
);

INVx1_ASAP7_75t_L g5864 ( 
.A(n_5249),
.Y(n_5864)
);

INVx1_ASAP7_75t_L g5865 ( 
.A(n_5608),
.Y(n_5865)
);

NAND2xp33_ASAP7_75t_R g5866 ( 
.A(n_5492),
.B(n_2911),
.Y(n_5866)
);

NOR2xp67_ASAP7_75t_L g5867 ( 
.A(n_5268),
.B(n_2912),
.Y(n_5867)
);

INVx1_ASAP7_75t_L g5868 ( 
.A(n_5610),
.Y(n_5868)
);

CKINVDCx5p33_ASAP7_75t_R g5869 ( 
.A(n_5499),
.Y(n_5869)
);

CKINVDCx5p33_ASAP7_75t_R g5870 ( 
.A(n_5514),
.Y(n_5870)
);

CKINVDCx5p33_ASAP7_75t_R g5871 ( 
.A(n_5518),
.Y(n_5871)
);

CKINVDCx20_ASAP7_75t_R g5872 ( 
.A(n_5596),
.Y(n_5872)
);

BUFx3_ASAP7_75t_L g5873 ( 
.A(n_5174),
.Y(n_5873)
);

INVx2_ASAP7_75t_L g5874 ( 
.A(n_5266),
.Y(n_5874)
);

INVx3_ASAP7_75t_L g5875 ( 
.A(n_5147),
.Y(n_5875)
);

CKINVDCx5p33_ASAP7_75t_R g5876 ( 
.A(n_5521),
.Y(n_5876)
);

AOI22xp5_ASAP7_75t_L g5877 ( 
.A1(n_5208),
.A2(n_3948),
.B1(n_4019),
.B2(n_3934),
.Y(n_5877)
);

INVx1_ASAP7_75t_SL g5878 ( 
.A(n_5206),
.Y(n_5878)
);

INVx2_ASAP7_75t_L g5879 ( 
.A(n_5270),
.Y(n_5879)
);

CKINVDCx20_ASAP7_75t_R g5880 ( 
.A(n_5434),
.Y(n_5880)
);

CKINVDCx20_ASAP7_75t_R g5881 ( 
.A(n_5457),
.Y(n_5881)
);

CKINVDCx11_ASAP7_75t_R g5882 ( 
.A(n_5587),
.Y(n_5882)
);

CKINVDCx5p33_ASAP7_75t_R g5883 ( 
.A(n_5522),
.Y(n_5883)
);

INVx1_ASAP7_75t_L g5884 ( 
.A(n_5613),
.Y(n_5884)
);

INVxp33_ASAP7_75t_SL g5885 ( 
.A(n_5592),
.Y(n_5885)
);

CKINVDCx5p33_ASAP7_75t_R g5886 ( 
.A(n_5523),
.Y(n_5886)
);

CKINVDCx5p33_ASAP7_75t_R g5887 ( 
.A(n_5524),
.Y(n_5887)
);

INVxp33_ASAP7_75t_SL g5888 ( 
.A(n_5520),
.Y(n_5888)
);

CKINVDCx5p33_ASAP7_75t_R g5889 ( 
.A(n_5543),
.Y(n_5889)
);

INVx1_ASAP7_75t_L g5890 ( 
.A(n_5616),
.Y(n_5890)
);

INVx1_ASAP7_75t_L g5891 ( 
.A(n_5620),
.Y(n_5891)
);

CKINVDCx5p33_ASAP7_75t_R g5892 ( 
.A(n_5560),
.Y(n_5892)
);

CKINVDCx5p33_ASAP7_75t_R g5893 ( 
.A(n_5562),
.Y(n_5893)
);

OAI22xp33_ASAP7_75t_L g5894 ( 
.A1(n_5600),
.A2(n_4033),
.B1(n_4035),
.B2(n_4032),
.Y(n_5894)
);

CKINVDCx20_ASAP7_75t_R g5895 ( 
.A(n_5213),
.Y(n_5895)
);

CKINVDCx5p33_ASAP7_75t_R g5896 ( 
.A(n_5567),
.Y(n_5896)
);

INVx1_ASAP7_75t_L g5897 ( 
.A(n_5622),
.Y(n_5897)
);

CKINVDCx20_ASAP7_75t_R g5898 ( 
.A(n_5491),
.Y(n_5898)
);

NOR2xp67_ASAP7_75t_L g5899 ( 
.A(n_5549),
.B(n_2915),
.Y(n_5899)
);

CKINVDCx20_ASAP7_75t_R g5900 ( 
.A(n_5515),
.Y(n_5900)
);

INVx1_ASAP7_75t_L g5901 ( 
.A(n_5625),
.Y(n_5901)
);

CKINVDCx5p33_ASAP7_75t_R g5902 ( 
.A(n_5568),
.Y(n_5902)
);

CKINVDCx5p33_ASAP7_75t_R g5903 ( 
.A(n_5571),
.Y(n_5903)
);

CKINVDCx5p33_ASAP7_75t_R g5904 ( 
.A(n_5574),
.Y(n_5904)
);

INVx1_ASAP7_75t_L g5905 ( 
.A(n_5626),
.Y(n_5905)
);

NOR2xp33_ASAP7_75t_L g5906 ( 
.A(n_5217),
.B(n_2916),
.Y(n_5906)
);

BUFx2_ASAP7_75t_L g5907 ( 
.A(n_5129),
.Y(n_5907)
);

INVx1_ASAP7_75t_L g5908 ( 
.A(n_5635),
.Y(n_5908)
);

NOR2xp33_ASAP7_75t_R g5909 ( 
.A(n_5644),
.B(n_4040),
.Y(n_5909)
);

CKINVDCx20_ASAP7_75t_R g5910 ( 
.A(n_5591),
.Y(n_5910)
);

BUFx10_ASAP7_75t_L g5911 ( 
.A(n_5449),
.Y(n_5911)
);

NOR2xp33_ASAP7_75t_R g5912 ( 
.A(n_5577),
.B(n_4052),
.Y(n_5912)
);

CKINVDCx20_ASAP7_75t_R g5913 ( 
.A(n_5584),
.Y(n_5913)
);

NOR2xp33_ASAP7_75t_R g5914 ( 
.A(n_5579),
.B(n_4063),
.Y(n_5914)
);

BUFx2_ASAP7_75t_L g5915 ( 
.A(n_5246),
.Y(n_5915)
);

CKINVDCx5p33_ASAP7_75t_R g5916 ( 
.A(n_5443),
.Y(n_5916)
);

CKINVDCx5p33_ASAP7_75t_R g5917 ( 
.A(n_5598),
.Y(n_5917)
);

CKINVDCx20_ASAP7_75t_R g5918 ( 
.A(n_5586),
.Y(n_5918)
);

CKINVDCx5p33_ASAP7_75t_R g5919 ( 
.A(n_5599),
.Y(n_5919)
);

INVxp67_ASAP7_75t_L g5920 ( 
.A(n_5123),
.Y(n_5920)
);

INVx2_ASAP7_75t_L g5921 ( 
.A(n_5271),
.Y(n_5921)
);

INVx2_ASAP7_75t_L g5922 ( 
.A(n_5275),
.Y(n_5922)
);

INVx3_ASAP7_75t_L g5923 ( 
.A(n_5182),
.Y(n_5923)
);

INVx2_ASAP7_75t_L g5924 ( 
.A(n_5282),
.Y(n_5924)
);

CKINVDCx5p33_ASAP7_75t_R g5925 ( 
.A(n_5595),
.Y(n_5925)
);

CKINVDCx5p33_ASAP7_75t_R g5926 ( 
.A(n_5564),
.Y(n_5926)
);

BUFx6f_ASAP7_75t_L g5927 ( 
.A(n_5623),
.Y(n_5927)
);

CKINVDCx20_ASAP7_75t_R g5928 ( 
.A(n_5488),
.Y(n_5928)
);

INVx1_ASAP7_75t_L g5929 ( 
.A(n_5636),
.Y(n_5929)
);

INVx1_ASAP7_75t_L g5930 ( 
.A(n_5643),
.Y(n_5930)
);

CKINVDCx5p33_ASAP7_75t_R g5931 ( 
.A(n_5155),
.Y(n_5931)
);

CKINVDCx20_ASAP7_75t_R g5932 ( 
.A(n_5458),
.Y(n_5932)
);

CKINVDCx5p33_ASAP7_75t_R g5933 ( 
.A(n_5176),
.Y(n_5933)
);

CKINVDCx20_ASAP7_75t_R g5934 ( 
.A(n_5288),
.Y(n_5934)
);

BUFx2_ASAP7_75t_L g5935 ( 
.A(n_5246),
.Y(n_5935)
);

CKINVDCx5p33_ASAP7_75t_R g5936 ( 
.A(n_5171),
.Y(n_5936)
);

CKINVDCx5p33_ASAP7_75t_R g5937 ( 
.A(n_5171),
.Y(n_5937)
);

CKINVDCx20_ASAP7_75t_R g5938 ( 
.A(n_5388),
.Y(n_5938)
);

NOR2xp33_ASAP7_75t_R g5939 ( 
.A(n_5429),
.B(n_4085),
.Y(n_5939)
);

CKINVDCx20_ASAP7_75t_R g5940 ( 
.A(n_5597),
.Y(n_5940)
);

AND3x2_ASAP7_75t_L g5941 ( 
.A(n_5166),
.B(n_3201),
.C(n_3188),
.Y(n_5941)
);

INVx1_ASAP7_75t_L g5942 ( 
.A(n_5658),
.Y(n_5942)
);

INVx1_ASAP7_75t_L g5943 ( 
.A(n_5659),
.Y(n_5943)
);

BUFx10_ASAP7_75t_L g5944 ( 
.A(n_5534),
.Y(n_5944)
);

CKINVDCx6p67_ASAP7_75t_R g5945 ( 
.A(n_5446),
.Y(n_5945)
);

CKINVDCx5p33_ASAP7_75t_R g5946 ( 
.A(n_5556),
.Y(n_5946)
);

CKINVDCx20_ASAP7_75t_R g5947 ( 
.A(n_5383),
.Y(n_5947)
);

CKINVDCx5p33_ASAP7_75t_R g5948 ( 
.A(n_5556),
.Y(n_5948)
);

CKINVDCx5p33_ASAP7_75t_R g5949 ( 
.A(n_5161),
.Y(n_5949)
);

INVx1_ASAP7_75t_L g5950 ( 
.A(n_5661),
.Y(n_5950)
);

INVx1_ASAP7_75t_L g5951 ( 
.A(n_5662),
.Y(n_5951)
);

INVx1_ASAP7_75t_L g5952 ( 
.A(n_5665),
.Y(n_5952)
);

HB1xp67_ASAP7_75t_L g5953 ( 
.A(n_5605),
.Y(n_5953)
);

INVx2_ASAP7_75t_L g5954 ( 
.A(n_5283),
.Y(n_5954)
);

INVx2_ASAP7_75t_L g5955 ( 
.A(n_5307),
.Y(n_5955)
);

NAND2xp5_ASAP7_75t_L g5956 ( 
.A(n_5132),
.B(n_2918),
.Y(n_5956)
);

CKINVDCx5p33_ASAP7_75t_R g5957 ( 
.A(n_5261),
.Y(n_5957)
);

INVx2_ASAP7_75t_L g5958 ( 
.A(n_5308),
.Y(n_5958)
);

BUFx3_ASAP7_75t_L g5959 ( 
.A(n_5242),
.Y(n_5959)
);

INVx3_ASAP7_75t_L g5960 ( 
.A(n_5444),
.Y(n_5960)
);

INVx1_ASAP7_75t_L g5961 ( 
.A(n_5666),
.Y(n_5961)
);

INVx1_ASAP7_75t_L g5962 ( 
.A(n_5669),
.Y(n_5962)
);

CKINVDCx5p33_ASAP7_75t_R g5963 ( 
.A(n_5628),
.Y(n_5963)
);

INVx1_ASAP7_75t_L g5964 ( 
.A(n_5673),
.Y(n_5964)
);

INVx1_ASAP7_75t_L g5965 ( 
.A(n_5675),
.Y(n_5965)
);

CKINVDCx5p33_ASAP7_75t_R g5966 ( 
.A(n_5628),
.Y(n_5966)
);

INVx1_ASAP7_75t_L g5967 ( 
.A(n_5679),
.Y(n_5967)
);

INVx1_ASAP7_75t_L g5968 ( 
.A(n_5427),
.Y(n_5968)
);

CKINVDCx5p33_ASAP7_75t_R g5969 ( 
.A(n_5446),
.Y(n_5969)
);

INVx1_ASAP7_75t_L g5970 ( 
.A(n_5436),
.Y(n_5970)
);

CKINVDCx5p33_ASAP7_75t_R g5971 ( 
.A(n_5236),
.Y(n_5971)
);

CKINVDCx5p33_ASAP7_75t_R g5972 ( 
.A(n_5260),
.Y(n_5972)
);

CKINVDCx20_ASAP7_75t_R g5973 ( 
.A(n_5456),
.Y(n_5973)
);

NOR2xp33_ASAP7_75t_R g5974 ( 
.A(n_5505),
.B(n_4114),
.Y(n_5974)
);

CKINVDCx5p33_ASAP7_75t_R g5975 ( 
.A(n_5450),
.Y(n_5975)
);

INVx1_ASAP7_75t_L g5976 ( 
.A(n_5289),
.Y(n_5976)
);

INVx1_ASAP7_75t_L g5977 ( 
.A(n_5290),
.Y(n_5977)
);

INVx1_ASAP7_75t_L g5978 ( 
.A(n_5294),
.Y(n_5978)
);

INVx1_ASAP7_75t_L g5979 ( 
.A(n_5301),
.Y(n_5979)
);

HB1xp67_ASAP7_75t_L g5980 ( 
.A(n_5672),
.Y(n_5980)
);

NOR2xp33_ASAP7_75t_L g5981 ( 
.A(n_5225),
.B(n_2922),
.Y(n_5981)
);

CKINVDCx20_ASAP7_75t_R g5982 ( 
.A(n_5607),
.Y(n_5982)
);

CKINVDCx5p33_ASAP7_75t_R g5983 ( 
.A(n_5263),
.Y(n_5983)
);

CKINVDCx5p33_ASAP7_75t_R g5984 ( 
.A(n_5369),
.Y(n_5984)
);

NOR2xp33_ASAP7_75t_L g5985 ( 
.A(n_5226),
.B(n_2924),
.Y(n_5985)
);

INVx1_ASAP7_75t_L g5986 ( 
.A(n_5311),
.Y(n_5986)
);

NOR2xp67_ASAP7_75t_L g5987 ( 
.A(n_5254),
.B(n_2928),
.Y(n_5987)
);

CKINVDCx20_ASAP7_75t_R g5988 ( 
.A(n_5617),
.Y(n_5988)
);

CKINVDCx5p33_ASAP7_75t_R g5989 ( 
.A(n_5428),
.Y(n_5989)
);

CKINVDCx5p33_ASAP7_75t_R g5990 ( 
.A(n_5252),
.Y(n_5990)
);

INVx1_ASAP7_75t_L g5991 ( 
.A(n_5326),
.Y(n_5991)
);

CKINVDCx5p33_ASAP7_75t_R g5992 ( 
.A(n_5397),
.Y(n_5992)
);

AOI22xp5_ASAP7_75t_L g5993 ( 
.A1(n_5209),
.A2(n_4136),
.B1(n_4197),
.B2(n_4121),
.Y(n_5993)
);

NAND2xp5_ASAP7_75t_L g5994 ( 
.A(n_5611),
.B(n_2930),
.Y(n_5994)
);

CKINVDCx20_ASAP7_75t_R g5995 ( 
.A(n_5650),
.Y(n_5995)
);

CKINVDCx5p33_ASAP7_75t_R g5996 ( 
.A(n_5441),
.Y(n_5996)
);

INVx2_ASAP7_75t_L g5997 ( 
.A(n_5310),
.Y(n_5997)
);

CKINVDCx5p33_ASAP7_75t_R g5998 ( 
.A(n_5447),
.Y(n_5998)
);

XOR2xp5_ASAP7_75t_L g5999 ( 
.A(n_5189),
.B(n_2934),
.Y(n_5999)
);

CKINVDCx5p33_ASAP7_75t_R g6000 ( 
.A(n_5448),
.Y(n_6000)
);

AND2x2_ASAP7_75t_L g6001 ( 
.A(n_5269),
.B(n_2935),
.Y(n_6001)
);

CKINVDCx5p33_ASAP7_75t_R g6002 ( 
.A(n_5642),
.Y(n_6002)
);

CKINVDCx5p33_ASAP7_75t_R g6003 ( 
.A(n_5694),
.Y(n_6003)
);

CKINVDCx5p33_ASAP7_75t_R g6004 ( 
.A(n_5232),
.Y(n_6004)
);

INVx1_ASAP7_75t_L g6005 ( 
.A(n_5349),
.Y(n_6005)
);

INVx3_ASAP7_75t_L g6006 ( 
.A(n_5184),
.Y(n_6006)
);

CKINVDCx5p33_ASAP7_75t_R g6007 ( 
.A(n_5232),
.Y(n_6007)
);

NOR2xp33_ASAP7_75t_R g6008 ( 
.A(n_5508),
.B(n_2938),
.Y(n_6008)
);

INVx1_ASAP7_75t_L g6009 ( 
.A(n_5350),
.Y(n_6009)
);

CKINVDCx5p33_ASAP7_75t_R g6010 ( 
.A(n_5229),
.Y(n_6010)
);

CKINVDCx5p33_ASAP7_75t_R g6011 ( 
.A(n_5201),
.Y(n_6011)
);

CKINVDCx5p33_ASAP7_75t_R g6012 ( 
.A(n_5327),
.Y(n_6012)
);

BUFx2_ASAP7_75t_L g6013 ( 
.A(n_5470),
.Y(n_6013)
);

CKINVDCx5p33_ASAP7_75t_R g6014 ( 
.A(n_5327),
.Y(n_6014)
);

CKINVDCx5p33_ASAP7_75t_R g6015 ( 
.A(n_5594),
.Y(n_6015)
);

CKINVDCx5p33_ASAP7_75t_R g6016 ( 
.A(n_5339),
.Y(n_6016)
);

INVx2_ASAP7_75t_L g6017 ( 
.A(n_5313),
.Y(n_6017)
);

CKINVDCx5p33_ASAP7_75t_R g6018 ( 
.A(n_5409),
.Y(n_6018)
);

INVx2_ASAP7_75t_L g6019 ( 
.A(n_5314),
.Y(n_6019)
);

CKINVDCx5p33_ASAP7_75t_R g6020 ( 
.A(n_5566),
.Y(n_6020)
);

NOR2xp33_ASAP7_75t_R g6021 ( 
.A(n_5511),
.B(n_2940),
.Y(n_6021)
);

BUFx6f_ASAP7_75t_L g6022 ( 
.A(n_5648),
.Y(n_6022)
);

AND2x6_ASAP7_75t_L g6023 ( 
.A(n_5136),
.B(n_3204),
.Y(n_6023)
);

NAND2xp33_ASAP7_75t_R g6024 ( 
.A(n_5498),
.B(n_2941),
.Y(n_6024)
);

CKINVDCx5p33_ASAP7_75t_R g6025 ( 
.A(n_5572),
.Y(n_6025)
);

OAI22xp5_ASAP7_75t_SL g6026 ( 
.A1(n_5141),
.A2(n_2944),
.B1(n_2948),
.B2(n_2942),
.Y(n_6026)
);

AND2x2_ASAP7_75t_L g6027 ( 
.A(n_5689),
.B(n_2952),
.Y(n_6027)
);

NAND2xp33_ASAP7_75t_L g6028 ( 
.A(n_5262),
.B(n_2953),
.Y(n_6028)
);

CKINVDCx5p33_ASAP7_75t_R g6029 ( 
.A(n_5575),
.Y(n_6029)
);

CKINVDCx5p33_ASAP7_75t_R g6030 ( 
.A(n_5580),
.Y(n_6030)
);

HB1xp67_ASAP7_75t_L g6031 ( 
.A(n_5481),
.Y(n_6031)
);

XNOR2xp5_ASAP7_75t_L g6032 ( 
.A(n_5264),
.B(n_2955),
.Y(n_6032)
);

CKINVDCx16_ASAP7_75t_R g6033 ( 
.A(n_5280),
.Y(n_6033)
);

CKINVDCx5p33_ASAP7_75t_R g6034 ( 
.A(n_5535),
.Y(n_6034)
);

CKINVDCx5p33_ASAP7_75t_R g6035 ( 
.A(n_5544),
.Y(n_6035)
);

CKINVDCx5p33_ASAP7_75t_R g6036 ( 
.A(n_5506),
.Y(n_6036)
);

INVx1_ASAP7_75t_L g6037 ( 
.A(n_5352),
.Y(n_6037)
);

CKINVDCx20_ASAP7_75t_R g6038 ( 
.A(n_5653),
.Y(n_6038)
);

CKINVDCx5p33_ASAP7_75t_R g6039 ( 
.A(n_5517),
.Y(n_6039)
);

NOR2xp67_ASAP7_75t_L g6040 ( 
.A(n_5503),
.B(n_2957),
.Y(n_6040)
);

NOR2xp33_ASAP7_75t_R g6041 ( 
.A(n_5493),
.B(n_2960),
.Y(n_6041)
);

INVx2_ASAP7_75t_L g6042 ( 
.A(n_5317),
.Y(n_6042)
);

HB1xp67_ASAP7_75t_L g6043 ( 
.A(n_5483),
.Y(n_6043)
);

INVxp33_ASAP7_75t_SL g6044 ( 
.A(n_5526),
.Y(n_6044)
);

BUFx3_ASAP7_75t_L g6045 ( 
.A(n_5654),
.Y(n_6045)
);

CKINVDCx5p33_ASAP7_75t_R g6046 ( 
.A(n_5542),
.Y(n_6046)
);

NAND2xp33_ASAP7_75t_R g6047 ( 
.A(n_5463),
.B(n_2961),
.Y(n_6047)
);

INVx1_ASAP7_75t_L g6048 ( 
.A(n_5354),
.Y(n_6048)
);

NAND2xp33_ASAP7_75t_R g6049 ( 
.A(n_5465),
.B(n_2962),
.Y(n_6049)
);

NOR2xp33_ASAP7_75t_R g6050 ( 
.A(n_5496),
.B(n_2963),
.Y(n_6050)
);

NAND2xp5_ASAP7_75t_SL g6051 ( 
.A(n_5391),
.B(n_2964),
.Y(n_6051)
);

NOR2xp33_ASAP7_75t_R g6052 ( 
.A(n_5500),
.B(n_2967),
.Y(n_6052)
);

CKINVDCx5p33_ASAP7_75t_R g6053 ( 
.A(n_5295),
.Y(n_6053)
);

CKINVDCx5p33_ASAP7_75t_R g6054 ( 
.A(n_5295),
.Y(n_6054)
);

AND2x4_ASAP7_75t_L g6055 ( 
.A(n_5404),
.B(n_3226),
.Y(n_6055)
);

OR2x2_ASAP7_75t_L g6056 ( 
.A(n_5621),
.B(n_5285),
.Y(n_6056)
);

CKINVDCx20_ASAP7_75t_R g6057 ( 
.A(n_5489),
.Y(n_6057)
);

CKINVDCx5p33_ASAP7_75t_R g6058 ( 
.A(n_5286),
.Y(n_6058)
);

CKINVDCx5p33_ASAP7_75t_R g6059 ( 
.A(n_5286),
.Y(n_6059)
);

BUFx6f_ASAP7_75t_L g6060 ( 
.A(n_5656),
.Y(n_6060)
);

NOR2xp33_ASAP7_75t_L g6061 ( 
.A(n_5214),
.B(n_2969),
.Y(n_6061)
);

AOI21x1_ASAP7_75t_L g6062 ( 
.A1(n_5340),
.A2(n_3239),
.B(n_3236),
.Y(n_6062)
);

INVx1_ASAP7_75t_L g6063 ( 
.A(n_5359),
.Y(n_6063)
);

CKINVDCx5p33_ASAP7_75t_R g6064 ( 
.A(n_5527),
.Y(n_6064)
);

CKINVDCx5p33_ASAP7_75t_R g6065 ( 
.A(n_5538),
.Y(n_6065)
);

CKINVDCx5p33_ASAP7_75t_R g6066 ( 
.A(n_5158),
.Y(n_6066)
);

CKINVDCx5p33_ASAP7_75t_R g6067 ( 
.A(n_5494),
.Y(n_6067)
);

NAND2xp5_ASAP7_75t_L g6068 ( 
.A(n_5631),
.B(n_2970),
.Y(n_6068)
);

CKINVDCx5p33_ASAP7_75t_R g6069 ( 
.A(n_5528),
.Y(n_6069)
);

CKINVDCx20_ASAP7_75t_R g6070 ( 
.A(n_5554),
.Y(n_6070)
);

CKINVDCx20_ASAP7_75t_R g6071 ( 
.A(n_5469),
.Y(n_6071)
);

AND2x2_ASAP7_75t_L g6072 ( 
.A(n_5222),
.B(n_2971),
.Y(n_6072)
);

CKINVDCx5p33_ASAP7_75t_R g6073 ( 
.A(n_5430),
.Y(n_6073)
);

CKINVDCx20_ASAP7_75t_R g6074 ( 
.A(n_5471),
.Y(n_6074)
);

HB1xp67_ASAP7_75t_L g6075 ( 
.A(n_5169),
.Y(n_6075)
);

AOI21x1_ASAP7_75t_L g6076 ( 
.A1(n_5633),
.A2(n_3245),
.B(n_3243),
.Y(n_6076)
);

CKINVDCx5p33_ASAP7_75t_R g6077 ( 
.A(n_5437),
.Y(n_6077)
);

CKINVDCx5p33_ASAP7_75t_R g6078 ( 
.A(n_5472),
.Y(n_6078)
);

CKINVDCx20_ASAP7_75t_R g6079 ( 
.A(n_5475),
.Y(n_6079)
);

INVx1_ASAP7_75t_L g6080 ( 
.A(n_5364),
.Y(n_6080)
);

NOR2xp33_ASAP7_75t_L g6081 ( 
.A(n_5637),
.B(n_2976),
.Y(n_6081)
);

NAND2xp5_ASAP7_75t_L g6082 ( 
.A(n_5638),
.B(n_2977),
.Y(n_6082)
);

CKINVDCx5p33_ASAP7_75t_R g6083 ( 
.A(n_5476),
.Y(n_6083)
);

INVx1_ASAP7_75t_L g6084 ( 
.A(n_5372),
.Y(n_6084)
);

INVx1_ASAP7_75t_L g6085 ( 
.A(n_5385),
.Y(n_6085)
);

INVx1_ASAP7_75t_L g6086 ( 
.A(n_5386),
.Y(n_6086)
);

CKINVDCx5p33_ASAP7_75t_R g6087 ( 
.A(n_5479),
.Y(n_6087)
);

CKINVDCx5p33_ASAP7_75t_R g6088 ( 
.A(n_5482),
.Y(n_6088)
);

NOR2xp33_ASAP7_75t_R g6089 ( 
.A(n_5440),
.B(n_2979),
.Y(n_6089)
);

INVx1_ASAP7_75t_L g6090 ( 
.A(n_5387),
.Y(n_6090)
);

NOR2xp33_ASAP7_75t_R g6091 ( 
.A(n_5485),
.B(n_2989),
.Y(n_6091)
);

OA22x2_ASAP7_75t_L g6092 ( 
.A1(n_5196),
.A2(n_2991),
.B1(n_2992),
.B2(n_2990),
.Y(n_6092)
);

CKINVDCx5p33_ASAP7_75t_R g6093 ( 
.A(n_5603),
.Y(n_6093)
);

CKINVDCx5p33_ASAP7_75t_R g6094 ( 
.A(n_5615),
.Y(n_6094)
);

INVx2_ASAP7_75t_L g6095 ( 
.A(n_5321),
.Y(n_6095)
);

INVx1_ASAP7_75t_L g6096 ( 
.A(n_5389),
.Y(n_6096)
);

NAND2xp33_ASAP7_75t_SL g6097 ( 
.A(n_5318),
.B(n_2997),
.Y(n_6097)
);

HB1xp67_ASAP7_75t_L g6098 ( 
.A(n_5335),
.Y(n_6098)
);

CKINVDCx5p33_ASAP7_75t_R g6099 ( 
.A(n_5618),
.Y(n_6099)
);

CKINVDCx5p33_ASAP7_75t_R g6100 ( 
.A(n_5667),
.Y(n_6100)
);

CKINVDCx20_ASAP7_75t_R g6101 ( 
.A(n_5175),
.Y(n_6101)
);

INVx1_ASAP7_75t_L g6102 ( 
.A(n_5393),
.Y(n_6102)
);

CKINVDCx5p33_ASAP7_75t_R g6103 ( 
.A(n_5674),
.Y(n_6103)
);

NOR2xp33_ASAP7_75t_R g6104 ( 
.A(n_5423),
.B(n_2998),
.Y(n_6104)
);

CKINVDCx5p33_ASAP7_75t_R g6105 ( 
.A(n_5677),
.Y(n_6105)
);

INVx1_ASAP7_75t_L g6106 ( 
.A(n_5398),
.Y(n_6106)
);

CKINVDCx5p33_ASAP7_75t_R g6107 ( 
.A(n_5330),
.Y(n_6107)
);

NOR2xp67_ASAP7_75t_L g6108 ( 
.A(n_5433),
.B(n_3001),
.Y(n_6108)
);

NOR2xp33_ASAP7_75t_R g6109 ( 
.A(n_5425),
.B(n_3003),
.Y(n_6109)
);

CKINVDCx5p33_ASAP7_75t_R g6110 ( 
.A(n_5555),
.Y(n_6110)
);

CKINVDCx5p33_ASAP7_75t_R g6111 ( 
.A(n_5563),
.Y(n_6111)
);

INVx1_ASAP7_75t_L g6112 ( 
.A(n_5401),
.Y(n_6112)
);

CKINVDCx5p33_ASAP7_75t_R g6113 ( 
.A(n_5149),
.Y(n_6113)
);

INVx2_ASAP7_75t_L g6114 ( 
.A(n_5322),
.Y(n_6114)
);

CKINVDCx5p33_ASAP7_75t_R g6115 ( 
.A(n_5435),
.Y(n_6115)
);

CKINVDCx5p33_ASAP7_75t_R g6116 ( 
.A(n_5186),
.Y(n_6116)
);

CKINVDCx5p33_ASAP7_75t_R g6117 ( 
.A(n_5194),
.Y(n_6117)
);

BUFx3_ASAP7_75t_L g6118 ( 
.A(n_5670),
.Y(n_6118)
);

NAND2xp5_ASAP7_75t_L g6119 ( 
.A(n_5645),
.B(n_3004),
.Y(n_6119)
);

INVx1_ASAP7_75t_L g6120 ( 
.A(n_5402),
.Y(n_6120)
);

CKINVDCx5p33_ASAP7_75t_R g6121 ( 
.A(n_5210),
.Y(n_6121)
);

INVx1_ASAP7_75t_L g6122 ( 
.A(n_5403),
.Y(n_6122)
);

NOR2xp33_ASAP7_75t_R g6123 ( 
.A(n_5344),
.B(n_3006),
.Y(n_6123)
);

INVx1_ASAP7_75t_L g6124 ( 
.A(n_5413),
.Y(n_6124)
);

INVx1_ASAP7_75t_L g6125 ( 
.A(n_5414),
.Y(n_6125)
);

NOR2xp33_ASAP7_75t_R g6126 ( 
.A(n_5346),
.B(n_3015),
.Y(n_6126)
);

CKINVDCx5p33_ASAP7_75t_R g6127 ( 
.A(n_5259),
.Y(n_6127)
);

INVx1_ASAP7_75t_L g6128 ( 
.A(n_5312),
.Y(n_6128)
);

CKINVDCx5p33_ASAP7_75t_R g6129 ( 
.A(n_5302),
.Y(n_6129)
);

AND2x2_ASAP7_75t_L g6130 ( 
.A(n_5223),
.B(n_3016),
.Y(n_6130)
);

CKINVDCx5p33_ASAP7_75t_R g6131 ( 
.A(n_5394),
.Y(n_6131)
);

CKINVDCx5p33_ASAP7_75t_R g6132 ( 
.A(n_5478),
.Y(n_6132)
);

CKINVDCx5p33_ASAP7_75t_R g6133 ( 
.A(n_5487),
.Y(n_6133)
);

INVx1_ASAP7_75t_L g6134 ( 
.A(n_5296),
.Y(n_6134)
);

CKINVDCx5p33_ASAP7_75t_R g6135 ( 
.A(n_5495),
.Y(n_6135)
);

BUFx6f_ASAP7_75t_L g6136 ( 
.A(n_5686),
.Y(n_6136)
);

INVx1_ASAP7_75t_L g6137 ( 
.A(n_5300),
.Y(n_6137)
);

CKINVDCx5p33_ASAP7_75t_R g6138 ( 
.A(n_5381),
.Y(n_6138)
);

CKINVDCx20_ASAP7_75t_R g6139 ( 
.A(n_5204),
.Y(n_6139)
);

INVx2_ASAP7_75t_L g6140 ( 
.A(n_5337),
.Y(n_6140)
);

CKINVDCx5p33_ASAP7_75t_R g6141 ( 
.A(n_5395),
.Y(n_6141)
);

AND2x2_ASAP7_75t_L g6142 ( 
.A(n_5243),
.B(n_3021),
.Y(n_6142)
);

CKINVDCx5p33_ASAP7_75t_R g6143 ( 
.A(n_5399),
.Y(n_6143)
);

AND2x2_ASAP7_75t_L g6144 ( 
.A(n_5274),
.B(n_3023),
.Y(n_6144)
);

CKINVDCx5p33_ASAP7_75t_R g6145 ( 
.A(n_5418),
.Y(n_6145)
);

HB1xp67_ASAP7_75t_L g6146 ( 
.A(n_5144),
.Y(n_6146)
);

CKINVDCx20_ASAP7_75t_R g6147 ( 
.A(n_5267),
.Y(n_6147)
);

NAND2xp33_ASAP7_75t_SL g6148 ( 
.A(n_5373),
.B(n_3025),
.Y(n_6148)
);

BUFx3_ASAP7_75t_L g6149 ( 
.A(n_5368),
.Y(n_6149)
);

BUFx6f_ASAP7_75t_SL g6150 ( 
.A(n_5347),
.Y(n_6150)
);

CKINVDCx5p33_ASAP7_75t_R g6151 ( 
.A(n_5432),
.Y(n_6151)
);

CKINVDCx20_ASAP7_75t_R g6152 ( 
.A(n_5199),
.Y(n_6152)
);

CKINVDCx5p33_ASAP7_75t_R g6153 ( 
.A(n_5241),
.Y(n_6153)
);

CKINVDCx5p33_ASAP7_75t_R g6154 ( 
.A(n_5451),
.Y(n_6154)
);

INVx2_ASAP7_75t_L g6155 ( 
.A(n_5338),
.Y(n_6155)
);

INVx2_ASAP7_75t_L g6156 ( 
.A(n_5342),
.Y(n_6156)
);

OR2x6_ASAP7_75t_L g6157 ( 
.A(n_5578),
.B(n_3267),
.Y(n_6157)
);

INVx1_ASAP7_75t_L g6158 ( 
.A(n_5343),
.Y(n_6158)
);

CKINVDCx5p33_ASAP7_75t_R g6159 ( 
.A(n_5460),
.Y(n_6159)
);

BUFx6f_ASAP7_75t_L g6160 ( 
.A(n_5227),
.Y(n_6160)
);

AO21x2_ASAP7_75t_L g6161 ( 
.A1(n_5531),
.A2(n_3280),
.B(n_3277),
.Y(n_6161)
);

NOR2xp33_ASAP7_75t_L g6162 ( 
.A(n_5652),
.B(n_3027),
.Y(n_6162)
);

CKINVDCx5p33_ASAP7_75t_R g6163 ( 
.A(n_5374),
.Y(n_6163)
);

CKINVDCx5p33_ASAP7_75t_R g6164 ( 
.A(n_5374),
.Y(n_6164)
);

CKINVDCx5p33_ASAP7_75t_R g6165 ( 
.A(n_5207),
.Y(n_6165)
);

CKINVDCx20_ASAP7_75t_R g6166 ( 
.A(n_5454),
.Y(n_6166)
);

BUFx6f_ASAP7_75t_L g6167 ( 
.A(n_5228),
.Y(n_6167)
);

CKINVDCx5p33_ASAP7_75t_R g6168 ( 
.A(n_5239),
.Y(n_6168)
);

BUFx6f_ASAP7_75t_L g6169 ( 
.A(n_5218),
.Y(n_6169)
);

CKINVDCx5p33_ASAP7_75t_R g6170 ( 
.A(n_5347),
.Y(n_6170)
);

CKINVDCx5p33_ASAP7_75t_R g6171 ( 
.A(n_5445),
.Y(n_6171)
);

CKINVDCx5p33_ASAP7_75t_R g6172 ( 
.A(n_5421),
.Y(n_6172)
);

CKINVDCx5p33_ASAP7_75t_R g6173 ( 
.A(n_5664),
.Y(n_6173)
);

NOR2xp33_ASAP7_75t_R g6174 ( 
.A(n_5348),
.B(n_3028),
.Y(n_6174)
);

CKINVDCx20_ASAP7_75t_R g6175 ( 
.A(n_5680),
.Y(n_6175)
);

OAI21x1_ASAP7_75t_L g6176 ( 
.A1(n_5205),
.A2(n_3285),
.B(n_3282),
.Y(n_6176)
);

CKINVDCx5p33_ASAP7_75t_R g6177 ( 
.A(n_5698),
.Y(n_6177)
);

INVx2_ASAP7_75t_L g6178 ( 
.A(n_5355),
.Y(n_6178)
);

INVx2_ASAP7_75t_L g6179 ( 
.A(n_5356),
.Y(n_6179)
);

CKINVDCx20_ASAP7_75t_R g6180 ( 
.A(n_5202),
.Y(n_6180)
);

INVx2_ASAP7_75t_L g6181 ( 
.A(n_5358),
.Y(n_6181)
);

NOR2xp33_ASAP7_75t_R g6182 ( 
.A(n_5353),
.B(n_3030),
.Y(n_6182)
);

INVx3_ASAP7_75t_L g6183 ( 
.A(n_5365),
.Y(n_6183)
);

INVx1_ASAP7_75t_L g6184 ( 
.A(n_5377),
.Y(n_6184)
);

CKINVDCx5p33_ASAP7_75t_R g6185 ( 
.A(n_5234),
.Y(n_6185)
);

CKINVDCx5p33_ASAP7_75t_R g6186 ( 
.A(n_5293),
.Y(n_6186)
);

CKINVDCx5p33_ASAP7_75t_R g6187 ( 
.A(n_5297),
.Y(n_6187)
);

CKINVDCx5p33_ASAP7_75t_R g6188 ( 
.A(n_5323),
.Y(n_6188)
);

CKINVDCx5p33_ASAP7_75t_R g6189 ( 
.A(n_5247),
.Y(n_6189)
);

CKINVDCx5p33_ASAP7_75t_R g6190 ( 
.A(n_5258),
.Y(n_6190)
);

INVx2_ASAP7_75t_L g6191 ( 
.A(n_5122),
.Y(n_6191)
);

CKINVDCx20_ASAP7_75t_R g6192 ( 
.A(n_5151),
.Y(n_6192)
);

BUFx6f_ASAP7_75t_L g6193 ( 
.A(n_5272),
.Y(n_6193)
);

CKINVDCx20_ASAP7_75t_R g6194 ( 
.A(n_5150),
.Y(n_6194)
);

CKINVDCx5p33_ASAP7_75t_R g6195 ( 
.A(n_5287),
.Y(n_6195)
);

CKINVDCx16_ASAP7_75t_R g6196 ( 
.A(n_5532),
.Y(n_6196)
);

CKINVDCx5p33_ASAP7_75t_R g6197 ( 
.A(n_5298),
.Y(n_6197)
);

CKINVDCx20_ASAP7_75t_R g6198 ( 
.A(n_5277),
.Y(n_6198)
);

CKINVDCx5p33_ASAP7_75t_R g6199 ( 
.A(n_5324),
.Y(n_6199)
);

NOR2xp33_ASAP7_75t_L g6200 ( 
.A(n_5255),
.B(n_3031),
.Y(n_6200)
);

NOR2xp33_ASAP7_75t_L g6201 ( 
.A(n_5279),
.B(n_3036),
.Y(n_6201)
);

BUFx3_ASAP7_75t_L g6202 ( 
.A(n_5606),
.Y(n_6202)
);

CKINVDCx20_ASAP7_75t_R g6203 ( 
.A(n_5291),
.Y(n_6203)
);

INVx1_ASAP7_75t_L g6204 ( 
.A(n_5126),
.Y(n_6204)
);

CKINVDCx5p33_ASAP7_75t_R g6205 ( 
.A(n_5341),
.Y(n_6205)
);

AND2x2_ASAP7_75t_L g6206 ( 
.A(n_5303),
.B(n_3037),
.Y(n_6206)
);

INVx3_ASAP7_75t_L g6207 ( 
.A(n_5305),
.Y(n_6207)
);

NAND2xp5_ASAP7_75t_L g6208 ( 
.A(n_5245),
.B(n_3038),
.Y(n_6208)
);

CKINVDCx5p33_ASAP7_75t_R g6209 ( 
.A(n_5367),
.Y(n_6209)
);

CKINVDCx5p33_ASAP7_75t_R g6210 ( 
.A(n_5370),
.Y(n_6210)
);

INVxp67_ASAP7_75t_SL g6211 ( 
.A(n_5361),
.Y(n_6211)
);

INVx1_ASAP7_75t_L g6212 ( 
.A(n_5609),
.Y(n_6212)
);

OR2x2_ASAP7_75t_L g6213 ( 
.A(n_5334),
.B(n_3040),
.Y(n_6213)
);

INVx2_ASAP7_75t_SL g6214 ( 
.A(n_5400),
.Y(n_6214)
);

CKINVDCx5p33_ASAP7_75t_R g6215 ( 
.A(n_5382),
.Y(n_6215)
);

BUFx2_ASAP7_75t_L g6216 ( 
.A(n_5651),
.Y(n_6216)
);

BUFx10_ASAP7_75t_L g6217 ( 
.A(n_5640),
.Y(n_6217)
);

CKINVDCx5p33_ASAP7_75t_R g6218 ( 
.A(n_5212),
.Y(n_6218)
);

INVx2_ASAP7_75t_L g6219 ( 
.A(n_5614),
.Y(n_6219)
);

CKINVDCx5p33_ASAP7_75t_R g6220 ( 
.A(n_5220),
.Y(n_6220)
);

CKINVDCx5p33_ASAP7_75t_R g6221 ( 
.A(n_5336),
.Y(n_6221)
);

INVx2_ASAP7_75t_L g6222 ( 
.A(n_5619),
.Y(n_6222)
);

CKINVDCx5p33_ASAP7_75t_R g6223 ( 
.A(n_5250),
.Y(n_6223)
);

INVx2_ASAP7_75t_L g6224 ( 
.A(n_5629),
.Y(n_6224)
);

NAND2xp33_ASAP7_75t_R g6225 ( 
.A(n_5453),
.B(n_3046),
.Y(n_6225)
);

CKINVDCx5p33_ASAP7_75t_R g6226 ( 
.A(n_5284),
.Y(n_6226)
);

INVx1_ASAP7_75t_L g6227 ( 
.A(n_5632),
.Y(n_6227)
);

NAND2xp5_ASAP7_75t_L g6228 ( 
.A(n_5138),
.B(n_3048),
.Y(n_6228)
);

INVx2_ASAP7_75t_L g6229 ( 
.A(n_5634),
.Y(n_6229)
);

CKINVDCx5p33_ASAP7_75t_R g6230 ( 
.A(n_5306),
.Y(n_6230)
);

INVx1_ASAP7_75t_L g6231 ( 
.A(n_5649),
.Y(n_6231)
);

CKINVDCx5p33_ASAP7_75t_R g6232 ( 
.A(n_5309),
.Y(n_6232)
);

INVx2_ASAP7_75t_L g6233 ( 
.A(n_5663),
.Y(n_6233)
);

HB1xp67_ASAP7_75t_L g6234 ( 
.A(n_5455),
.Y(n_6234)
);

INVx1_ASAP7_75t_L g6235 ( 
.A(n_5671),
.Y(n_6235)
);

CKINVDCx5p33_ASAP7_75t_R g6236 ( 
.A(n_5316),
.Y(n_6236)
);

CKINVDCx20_ASAP7_75t_R g6237 ( 
.A(n_5408),
.Y(n_6237)
);

CKINVDCx5p33_ASAP7_75t_R g6238 ( 
.A(n_5333),
.Y(n_6238)
);

CKINVDCx5p33_ASAP7_75t_R g6239 ( 
.A(n_5363),
.Y(n_6239)
);

CKINVDCx5p33_ASAP7_75t_R g6240 ( 
.A(n_5366),
.Y(n_6240)
);

CKINVDCx5p33_ASAP7_75t_R g6241 ( 
.A(n_5384),
.Y(n_6241)
);

INVx2_ASAP7_75t_L g6242 ( 
.A(n_5684),
.Y(n_6242)
);

INVx1_ASAP7_75t_L g6243 ( 
.A(n_5329),
.Y(n_6243)
);

NAND2xp5_ASAP7_75t_L g6244 ( 
.A(n_5497),
.B(n_3049),
.Y(n_6244)
);

BUFx2_ASAP7_75t_L g6245 ( 
.A(n_5668),
.Y(n_6245)
);

NOR2xp33_ASAP7_75t_R g6246 ( 
.A(n_5655),
.B(n_3054),
.Y(n_6246)
);

OR2x2_ASAP7_75t_L g6247 ( 
.A(n_5420),
.B(n_3064),
.Y(n_6247)
);

INVxp67_ASAP7_75t_SL g6248 ( 
.A(n_5681),
.Y(n_6248)
);

NOR2xp33_ASAP7_75t_R g6249 ( 
.A(n_5257),
.B(n_3066),
.Y(n_6249)
);

CKINVDCx5p33_ASAP7_75t_R g6250 ( 
.A(n_5688),
.Y(n_6250)
);

NOR2xp33_ASAP7_75t_R g6251 ( 
.A(n_5278),
.B(n_3067),
.Y(n_6251)
);

INVx1_ASAP7_75t_L g6252 ( 
.A(n_5357),
.Y(n_6252)
);

BUFx16f_ASAP7_75t_R g6253 ( 
.A(n_5695),
.Y(n_6253)
);

CKINVDCx20_ASAP7_75t_R g6254 ( 
.A(n_5422),
.Y(n_6254)
);

INVx1_ASAP7_75t_L g6255 ( 
.A(n_5304),
.Y(n_6255)
);

CKINVDCx5p33_ASAP7_75t_R g6256 ( 
.A(n_5697),
.Y(n_6256)
);

INVx2_ASAP7_75t_L g6257 ( 
.A(n_5320),
.Y(n_6257)
);

CKINVDCx5p33_ASAP7_75t_R g6258 ( 
.A(n_5431),
.Y(n_6258)
);

NAND2xp5_ASAP7_75t_SL g6259 ( 
.A(n_6173),
.B(n_5416),
.Y(n_6259)
);

NOR2xp33_ASAP7_75t_L g6260 ( 
.A(n_6172),
.B(n_6209),
.Y(n_6260)
);

BUFx3_ASAP7_75t_L g6261 ( 
.A(n_6116),
.Y(n_6261)
);

INVx4_ASAP7_75t_L g6262 ( 
.A(n_5807),
.Y(n_6262)
);

BUFx3_ASAP7_75t_L g6263 ( 
.A(n_6117),
.Y(n_6263)
);

INVx2_ASAP7_75t_L g6264 ( 
.A(n_5708),
.Y(n_6264)
);

INVx1_ASAP7_75t_L g6265 ( 
.A(n_5700),
.Y(n_6265)
);

INVx3_ASAP7_75t_L g6266 ( 
.A(n_6149),
.Y(n_6266)
);

BUFx6f_ASAP7_75t_L g6267 ( 
.A(n_5716),
.Y(n_6267)
);

NAND2xp5_ASAP7_75t_L g6268 ( 
.A(n_6177),
.B(n_5438),
.Y(n_6268)
);

INVx1_ASAP7_75t_SL g6269 ( 
.A(n_5704),
.Y(n_6269)
);

INVx2_ASAP7_75t_L g6270 ( 
.A(n_5711),
.Y(n_6270)
);

NAND2xp5_ASAP7_75t_SL g6271 ( 
.A(n_6210),
.B(n_5183),
.Y(n_6271)
);

INVx4_ASAP7_75t_L g6272 ( 
.A(n_6073),
.Y(n_6272)
);

NAND2xp5_ASAP7_75t_SL g6273 ( 
.A(n_6215),
.B(n_5281),
.Y(n_6273)
);

AOI22xp33_ASAP7_75t_L g6274 ( 
.A1(n_6234),
.A2(n_5375),
.B1(n_5411),
.B2(n_5378),
.Y(n_6274)
);

AOI22xp33_ASAP7_75t_SL g6275 ( 
.A1(n_5885),
.A2(n_5462),
.B1(n_5461),
.B2(n_3079),
.Y(n_6275)
);

BUFx6f_ASAP7_75t_L g6276 ( 
.A(n_5716),
.Y(n_6276)
);

AND2x6_ASAP7_75t_L g6277 ( 
.A(n_6134),
.B(n_5362),
.Y(n_6277)
);

INVx1_ASAP7_75t_L g6278 ( 
.A(n_5705),
.Y(n_6278)
);

INVx1_ASAP7_75t_L g6279 ( 
.A(n_5706),
.Y(n_6279)
);

AND2x2_ASAP7_75t_L g6280 ( 
.A(n_5878),
.B(n_5325),
.Y(n_6280)
);

INVx3_ASAP7_75t_L g6281 ( 
.A(n_6160),
.Y(n_6281)
);

INVx2_ASAP7_75t_L g6282 ( 
.A(n_5715),
.Y(n_6282)
);

INVx4_ASAP7_75t_L g6283 ( 
.A(n_6077),
.Y(n_6283)
);

NOR2xp33_ASAP7_75t_SL g6284 ( 
.A(n_5710),
.B(n_3071),
.Y(n_6284)
);

NAND2xp5_ASAP7_75t_L g6285 ( 
.A(n_5818),
.B(n_5332),
.Y(n_6285)
);

AOI22xp33_ASAP7_75t_L g6286 ( 
.A1(n_5906),
.A2(n_5371),
.B1(n_5390),
.B2(n_5331),
.Y(n_6286)
);

INVx1_ASAP7_75t_L g6287 ( 
.A(n_5719),
.Y(n_6287)
);

INVx3_ASAP7_75t_L g6288 ( 
.A(n_6160),
.Y(n_6288)
);

INVx1_ASAP7_75t_L g6289 ( 
.A(n_5721),
.Y(n_6289)
);

NAND2xp5_ASAP7_75t_L g6290 ( 
.A(n_6081),
.B(n_5396),
.Y(n_6290)
);

OR2x2_ASAP7_75t_L g6291 ( 
.A(n_5757),
.B(n_5781),
.Y(n_6291)
);

OR2x2_ASAP7_75t_L g6292 ( 
.A(n_5755),
.B(n_5417),
.Y(n_6292)
);

INVx3_ASAP7_75t_L g6293 ( 
.A(n_6160),
.Y(n_6293)
);

INVx1_ASAP7_75t_L g6294 ( 
.A(n_5731),
.Y(n_6294)
);

INVx5_ASAP7_75t_L g6295 ( 
.A(n_5944),
.Y(n_6295)
);

BUFx10_ASAP7_75t_L g6296 ( 
.A(n_6150),
.Y(n_6296)
);

BUFx6f_ASAP7_75t_L g6297 ( 
.A(n_5716),
.Y(n_6297)
);

INVx1_ASAP7_75t_L g6298 ( 
.A(n_5747),
.Y(n_6298)
);

HB1xp67_ASAP7_75t_L g6299 ( 
.A(n_5723),
.Y(n_6299)
);

AOI22xp33_ASAP7_75t_L g6300 ( 
.A1(n_6056),
.A2(n_5657),
.B1(n_5412),
.B2(n_5376),
.Y(n_6300)
);

INVx2_ASAP7_75t_L g6301 ( 
.A(n_5720),
.Y(n_6301)
);

INVx1_ASAP7_75t_L g6302 ( 
.A(n_5760),
.Y(n_6302)
);

NAND2xp5_ASAP7_75t_L g6303 ( 
.A(n_6162),
.B(n_5468),
.Y(n_6303)
);

INVx5_ASAP7_75t_L g6304 ( 
.A(n_5944),
.Y(n_6304)
);

INVx1_ASAP7_75t_L g6305 ( 
.A(n_5762),
.Y(n_6305)
);

NOR2xp33_ASAP7_75t_L g6306 ( 
.A(n_6020),
.B(n_3080),
.Y(n_6306)
);

NOR2xp33_ASAP7_75t_L g6307 ( 
.A(n_6025),
.B(n_3081),
.Y(n_6307)
);

INVx2_ASAP7_75t_SL g6308 ( 
.A(n_5730),
.Y(n_6308)
);

BUFx4f_ASAP7_75t_L g6309 ( 
.A(n_5752),
.Y(n_6309)
);

NAND2xp5_ASAP7_75t_SL g6310 ( 
.A(n_6185),
.B(n_5477),
.Y(n_6310)
);

INVx2_ASAP7_75t_L g6311 ( 
.A(n_5733),
.Y(n_6311)
);

INVx1_ASAP7_75t_L g6312 ( 
.A(n_5765),
.Y(n_6312)
);

AND2x2_ASAP7_75t_L g6313 ( 
.A(n_6072),
.B(n_5490),
.Y(n_6313)
);

NAND2xp5_ASAP7_75t_SL g6314 ( 
.A(n_6186),
.B(n_3083),
.Y(n_6314)
);

INVxp33_ASAP7_75t_SL g6315 ( 
.A(n_5848),
.Y(n_6315)
);

INVx1_ASAP7_75t_SL g6316 ( 
.A(n_5992),
.Y(n_6316)
);

NAND2xp33_ASAP7_75t_L g6317 ( 
.A(n_5751),
.B(n_3086),
.Y(n_6317)
);

NAND2xp5_ASAP7_75t_L g6318 ( 
.A(n_5981),
.B(n_3087),
.Y(n_6318)
);

BUFx6f_ASAP7_75t_L g6319 ( 
.A(n_5764),
.Y(n_6319)
);

INVx1_ASAP7_75t_L g6320 ( 
.A(n_5774),
.Y(n_6320)
);

BUFx3_ASAP7_75t_L g6321 ( 
.A(n_6121),
.Y(n_6321)
);

INVx2_ASAP7_75t_L g6322 ( 
.A(n_5714),
.Y(n_6322)
);

AND2x4_ASAP7_75t_L g6323 ( 
.A(n_5823),
.B(n_3298),
.Y(n_6323)
);

INVx3_ASAP7_75t_L g6324 ( 
.A(n_6167),
.Y(n_6324)
);

NAND2xp5_ASAP7_75t_SL g6325 ( 
.A(n_6187),
.B(n_3089),
.Y(n_6325)
);

INVx2_ASAP7_75t_SL g6326 ( 
.A(n_6154),
.Y(n_6326)
);

NOR2xp33_ASAP7_75t_L g6327 ( 
.A(n_6029),
.B(n_3091),
.Y(n_6327)
);

BUFx3_ASAP7_75t_L g6328 ( 
.A(n_6138),
.Y(n_6328)
);

INVx1_ASAP7_75t_L g6329 ( 
.A(n_5779),
.Y(n_6329)
);

CKINVDCx5p33_ASAP7_75t_R g6330 ( 
.A(n_5713),
.Y(n_6330)
);

NOR2xp33_ASAP7_75t_SL g6331 ( 
.A(n_5718),
.B(n_3092),
.Y(n_6331)
);

NAND2xp5_ASAP7_75t_SL g6332 ( 
.A(n_6188),
.B(n_3097),
.Y(n_6332)
);

NOR2xp33_ASAP7_75t_L g6333 ( 
.A(n_6030),
.B(n_3099),
.Y(n_6333)
);

NAND2xp5_ASAP7_75t_SL g6334 ( 
.A(n_6036),
.B(n_3100),
.Y(n_6334)
);

INVx1_ASAP7_75t_L g6335 ( 
.A(n_5790),
.Y(n_6335)
);

NAND2xp5_ASAP7_75t_L g6336 ( 
.A(n_5985),
.B(n_3102),
.Y(n_6336)
);

INVx3_ASAP7_75t_L g6337 ( 
.A(n_6167),
.Y(n_6337)
);

BUFx3_ASAP7_75t_L g6338 ( 
.A(n_6141),
.Y(n_6338)
);

INVx2_ASAP7_75t_L g6339 ( 
.A(n_5714),
.Y(n_6339)
);

INVx2_ASAP7_75t_L g6340 ( 
.A(n_5798),
.Y(n_6340)
);

NAND2xp5_ASAP7_75t_L g6341 ( 
.A(n_6039),
.B(n_3104),
.Y(n_6341)
);

BUFx8_ASAP7_75t_SL g6342 ( 
.A(n_5712),
.Y(n_6342)
);

INVx4_ASAP7_75t_L g6343 ( 
.A(n_6143),
.Y(n_6343)
);

INVx4_ASAP7_75t_L g6344 ( 
.A(n_6145),
.Y(n_6344)
);

AND2x2_ASAP7_75t_L g6345 ( 
.A(n_5758),
.B(n_3105),
.Y(n_6345)
);

NAND2xp5_ASAP7_75t_L g6346 ( 
.A(n_6046),
.B(n_3107),
.Y(n_6346)
);

NAND2xp5_ASAP7_75t_SL g6347 ( 
.A(n_5776),
.B(n_3109),
.Y(n_6347)
);

NAND2xp33_ASAP7_75t_L g6348 ( 
.A(n_5780),
.B(n_3110),
.Y(n_6348)
);

OR2x6_ASAP7_75t_L g6349 ( 
.A(n_5794),
.B(n_3301),
.Y(n_6349)
);

NAND2xp5_ASAP7_75t_L g6350 ( 
.A(n_6061),
.B(n_3114),
.Y(n_6350)
);

INVxp67_ASAP7_75t_SL g6351 ( 
.A(n_6031),
.Y(n_6351)
);

INVx1_ASAP7_75t_L g6352 ( 
.A(n_5799),
.Y(n_6352)
);

INVx3_ASAP7_75t_L g6353 ( 
.A(n_6167),
.Y(n_6353)
);

AND2x2_ASAP7_75t_SL g6354 ( 
.A(n_6033),
.B(n_3304),
.Y(n_6354)
);

INVx5_ASAP7_75t_L g6355 ( 
.A(n_5764),
.Y(n_6355)
);

BUFx3_ASAP7_75t_L g6356 ( 
.A(n_6168),
.Y(n_6356)
);

BUFx6f_ASAP7_75t_L g6357 ( 
.A(n_5764),
.Y(n_6357)
);

INVx1_ASAP7_75t_L g6358 ( 
.A(n_5805),
.Y(n_6358)
);

BUFx3_ASAP7_75t_L g6359 ( 
.A(n_6189),
.Y(n_6359)
);

NOR2xp33_ASAP7_75t_L g6360 ( 
.A(n_5863),
.B(n_3119),
.Y(n_6360)
);

BUFx3_ASAP7_75t_L g6361 ( 
.A(n_6190),
.Y(n_6361)
);

AOI22xp33_ASAP7_75t_L g6362 ( 
.A1(n_6243),
.A2(n_3316),
.B1(n_3317),
.B2(n_3307),
.Y(n_6362)
);

INVxp67_ASAP7_75t_SL g6363 ( 
.A(n_6043),
.Y(n_6363)
);

INVx3_ASAP7_75t_L g6364 ( 
.A(n_6193),
.Y(n_6364)
);

NOR2xp33_ASAP7_75t_L g6365 ( 
.A(n_5869),
.B(n_3122),
.Y(n_6365)
);

INVx1_ASAP7_75t_L g6366 ( 
.A(n_5814),
.Y(n_6366)
);

INVx1_ASAP7_75t_L g6367 ( 
.A(n_5820),
.Y(n_6367)
);

INVx2_ASAP7_75t_L g6368 ( 
.A(n_5830),
.Y(n_6368)
);

INVx2_ASAP7_75t_L g6369 ( 
.A(n_5835),
.Y(n_6369)
);

INVx2_ASAP7_75t_L g6370 ( 
.A(n_5836),
.Y(n_6370)
);

BUFx4f_ASAP7_75t_L g6371 ( 
.A(n_5945),
.Y(n_6371)
);

INVx6_ASAP7_75t_L g6372 ( 
.A(n_5717),
.Y(n_6372)
);

INVx1_ASAP7_75t_L g6373 ( 
.A(n_5847),
.Y(n_6373)
);

AND2x2_ASAP7_75t_L g6374 ( 
.A(n_6001),
.B(n_3123),
.Y(n_6374)
);

INVx1_ASAP7_75t_L g6375 ( 
.A(n_5856),
.Y(n_6375)
);

INVx1_ASAP7_75t_L g6376 ( 
.A(n_5861),
.Y(n_6376)
);

NAND2xp5_ASAP7_75t_L g6377 ( 
.A(n_6211),
.B(n_3124),
.Y(n_6377)
);

INVx3_ASAP7_75t_L g6378 ( 
.A(n_6193),
.Y(n_6378)
);

AND2x2_ASAP7_75t_L g6379 ( 
.A(n_6144),
.B(n_6206),
.Y(n_6379)
);

BUFx6f_ASAP7_75t_L g6380 ( 
.A(n_5767),
.Y(n_6380)
);

INVx4_ASAP7_75t_L g6381 ( 
.A(n_5734),
.Y(n_6381)
);

NAND2xp5_ASAP7_75t_L g6382 ( 
.A(n_5994),
.B(n_3127),
.Y(n_6382)
);

INVx3_ASAP7_75t_L g6383 ( 
.A(n_6193),
.Y(n_6383)
);

AND2x2_ASAP7_75t_L g6384 ( 
.A(n_5748),
.B(n_3128),
.Y(n_6384)
);

CKINVDCx20_ASAP7_75t_R g6385 ( 
.A(n_5701),
.Y(n_6385)
);

INVx1_ASAP7_75t_L g6386 ( 
.A(n_5864),
.Y(n_6386)
);

INVx2_ASAP7_75t_L g6387 ( 
.A(n_5865),
.Y(n_6387)
);

NOR2xp33_ASAP7_75t_L g6388 ( 
.A(n_5750),
.B(n_3130),
.Y(n_6388)
);

NAND2xp5_ASAP7_75t_SL g6389 ( 
.A(n_6159),
.B(n_3132),
.Y(n_6389)
);

NAND2xp5_ASAP7_75t_L g6390 ( 
.A(n_6068),
.B(n_3134),
.Y(n_6390)
);

INVx1_ASAP7_75t_L g6391 ( 
.A(n_5868),
.Y(n_6391)
);

NAND2xp5_ASAP7_75t_L g6392 ( 
.A(n_6082),
.B(n_3137),
.Y(n_6392)
);

INVx2_ASAP7_75t_SL g6393 ( 
.A(n_6016),
.Y(n_6393)
);

AND2x2_ASAP7_75t_L g6394 ( 
.A(n_6130),
.B(n_3139),
.Y(n_6394)
);

NAND2xp5_ASAP7_75t_SL g6395 ( 
.A(n_6018),
.B(n_3141),
.Y(n_6395)
);

INVx2_ASAP7_75t_L g6396 ( 
.A(n_5884),
.Y(n_6396)
);

NAND2xp5_ASAP7_75t_L g6397 ( 
.A(n_6119),
.B(n_3151),
.Y(n_6397)
);

INVx1_ASAP7_75t_L g6398 ( 
.A(n_5890),
.Y(n_6398)
);

BUFx6f_ASAP7_75t_L g6399 ( 
.A(n_5767),
.Y(n_6399)
);

INVx2_ASAP7_75t_L g6400 ( 
.A(n_5891),
.Y(n_6400)
);

NOR2xp33_ASAP7_75t_L g6401 ( 
.A(n_5920),
.B(n_3154),
.Y(n_6401)
);

BUFx3_ASAP7_75t_L g6402 ( 
.A(n_6195),
.Y(n_6402)
);

INVx1_ASAP7_75t_SL g6403 ( 
.A(n_5932),
.Y(n_6403)
);

HB1xp67_ASAP7_75t_L g6404 ( 
.A(n_6098),
.Y(n_6404)
);

NAND2xp5_ASAP7_75t_SL g6405 ( 
.A(n_6214),
.B(n_3155),
.Y(n_6405)
);

BUFx3_ASAP7_75t_L g6406 ( 
.A(n_6197),
.Y(n_6406)
);

INVx6_ASAP7_75t_L g6407 ( 
.A(n_5767),
.Y(n_6407)
);

INVx1_ASAP7_75t_L g6408 ( 
.A(n_5897),
.Y(n_6408)
);

INVx2_ASAP7_75t_L g6409 ( 
.A(n_5901),
.Y(n_6409)
);

NAND2xp5_ASAP7_75t_SL g6410 ( 
.A(n_6239),
.B(n_3158),
.Y(n_6410)
);

INVx1_ASAP7_75t_L g6411 ( 
.A(n_5905),
.Y(n_6411)
);

OR2x6_ASAP7_75t_L g6412 ( 
.A(n_5822),
.B(n_3321),
.Y(n_6412)
);

NOR2xp33_ASAP7_75t_L g6413 ( 
.A(n_5953),
.B(n_3159),
.Y(n_6413)
);

INVx1_ASAP7_75t_L g6414 ( 
.A(n_5908),
.Y(n_6414)
);

NAND2xp5_ASAP7_75t_L g6415 ( 
.A(n_6200),
.B(n_3160),
.Y(n_6415)
);

AND2x2_ASAP7_75t_L g6416 ( 
.A(n_6142),
.B(n_3161),
.Y(n_6416)
);

INVx5_ASAP7_75t_L g6417 ( 
.A(n_5782),
.Y(n_6417)
);

INVx1_ASAP7_75t_L g6418 ( 
.A(n_5929),
.Y(n_6418)
);

INVx2_ASAP7_75t_L g6419 ( 
.A(n_5930),
.Y(n_6419)
);

BUFx3_ASAP7_75t_L g6420 ( 
.A(n_6199),
.Y(n_6420)
);

INVx1_ASAP7_75t_L g6421 ( 
.A(n_5942),
.Y(n_6421)
);

INVxp33_ASAP7_75t_L g6422 ( 
.A(n_5808),
.Y(n_6422)
);

INVx3_ASAP7_75t_L g6423 ( 
.A(n_6169),
.Y(n_6423)
);

INVx3_ASAP7_75t_L g6424 ( 
.A(n_6169),
.Y(n_6424)
);

BUFx10_ASAP7_75t_L g6425 ( 
.A(n_6150),
.Y(n_6425)
);

AND2x2_ASAP7_75t_SL g6426 ( 
.A(n_5877),
.B(n_3325),
.Y(n_6426)
);

INVx5_ASAP7_75t_L g6427 ( 
.A(n_5782),
.Y(n_6427)
);

OR2x6_ASAP7_75t_L g6428 ( 
.A(n_5907),
.B(n_3336),
.Y(n_6428)
);

INVx2_ASAP7_75t_L g6429 ( 
.A(n_5943),
.Y(n_6429)
);

BUFx3_ASAP7_75t_L g6430 ( 
.A(n_6205),
.Y(n_6430)
);

HB1xp67_ASAP7_75t_L g6431 ( 
.A(n_5980),
.Y(n_6431)
);

CKINVDCx5p33_ASAP7_75t_R g6432 ( 
.A(n_5724),
.Y(n_6432)
);

INVx4_ASAP7_75t_L g6433 ( 
.A(n_5736),
.Y(n_6433)
);

BUFx4f_ASAP7_75t_L g6434 ( 
.A(n_6023),
.Y(n_6434)
);

NOR2xp33_ASAP7_75t_L g6435 ( 
.A(n_5727),
.B(n_3162),
.Y(n_6435)
);

NAND2xp33_ASAP7_75t_L g6436 ( 
.A(n_5792),
.B(n_3163),
.Y(n_6436)
);

NOR2x1p5_ASAP7_75t_L g6437 ( 
.A(n_5851),
.B(n_3164),
.Y(n_6437)
);

INVx2_ASAP7_75t_L g6438 ( 
.A(n_5950),
.Y(n_6438)
);

BUFx3_ASAP7_75t_L g6439 ( 
.A(n_5784),
.Y(n_6439)
);

INVx3_ASAP7_75t_L g6440 ( 
.A(n_6169),
.Y(n_6440)
);

INVx2_ASAP7_75t_L g6441 ( 
.A(n_5951),
.Y(n_6441)
);

INVx4_ASAP7_75t_L g6442 ( 
.A(n_5737),
.Y(n_6442)
);

NAND2xp5_ASAP7_75t_SL g6443 ( 
.A(n_6240),
.B(n_3166),
.Y(n_6443)
);

NAND2xp5_ASAP7_75t_L g6444 ( 
.A(n_6201),
.B(n_3169),
.Y(n_6444)
);

INVxp67_ASAP7_75t_SL g6445 ( 
.A(n_6183),
.Y(n_6445)
);

NAND2xp5_ASAP7_75t_L g6446 ( 
.A(n_5952),
.B(n_3170),
.Y(n_6446)
);

NAND2xp5_ASAP7_75t_L g6447 ( 
.A(n_5961),
.B(n_5962),
.Y(n_6447)
);

BUFx4f_ASAP7_75t_L g6448 ( 
.A(n_6023),
.Y(n_6448)
);

OAI22xp5_ASAP7_75t_L g6449 ( 
.A1(n_6093),
.A2(n_6099),
.B1(n_6100),
.B2(n_6094),
.Y(n_6449)
);

INVx2_ASAP7_75t_L g6450 ( 
.A(n_5964),
.Y(n_6450)
);

AND2x2_ASAP7_75t_L g6451 ( 
.A(n_6027),
.B(n_3172),
.Y(n_6451)
);

NAND2xp5_ASAP7_75t_SL g6452 ( 
.A(n_6241),
.B(n_3173),
.Y(n_6452)
);

INVx1_ASAP7_75t_L g6453 ( 
.A(n_5965),
.Y(n_6453)
);

NAND2xp5_ASAP7_75t_SL g6454 ( 
.A(n_6258),
.B(n_3174),
.Y(n_6454)
);

NOR2xp33_ASAP7_75t_L g6455 ( 
.A(n_6216),
.B(n_3175),
.Y(n_6455)
);

INVx4_ASAP7_75t_L g6456 ( 
.A(n_5739),
.Y(n_6456)
);

NAND2xp5_ASAP7_75t_L g6457 ( 
.A(n_5967),
.B(n_3177),
.Y(n_6457)
);

INVx4_ASAP7_75t_L g6458 ( 
.A(n_5740),
.Y(n_6458)
);

INVx1_ASAP7_75t_L g6459 ( 
.A(n_5976),
.Y(n_6459)
);

BUFx6f_ASAP7_75t_L g6460 ( 
.A(n_5782),
.Y(n_6460)
);

NAND2xp5_ASAP7_75t_L g6461 ( 
.A(n_5977),
.B(n_3178),
.Y(n_6461)
);

NAND2xp5_ASAP7_75t_SL g6462 ( 
.A(n_5996),
.B(n_3182),
.Y(n_6462)
);

INVx3_ASAP7_75t_L g6463 ( 
.A(n_5810),
.Y(n_6463)
);

BUFx2_ASAP7_75t_L g6464 ( 
.A(n_5825),
.Y(n_6464)
);

NAND2xp5_ASAP7_75t_SL g6465 ( 
.A(n_5998),
.B(n_3186),
.Y(n_6465)
);

INVx1_ASAP7_75t_L g6466 ( 
.A(n_5978),
.Y(n_6466)
);

AND2x2_ASAP7_75t_L g6467 ( 
.A(n_6146),
.B(n_3187),
.Y(n_6467)
);

AOI22xp33_ASAP7_75t_L g6468 ( 
.A1(n_6252),
.A2(n_3342),
.B1(n_3352),
.B2(n_3339),
.Y(n_6468)
);

INVx1_ASAP7_75t_L g6469 ( 
.A(n_5979),
.Y(n_6469)
);

NAND2xp5_ASAP7_75t_L g6470 ( 
.A(n_5986),
.B(n_3189),
.Y(n_6470)
);

AOI22xp33_ASAP7_75t_L g6471 ( 
.A1(n_6137),
.A2(n_3374),
.B1(n_3377),
.B2(n_3363),
.Y(n_6471)
);

NAND2xp5_ASAP7_75t_L g6472 ( 
.A(n_5991),
.B(n_3191),
.Y(n_6472)
);

INVx1_ASAP7_75t_L g6473 ( 
.A(n_6005),
.Y(n_6473)
);

INVx5_ASAP7_75t_L g6474 ( 
.A(n_5810),
.Y(n_6474)
);

INVx2_ASAP7_75t_L g6475 ( 
.A(n_6009),
.Y(n_6475)
);

NOR2xp33_ASAP7_75t_L g6476 ( 
.A(n_5804),
.B(n_3194),
.Y(n_6476)
);

INVx3_ASAP7_75t_L g6477 ( 
.A(n_5810),
.Y(n_6477)
);

INVx1_ASAP7_75t_L g6478 ( 
.A(n_6037),
.Y(n_6478)
);

OAI22xp33_ASAP7_75t_L g6479 ( 
.A1(n_6103),
.A2(n_3197),
.B1(n_3198),
.B2(n_3195),
.Y(n_6479)
);

NOR2xp33_ASAP7_75t_SL g6480 ( 
.A(n_5853),
.B(n_3199),
.Y(n_6480)
);

NOR2xp33_ASAP7_75t_L g6481 ( 
.A(n_5804),
.B(n_3200),
.Y(n_6481)
);

OR2x2_ASAP7_75t_L g6482 ( 
.A(n_6247),
.B(n_3203),
.Y(n_6482)
);

NAND2xp5_ASAP7_75t_SL g6483 ( 
.A(n_6000),
.B(n_3205),
.Y(n_6483)
);

INVx1_ASAP7_75t_L g6484 ( 
.A(n_6048),
.Y(n_6484)
);

OR2x2_ASAP7_75t_L g6485 ( 
.A(n_5993),
.B(n_3210),
.Y(n_6485)
);

NOR2xp33_ASAP7_75t_L g6486 ( 
.A(n_5911),
.B(n_3211),
.Y(n_6486)
);

INVx1_ASAP7_75t_L g6487 ( 
.A(n_6063),
.Y(n_6487)
);

AO22x2_ASAP7_75t_L g6488 ( 
.A1(n_5999),
.A2(n_3378),
.B1(n_3383),
.B2(n_3380),
.Y(n_6488)
);

INVx4_ASAP7_75t_L g6489 ( 
.A(n_5742),
.Y(n_6489)
);

INVx1_ASAP7_75t_L g6490 ( 
.A(n_6080),
.Y(n_6490)
);

INVx1_ASAP7_75t_L g6491 ( 
.A(n_6084),
.Y(n_6491)
);

INVx2_ASAP7_75t_L g6492 ( 
.A(n_6085),
.Y(n_6492)
);

AND2x4_ASAP7_75t_L g6493 ( 
.A(n_5873),
.B(n_3386),
.Y(n_6493)
);

NAND2xp33_ASAP7_75t_L g6494 ( 
.A(n_5797),
.B(n_3212),
.Y(n_6494)
);

INVx3_ASAP7_75t_L g6495 ( 
.A(n_5927),
.Y(n_6495)
);

BUFx6f_ASAP7_75t_L g6496 ( 
.A(n_5927),
.Y(n_6496)
);

INVx1_ASAP7_75t_L g6497 ( 
.A(n_6086),
.Y(n_6497)
);

INVx1_ASAP7_75t_L g6498 ( 
.A(n_6090),
.Y(n_6498)
);

AND2x4_ASAP7_75t_L g6499 ( 
.A(n_5959),
.B(n_3390),
.Y(n_6499)
);

INVx1_ASAP7_75t_L g6500 ( 
.A(n_6096),
.Y(n_6500)
);

INVx1_ASAP7_75t_L g6501 ( 
.A(n_6102),
.Y(n_6501)
);

NAND2xp5_ASAP7_75t_L g6502 ( 
.A(n_6106),
.B(n_3214),
.Y(n_6502)
);

NAND2xp5_ASAP7_75t_SL g6503 ( 
.A(n_5838),
.B(n_3215),
.Y(n_6503)
);

INVx2_ASAP7_75t_SL g6504 ( 
.A(n_6013),
.Y(n_6504)
);

INVx2_ASAP7_75t_L g6505 ( 
.A(n_6112),
.Y(n_6505)
);

INVx4_ASAP7_75t_L g6506 ( 
.A(n_5800),
.Y(n_6506)
);

INVx1_ASAP7_75t_L g6507 ( 
.A(n_6120),
.Y(n_6507)
);

NAND2xp5_ASAP7_75t_L g6508 ( 
.A(n_6122),
.B(n_3216),
.Y(n_6508)
);

NAND2xp5_ASAP7_75t_L g6509 ( 
.A(n_6124),
.B(n_3219),
.Y(n_6509)
);

INVx1_ASAP7_75t_L g6510 ( 
.A(n_6125),
.Y(n_6510)
);

NAND2xp5_ASAP7_75t_SL g6511 ( 
.A(n_5839),
.B(n_3222),
.Y(n_6511)
);

AOI22xp33_ASAP7_75t_L g6512 ( 
.A1(n_6228),
.A2(n_3400),
.B1(n_3405),
.B2(n_3396),
.Y(n_6512)
);

BUFx4f_ASAP7_75t_L g6513 ( 
.A(n_6023),
.Y(n_6513)
);

BUFx3_ASAP7_75t_L g6514 ( 
.A(n_5827),
.Y(n_6514)
);

CKINVDCx20_ASAP7_75t_R g6515 ( 
.A(n_5735),
.Y(n_6515)
);

NAND2xp5_ASAP7_75t_SL g6516 ( 
.A(n_5840),
.B(n_3225),
.Y(n_6516)
);

INVx1_ASAP7_75t_L g6517 ( 
.A(n_5968),
.Y(n_6517)
);

AND2x2_ASAP7_75t_L g6518 ( 
.A(n_5916),
.B(n_3229),
.Y(n_6518)
);

INVx2_ASAP7_75t_L g6519 ( 
.A(n_5970),
.Y(n_6519)
);

INVx1_ASAP7_75t_L g6520 ( 
.A(n_6158),
.Y(n_6520)
);

AND2x2_ASAP7_75t_L g6521 ( 
.A(n_6221),
.B(n_3231),
.Y(n_6521)
);

BUFx10_ASAP7_75t_L g6522 ( 
.A(n_5729),
.Y(n_6522)
);

AND2x6_ASAP7_75t_L g6523 ( 
.A(n_6128),
.B(n_5787),
.Y(n_6523)
);

NAND2xp5_ASAP7_75t_L g6524 ( 
.A(n_5956),
.B(n_3232),
.Y(n_6524)
);

INVx1_ASAP7_75t_L g6525 ( 
.A(n_6184),
.Y(n_6525)
);

INVx2_ASAP7_75t_L g6526 ( 
.A(n_5743),
.Y(n_6526)
);

BUFx3_ASAP7_75t_L g6527 ( 
.A(n_5828),
.Y(n_6527)
);

INVx1_ASAP7_75t_L g6528 ( 
.A(n_5749),
.Y(n_6528)
);

AND2x2_ASAP7_75t_L g6529 ( 
.A(n_6171),
.B(n_5741),
.Y(n_6529)
);

AO21x1_ASAP7_75t_L g6530 ( 
.A1(n_6244),
.A2(n_3411),
.B(n_3408),
.Y(n_6530)
);

INVxp33_ASAP7_75t_L g6531 ( 
.A(n_5974),
.Y(n_6531)
);

BUFx3_ASAP7_75t_L g6532 ( 
.A(n_5829),
.Y(n_6532)
);

AOI22xp5_ASAP7_75t_L g6533 ( 
.A1(n_6192),
.A2(n_3234),
.B1(n_3238),
.B2(n_3233),
.Y(n_6533)
);

INVx4_ASAP7_75t_L g6534 ( 
.A(n_5744),
.Y(n_6534)
);

NAND2xp5_ASAP7_75t_SL g6535 ( 
.A(n_5846),
.B(n_3240),
.Y(n_6535)
);

INVx1_ASAP7_75t_L g6536 ( 
.A(n_5778),
.Y(n_6536)
);

INVx4_ASAP7_75t_L g6537 ( 
.A(n_5746),
.Y(n_6537)
);

INVx1_ASAP7_75t_L g6538 ( 
.A(n_5789),
.Y(n_6538)
);

INVx1_ASAP7_75t_L g6539 ( 
.A(n_5796),
.Y(n_6539)
);

INVx2_ASAP7_75t_L g6540 ( 
.A(n_5801),
.Y(n_6540)
);

CKINVDCx6p67_ASAP7_75t_R g6541 ( 
.A(n_5895),
.Y(n_6541)
);

OR2x2_ASAP7_75t_L g6542 ( 
.A(n_6196),
.B(n_3241),
.Y(n_6542)
);

AND2x4_ASAP7_75t_L g6543 ( 
.A(n_6202),
.B(n_3414),
.Y(n_6543)
);

NAND2xp5_ASAP7_75t_L g6544 ( 
.A(n_6208),
.B(n_3242),
.Y(n_6544)
);

AOI22xp33_ASAP7_75t_L g6545 ( 
.A1(n_6207),
.A2(n_3426),
.B1(n_3428),
.B2(n_3425),
.Y(n_6545)
);

BUFx3_ASAP7_75t_L g6546 ( 
.A(n_6045),
.Y(n_6546)
);

INVx1_ASAP7_75t_L g6547 ( 
.A(n_5806),
.Y(n_6547)
);

INVx2_ASAP7_75t_L g6548 ( 
.A(n_5816),
.Y(n_6548)
);

HB1xp67_ASAP7_75t_L g6549 ( 
.A(n_6067),
.Y(n_6549)
);

INVx1_ASAP7_75t_SL g6550 ( 
.A(n_6115),
.Y(n_6550)
);

INVx1_ASAP7_75t_L g6551 ( 
.A(n_5817),
.Y(n_6551)
);

INVx2_ASAP7_75t_L g6552 ( 
.A(n_5833),
.Y(n_6552)
);

INVx1_ASAP7_75t_L g6553 ( 
.A(n_5837),
.Y(n_6553)
);

INVx1_ASAP7_75t_L g6554 ( 
.A(n_5862),
.Y(n_6554)
);

NAND2xp5_ASAP7_75t_L g6555 ( 
.A(n_5702),
.B(n_3244),
.Y(n_6555)
);

OA22x2_ASAP7_75t_L g6556 ( 
.A1(n_5957),
.A2(n_3248),
.B1(n_3252),
.B2(n_3246),
.Y(n_6556)
);

NAND2xp5_ASAP7_75t_L g6557 ( 
.A(n_5702),
.B(n_3253),
.Y(n_6557)
);

INVx2_ASAP7_75t_L g6558 ( 
.A(n_5874),
.Y(n_6558)
);

NAND2xp5_ASAP7_75t_L g6559 ( 
.A(n_5707),
.B(n_3254),
.Y(n_6559)
);

INVx2_ASAP7_75t_SL g6560 ( 
.A(n_5927),
.Y(n_6560)
);

NAND2xp5_ASAP7_75t_L g6561 ( 
.A(n_5707),
.B(n_3257),
.Y(n_6561)
);

NOR2xp33_ASAP7_75t_L g6562 ( 
.A(n_5911),
.B(n_3258),
.Y(n_6562)
);

INVxp67_ASAP7_75t_L g6563 ( 
.A(n_6047),
.Y(n_6563)
);

NAND2xp5_ASAP7_75t_L g6564 ( 
.A(n_5834),
.B(n_3260),
.Y(n_6564)
);

INVx1_ASAP7_75t_L g6565 ( 
.A(n_5879),
.Y(n_6565)
);

INVx4_ASAP7_75t_SL g6566 ( 
.A(n_6023),
.Y(n_6566)
);

INVx2_ASAP7_75t_L g6567 ( 
.A(n_5921),
.Y(n_6567)
);

CKINVDCx20_ASAP7_75t_R g6568 ( 
.A(n_5795),
.Y(n_6568)
);

NOR2xp33_ASAP7_75t_L g6569 ( 
.A(n_5975),
.B(n_3263),
.Y(n_6569)
);

NAND2xp5_ASAP7_75t_L g6570 ( 
.A(n_5922),
.B(n_3268),
.Y(n_6570)
);

INVx2_ASAP7_75t_SL g6571 ( 
.A(n_6022),
.Y(n_6571)
);

BUFx6f_ASAP7_75t_L g6572 ( 
.A(n_6022),
.Y(n_6572)
);

OR2x6_ASAP7_75t_L g6573 ( 
.A(n_6157),
.B(n_3435),
.Y(n_6573)
);

NAND2xp5_ASAP7_75t_L g6574 ( 
.A(n_5924),
.B(n_3271),
.Y(n_6574)
);

NAND2xp5_ASAP7_75t_SL g6575 ( 
.A(n_5858),
.B(n_3274),
.Y(n_6575)
);

INVx1_ASAP7_75t_L g6576 ( 
.A(n_5954),
.Y(n_6576)
);

AOI22xp33_ASAP7_75t_L g6577 ( 
.A1(n_6207),
.A2(n_5894),
.B1(n_6044),
.B2(n_5787),
.Y(n_6577)
);

INVx1_ASAP7_75t_L g6578 ( 
.A(n_5955),
.Y(n_6578)
);

INVx1_ASAP7_75t_L g6579 ( 
.A(n_5958),
.Y(n_6579)
);

INVxp67_ASAP7_75t_SL g6580 ( 
.A(n_6183),
.Y(n_6580)
);

BUFx6f_ASAP7_75t_L g6581 ( 
.A(n_6022),
.Y(n_6581)
);

INVx4_ASAP7_75t_L g6582 ( 
.A(n_5854),
.Y(n_6582)
);

INVx1_ASAP7_75t_L g6583 ( 
.A(n_5997),
.Y(n_6583)
);

AND2x6_ASAP7_75t_L g6584 ( 
.A(n_6006),
.B(n_3437),
.Y(n_6584)
);

NAND2xp5_ASAP7_75t_L g6585 ( 
.A(n_6017),
.B(n_3279),
.Y(n_6585)
);

OAI221xp5_ASAP7_75t_L g6586 ( 
.A1(n_6213),
.A2(n_3452),
.B1(n_3457),
.B2(n_3447),
.C(n_3440),
.Y(n_6586)
);

INVx1_ASAP7_75t_L g6587 ( 
.A(n_6019),
.Y(n_6587)
);

INVx1_ASAP7_75t_L g6588 ( 
.A(n_6042),
.Y(n_6588)
);

AND2x4_ASAP7_75t_L g6589 ( 
.A(n_6118),
.B(n_3468),
.Y(n_6589)
);

AND2x2_ASAP7_75t_L g6590 ( 
.A(n_5926),
.B(n_3289),
.Y(n_6590)
);

BUFx10_ASAP7_75t_L g6591 ( 
.A(n_5726),
.Y(n_6591)
);

BUFx6f_ASAP7_75t_L g6592 ( 
.A(n_6060),
.Y(n_6592)
);

INVx2_ASAP7_75t_L g6593 ( 
.A(n_6095),
.Y(n_6593)
);

AND2x4_ASAP7_75t_L g6594 ( 
.A(n_6245),
.B(n_3485),
.Y(n_6594)
);

CKINVDCx20_ASAP7_75t_R g6595 ( 
.A(n_5722),
.Y(n_6595)
);

INVx1_ASAP7_75t_L g6596 ( 
.A(n_6114),
.Y(n_6596)
);

INVx3_ASAP7_75t_L g6597 ( 
.A(n_6060),
.Y(n_6597)
);

NOR2xp33_ASAP7_75t_L g6598 ( 
.A(n_5983),
.B(n_3292),
.Y(n_6598)
);

CKINVDCx5p33_ASAP7_75t_R g6599 ( 
.A(n_5725),
.Y(n_6599)
);

NAND2xp5_ASAP7_75t_SL g6600 ( 
.A(n_5859),
.B(n_3293),
.Y(n_6600)
);

BUFx2_ASAP7_75t_L g6601 ( 
.A(n_5824),
.Y(n_6601)
);

NAND3xp33_ASAP7_75t_L g6602 ( 
.A(n_5728),
.B(n_3297),
.C(n_3294),
.Y(n_6602)
);

NOR2xp33_ASAP7_75t_L g6603 ( 
.A(n_5984),
.B(n_3300),
.Y(n_6603)
);

BUFx4f_ASAP7_75t_L g6604 ( 
.A(n_6157),
.Y(n_6604)
);

OR2x6_ASAP7_75t_L g6605 ( 
.A(n_5915),
.B(n_3486),
.Y(n_6605)
);

INVx3_ASAP7_75t_L g6606 ( 
.A(n_6060),
.Y(n_6606)
);

CKINVDCx11_ASAP7_75t_R g6607 ( 
.A(n_6152),
.Y(n_6607)
);

INVx2_ASAP7_75t_L g6608 ( 
.A(n_6140),
.Y(n_6608)
);

NAND2xp5_ASAP7_75t_L g6609 ( 
.A(n_6155),
.B(n_3306),
.Y(n_6609)
);

INVx1_ASAP7_75t_L g6610 ( 
.A(n_6156),
.Y(n_6610)
);

NAND2xp5_ASAP7_75t_SL g6611 ( 
.A(n_5860),
.B(n_3308),
.Y(n_6611)
);

INVx2_ASAP7_75t_L g6612 ( 
.A(n_6178),
.Y(n_6612)
);

INVx5_ASAP7_75t_L g6613 ( 
.A(n_6136),
.Y(n_6613)
);

BUFx6f_ASAP7_75t_L g6614 ( 
.A(n_6136),
.Y(n_6614)
);

INVx2_ASAP7_75t_L g6615 ( 
.A(n_6179),
.Y(n_6615)
);

NAND2xp5_ASAP7_75t_L g6616 ( 
.A(n_6181),
.B(n_3310),
.Y(n_6616)
);

INVx2_ASAP7_75t_L g6617 ( 
.A(n_5756),
.Y(n_6617)
);

INVx1_ASAP7_75t_L g6618 ( 
.A(n_5763),
.Y(n_6618)
);

BUFx4f_ASAP7_75t_L g6619 ( 
.A(n_6136),
.Y(n_6619)
);

INVx1_ASAP7_75t_L g6620 ( 
.A(n_5770),
.Y(n_6620)
);

INVx5_ASAP7_75t_L g6621 ( 
.A(n_6217),
.Y(n_6621)
);

BUFx4f_ASAP7_75t_L g6622 ( 
.A(n_5935),
.Y(n_6622)
);

INVx1_ASAP7_75t_L g6623 ( 
.A(n_5772),
.Y(n_6623)
);

INVx1_ASAP7_75t_L g6624 ( 
.A(n_6204),
.Y(n_6624)
);

INVx2_ASAP7_75t_L g6625 ( 
.A(n_6191),
.Y(n_6625)
);

INVx4_ASAP7_75t_L g6626 ( 
.A(n_5855),
.Y(n_6626)
);

INVx1_ASAP7_75t_L g6627 ( 
.A(n_6212),
.Y(n_6627)
);

INVx1_ASAP7_75t_L g6628 ( 
.A(n_6227),
.Y(n_6628)
);

NOR3xp33_ASAP7_75t_L g6629 ( 
.A(n_6026),
.B(n_3314),
.C(n_3311),
.Y(n_6629)
);

INVx2_ASAP7_75t_SL g6630 ( 
.A(n_6075),
.Y(n_6630)
);

INVx2_ASAP7_75t_L g6631 ( 
.A(n_6219),
.Y(n_6631)
);

AND2x2_ASAP7_75t_L g6632 ( 
.A(n_5841),
.B(n_3318),
.Y(n_6632)
);

NAND2xp5_ASAP7_75t_L g6633 ( 
.A(n_6055),
.B(n_3319),
.Y(n_6633)
);

CKINVDCx5p33_ASAP7_75t_R g6634 ( 
.A(n_5699),
.Y(n_6634)
);

AOI22xp33_ASAP7_75t_L g6635 ( 
.A1(n_5888),
.A2(n_3491),
.B1(n_3492),
.B2(n_3487),
.Y(n_6635)
);

INVx2_ASAP7_75t_L g6636 ( 
.A(n_6222),
.Y(n_6636)
);

OR2x6_ASAP7_75t_L g6637 ( 
.A(n_5738),
.B(n_3493),
.Y(n_6637)
);

INVx1_ASAP7_75t_L g6638 ( 
.A(n_6231),
.Y(n_6638)
);

INVx1_ASAP7_75t_L g6639 ( 
.A(n_6235),
.Y(n_6639)
);

NOR2xp33_ASAP7_75t_L g6640 ( 
.A(n_5989),
.B(n_6175),
.Y(n_6640)
);

CKINVDCx16_ASAP7_75t_R g6641 ( 
.A(n_5753),
.Y(n_6641)
);

INVx1_ASAP7_75t_L g6642 ( 
.A(n_6224),
.Y(n_6642)
);

INVx2_ASAP7_75t_L g6643 ( 
.A(n_6229),
.Y(n_6643)
);

INVx2_ASAP7_75t_L g6644 ( 
.A(n_6233),
.Y(n_6644)
);

OR2x2_ASAP7_75t_L g6645 ( 
.A(n_5788),
.B(n_3320),
.Y(n_6645)
);

NAND2xp33_ASAP7_75t_L g6646 ( 
.A(n_5754),
.B(n_3322),
.Y(n_6646)
);

INVx1_ASAP7_75t_L g6647 ( 
.A(n_6242),
.Y(n_6647)
);

INVx2_ASAP7_75t_L g6648 ( 
.A(n_5793),
.Y(n_6648)
);

NAND2xp5_ASAP7_75t_L g6649 ( 
.A(n_6055),
.B(n_6255),
.Y(n_6649)
);

INVx3_ASAP7_75t_L g6650 ( 
.A(n_6217),
.Y(n_6650)
);

NAND2xp5_ASAP7_75t_SL g6651 ( 
.A(n_6153),
.B(n_3324),
.Y(n_6651)
);

INVx1_ASAP7_75t_SL g6652 ( 
.A(n_5831),
.Y(n_6652)
);

NAND2xp5_ASAP7_75t_SL g6653 ( 
.A(n_5949),
.B(n_3326),
.Y(n_6653)
);

INVx1_ASAP7_75t_L g6654 ( 
.A(n_5793),
.Y(n_6654)
);

BUFx3_ASAP7_75t_L g6655 ( 
.A(n_5931),
.Y(n_6655)
);

INVx1_ASAP7_75t_L g6656 ( 
.A(n_5826),
.Y(n_6656)
);

INVxp67_ASAP7_75t_L g6657 ( 
.A(n_6049),
.Y(n_6657)
);

BUFx2_ASAP7_75t_L g6658 ( 
.A(n_5832),
.Y(n_6658)
);

INVx1_ASAP7_75t_L g6659 ( 
.A(n_5826),
.Y(n_6659)
);

INVx2_ASAP7_75t_L g6660 ( 
.A(n_5849),
.Y(n_6660)
);

NAND2xp5_ASAP7_75t_SL g6661 ( 
.A(n_5870),
.B(n_3332),
.Y(n_6661)
);

INVx2_ASAP7_75t_L g6662 ( 
.A(n_5849),
.Y(n_6662)
);

NAND2xp5_ASAP7_75t_L g6663 ( 
.A(n_5850),
.B(n_3333),
.Y(n_6663)
);

NAND2xp5_ASAP7_75t_SL g6664 ( 
.A(n_5871),
.B(n_3334),
.Y(n_6664)
);

INVx2_ASAP7_75t_L g6665 ( 
.A(n_5875),
.Y(n_6665)
);

NAND2xp5_ASAP7_75t_L g6666 ( 
.A(n_5867),
.B(n_3335),
.Y(n_6666)
);

INVx1_ASAP7_75t_L g6667 ( 
.A(n_5875),
.Y(n_6667)
);

BUFx10_ASAP7_75t_L g6668 ( 
.A(n_5785),
.Y(n_6668)
);

AND2x2_ASAP7_75t_L g6669 ( 
.A(n_6064),
.B(n_3338),
.Y(n_6669)
);

INVx2_ASAP7_75t_L g6670 ( 
.A(n_5923),
.Y(n_6670)
);

INVx2_ASAP7_75t_L g6671 ( 
.A(n_5923),
.Y(n_6671)
);

NAND2xp5_ASAP7_75t_SL g6672 ( 
.A(n_5876),
.B(n_5883),
.Y(n_6672)
);

NOR2xp33_ASAP7_75t_L g6673 ( 
.A(n_5783),
.B(n_3340),
.Y(n_6673)
);

NAND2xp5_ASAP7_75t_L g6674 ( 
.A(n_6257),
.B(n_3341),
.Y(n_6674)
);

NAND2xp5_ASAP7_75t_SL g6675 ( 
.A(n_5886),
.B(n_3347),
.Y(n_6675)
);

BUFx4f_ASAP7_75t_L g6676 ( 
.A(n_6253),
.Y(n_6676)
);

BUFx3_ASAP7_75t_L g6677 ( 
.A(n_5933),
.Y(n_6677)
);

AND2x2_ASAP7_75t_L g6678 ( 
.A(n_6065),
.B(n_3348),
.Y(n_6678)
);

NAND2xp5_ASAP7_75t_L g6679 ( 
.A(n_6248),
.B(n_3356),
.Y(n_6679)
);

INVx2_ASAP7_75t_L g6680 ( 
.A(n_6062),
.Y(n_6680)
);

OR2x2_ASAP7_75t_L g6681 ( 
.A(n_5791),
.B(n_3358),
.Y(n_6681)
);

INVx1_ASAP7_75t_L g6682 ( 
.A(n_6076),
.Y(n_6682)
);

NAND2xp5_ASAP7_75t_L g6683 ( 
.A(n_5987),
.B(n_3359),
.Y(n_6683)
);

NOR2xp33_ASAP7_75t_L g6684 ( 
.A(n_5783),
.B(n_3361),
.Y(n_6684)
);

INVx1_ASAP7_75t_L g6685 ( 
.A(n_6176),
.Y(n_6685)
);

HB1xp67_ASAP7_75t_L g6686 ( 
.A(n_5917),
.Y(n_6686)
);

BUFx2_ASAP7_75t_L g6687 ( 
.A(n_5844),
.Y(n_6687)
);

AND2x4_ASAP7_75t_L g6688 ( 
.A(n_5872),
.B(n_3495),
.Y(n_6688)
);

INVx3_ASAP7_75t_L g6689 ( 
.A(n_5786),
.Y(n_6689)
);

NAND2xp5_ASAP7_75t_L g6690 ( 
.A(n_6040),
.B(n_3362),
.Y(n_6690)
);

AND2x4_ASAP7_75t_L g6691 ( 
.A(n_5745),
.B(n_3499),
.Y(n_6691)
);

BUFx6f_ASAP7_75t_L g6692 ( 
.A(n_5882),
.Y(n_6692)
);

INVx1_ASAP7_75t_L g6693 ( 
.A(n_6161),
.Y(n_6693)
);

NAND2xp5_ASAP7_75t_SL g6694 ( 
.A(n_5887),
.B(n_3364),
.Y(n_6694)
);

INVx1_ASAP7_75t_L g6695 ( 
.A(n_6161),
.Y(n_6695)
);

INVx1_ASAP7_75t_SL g6696 ( 
.A(n_5852),
.Y(n_6696)
);

NAND2xp33_ASAP7_75t_L g6697 ( 
.A(n_5963),
.B(n_3367),
.Y(n_6697)
);

INVx1_ASAP7_75t_L g6698 ( 
.A(n_6006),
.Y(n_6698)
);

AND2x6_ASAP7_75t_L g6699 ( 
.A(n_5960),
.B(n_3502),
.Y(n_6699)
);

AOI22xp33_ASAP7_75t_L g6700 ( 
.A1(n_6105),
.A2(n_3513),
.B1(n_3517),
.B2(n_3506),
.Y(n_6700)
);

INVx1_ASAP7_75t_L g6701 ( 
.A(n_5960),
.Y(n_6701)
);

INVx1_ASAP7_75t_L g6702 ( 
.A(n_6108),
.Y(n_6702)
);

OR2x2_ASAP7_75t_L g6703 ( 
.A(n_6002),
.B(n_3370),
.Y(n_6703)
);

INVx1_ASAP7_75t_SL g6704 ( 
.A(n_5880),
.Y(n_6704)
);

OR2x6_ASAP7_75t_L g6705 ( 
.A(n_6092),
.B(n_3518),
.Y(n_6705)
);

NAND2xp5_ASAP7_75t_L g6706 ( 
.A(n_5899),
.B(n_3371),
.Y(n_6706)
);

INVx1_ASAP7_75t_SL g6707 ( 
.A(n_5881),
.Y(n_6707)
);

INVx1_ASAP7_75t_L g6708 ( 
.A(n_6028),
.Y(n_6708)
);

INVx1_ASAP7_75t_L g6709 ( 
.A(n_6051),
.Y(n_6709)
);

BUFx3_ASAP7_75t_L g6710 ( 
.A(n_5761),
.Y(n_6710)
);

AND2x2_ASAP7_75t_L g6711 ( 
.A(n_5766),
.B(n_3372),
.Y(n_6711)
);

NAND2xp5_ASAP7_75t_SL g6712 ( 
.A(n_5889),
.B(n_3375),
.Y(n_6712)
);

INVx5_ASAP7_75t_L g6713 ( 
.A(n_5842),
.Y(n_6713)
);

AOI22xp33_ASAP7_75t_L g6714 ( 
.A1(n_6151),
.A2(n_3530),
.B1(n_3531),
.B2(n_3526),
.Y(n_6714)
);

NOR2xp33_ASAP7_75t_L g6715 ( 
.A(n_6127),
.B(n_3376),
.Y(n_6715)
);

INVx1_ASAP7_75t_L g6716 ( 
.A(n_6226),
.Y(n_6716)
);

INVx1_ASAP7_75t_L g6717 ( 
.A(n_6230),
.Y(n_6717)
);

INVx2_ASAP7_75t_L g6718 ( 
.A(n_6194),
.Y(n_6718)
);

NOR2xp33_ASAP7_75t_L g6719 ( 
.A(n_6129),
.B(n_3384),
.Y(n_6719)
);

NOR2xp33_ASAP7_75t_L g6720 ( 
.A(n_6131),
.B(n_3388),
.Y(n_6720)
);

AOI22xp33_ASAP7_75t_L g6721 ( 
.A1(n_6107),
.A2(n_3534),
.B1(n_3540),
.B2(n_3533),
.Y(n_6721)
);

AND2x4_ASAP7_75t_L g6722 ( 
.A(n_6250),
.B(n_3543),
.Y(n_6722)
);

NAND2xp5_ASAP7_75t_SL g6723 ( 
.A(n_5892),
.B(n_3394),
.Y(n_6723)
);

NAND2xp5_ASAP7_75t_L g6724 ( 
.A(n_6034),
.B(n_3395),
.Y(n_6724)
);

INVx2_ASAP7_75t_SL g6725 ( 
.A(n_5941),
.Y(n_6725)
);

AND2x6_ASAP7_75t_L g6726 ( 
.A(n_6225),
.B(n_3549),
.Y(n_6726)
);

INVx1_ASAP7_75t_L g6727 ( 
.A(n_6232),
.Y(n_6727)
);

NAND2xp5_ASAP7_75t_SL g6728 ( 
.A(n_5893),
.B(n_3399),
.Y(n_6728)
);

INVx1_ASAP7_75t_L g6729 ( 
.A(n_6236),
.Y(n_6729)
);

INVx2_ASAP7_75t_L g6730 ( 
.A(n_6238),
.Y(n_6730)
);

INVx4_ASAP7_75t_SL g6731 ( 
.A(n_6032),
.Y(n_6731)
);

OR2x6_ASAP7_75t_L g6732 ( 
.A(n_5768),
.B(n_3555),
.Y(n_6732)
);

INVx1_ASAP7_75t_SL g6733 ( 
.A(n_6198),
.Y(n_6733)
);

INVx1_ASAP7_75t_L g6734 ( 
.A(n_5919),
.Y(n_6734)
);

INVx3_ASAP7_75t_L g6735 ( 
.A(n_5769),
.Y(n_6735)
);

NAND2xp5_ASAP7_75t_L g6736 ( 
.A(n_6035),
.B(n_6123),
.Y(n_6736)
);

INVx2_ASAP7_75t_L g6737 ( 
.A(n_6180),
.Y(n_6737)
);

INVx1_ASAP7_75t_L g6738 ( 
.A(n_6218),
.Y(n_6738)
);

NOR2xp33_ASAP7_75t_L g6739 ( 
.A(n_6132),
.B(n_3402),
.Y(n_6739)
);

INVx2_ASAP7_75t_L g6740 ( 
.A(n_6166),
.Y(n_6740)
);

AND2x4_ASAP7_75t_L g6741 ( 
.A(n_6256),
.B(n_6071),
.Y(n_6741)
);

NAND2xp5_ASAP7_75t_L g6742 ( 
.A(n_6126),
.B(n_3407),
.Y(n_6742)
);

INVxp33_ASAP7_75t_L g6743 ( 
.A(n_6089),
.Y(n_6743)
);

NOR2xp33_ASAP7_75t_L g6744 ( 
.A(n_6133),
.B(n_3410),
.Y(n_6744)
);

INVx4_ASAP7_75t_L g6745 ( 
.A(n_5771),
.Y(n_6745)
);

NAND2x1p5_ASAP7_75t_L g6746 ( 
.A(n_5773),
.B(n_3565),
.Y(n_6746)
);

AND2x4_ASAP7_75t_L g6747 ( 
.A(n_6074),
.B(n_3569),
.Y(n_6747)
);

INVx1_ASAP7_75t_L g6748 ( 
.A(n_6220),
.Y(n_6748)
);

AOI22xp33_ASAP7_75t_L g6749 ( 
.A1(n_6069),
.A2(n_3585),
.B1(n_3601),
.B2(n_3584),
.Y(n_6749)
);

NAND2xp5_ASAP7_75t_SL g6750 ( 
.A(n_5896),
.B(n_3412),
.Y(n_6750)
);

NAND2xp5_ASAP7_75t_L g6751 ( 
.A(n_6174),
.B(n_6182),
.Y(n_6751)
);

INVx4_ASAP7_75t_L g6752 ( 
.A(n_5775),
.Y(n_6752)
);

HB1xp67_ASAP7_75t_L g6753 ( 
.A(n_6165),
.Y(n_6753)
);

INVxp67_ASAP7_75t_L g6754 ( 
.A(n_5709),
.Y(n_6754)
);

NOR2xp33_ASAP7_75t_L g6755 ( 
.A(n_6135),
.B(n_3418),
.Y(n_6755)
);

INVx1_ASAP7_75t_L g6756 ( 
.A(n_6249),
.Y(n_6756)
);

INVx1_ASAP7_75t_L g6757 ( 
.A(n_6251),
.Y(n_6757)
);

NAND2xp5_ASAP7_75t_L g6758 ( 
.A(n_5909),
.B(n_5939),
.Y(n_6758)
);

BUFx6f_ASAP7_75t_L g6759 ( 
.A(n_5857),
.Y(n_6759)
);

INVx2_ASAP7_75t_L g6760 ( 
.A(n_5902),
.Y(n_6760)
);

INVx1_ASAP7_75t_L g6761 ( 
.A(n_5903),
.Y(n_6761)
);

INVx2_ASAP7_75t_L g6762 ( 
.A(n_5904),
.Y(n_6762)
);

NAND2xp5_ASAP7_75t_L g6763 ( 
.A(n_6010),
.B(n_3419),
.Y(n_6763)
);

INVx3_ASAP7_75t_L g6764 ( 
.A(n_5777),
.Y(n_6764)
);

OR2x2_ASAP7_75t_L g6765 ( 
.A(n_6003),
.B(n_3424),
.Y(n_6765)
);

CKINVDCx5p33_ASAP7_75t_R g6766 ( 
.A(n_5732),
.Y(n_6766)
);

NAND2xp5_ASAP7_75t_L g6767 ( 
.A(n_6015),
.B(n_3427),
.Y(n_6767)
);

AND2x2_ASAP7_75t_L g6768 ( 
.A(n_6110),
.B(n_3430),
.Y(n_6768)
);

INVx2_ASAP7_75t_L g6769 ( 
.A(n_6113),
.Y(n_6769)
);

NOR2xp33_ASAP7_75t_L g6770 ( 
.A(n_5819),
.B(n_3431),
.Y(n_6770)
);

INVx2_ASAP7_75t_L g6771 ( 
.A(n_6223),
.Y(n_6771)
);

INVx2_ASAP7_75t_L g6772 ( 
.A(n_6203),
.Y(n_6772)
);

INVx1_ASAP7_75t_L g6773 ( 
.A(n_6246),
.Y(n_6773)
);

INVx3_ASAP7_75t_L g6774 ( 
.A(n_6111),
.Y(n_6774)
);

INVx1_ASAP7_75t_L g6775 ( 
.A(n_5803),
.Y(n_6775)
);

BUFx3_ASAP7_75t_L g6776 ( 
.A(n_5759),
.Y(n_6776)
);

AOI22xp33_ASAP7_75t_L g6777 ( 
.A1(n_6097),
.A2(n_3607),
.B1(n_3622),
.B2(n_3603),
.Y(n_6777)
);

AND2x2_ASAP7_75t_L g6778 ( 
.A(n_5821),
.B(n_3432),
.Y(n_6778)
);

CKINVDCx5p33_ASAP7_75t_R g6779 ( 
.A(n_5811),
.Y(n_6779)
);

NOR2xp33_ASAP7_75t_L g6780 ( 
.A(n_6011),
.B(n_3436),
.Y(n_6780)
);

NOR2x1p5_ASAP7_75t_L g6781 ( 
.A(n_5809),
.B(n_3443),
.Y(n_6781)
);

INVx1_ASAP7_75t_L g6782 ( 
.A(n_6078),
.Y(n_6782)
);

BUFx2_ASAP7_75t_L g6783 ( 
.A(n_6079),
.Y(n_6783)
);

AND2x2_ASAP7_75t_SL g6784 ( 
.A(n_5947),
.B(n_3623),
.Y(n_6784)
);

NAND2xp5_ASAP7_75t_L g6785 ( 
.A(n_6104),
.B(n_3445),
.Y(n_6785)
);

OR2x2_ASAP7_75t_L g6786 ( 
.A(n_5972),
.B(n_3446),
.Y(n_6786)
);

INVx2_ASAP7_75t_L g6787 ( 
.A(n_6237),
.Y(n_6787)
);

NAND2xp5_ASAP7_75t_SL g6788 ( 
.A(n_5966),
.B(n_3449),
.Y(n_6788)
);

CKINVDCx11_ASAP7_75t_R g6789 ( 
.A(n_5928),
.Y(n_6789)
);

NOR2xp33_ASAP7_75t_L g6790 ( 
.A(n_5990),
.B(n_3450),
.Y(n_6790)
);

NAND2xp5_ASAP7_75t_L g6791 ( 
.A(n_6109),
.B(n_3451),
.Y(n_6791)
);

OR2x2_ASAP7_75t_L g6792 ( 
.A(n_5843),
.B(n_6083),
.Y(n_6792)
);

AOI22xp33_ASAP7_75t_L g6793 ( 
.A1(n_6148),
.A2(n_3628),
.B1(n_3646),
.B2(n_3625),
.Y(n_6793)
);

INVx1_ASAP7_75t_L g6794 ( 
.A(n_6087),
.Y(n_6794)
);

AO22x2_ASAP7_75t_L g6795 ( 
.A1(n_5973),
.A2(n_5938),
.B1(n_5934),
.B2(n_6066),
.Y(n_6795)
);

INVx4_ASAP7_75t_L g6796 ( 
.A(n_6088),
.Y(n_6796)
);

NAND2xp5_ASAP7_75t_SL g6797 ( 
.A(n_5912),
.B(n_3455),
.Y(n_6797)
);

INVx1_ASAP7_75t_L g6798 ( 
.A(n_6254),
.Y(n_6798)
);

NOR2xp33_ASAP7_75t_L g6799 ( 
.A(n_6004),
.B(n_3456),
.Y(n_6799)
);

NAND2xp5_ASAP7_75t_L g6800 ( 
.A(n_6008),
.B(n_3459),
.Y(n_6800)
);

INVx1_ASAP7_75t_L g6801 ( 
.A(n_5925),
.Y(n_6801)
);

CKINVDCx20_ASAP7_75t_R g6802 ( 
.A(n_6147),
.Y(n_6802)
);

INVx4_ASAP7_75t_L g6803 ( 
.A(n_5812),
.Y(n_6803)
);

NOR2xp33_ASAP7_75t_L g6804 ( 
.A(n_6007),
.B(n_3460),
.Y(n_6804)
);

NOR2xp33_ASAP7_75t_L g6805 ( 
.A(n_6101),
.B(n_3461),
.Y(n_6805)
);

INVx2_ASAP7_75t_L g6806 ( 
.A(n_6057),
.Y(n_6806)
);

NAND2xp33_ASAP7_75t_L g6807 ( 
.A(n_5946),
.B(n_3462),
.Y(n_6807)
);

INVx1_ASAP7_75t_L g6808 ( 
.A(n_6265),
.Y(n_6808)
);

NAND2xp5_ASAP7_75t_SL g6809 ( 
.A(n_6268),
.B(n_5914),
.Y(n_6809)
);

INVx1_ASAP7_75t_L g6810 ( 
.A(n_6278),
.Y(n_6810)
);

INVx2_ASAP7_75t_L g6811 ( 
.A(n_6340),
.Y(n_6811)
);

NAND2xp5_ASAP7_75t_L g6812 ( 
.A(n_6290),
.B(n_6012),
.Y(n_6812)
);

NAND2xp5_ASAP7_75t_L g6813 ( 
.A(n_6303),
.B(n_6014),
.Y(n_6813)
);

NAND2xp5_ASAP7_75t_SL g6814 ( 
.A(n_6713),
.B(n_6379),
.Y(n_6814)
);

INVx2_ASAP7_75t_L g6815 ( 
.A(n_6368),
.Y(n_6815)
);

INVxp67_ASAP7_75t_SL g6816 ( 
.A(n_6504),
.Y(n_6816)
);

NAND2xp5_ASAP7_75t_L g6817 ( 
.A(n_6313),
.B(n_6021),
.Y(n_6817)
);

NAND2xp5_ASAP7_75t_SL g6818 ( 
.A(n_6713),
.B(n_6053),
.Y(n_6818)
);

NOR2xp33_ASAP7_75t_L g6819 ( 
.A(n_6260),
.B(n_6070),
.Y(n_6819)
);

NAND2xp33_ASAP7_75t_L g6820 ( 
.A(n_6758),
.B(n_5948),
.Y(n_6820)
);

NAND2xp5_ASAP7_75t_L g6821 ( 
.A(n_6318),
.B(n_6054),
.Y(n_6821)
);

NAND2xp5_ASAP7_75t_SL g6822 ( 
.A(n_6736),
.B(n_6058),
.Y(n_6822)
);

INVx1_ASAP7_75t_L g6823 ( 
.A(n_6279),
.Y(n_6823)
);

AOI22xp33_ASAP7_75t_L g6824 ( 
.A1(n_6426),
.A2(n_5988),
.B1(n_5995),
.B2(n_5982),
.Y(n_6824)
);

INVx1_ASAP7_75t_L g6825 ( 
.A(n_6287),
.Y(n_6825)
);

NAND2xp5_ASAP7_75t_L g6826 ( 
.A(n_6336),
.B(n_6059),
.Y(n_6826)
);

A2O1A1Ixp33_ASAP7_75t_L g6827 ( 
.A1(n_6435),
.A2(n_5937),
.B(n_5936),
.C(n_6139),
.Y(n_6827)
);

NOR2xp33_ASAP7_75t_L g6828 ( 
.A(n_6763),
.B(n_6163),
.Y(n_6828)
);

INVx1_ASAP7_75t_L g6829 ( 
.A(n_6289),
.Y(n_6829)
);

NAND2xp5_ASAP7_75t_L g6830 ( 
.A(n_6285),
.B(n_6280),
.Y(n_6830)
);

NAND2xp5_ASAP7_75t_L g6831 ( 
.A(n_6350),
.B(n_6164),
.Y(n_6831)
);

NAND2xp5_ASAP7_75t_L g6832 ( 
.A(n_6415),
.B(n_6170),
.Y(n_6832)
);

NAND2xp5_ASAP7_75t_L g6833 ( 
.A(n_6444),
.B(n_6041),
.Y(n_6833)
);

NOR2xp33_ASAP7_75t_L g6834 ( 
.A(n_6790),
.B(n_5910),
.Y(n_6834)
);

NOR2xp33_ASAP7_75t_L g6835 ( 
.A(n_6767),
.B(n_5913),
.Y(n_6835)
);

BUFx6f_ASAP7_75t_SL g6836 ( 
.A(n_6692),
.Y(n_6836)
);

NAND2xp5_ASAP7_75t_SL g6837 ( 
.A(n_6326),
.B(n_5969),
.Y(n_6837)
);

NAND2xp5_ASAP7_75t_SL g6838 ( 
.A(n_6760),
.B(n_5940),
.Y(n_6838)
);

NAND2xp5_ASAP7_75t_SL g6839 ( 
.A(n_6762),
.B(n_6050),
.Y(n_6839)
);

NAND2xp5_ASAP7_75t_SL g6840 ( 
.A(n_6761),
.B(n_6052),
.Y(n_6840)
);

NAND2xp5_ASAP7_75t_L g6841 ( 
.A(n_6382),
.B(n_6091),
.Y(n_6841)
);

NOR2xp33_ASAP7_75t_L g6842 ( 
.A(n_6715),
.B(n_5918),
.Y(n_6842)
);

NOR2xp33_ASAP7_75t_L g6843 ( 
.A(n_6719),
.B(n_6038),
.Y(n_6843)
);

NOR2xp33_ASAP7_75t_L g6844 ( 
.A(n_6720),
.B(n_5898),
.Y(n_6844)
);

INVx1_ASAP7_75t_L g6845 ( 
.A(n_6294),
.Y(n_6845)
);

NAND2xp5_ASAP7_75t_L g6846 ( 
.A(n_6390),
.B(n_5971),
.Y(n_6846)
);

INVx1_ASAP7_75t_L g6847 ( 
.A(n_6298),
.Y(n_6847)
);

INVx1_ASAP7_75t_L g6848 ( 
.A(n_6302),
.Y(n_6848)
);

AND2x4_ASAP7_75t_L g6849 ( 
.A(n_6439),
.B(n_5900),
.Y(n_6849)
);

INVx2_ASAP7_75t_SL g6850 ( 
.A(n_6291),
.Y(n_6850)
);

NAND3xp33_ASAP7_75t_L g6851 ( 
.A(n_6739),
.B(n_5703),
.C(n_5802),
.Y(n_6851)
);

INVxp67_ASAP7_75t_L g6852 ( 
.A(n_6431),
.Y(n_6852)
);

NAND2xp33_ASAP7_75t_L g6853 ( 
.A(n_6751),
.B(n_5813),
.Y(n_6853)
);

INVx2_ASAP7_75t_L g6854 ( 
.A(n_6369),
.Y(n_6854)
);

INVx2_ASAP7_75t_SL g6855 ( 
.A(n_6269),
.Y(n_6855)
);

INVx1_ASAP7_75t_L g6856 ( 
.A(n_6305),
.Y(n_6856)
);

INVxp67_ASAP7_75t_L g6857 ( 
.A(n_6549),
.Y(n_6857)
);

AND2x2_ASAP7_75t_L g6858 ( 
.A(n_6744),
.B(n_3464),
.Y(n_6858)
);

NAND2xp5_ASAP7_75t_L g6859 ( 
.A(n_6392),
.B(n_3465),
.Y(n_6859)
);

INVx2_ASAP7_75t_L g6860 ( 
.A(n_6370),
.Y(n_6860)
);

NOR3xp33_ASAP7_75t_L g6861 ( 
.A(n_6449),
.B(n_5815),
.C(n_3471),
.Y(n_6861)
);

O2A1O1Ixp33_ASAP7_75t_L g6862 ( 
.A1(n_6259),
.A2(n_3656),
.B(n_3659),
.C(n_3657),
.Y(n_6862)
);

NAND2xp5_ASAP7_75t_SL g6863 ( 
.A(n_6563),
.B(n_5845),
.Y(n_6863)
);

NAND2xp33_ASAP7_75t_SL g6864 ( 
.A(n_6743),
.B(n_5866),
.Y(n_6864)
);

NAND2xp5_ASAP7_75t_L g6865 ( 
.A(n_6397),
.B(n_3470),
.Y(n_6865)
);

BUFx3_ASAP7_75t_L g6866 ( 
.A(n_6328),
.Y(n_6866)
);

NOR2xp33_ASAP7_75t_L g6867 ( 
.A(n_6755),
.B(n_3472),
.Y(n_6867)
);

INVx2_ASAP7_75t_L g6868 ( 
.A(n_6387),
.Y(n_6868)
);

INVx2_ASAP7_75t_L g6869 ( 
.A(n_6396),
.Y(n_6869)
);

NOR2xp33_ASAP7_75t_SL g6870 ( 
.A(n_6315),
.B(n_3474),
.Y(n_6870)
);

INVx1_ASAP7_75t_L g6871 ( 
.A(n_6312),
.Y(n_6871)
);

NAND3xp33_ASAP7_75t_L g6872 ( 
.A(n_6306),
.B(n_6024),
.C(n_3476),
.Y(n_6872)
);

INVx2_ASAP7_75t_L g6873 ( 
.A(n_6400),
.Y(n_6873)
);

NAND3xp33_ASAP7_75t_L g6874 ( 
.A(n_6307),
.B(n_3479),
.C(n_3475),
.Y(n_6874)
);

OAI22xp5_ASAP7_75t_L g6875 ( 
.A1(n_6577),
.A2(n_3481),
.B1(n_3498),
.B2(n_3483),
.Y(n_6875)
);

NAND2xp5_ASAP7_75t_L g6876 ( 
.A(n_6447),
.B(n_3503),
.Y(n_6876)
);

NAND2xp5_ASAP7_75t_L g6877 ( 
.A(n_6544),
.B(n_3508),
.Y(n_6877)
);

NAND2xp5_ASAP7_75t_L g6878 ( 
.A(n_6320),
.B(n_3514),
.Y(n_6878)
);

INVxp67_ASAP7_75t_L g6879 ( 
.A(n_6686),
.Y(n_6879)
);

NAND2xp5_ASAP7_75t_L g6880 ( 
.A(n_6329),
.B(n_6335),
.Y(n_6880)
);

NAND2xp5_ASAP7_75t_L g6881 ( 
.A(n_6352),
.B(n_3515),
.Y(n_6881)
);

INVx2_ASAP7_75t_L g6882 ( 
.A(n_6409),
.Y(n_6882)
);

BUFx5_ASAP7_75t_L g6883 ( 
.A(n_6523),
.Y(n_6883)
);

NAND2xp5_ASAP7_75t_L g6884 ( 
.A(n_6358),
.B(n_3516),
.Y(n_6884)
);

BUFx6f_ASAP7_75t_L g6885 ( 
.A(n_6267),
.Y(n_6885)
);

NAND2xp5_ASAP7_75t_L g6886 ( 
.A(n_6366),
.B(n_3521),
.Y(n_6886)
);

NAND2xp5_ASAP7_75t_SL g6887 ( 
.A(n_6657),
.B(n_3522),
.Y(n_6887)
);

NOR2xp33_ASAP7_75t_L g6888 ( 
.A(n_6724),
.B(n_3524),
.Y(n_6888)
);

NAND2xp5_ASAP7_75t_SL g6889 ( 
.A(n_6550),
.B(n_3525),
.Y(n_6889)
);

INVx1_ASAP7_75t_L g6890 ( 
.A(n_6367),
.Y(n_6890)
);

NAND2xp5_ASAP7_75t_L g6891 ( 
.A(n_6373),
.B(n_3528),
.Y(n_6891)
);

NOR2xp33_ASAP7_75t_L g6892 ( 
.A(n_6360),
.B(n_3532),
.Y(n_6892)
);

NAND2xp5_ASAP7_75t_L g6893 ( 
.A(n_6375),
.B(n_3535),
.Y(n_6893)
);

INVx2_ASAP7_75t_SL g6894 ( 
.A(n_6407),
.Y(n_6894)
);

NOR2xp33_ASAP7_75t_SL g6895 ( 
.A(n_6330),
.B(n_3536),
.Y(n_6895)
);

NAND2xp5_ASAP7_75t_L g6896 ( 
.A(n_6376),
.B(n_3537),
.Y(n_6896)
);

INVx2_ASAP7_75t_L g6897 ( 
.A(n_6419),
.Y(n_6897)
);

INVx2_ASAP7_75t_L g6898 ( 
.A(n_6429),
.Y(n_6898)
);

NAND2xp5_ASAP7_75t_L g6899 ( 
.A(n_6386),
.B(n_3539),
.Y(n_6899)
);

NAND2xp5_ASAP7_75t_L g6900 ( 
.A(n_6391),
.B(n_3542),
.Y(n_6900)
);

HB1xp67_ASAP7_75t_L g6901 ( 
.A(n_6299),
.Y(n_6901)
);

INVx2_ASAP7_75t_SL g6902 ( 
.A(n_6619),
.Y(n_6902)
);

NAND2xp5_ASAP7_75t_L g6903 ( 
.A(n_6398),
.B(n_3544),
.Y(n_6903)
);

NAND3xp33_ASAP7_75t_L g6904 ( 
.A(n_6327),
.B(n_3547),
.C(n_3546),
.Y(n_6904)
);

INVx1_ASAP7_75t_L g6905 ( 
.A(n_6408),
.Y(n_6905)
);

NOR2xp33_ASAP7_75t_L g6906 ( 
.A(n_6365),
.B(n_3551),
.Y(n_6906)
);

NOR2xp33_ASAP7_75t_L g6907 ( 
.A(n_6754),
.B(n_3552),
.Y(n_6907)
);

NAND2xp5_ASAP7_75t_L g6908 ( 
.A(n_6411),
.B(n_3554),
.Y(n_6908)
);

BUFx6f_ASAP7_75t_L g6909 ( 
.A(n_6267),
.Y(n_6909)
);

NAND2xp5_ASAP7_75t_L g6910 ( 
.A(n_6414),
.B(n_3556),
.Y(n_6910)
);

BUFx6f_ASAP7_75t_L g6911 ( 
.A(n_6276),
.Y(n_6911)
);

NAND2xp5_ASAP7_75t_L g6912 ( 
.A(n_6418),
.B(n_6421),
.Y(n_6912)
);

INVx2_ASAP7_75t_L g6913 ( 
.A(n_6438),
.Y(n_6913)
);

NAND2xp5_ASAP7_75t_L g6914 ( 
.A(n_6453),
.B(n_3559),
.Y(n_6914)
);

NOR2xp33_ASAP7_75t_L g6915 ( 
.A(n_6333),
.B(n_3560),
.Y(n_6915)
);

NAND2xp5_ASAP7_75t_L g6916 ( 
.A(n_6459),
.B(n_6466),
.Y(n_6916)
);

INVx1_ASAP7_75t_L g6917 ( 
.A(n_6469),
.Y(n_6917)
);

NAND2xp5_ASAP7_75t_L g6918 ( 
.A(n_6473),
.B(n_3561),
.Y(n_6918)
);

NAND2xp5_ASAP7_75t_L g6919 ( 
.A(n_6478),
.B(n_3564),
.Y(n_6919)
);

NOR2xp33_ASAP7_75t_L g6920 ( 
.A(n_6780),
.B(n_3566),
.Y(n_6920)
);

INVxp67_ASAP7_75t_L g6921 ( 
.A(n_6404),
.Y(n_6921)
);

BUFx3_ASAP7_75t_L g6922 ( 
.A(n_6338),
.Y(n_6922)
);

BUFx5_ASAP7_75t_L g6923 ( 
.A(n_6523),
.Y(n_6923)
);

INVx1_ASAP7_75t_L g6924 ( 
.A(n_6484),
.Y(n_6924)
);

INVx2_ASAP7_75t_L g6925 ( 
.A(n_6441),
.Y(n_6925)
);

INVx1_ASAP7_75t_L g6926 ( 
.A(n_6487),
.Y(n_6926)
);

NAND2x1p5_ASAP7_75t_L g6927 ( 
.A(n_6355),
.B(n_3669),
.Y(n_6927)
);

NAND2xp5_ASAP7_75t_L g6928 ( 
.A(n_6490),
.B(n_3567),
.Y(n_6928)
);

NAND2xp5_ASAP7_75t_SL g6929 ( 
.A(n_6734),
.B(n_3570),
.Y(n_6929)
);

NAND2xp5_ASAP7_75t_L g6930 ( 
.A(n_6491),
.B(n_3571),
.Y(n_6930)
);

NOR2xp67_ASAP7_75t_L g6931 ( 
.A(n_6796),
.B(n_3572),
.Y(n_6931)
);

INVx1_ASAP7_75t_L g6932 ( 
.A(n_6497),
.Y(n_6932)
);

NAND2xp5_ASAP7_75t_L g6933 ( 
.A(n_6498),
.B(n_6500),
.Y(n_6933)
);

INVx1_ASAP7_75t_L g6934 ( 
.A(n_6501),
.Y(n_6934)
);

NAND2xp5_ASAP7_75t_L g6935 ( 
.A(n_6507),
.B(n_3574),
.Y(n_6935)
);

OR2x6_ASAP7_75t_L g6936 ( 
.A(n_6262),
.B(n_3670),
.Y(n_6936)
);

NAND2xp5_ASAP7_75t_L g6937 ( 
.A(n_6510),
.B(n_3575),
.Y(n_6937)
);

NOR2xp33_ASAP7_75t_L g6938 ( 
.A(n_6598),
.B(n_3576),
.Y(n_6938)
);

NAND2xp5_ASAP7_75t_L g6939 ( 
.A(n_6524),
.B(n_3588),
.Y(n_6939)
);

INVx2_ASAP7_75t_L g6940 ( 
.A(n_6450),
.Y(n_6940)
);

NAND2xp5_ASAP7_75t_SL g6941 ( 
.A(n_6292),
.B(n_3589),
.Y(n_6941)
);

NAND2xp5_ASAP7_75t_L g6942 ( 
.A(n_6475),
.B(n_3591),
.Y(n_6942)
);

NAND2xp5_ASAP7_75t_L g6943 ( 
.A(n_6492),
.B(n_3594),
.Y(n_6943)
);

OR2x6_ASAP7_75t_L g6944 ( 
.A(n_6381),
.B(n_3671),
.Y(n_6944)
);

OAI22xp5_ASAP7_75t_L g6945 ( 
.A1(n_6445),
.A2(n_3596),
.B1(n_3608),
.B2(n_3599),
.Y(n_6945)
);

NAND2xp5_ASAP7_75t_L g6946 ( 
.A(n_6505),
.B(n_3609),
.Y(n_6946)
);

NAND2xp5_ASAP7_75t_L g6947 ( 
.A(n_6451),
.B(n_6286),
.Y(n_6947)
);

INVx2_ASAP7_75t_L g6948 ( 
.A(n_6264),
.Y(n_6948)
);

BUFx5_ASAP7_75t_L g6949 ( 
.A(n_6523),
.Y(n_6949)
);

BUFx6f_ASAP7_75t_L g6950 ( 
.A(n_6276),
.Y(n_6950)
);

INVx2_ASAP7_75t_L g6951 ( 
.A(n_6270),
.Y(n_6951)
);

NOR2xp33_ASAP7_75t_L g6952 ( 
.A(n_6603),
.B(n_3611),
.Y(n_6952)
);

OR2x6_ASAP7_75t_L g6953 ( 
.A(n_6433),
.B(n_3674),
.Y(n_6953)
);

AND2x2_ASAP7_75t_SL g6954 ( 
.A(n_6641),
.B(n_6354),
.Y(n_6954)
);

INVx2_ASAP7_75t_L g6955 ( 
.A(n_6282),
.Y(n_6955)
);

NOR2xp33_ASAP7_75t_L g6956 ( 
.A(n_6341),
.B(n_3612),
.Y(n_6956)
);

NAND2xp5_ASAP7_75t_L g6957 ( 
.A(n_6374),
.B(n_3613),
.Y(n_6957)
);

AND2x2_ASAP7_75t_L g6958 ( 
.A(n_6590),
.B(n_3615),
.Y(n_6958)
);

CKINVDCx5p33_ASAP7_75t_R g6959 ( 
.A(n_6342),
.Y(n_6959)
);

BUFx12f_ASAP7_75t_L g6960 ( 
.A(n_6607),
.Y(n_6960)
);

NAND2xp5_ASAP7_75t_L g6961 ( 
.A(n_6394),
.B(n_6416),
.Y(n_6961)
);

NAND2xp5_ASAP7_75t_L g6962 ( 
.A(n_6564),
.B(n_3616),
.Y(n_6962)
);

AOI22xp5_ASAP7_75t_L g6963 ( 
.A1(n_6726),
.A2(n_3624),
.B1(n_3630),
.B2(n_3626),
.Y(n_6963)
);

INVx1_ASAP7_75t_L g6964 ( 
.A(n_6517),
.Y(n_6964)
);

INVx1_ASAP7_75t_L g6965 ( 
.A(n_6520),
.Y(n_6965)
);

NAND2xp5_ASAP7_75t_L g6966 ( 
.A(n_6709),
.B(n_3634),
.Y(n_6966)
);

AOI22xp5_ASAP7_75t_L g6967 ( 
.A1(n_6726),
.A2(n_3635),
.B1(n_3638),
.B2(n_3637),
.Y(n_6967)
);

NAND2xp5_ASAP7_75t_L g6968 ( 
.A(n_6346),
.B(n_3639),
.Y(n_6968)
);

NAND2xp5_ASAP7_75t_L g6969 ( 
.A(n_6580),
.B(n_3641),
.Y(n_6969)
);

NAND2xp5_ASAP7_75t_L g6970 ( 
.A(n_6778),
.B(n_3642),
.Y(n_6970)
);

OR2x6_ASAP7_75t_L g6971 ( 
.A(n_6442),
.B(n_6456),
.Y(n_6971)
);

INVx2_ASAP7_75t_L g6972 ( 
.A(n_6301),
.Y(n_6972)
);

INVx1_ASAP7_75t_L g6973 ( 
.A(n_6525),
.Y(n_6973)
);

AND2x6_ASAP7_75t_L g6974 ( 
.A(n_6708),
.B(n_3677),
.Y(n_6974)
);

INVx1_ASAP7_75t_L g6975 ( 
.A(n_6624),
.Y(n_6975)
);

INVx1_ASAP7_75t_L g6976 ( 
.A(n_6627),
.Y(n_6976)
);

NAND2xp5_ASAP7_75t_L g6977 ( 
.A(n_6384),
.B(n_3643),
.Y(n_6977)
);

INVx1_ASAP7_75t_L g6978 ( 
.A(n_6628),
.Y(n_6978)
);

INVx1_ASAP7_75t_L g6979 ( 
.A(n_6638),
.Y(n_6979)
);

NAND2xp5_ASAP7_75t_SL g6980 ( 
.A(n_6782),
.B(n_6794),
.Y(n_6980)
);

NAND2xp5_ASAP7_75t_SL g6981 ( 
.A(n_6801),
.B(n_3647),
.Y(n_6981)
);

NAND2xp33_ASAP7_75t_SL g6982 ( 
.A(n_6531),
.B(n_3648),
.Y(n_6982)
);

AND2x2_ASAP7_75t_SL g6983 ( 
.A(n_6784),
.B(n_3679),
.Y(n_6983)
);

INVx1_ASAP7_75t_L g6984 ( 
.A(n_6639),
.Y(n_6984)
);

INVx1_ASAP7_75t_L g6985 ( 
.A(n_6528),
.Y(n_6985)
);

NOR2xp33_ASAP7_75t_L g6986 ( 
.A(n_6703),
.B(n_3649),
.Y(n_6986)
);

NOR2xp33_ASAP7_75t_L g6987 ( 
.A(n_6765),
.B(n_6786),
.Y(n_6987)
);

INVx8_ASAP7_75t_L g6988 ( 
.A(n_6355),
.Y(n_6988)
);

NAND2xp5_ASAP7_75t_L g6989 ( 
.A(n_6377),
.B(n_6726),
.Y(n_6989)
);

NAND2xp5_ASAP7_75t_L g6990 ( 
.A(n_6519),
.B(n_6512),
.Y(n_6990)
);

NAND2xp5_ASAP7_75t_SL g6991 ( 
.A(n_6393),
.B(n_3650),
.Y(n_6991)
);

INVxp67_ASAP7_75t_L g6992 ( 
.A(n_6351),
.Y(n_6992)
);

NAND2xp33_ASAP7_75t_SL g6993 ( 
.A(n_6756),
.B(n_3651),
.Y(n_6993)
);

CKINVDCx20_ASAP7_75t_R g6994 ( 
.A(n_6568),
.Y(n_6994)
);

NAND2xp5_ASAP7_75t_SL g6995 ( 
.A(n_6757),
.B(n_3654),
.Y(n_6995)
);

NAND2xp5_ASAP7_75t_L g6996 ( 
.A(n_6310),
.B(n_3660),
.Y(n_6996)
);

NAND2xp5_ASAP7_75t_L g6997 ( 
.A(n_6455),
.B(n_3662),
.Y(n_6997)
);

NAND2xp5_ASAP7_75t_L g6998 ( 
.A(n_6526),
.B(n_3663),
.Y(n_6998)
);

AND2x2_ASAP7_75t_L g6999 ( 
.A(n_6669),
.B(n_3664),
.Y(n_6999)
);

BUFx6f_ASAP7_75t_SL g7000 ( 
.A(n_6692),
.Y(n_7000)
);

AOI22xp5_ASAP7_75t_L g7001 ( 
.A1(n_6347),
.A2(n_3666),
.B1(n_3672),
.B2(n_3667),
.Y(n_7001)
);

NOR2xp33_ASAP7_75t_L g7002 ( 
.A(n_6569),
.B(n_3673),
.Y(n_7002)
);

AOI22xp33_ASAP7_75t_L g7003 ( 
.A1(n_6530),
.A2(n_3686),
.B1(n_3689),
.B2(n_3684),
.Y(n_7003)
);

NAND2xp5_ASAP7_75t_L g7004 ( 
.A(n_6540),
.B(n_3675),
.Y(n_7004)
);

NOR2xp33_ASAP7_75t_L g7005 ( 
.A(n_6805),
.B(n_6672),
.Y(n_7005)
);

NAND2xp5_ASAP7_75t_L g7006 ( 
.A(n_6548),
.B(n_3678),
.Y(n_7006)
);

NAND2xp5_ASAP7_75t_SL g7007 ( 
.A(n_6275),
.B(n_3682),
.Y(n_7007)
);

NOR2xp33_ASAP7_75t_L g7008 ( 
.A(n_6422),
.B(n_3683),
.Y(n_7008)
);

NAND2x1_ASAP7_75t_L g7009 ( 
.A(n_6698),
.B(n_3290),
.Y(n_7009)
);

BUFx6f_ASAP7_75t_L g7010 ( 
.A(n_6297),
.Y(n_7010)
);

INVx1_ASAP7_75t_L g7011 ( 
.A(n_6536),
.Y(n_7011)
);

NAND2xp5_ASAP7_75t_L g7012 ( 
.A(n_6552),
.B(n_3685),
.Y(n_7012)
);

NAND2xp5_ASAP7_75t_L g7013 ( 
.A(n_6558),
.B(n_3694),
.Y(n_7013)
);

AOI22xp5_ASAP7_75t_L g7014 ( 
.A1(n_6702),
.A2(n_3697),
.B1(n_3699),
.B2(n_3695),
.Y(n_7014)
);

NOR2xp33_ASAP7_75t_L g7015 ( 
.A(n_6316),
.B(n_3700),
.Y(n_7015)
);

NAND2xp5_ASAP7_75t_SL g7016 ( 
.A(n_6773),
.B(n_3709),
.Y(n_7016)
);

NAND2xp5_ASAP7_75t_L g7017 ( 
.A(n_6567),
.B(n_3710),
.Y(n_7017)
);

NAND2xp5_ASAP7_75t_L g7018 ( 
.A(n_6593),
.B(n_3713),
.Y(n_7018)
);

NOR2xp33_ASAP7_75t_L g7019 ( 
.A(n_6363),
.B(n_6770),
.Y(n_7019)
);

NAND2xp5_ASAP7_75t_L g7020 ( 
.A(n_6608),
.B(n_3714),
.Y(n_7020)
);

INVx2_ASAP7_75t_L g7021 ( 
.A(n_6311),
.Y(n_7021)
);

NAND2xp5_ASAP7_75t_L g7022 ( 
.A(n_6612),
.B(n_3715),
.Y(n_7022)
);

AOI22xp33_ASAP7_75t_L g7023 ( 
.A1(n_6586),
.A2(n_3692),
.B1(n_3704),
.B2(n_3691),
.Y(n_7023)
);

NAND2xp5_ASAP7_75t_L g7024 ( 
.A(n_6615),
.B(n_3716),
.Y(n_7024)
);

AND2x4_ASAP7_75t_L g7025 ( 
.A(n_6261),
.B(n_3717),
.Y(n_7025)
);

INVx2_ASAP7_75t_L g7026 ( 
.A(n_6617),
.Y(n_7026)
);

NAND2xp5_ASAP7_75t_SL g7027 ( 
.A(n_6735),
.B(n_3718),
.Y(n_7027)
);

INVx8_ASAP7_75t_L g7028 ( 
.A(n_6417),
.Y(n_7028)
);

AOI22xp33_ASAP7_75t_L g7029 ( 
.A1(n_6545),
.A2(n_6539),
.B1(n_6547),
.B2(n_6538),
.Y(n_7029)
);

AND2x2_ASAP7_75t_L g7030 ( 
.A(n_6678),
.B(n_3719),
.Y(n_7030)
);

INVx1_ASAP7_75t_L g7031 ( 
.A(n_6551),
.Y(n_7031)
);

NAND2xp5_ASAP7_75t_L g7032 ( 
.A(n_6553),
.B(n_3720),
.Y(n_7032)
);

INVx1_ASAP7_75t_L g7033 ( 
.A(n_6554),
.Y(n_7033)
);

NAND2xp5_ASAP7_75t_L g7034 ( 
.A(n_6565),
.B(n_3723),
.Y(n_7034)
);

INVxp33_ASAP7_75t_L g7035 ( 
.A(n_6529),
.Y(n_7035)
);

NAND2xp5_ASAP7_75t_L g7036 ( 
.A(n_6576),
.B(n_3725),
.Y(n_7036)
);

AND2x2_ASAP7_75t_L g7037 ( 
.A(n_6768),
.B(n_3726),
.Y(n_7037)
);

INVx1_ASAP7_75t_L g7038 ( 
.A(n_6578),
.Y(n_7038)
);

INVx1_ASAP7_75t_L g7039 ( 
.A(n_6579),
.Y(n_7039)
);

INVx1_ASAP7_75t_SL g7040 ( 
.A(n_6783),
.Y(n_7040)
);

INVx1_ASAP7_75t_L g7041 ( 
.A(n_6583),
.Y(n_7041)
);

AOI221xp5_ASAP7_75t_L g7042 ( 
.A1(n_6479),
.A2(n_3735),
.B1(n_3741),
.B2(n_3722),
.C(n_3721),
.Y(n_7042)
);

NAND2xp5_ASAP7_75t_SL g7043 ( 
.A(n_6764),
.B(n_3732),
.Y(n_7043)
);

HB1xp67_ASAP7_75t_L g7044 ( 
.A(n_6417),
.Y(n_7044)
);

NAND2xp5_ASAP7_75t_L g7045 ( 
.A(n_6587),
.B(n_3733),
.Y(n_7045)
);

BUFx3_ASAP7_75t_L g7046 ( 
.A(n_6356),
.Y(n_7046)
);

NAND2xp5_ASAP7_75t_L g7047 ( 
.A(n_6588),
.B(n_3736),
.Y(n_7047)
);

INVx2_ASAP7_75t_L g7048 ( 
.A(n_6625),
.Y(n_7048)
);

OR2x2_ASAP7_75t_L g7049 ( 
.A(n_6403),
.B(n_3738),
.Y(n_7049)
);

AND2x2_ASAP7_75t_L g7050 ( 
.A(n_6518),
.B(n_6711),
.Y(n_7050)
);

NAND2xp5_ASAP7_75t_L g7051 ( 
.A(n_6596),
.B(n_3739),
.Y(n_7051)
);

NAND2xp5_ASAP7_75t_L g7052 ( 
.A(n_6610),
.B(n_3740),
.Y(n_7052)
);

NAND2xp5_ASAP7_75t_SL g7053 ( 
.A(n_6284),
.B(n_3746),
.Y(n_7053)
);

OAI221xp5_ASAP7_75t_L g7054 ( 
.A1(n_6700),
.A2(n_3747),
.B1(n_3751),
.B2(n_3750),
.C(n_3748),
.Y(n_7054)
);

NAND2xp5_ASAP7_75t_L g7055 ( 
.A(n_6618),
.B(n_3757),
.Y(n_7055)
);

NOR2xp33_ASAP7_75t_L g7056 ( 
.A(n_6486),
.B(n_3758),
.Y(n_7056)
);

NAND2xp5_ASAP7_75t_L g7057 ( 
.A(n_6620),
.B(n_6623),
.Y(n_7057)
);

NAND2xp5_ASAP7_75t_SL g7058 ( 
.A(n_6331),
.B(n_3759),
.Y(n_7058)
);

INVx2_ASAP7_75t_SL g7059 ( 
.A(n_6427),
.Y(n_7059)
);

INVx1_ASAP7_75t_L g7060 ( 
.A(n_6642),
.Y(n_7060)
);

INVx2_ASAP7_75t_SL g7061 ( 
.A(n_6427),
.Y(n_7061)
);

INVx1_ASAP7_75t_L g7062 ( 
.A(n_6647),
.Y(n_7062)
);

INVx1_ASAP7_75t_L g7063 ( 
.A(n_6631),
.Y(n_7063)
);

NOR2xp33_ASAP7_75t_L g7064 ( 
.A(n_6562),
.B(n_3761),
.Y(n_7064)
);

AND2x2_ASAP7_75t_L g7065 ( 
.A(n_6345),
.B(n_3767),
.Y(n_7065)
);

NOR2xp33_ASAP7_75t_L g7066 ( 
.A(n_6673),
.B(n_3768),
.Y(n_7066)
);

NAND2xp33_ASAP7_75t_SL g7067 ( 
.A(n_6297),
.B(n_3772),
.Y(n_7067)
);

NOR2xp33_ASAP7_75t_L g7068 ( 
.A(n_6684),
.B(n_3775),
.Y(n_7068)
);

NAND2xp5_ASAP7_75t_SL g7069 ( 
.A(n_6308),
.B(n_3777),
.Y(n_7069)
);

INVx2_ASAP7_75t_L g7070 ( 
.A(n_6636),
.Y(n_7070)
);

NAND2xp5_ASAP7_75t_SL g7071 ( 
.A(n_6774),
.B(n_3778),
.Y(n_7071)
);

NAND2xp5_ASAP7_75t_L g7072 ( 
.A(n_6322),
.B(n_3779),
.Y(n_7072)
);

NAND2xp5_ASAP7_75t_L g7073 ( 
.A(n_6339),
.B(n_3780),
.Y(n_7073)
);

NAND2xp33_ASAP7_75t_L g7074 ( 
.A(n_6277),
.B(n_3781),
.Y(n_7074)
);

NOR2xp33_ASAP7_75t_L g7075 ( 
.A(n_6476),
.B(n_6481),
.Y(n_7075)
);

AND2x2_ASAP7_75t_L g7076 ( 
.A(n_6467),
.B(n_6632),
.Y(n_7076)
);

NOR2xp33_ASAP7_75t_L g7077 ( 
.A(n_6645),
.B(n_6681),
.Y(n_7077)
);

INVx2_ASAP7_75t_L g7078 ( 
.A(n_6643),
.Y(n_7078)
);

NAND2xp5_ASAP7_75t_L g7079 ( 
.A(n_6471),
.B(n_3783),
.Y(n_7079)
);

INVx2_ASAP7_75t_L g7080 ( 
.A(n_6644),
.Y(n_7080)
);

NAND2xp5_ASAP7_75t_L g7081 ( 
.A(n_6413),
.B(n_3784),
.Y(n_7081)
);

AO221x1_ASAP7_75t_L g7082 ( 
.A1(n_6488),
.A2(n_6682),
.B1(n_6695),
.B2(n_6693),
.C(n_6795),
.Y(n_7082)
);

INVx2_ASAP7_75t_L g7083 ( 
.A(n_6648),
.Y(n_7083)
);

NOR2x1p5_ASAP7_75t_L g7084 ( 
.A(n_6263),
.B(n_3786),
.Y(n_7084)
);

OR2x2_ASAP7_75t_L g7085 ( 
.A(n_6737),
.B(n_3789),
.Y(n_7085)
);

NAND2xp5_ASAP7_75t_L g7086 ( 
.A(n_6362),
.B(n_3791),
.Y(n_7086)
);

NOR2xp33_ASAP7_75t_L g7087 ( 
.A(n_6740),
.B(n_3792),
.Y(n_7087)
);

NAND2xp5_ASAP7_75t_SL g7088 ( 
.A(n_6689),
.B(n_3794),
.Y(n_7088)
);

NAND2xp5_ASAP7_75t_L g7089 ( 
.A(n_6468),
.B(n_3795),
.Y(n_7089)
);

NOR2xp33_ASAP7_75t_L g7090 ( 
.A(n_6718),
.B(n_3796),
.Y(n_7090)
);

NAND2xp5_ASAP7_75t_SL g7091 ( 
.A(n_6604),
.B(n_3800),
.Y(n_7091)
);

INVx2_ASAP7_75t_L g7092 ( 
.A(n_6660),
.Y(n_7092)
);

INVx2_ASAP7_75t_L g7093 ( 
.A(n_6662),
.Y(n_7093)
);

NAND2xp5_ASAP7_75t_SL g7094 ( 
.A(n_6710),
.B(n_3801),
.Y(n_7094)
);

NAND2xp5_ASAP7_75t_SL g7095 ( 
.A(n_6630),
.B(n_3803),
.Y(n_7095)
);

INVx2_ASAP7_75t_L g7096 ( 
.A(n_6665),
.Y(n_7096)
);

NAND2xp5_ASAP7_75t_L g7097 ( 
.A(n_6679),
.B(n_3807),
.Y(n_7097)
);

OR2x2_ASAP7_75t_L g7098 ( 
.A(n_6806),
.B(n_3812),
.Y(n_7098)
);

NOR3xp33_ASAP7_75t_L g7099 ( 
.A(n_6799),
.B(n_3816),
.C(n_3813),
.Y(n_7099)
);

NOR2xp33_ASAP7_75t_L g7100 ( 
.A(n_6314),
.B(n_3820),
.Y(n_7100)
);

OAI22xp5_ASAP7_75t_L g7101 ( 
.A1(n_6274),
.A2(n_3835),
.B1(n_3838),
.B2(n_3827),
.Y(n_7101)
);

INVxp33_ASAP7_75t_L g7102 ( 
.A(n_6521),
.Y(n_7102)
);

NAND2xp5_ASAP7_75t_L g7103 ( 
.A(n_6714),
.B(n_3841),
.Y(n_7103)
);

OAI221xp5_ASAP7_75t_L g7104 ( 
.A1(n_6749),
.A2(n_3846),
.B1(n_3847),
.B2(n_3844),
.C(n_3843),
.Y(n_7104)
);

NAND2xp5_ASAP7_75t_L g7105 ( 
.A(n_6721),
.B(n_3848),
.Y(n_7105)
);

NAND2xp5_ASAP7_75t_L g7106 ( 
.A(n_6401),
.B(n_3849),
.Y(n_7106)
);

AND2x2_ASAP7_75t_L g7107 ( 
.A(n_6388),
.B(n_6482),
.Y(n_7107)
);

NOR2xp33_ASAP7_75t_L g7108 ( 
.A(n_6325),
.B(n_3850),
.Y(n_7108)
);

AND2x6_ASAP7_75t_L g7109 ( 
.A(n_6701),
.B(n_3744),
.Y(n_7109)
);

NAND2xp5_ASAP7_75t_L g7110 ( 
.A(n_6446),
.B(n_3852),
.Y(n_7110)
);

INVxp67_ASAP7_75t_L g7111 ( 
.A(n_6601),
.Y(n_7111)
);

AND2x4_ASAP7_75t_SL g7112 ( 
.A(n_6458),
.B(n_6489),
.Y(n_7112)
);

BUFx6f_ASAP7_75t_L g7113 ( 
.A(n_6319),
.Y(n_7113)
);

INVx1_ASAP7_75t_L g7114 ( 
.A(n_6654),
.Y(n_7114)
);

AND2x2_ASAP7_75t_L g7115 ( 
.A(n_6747),
.B(n_3853),
.Y(n_7115)
);

NAND2xp5_ASAP7_75t_L g7116 ( 
.A(n_6457),
.B(n_3855),
.Y(n_7116)
);

INVx1_ASAP7_75t_L g7117 ( 
.A(n_6656),
.Y(n_7117)
);

NAND2xp5_ASAP7_75t_L g7118 ( 
.A(n_6461),
.B(n_3859),
.Y(n_7118)
);

NAND2xp5_ASAP7_75t_L g7119 ( 
.A(n_6470),
.B(n_3860),
.Y(n_7119)
);

INVx2_ASAP7_75t_L g7120 ( 
.A(n_6670),
.Y(n_7120)
);

NAND2xp5_ASAP7_75t_SL g7121 ( 
.A(n_6649),
.B(n_3861),
.Y(n_7121)
);

AOI22xp5_ASAP7_75t_L g7122 ( 
.A1(n_6683),
.A2(n_3863),
.B1(n_3868),
.B2(n_3862),
.Y(n_7122)
);

INVx2_ASAP7_75t_L g7123 ( 
.A(n_6671),
.Y(n_7123)
);

NOR3xp33_ASAP7_75t_L g7124 ( 
.A(n_6804),
.B(n_3871),
.C(n_3869),
.Y(n_7124)
);

NAND2xp5_ASAP7_75t_L g7125 ( 
.A(n_6472),
.B(n_3880),
.Y(n_7125)
);

NAND2xp5_ASAP7_75t_L g7126 ( 
.A(n_6502),
.B(n_3886),
.Y(n_7126)
);

NAND2xp5_ASAP7_75t_L g7127 ( 
.A(n_6508),
.B(n_3887),
.Y(n_7127)
);

NOR2xp33_ASAP7_75t_L g7128 ( 
.A(n_6332),
.B(n_3888),
.Y(n_7128)
);

INVx2_ASAP7_75t_L g7129 ( 
.A(n_6659),
.Y(n_7129)
);

NOR3xp33_ASAP7_75t_L g7130 ( 
.A(n_6602),
.B(n_3890),
.C(n_3889),
.Y(n_7130)
);

NAND2xp5_ASAP7_75t_L g7131 ( 
.A(n_6509),
.B(n_3894),
.Y(n_7131)
);

NAND2xp5_ASAP7_75t_L g7132 ( 
.A(n_6663),
.B(n_3895),
.Y(n_7132)
);

INVx2_ASAP7_75t_L g7133 ( 
.A(n_6667),
.Y(n_7133)
);

NAND2xp5_ASAP7_75t_SL g7134 ( 
.A(n_6582),
.B(n_3896),
.Y(n_7134)
);

OAI22xp33_ASAP7_75t_L g7135 ( 
.A1(n_6485),
.A2(n_3898),
.B1(n_3901),
.B2(n_3897),
.Y(n_7135)
);

INVx2_ASAP7_75t_SL g7136 ( 
.A(n_6474),
.Y(n_7136)
);

NOR3xp33_ASAP7_75t_L g7137 ( 
.A(n_6640),
.B(n_3908),
.C(n_3907),
.Y(n_7137)
);

INVx2_ASAP7_75t_L g7138 ( 
.A(n_6680),
.Y(n_7138)
);

OR2x2_ASAP7_75t_L g7139 ( 
.A(n_6733),
.B(n_3914),
.Y(n_7139)
);

CKINVDCx5p33_ASAP7_75t_R g7140 ( 
.A(n_6599),
.Y(n_7140)
);

NAND2xp5_ASAP7_75t_SL g7141 ( 
.A(n_6626),
.B(n_3915),
.Y(n_7141)
);

NOR2xp33_ASAP7_75t_L g7142 ( 
.A(n_6334),
.B(n_3917),
.Y(n_7142)
);

INVx1_ASAP7_75t_L g7143 ( 
.A(n_6570),
.Y(n_7143)
);

NAND2xp5_ASAP7_75t_L g7144 ( 
.A(n_6666),
.B(n_3922),
.Y(n_7144)
);

AND2x4_ASAP7_75t_L g7145 ( 
.A(n_6321),
.B(n_3749),
.Y(n_7145)
);

NAND2xp5_ASAP7_75t_L g7146 ( 
.A(n_6742),
.B(n_3928),
.Y(n_7146)
);

INVx3_ASAP7_75t_L g7147 ( 
.A(n_6359),
.Y(n_7147)
);

NAND2xp5_ASAP7_75t_L g7148 ( 
.A(n_6690),
.B(n_3930),
.Y(n_7148)
);

CKINVDCx5p33_ASAP7_75t_R g7149 ( 
.A(n_6432),
.Y(n_7149)
);

NAND2xp5_ASAP7_75t_L g7150 ( 
.A(n_6555),
.B(n_3931),
.Y(n_7150)
);

INVx1_ASAP7_75t_L g7151 ( 
.A(n_6574),
.Y(n_7151)
);

NAND2xp5_ASAP7_75t_SL g7152 ( 
.A(n_6706),
.B(n_3933),
.Y(n_7152)
);

INVx1_ASAP7_75t_L g7153 ( 
.A(n_6585),
.Y(n_7153)
);

INVx2_ASAP7_75t_L g7154 ( 
.A(n_6423),
.Y(n_7154)
);

NAND2xp5_ASAP7_75t_L g7155 ( 
.A(n_6557),
.B(n_3935),
.Y(n_7155)
);

AND2x2_ASAP7_75t_L g7156 ( 
.A(n_6746),
.B(n_3936),
.Y(n_7156)
);

NAND2xp5_ASAP7_75t_SL g7157 ( 
.A(n_6745),
.B(n_3937),
.Y(n_7157)
);

NAND2xp5_ASAP7_75t_L g7158 ( 
.A(n_6559),
.B(n_3938),
.Y(n_7158)
);

INVx2_ASAP7_75t_L g7159 ( 
.A(n_6424),
.Y(n_7159)
);

OAI22xp33_ASAP7_75t_L g7160 ( 
.A1(n_6785),
.A2(n_3945),
.B1(n_3946),
.B2(n_3944),
.Y(n_7160)
);

INVx1_ASAP7_75t_L g7161 ( 
.A(n_6609),
.Y(n_7161)
);

INVx1_ASAP7_75t_L g7162 ( 
.A(n_6616),
.Y(n_7162)
);

NAND2xp5_ASAP7_75t_L g7163 ( 
.A(n_6561),
.B(n_3954),
.Y(n_7163)
);

NAND2xp5_ASAP7_75t_SL g7164 ( 
.A(n_6752),
.B(n_3955),
.Y(n_7164)
);

NAND3xp33_ASAP7_75t_SL g7165 ( 
.A(n_6629),
.B(n_3958),
.C(n_3956),
.Y(n_7165)
);

INVx1_ASAP7_75t_L g7166 ( 
.A(n_6674),
.Y(n_7166)
);

INVx3_ASAP7_75t_L g7167 ( 
.A(n_6361),
.Y(n_7167)
);

NOR2xp33_ASAP7_75t_L g7168 ( 
.A(n_6653),
.B(n_3959),
.Y(n_7168)
);

INVx1_ASAP7_75t_L g7169 ( 
.A(n_6440),
.Y(n_7169)
);

BUFx6f_ASAP7_75t_L g7170 ( 
.A(n_6319),
.Y(n_7170)
);

INVxp67_ASAP7_75t_SL g7171 ( 
.A(n_6357),
.Y(n_7171)
);

INVx1_ASAP7_75t_L g7172 ( 
.A(n_6499),
.Y(n_7172)
);

INVx2_ASAP7_75t_SL g7173 ( 
.A(n_6474),
.Y(n_7173)
);

NAND2xp5_ASAP7_75t_SL g7174 ( 
.A(n_6655),
.B(n_3961),
.Y(n_7174)
);

NAND2xp5_ASAP7_75t_L g7175 ( 
.A(n_6791),
.B(n_3962),
.Y(n_7175)
);

INVxp67_ASAP7_75t_L g7176 ( 
.A(n_6464),
.Y(n_7176)
);

NAND2xp5_ASAP7_75t_SL g7177 ( 
.A(n_6677),
.B(n_3964),
.Y(n_7177)
);

OR2x2_ASAP7_75t_L g7178 ( 
.A(n_6792),
.B(n_3967),
.Y(n_7178)
);

INVx2_ASAP7_75t_L g7179 ( 
.A(n_6281),
.Y(n_7179)
);

NAND2xp5_ASAP7_75t_SL g7180 ( 
.A(n_6800),
.B(n_3968),
.Y(n_7180)
);

OR2x2_ASAP7_75t_L g7181 ( 
.A(n_6772),
.B(n_3973),
.Y(n_7181)
);

INVx2_ASAP7_75t_L g7182 ( 
.A(n_6288),
.Y(n_7182)
);

NAND2xp5_ASAP7_75t_L g7183 ( 
.A(n_6277),
.B(n_3982),
.Y(n_7183)
);

INVx1_ASAP7_75t_L g7184 ( 
.A(n_6463),
.Y(n_7184)
);

INVxp67_ASAP7_75t_L g7185 ( 
.A(n_6658),
.Y(n_7185)
);

AOI22xp5_ASAP7_75t_L g7186 ( 
.A1(n_6273),
.A2(n_3984),
.B1(n_3985),
.B2(n_3983),
.Y(n_7186)
);

AND2x4_ASAP7_75t_L g7187 ( 
.A(n_6402),
.B(n_3760),
.Y(n_7187)
);

INVx8_ASAP7_75t_L g7188 ( 
.A(n_6613),
.Y(n_7188)
);

NAND2xp5_ASAP7_75t_SL g7189 ( 
.A(n_6634),
.B(n_3987),
.Y(n_7189)
);

NAND2xp5_ASAP7_75t_L g7190 ( 
.A(n_6277),
.B(n_3991),
.Y(n_7190)
);

NAND2xp5_ASAP7_75t_SL g7191 ( 
.A(n_6434),
.B(n_3992),
.Y(n_7191)
);

NOR2xp33_ASAP7_75t_L g7192 ( 
.A(n_6542),
.B(n_3994),
.Y(n_7192)
);

NAND2xp5_ASAP7_75t_L g7193 ( 
.A(n_6635),
.B(n_3996),
.Y(n_7193)
);

AND2x4_ASAP7_75t_L g7194 ( 
.A(n_6406),
.B(n_3762),
.Y(n_7194)
);

INVx1_ASAP7_75t_L g7195 ( 
.A(n_6477),
.Y(n_7195)
);

INVx2_ASAP7_75t_L g7196 ( 
.A(n_6293),
.Y(n_7196)
);

AOI22xp5_ASAP7_75t_L g7197 ( 
.A1(n_6405),
.A2(n_4002),
.B1(n_4006),
.B2(n_3998),
.Y(n_7197)
);

NAND2xp5_ASAP7_75t_SL g7198 ( 
.A(n_6448),
.B(n_4008),
.Y(n_7198)
);

NOR2xp67_ASAP7_75t_L g7199 ( 
.A(n_6506),
.B(n_4013),
.Y(n_7199)
);

INVx1_ASAP7_75t_L g7200 ( 
.A(n_6495),
.Y(n_7200)
);

NAND2xp5_ASAP7_75t_L g7201 ( 
.A(n_6777),
.B(n_4014),
.Y(n_7201)
);

NAND2xp5_ASAP7_75t_L g7202 ( 
.A(n_6793),
.B(n_6584),
.Y(n_7202)
);

NAND2xp5_ASAP7_75t_L g7203 ( 
.A(n_6584),
.B(n_4015),
.Y(n_7203)
);

HB1xp67_ASAP7_75t_L g7204 ( 
.A(n_6613),
.Y(n_7204)
);

NAND2xp5_ASAP7_75t_L g7205 ( 
.A(n_6584),
.B(n_4017),
.Y(n_7205)
);

INVx1_ASAP7_75t_L g7206 ( 
.A(n_6597),
.Y(n_7206)
);

NOR2xp33_ASAP7_75t_L g7207 ( 
.A(n_6462),
.B(n_4027),
.Y(n_7207)
);

NOR2xp33_ASAP7_75t_L g7208 ( 
.A(n_6465),
.B(n_4028),
.Y(n_7208)
);

NAND2xp5_ASAP7_75t_L g7209 ( 
.A(n_6699),
.B(n_4029),
.Y(n_7209)
);

NOR2xp33_ASAP7_75t_L g7210 ( 
.A(n_6483),
.B(n_4031),
.Y(n_7210)
);

INVx5_ASAP7_75t_L g7211 ( 
.A(n_6372),
.Y(n_7211)
);

INVx1_ASAP7_75t_L g7212 ( 
.A(n_6606),
.Y(n_7212)
);

NAND2xp5_ASAP7_75t_L g7213 ( 
.A(n_6699),
.B(n_4036),
.Y(n_7213)
);

NOR2xp33_ASAP7_75t_L g7214 ( 
.A(n_6661),
.B(n_6664),
.Y(n_7214)
);

INVx2_ASAP7_75t_L g7215 ( 
.A(n_6324),
.Y(n_7215)
);

INVx2_ASAP7_75t_L g7216 ( 
.A(n_6337),
.Y(n_7216)
);

NOR3xp33_ASAP7_75t_L g7217 ( 
.A(n_6675),
.B(n_4043),
.C(n_4037),
.Y(n_7217)
);

AND2x2_ASAP7_75t_L g7218 ( 
.A(n_6594),
.B(n_4045),
.Y(n_7218)
);

NAND2xp33_ASAP7_75t_L g7219 ( 
.A(n_6699),
.B(n_4054),
.Y(n_7219)
);

INVx2_ASAP7_75t_L g7220 ( 
.A(n_6353),
.Y(n_7220)
);

NAND3xp33_ASAP7_75t_L g7221 ( 
.A(n_6533),
.B(n_6348),
.C(n_6317),
.Y(n_7221)
);

BUFx3_ASAP7_75t_L g7222 ( 
.A(n_6420),
.Y(n_7222)
);

INVxp67_ASAP7_75t_L g7223 ( 
.A(n_6687),
.Y(n_7223)
);

NAND2xp5_ASAP7_75t_L g7224 ( 
.A(n_6633),
.B(n_4057),
.Y(n_7224)
);

A2O1A1Ixp33_ASAP7_75t_L g7225 ( 
.A1(n_6513),
.A2(n_3763),
.B(n_3773),
.C(n_3771),
.Y(n_7225)
);

NAND2xp5_ASAP7_75t_SL g7226 ( 
.A(n_6266),
.B(n_4058),
.Y(n_7226)
);

CKINVDCx5p33_ASAP7_75t_R g7227 ( 
.A(n_6766),
.Y(n_7227)
);

NOR2xp33_ASAP7_75t_L g7228 ( 
.A(n_6694),
.B(n_6712),
.Y(n_7228)
);

CKINVDCx5p33_ASAP7_75t_R g7229 ( 
.A(n_6515),
.Y(n_7229)
);

INVx1_ASAP7_75t_L g7230 ( 
.A(n_6364),
.Y(n_7230)
);

INVx2_ASAP7_75t_L g7231 ( 
.A(n_6378),
.Y(n_7231)
);

NAND2xp5_ASAP7_75t_L g7232 ( 
.A(n_6383),
.B(n_4060),
.Y(n_7232)
);

HB1xp67_ASAP7_75t_L g7233 ( 
.A(n_6430),
.Y(n_7233)
);

NAND2xp33_ASAP7_75t_L g7234 ( 
.A(n_6357),
.B(n_4067),
.Y(n_7234)
);

INVx1_ASAP7_75t_L g7235 ( 
.A(n_6560),
.Y(n_7235)
);

NAND2xp5_ASAP7_75t_SL g7236 ( 
.A(n_6621),
.B(n_4068),
.Y(n_7236)
);

INVx1_ASAP7_75t_L g7237 ( 
.A(n_6571),
.Y(n_7237)
);

AOI221xp5_ASAP7_75t_L g7238 ( 
.A1(n_6723),
.A2(n_3793),
.B1(n_3802),
.B2(n_3797),
.C(n_3790),
.Y(n_7238)
);

BUFx6f_ASAP7_75t_L g7239 ( 
.A(n_6380),
.Y(n_7239)
);

BUFx6f_ASAP7_75t_SL g7240 ( 
.A(n_6296),
.Y(n_7240)
);

INVx1_ASAP7_75t_L g7241 ( 
.A(n_6493),
.Y(n_7241)
);

OAI22xp5_ASAP7_75t_L g7242 ( 
.A1(n_6300),
.A2(n_4072),
.B1(n_4073),
.B2(n_4071),
.Y(n_7242)
);

OAI22xp5_ASAP7_75t_L g7243 ( 
.A1(n_6775),
.A2(n_4075),
.B1(n_4078),
.B2(n_4074),
.Y(n_7243)
);

NAND2xp5_ASAP7_75t_L g7244 ( 
.A(n_6271),
.B(n_4081),
.Y(n_7244)
);

NAND2xp5_ASAP7_75t_SL g7245 ( 
.A(n_6621),
.B(n_6730),
.Y(n_7245)
);

INVx1_ASAP7_75t_L g7246 ( 
.A(n_6543),
.Y(n_7246)
);

NAND2xp5_ASAP7_75t_SL g7247 ( 
.A(n_6295),
.B(n_4083),
.Y(n_7247)
);

NAND2xp5_ASAP7_75t_L g7248 ( 
.A(n_6503),
.B(n_4084),
.Y(n_7248)
);

AOI22xp5_ASAP7_75t_L g7249 ( 
.A1(n_6511),
.A2(n_4091),
.B1(n_4095),
.B2(n_4090),
.Y(n_7249)
);

INVx2_ASAP7_75t_SL g7250 ( 
.A(n_6380),
.Y(n_7250)
);

NOR2xp33_ASAP7_75t_L g7251 ( 
.A(n_6728),
.B(n_4096),
.Y(n_7251)
);

INVx2_ASAP7_75t_L g7252 ( 
.A(n_6685),
.Y(n_7252)
);

NOR2xp33_ASAP7_75t_L g7253 ( 
.A(n_6750),
.B(n_4097),
.Y(n_7253)
);

NAND2xp5_ASAP7_75t_SL g7254 ( 
.A(n_6295),
.B(n_4099),
.Y(n_7254)
);

NAND2xp5_ASAP7_75t_L g7255 ( 
.A(n_6516),
.B(n_4100),
.Y(n_7255)
);

INVx1_ASAP7_75t_L g7256 ( 
.A(n_6399),
.Y(n_7256)
);

NAND2xp5_ASAP7_75t_SL g7257 ( 
.A(n_6304),
.B(n_4101),
.Y(n_7257)
);

BUFx5_ASAP7_75t_L g7258 ( 
.A(n_6514),
.Y(n_7258)
);

NOR2xp33_ASAP7_75t_L g7259 ( 
.A(n_6652),
.B(n_4102),
.Y(n_7259)
);

AND2x2_ASAP7_75t_L g7260 ( 
.A(n_6688),
.B(n_4103),
.Y(n_7260)
);

NAND2xp5_ASAP7_75t_SL g7261 ( 
.A(n_6304),
.B(n_4107),
.Y(n_7261)
);

NAND2xp5_ASAP7_75t_L g7262 ( 
.A(n_6535),
.B(n_6575),
.Y(n_7262)
);

NAND2xp5_ASAP7_75t_L g7263 ( 
.A(n_6600),
.B(n_4108),
.Y(n_7263)
);

NAND2xp5_ASAP7_75t_L g7264 ( 
.A(n_6611),
.B(n_4110),
.Y(n_7264)
);

NAND2xp33_ASAP7_75t_L g7265 ( 
.A(n_6399),
.B(n_4113),
.Y(n_7265)
);

OR2x6_ASAP7_75t_L g7266 ( 
.A(n_6272),
.B(n_3809),
.Y(n_7266)
);

INVx2_ASAP7_75t_L g7267 ( 
.A(n_6460),
.Y(n_7267)
);

NAND2xp5_ASAP7_75t_L g7268 ( 
.A(n_6436),
.B(n_4117),
.Y(n_7268)
);

INVx1_ASAP7_75t_L g7269 ( 
.A(n_6460),
.Y(n_7269)
);

INVx1_ASAP7_75t_SL g7270 ( 
.A(n_6696),
.Y(n_7270)
);

AND2x2_ASAP7_75t_SL g7271 ( 
.A(n_6676),
.B(n_3810),
.Y(n_7271)
);

AND2x2_ASAP7_75t_L g7272 ( 
.A(n_6769),
.B(n_4118),
.Y(n_7272)
);

INVxp33_ASAP7_75t_L g7273 ( 
.A(n_6741),
.Y(n_7273)
);

AND2x2_ASAP7_75t_SL g7274 ( 
.A(n_6622),
.B(n_3811),
.Y(n_7274)
);

NAND2xp5_ASAP7_75t_SL g7275 ( 
.A(n_6283),
.B(n_4119),
.Y(n_7275)
);

NAND2xp5_ASAP7_75t_L g7276 ( 
.A(n_6494),
.B(n_4122),
.Y(n_7276)
);

NAND2xp5_ASAP7_75t_L g7277 ( 
.A(n_6389),
.B(n_4124),
.Y(n_7277)
);

INVx1_ASAP7_75t_L g7278 ( 
.A(n_6496),
.Y(n_7278)
);

INVx2_ASAP7_75t_L g7279 ( 
.A(n_6496),
.Y(n_7279)
);

INVxp67_ASAP7_75t_L g7280 ( 
.A(n_6722),
.Y(n_7280)
);

NOR2xp33_ASAP7_75t_L g7281 ( 
.A(n_6704),
.B(n_4126),
.Y(n_7281)
);

NOR2xp33_ASAP7_75t_L g7282 ( 
.A(n_6707),
.B(n_4128),
.Y(n_7282)
);

AND2x4_ASAP7_75t_L g7283 ( 
.A(n_6546),
.B(n_3817),
.Y(n_7283)
);

INVx1_ASAP7_75t_L g7284 ( 
.A(n_6572),
.Y(n_7284)
);

INVx2_ASAP7_75t_L g7285 ( 
.A(n_6572),
.Y(n_7285)
);

AND2x2_ASAP7_75t_L g7286 ( 
.A(n_6771),
.B(n_4129),
.Y(n_7286)
);

INVx1_ASAP7_75t_L g7287 ( 
.A(n_6581),
.Y(n_7287)
);

INVxp33_ASAP7_75t_L g7288 ( 
.A(n_6753),
.Y(n_7288)
);

NAND2xp5_ASAP7_75t_L g7289 ( 
.A(n_6646),
.B(n_4130),
.Y(n_7289)
);

INVx2_ASAP7_75t_L g7290 ( 
.A(n_6581),
.Y(n_7290)
);

NOR2xp33_ASAP7_75t_L g7291 ( 
.A(n_6779),
.B(n_6395),
.Y(n_7291)
);

HB1xp67_ASAP7_75t_L g7292 ( 
.A(n_6592),
.Y(n_7292)
);

NAND2xp5_ASAP7_75t_L g7293 ( 
.A(n_6797),
.B(n_4132),
.Y(n_7293)
);

NAND2xp5_ASAP7_75t_L g7294 ( 
.A(n_6410),
.B(n_4135),
.Y(n_7294)
);

INVx2_ASAP7_75t_SL g7295 ( 
.A(n_6592),
.Y(n_7295)
);

INVx1_ASAP7_75t_L g7296 ( 
.A(n_6614),
.Y(n_7296)
);

INVx1_ASAP7_75t_L g7297 ( 
.A(n_6614),
.Y(n_7297)
);

OR2x6_ASAP7_75t_L g7298 ( 
.A(n_6343),
.B(n_3819),
.Y(n_7298)
);

NAND2xp5_ASAP7_75t_L g7299 ( 
.A(n_6443),
.B(n_4137),
.Y(n_7299)
);

NOR2xp33_ASAP7_75t_L g7300 ( 
.A(n_6454),
.B(n_4140),
.Y(n_7300)
);

INVx2_ASAP7_75t_L g7301 ( 
.A(n_6705),
.Y(n_7301)
);

INVx1_ASAP7_75t_L g7302 ( 
.A(n_6705),
.Y(n_7302)
);

BUFx4_ASAP7_75t_L g7303 ( 
.A(n_6798),
.Y(n_7303)
);

NAND2xp5_ASAP7_75t_SL g7304 ( 
.A(n_6344),
.B(n_4142),
.Y(n_7304)
);

NAND2xp5_ASAP7_75t_L g7305 ( 
.A(n_6452),
.B(n_4143),
.Y(n_7305)
);

INVx1_ASAP7_75t_L g7306 ( 
.A(n_6589),
.Y(n_7306)
);

NAND2xp5_ASAP7_75t_SL g7307 ( 
.A(n_6480),
.B(n_4144),
.Y(n_7307)
);

NAND2xp5_ASAP7_75t_L g7308 ( 
.A(n_6323),
.B(n_4147),
.Y(n_7308)
);

INVx5_ASAP7_75t_L g7309 ( 
.A(n_6425),
.Y(n_7309)
);

NAND2xp5_ASAP7_75t_L g7310 ( 
.A(n_6697),
.B(n_4150),
.Y(n_7310)
);

INVx1_ASAP7_75t_L g7311 ( 
.A(n_6556),
.Y(n_7311)
);

AND2x4_ASAP7_75t_L g7312 ( 
.A(n_7211),
.B(n_6527),
.Y(n_7312)
);

NAND2x1p5_ASAP7_75t_L g7313 ( 
.A(n_7211),
.B(n_6532),
.Y(n_7313)
);

NAND2xp5_ASAP7_75t_SL g7314 ( 
.A(n_7019),
.B(n_6716),
.Y(n_7314)
);

INVx1_ASAP7_75t_L g7315 ( 
.A(n_6808),
.Y(n_7315)
);

INVx1_ASAP7_75t_SL g7316 ( 
.A(n_6855),
.Y(n_7316)
);

INVx1_ASAP7_75t_L g7317 ( 
.A(n_6810),
.Y(n_7317)
);

INVx1_ASAP7_75t_L g7318 ( 
.A(n_6823),
.Y(n_7318)
);

INVx1_ASAP7_75t_L g7319 ( 
.A(n_6825),
.Y(n_7319)
);

INVx2_ASAP7_75t_L g7320 ( 
.A(n_6829),
.Y(n_7320)
);

INVx1_ASAP7_75t_L g7321 ( 
.A(n_6845),
.Y(n_7321)
);

INVx2_ASAP7_75t_L g7322 ( 
.A(n_6847),
.Y(n_7322)
);

AO22x2_ASAP7_75t_L g7323 ( 
.A1(n_6851),
.A2(n_6731),
.B1(n_6566),
.B2(n_6787),
.Y(n_7323)
);

INVx1_ASAP7_75t_L g7324 ( 
.A(n_6848),
.Y(n_7324)
);

BUFx2_ASAP7_75t_L g7325 ( 
.A(n_6901),
.Y(n_7325)
);

BUFx6f_ASAP7_75t_SL g7326 ( 
.A(n_6866),
.Y(n_7326)
);

AOI22xp5_ASAP7_75t_L g7327 ( 
.A1(n_6867),
.A2(n_6717),
.B1(n_6729),
.B2(n_6727),
.Y(n_7327)
);

INVx2_ASAP7_75t_L g7328 ( 
.A(n_6856),
.Y(n_7328)
);

AND2x4_ASAP7_75t_L g7329 ( 
.A(n_6922),
.B(n_6534),
.Y(n_7329)
);

NOR2xp33_ASAP7_75t_L g7330 ( 
.A(n_7075),
.B(n_6537),
.Y(n_7330)
);

AND2x4_ASAP7_75t_L g7331 ( 
.A(n_7046),
.B(n_6650),
.Y(n_7331)
);

BUFx8_ASAP7_75t_L g7332 ( 
.A(n_6836),
.Y(n_7332)
);

INVx1_ASAP7_75t_L g7333 ( 
.A(n_6871),
.Y(n_7333)
);

AO22x1_ASAP7_75t_L g7334 ( 
.A1(n_6844),
.A2(n_6691),
.B1(n_6748),
.B2(n_6738),
.Y(n_7334)
);

INVx1_ASAP7_75t_L g7335 ( 
.A(n_6890),
.Y(n_7335)
);

OAI221xp5_ASAP7_75t_L g7336 ( 
.A1(n_7002),
.A2(n_6573),
.B1(n_6732),
.B2(n_6725),
.C(n_6651),
.Y(n_7336)
);

BUFx8_ASAP7_75t_L g7337 ( 
.A(n_7000),
.Y(n_7337)
);

INVx1_ASAP7_75t_L g7338 ( 
.A(n_6905),
.Y(n_7338)
);

INVx2_ASAP7_75t_L g7339 ( 
.A(n_6917),
.Y(n_7339)
);

INVx1_ASAP7_75t_L g7340 ( 
.A(n_6924),
.Y(n_7340)
);

INVx1_ASAP7_75t_L g7341 ( 
.A(n_6926),
.Y(n_7341)
);

INVx1_ASAP7_75t_L g7342 ( 
.A(n_6932),
.Y(n_7342)
);

AND2x2_ASAP7_75t_L g7343 ( 
.A(n_7050),
.B(n_6412),
.Y(n_7343)
);

CKINVDCx5p33_ASAP7_75t_R g7344 ( 
.A(n_7140),
.Y(n_7344)
);

NAND2xp5_ASAP7_75t_SL g7345 ( 
.A(n_7005),
.B(n_6776),
.Y(n_7345)
);

INVxp67_ASAP7_75t_L g7346 ( 
.A(n_6850),
.Y(n_7346)
);

NAND2x1p5_ASAP7_75t_L g7347 ( 
.A(n_7147),
.B(n_6309),
.Y(n_7347)
);

INVx2_ASAP7_75t_L g7348 ( 
.A(n_6934),
.Y(n_7348)
);

INVx1_ASAP7_75t_L g7349 ( 
.A(n_6880),
.Y(n_7349)
);

NAND2x1p5_ASAP7_75t_L g7350 ( 
.A(n_7167),
.B(n_6371),
.Y(n_7350)
);

INVx1_ASAP7_75t_L g7351 ( 
.A(n_6912),
.Y(n_7351)
);

NAND2xp5_ASAP7_75t_L g7352 ( 
.A(n_6830),
.B(n_6788),
.Y(n_7352)
);

INVx1_ASAP7_75t_L g7353 ( 
.A(n_6916),
.Y(n_7353)
);

AO22x2_ASAP7_75t_L g7354 ( 
.A1(n_6875),
.A2(n_3823),
.B1(n_3829),
.B2(n_3825),
.Y(n_7354)
);

OAI221xp5_ASAP7_75t_L g7355 ( 
.A1(n_6915),
.A2(n_6573),
.B1(n_6732),
.B2(n_6637),
.C(n_6412),
.Y(n_7355)
);

XNOR2xp5_ASAP7_75t_L g7356 ( 
.A(n_6994),
.B(n_6802),
.Y(n_7356)
);

INVx1_ASAP7_75t_L g7357 ( 
.A(n_6933),
.Y(n_7357)
);

INVx1_ASAP7_75t_L g7358 ( 
.A(n_6964),
.Y(n_7358)
);

INVx1_ASAP7_75t_L g7359 ( 
.A(n_6965),
.Y(n_7359)
);

NAND2xp5_ASAP7_75t_L g7360 ( 
.A(n_6812),
.B(n_6807),
.Y(n_7360)
);

AOI22xp33_ASAP7_75t_L g7361 ( 
.A1(n_6892),
.A2(n_6605),
.B1(n_6349),
.B2(n_6428),
.Y(n_7361)
);

INVx1_ASAP7_75t_L g7362 ( 
.A(n_6973),
.Y(n_7362)
);

AO22x2_ASAP7_75t_L g7363 ( 
.A1(n_6947),
.A2(n_3830),
.B1(n_3840),
.B2(n_3832),
.Y(n_7363)
);

NAND2xp5_ASAP7_75t_L g7364 ( 
.A(n_6813),
.B(n_6605),
.Y(n_7364)
);

OAI22xp33_ASAP7_75t_SL g7365 ( 
.A1(n_7056),
.A2(n_6349),
.B1(n_6637),
.B2(n_6428),
.Y(n_7365)
);

NAND2x1p5_ASAP7_75t_L g7366 ( 
.A(n_7222),
.B(n_6803),
.Y(n_7366)
);

CKINVDCx11_ASAP7_75t_R g7367 ( 
.A(n_6960),
.Y(n_7367)
);

INVx2_ASAP7_75t_L g7368 ( 
.A(n_6975),
.Y(n_7368)
);

INVx5_ASAP7_75t_L g7369 ( 
.A(n_6988),
.Y(n_7369)
);

INVx1_ASAP7_75t_L g7370 ( 
.A(n_6976),
.Y(n_7370)
);

AO22x2_ASAP7_75t_L g7371 ( 
.A1(n_6863),
.A2(n_3842),
.B1(n_3856),
.B2(n_3854),
.Y(n_7371)
);

INVx1_ASAP7_75t_L g7372 ( 
.A(n_6978),
.Y(n_7372)
);

OAI221xp5_ASAP7_75t_L g7373 ( 
.A1(n_6906),
.A2(n_6759),
.B1(n_3874),
.B2(n_3892),
.C(n_3882),
.Y(n_7373)
);

AO22x2_ASAP7_75t_L g7374 ( 
.A1(n_7311),
.A2(n_3867),
.B1(n_3903),
.B2(n_3900),
.Y(n_7374)
);

INVx1_ASAP7_75t_L g7375 ( 
.A(n_6979),
.Y(n_7375)
);

AND2x2_ASAP7_75t_L g7376 ( 
.A(n_6858),
.B(n_6437),
.Y(n_7376)
);

INVx2_ASAP7_75t_L g7377 ( 
.A(n_6984),
.Y(n_7377)
);

NAND2xp5_ASAP7_75t_L g7378 ( 
.A(n_6888),
.B(n_6541),
.Y(n_7378)
);

AOI22xp5_ASAP7_75t_L g7379 ( 
.A1(n_6843),
.A2(n_6595),
.B1(n_6789),
.B2(n_6385),
.Y(n_7379)
);

AO22x2_ASAP7_75t_L g7380 ( 
.A1(n_6872),
.A2(n_3906),
.B1(n_3923),
.B2(n_3913),
.Y(n_7380)
);

NAND2xp33_ASAP7_75t_L g7381 ( 
.A(n_7258),
.B(n_6759),
.Y(n_7381)
);

NAND2xp5_ASAP7_75t_L g7382 ( 
.A(n_7107),
.B(n_6781),
.Y(n_7382)
);

INVx3_ASAP7_75t_L g7383 ( 
.A(n_6988),
.Y(n_7383)
);

NAND2xp5_ASAP7_75t_L g7384 ( 
.A(n_7143),
.B(n_6668),
.Y(n_7384)
);

AO22x2_ASAP7_75t_L g7385 ( 
.A1(n_7221),
.A2(n_3924),
.B1(n_3932),
.B2(n_3927),
.Y(n_7385)
);

INVx3_ASAP7_75t_L g7386 ( 
.A(n_7028),
.Y(n_7386)
);

NAND2x1p5_ASAP7_75t_L g7387 ( 
.A(n_6885),
.B(n_6909),
.Y(n_7387)
);

INVx1_ASAP7_75t_L g7388 ( 
.A(n_7057),
.Y(n_7388)
);

INVx1_ASAP7_75t_L g7389 ( 
.A(n_6985),
.Y(n_7389)
);

AND2x2_ASAP7_75t_L g7390 ( 
.A(n_7065),
.B(n_6522),
.Y(n_7390)
);

AO22x2_ASAP7_75t_L g7391 ( 
.A1(n_7007),
.A2(n_3950),
.B1(n_3960),
.B2(n_3957),
.Y(n_7391)
);

AO22x2_ASAP7_75t_L g7392 ( 
.A1(n_7165),
.A2(n_3963),
.B1(n_3974),
.B2(n_3970),
.Y(n_7392)
);

INVx1_ASAP7_75t_L g7393 ( 
.A(n_7011),
.Y(n_7393)
);

INVxp67_ASAP7_75t_L g7394 ( 
.A(n_7049),
.Y(n_7394)
);

CKINVDCx5p33_ASAP7_75t_R g7395 ( 
.A(n_7149),
.Y(n_7395)
);

AO22x2_ASAP7_75t_L g7396 ( 
.A1(n_7302),
.A2(n_3975),
.B1(n_3988),
.B2(n_3976),
.Y(n_7396)
);

AND2x4_ASAP7_75t_L g7397 ( 
.A(n_7112),
.B(n_6816),
.Y(n_7397)
);

NAND2xp5_ASAP7_75t_L g7398 ( 
.A(n_7151),
.B(n_4000),
.Y(n_7398)
);

HB1xp67_ASAP7_75t_L g7399 ( 
.A(n_6852),
.Y(n_7399)
);

AO22x2_ASAP7_75t_L g7400 ( 
.A1(n_7242),
.A2(n_6809),
.B1(n_7082),
.B2(n_6814),
.Y(n_7400)
);

NAND2xp5_ASAP7_75t_L g7401 ( 
.A(n_7153),
.B(n_4001),
.Y(n_7401)
);

CKINVDCx5p33_ASAP7_75t_R g7402 ( 
.A(n_7227),
.Y(n_7402)
);

AND2x4_ASAP7_75t_L g7403 ( 
.A(n_7233),
.B(n_6591),
.Y(n_7403)
);

INVx2_ASAP7_75t_L g7404 ( 
.A(n_6811),
.Y(n_7404)
);

INVx1_ASAP7_75t_L g7405 ( 
.A(n_7031),
.Y(n_7405)
);

INVx1_ASAP7_75t_L g7406 ( 
.A(n_7033),
.Y(n_7406)
);

INVx1_ASAP7_75t_L g7407 ( 
.A(n_7038),
.Y(n_7407)
);

NAND2x1p5_ASAP7_75t_L g7408 ( 
.A(n_6885),
.B(n_4003),
.Y(n_7408)
);

AND2x4_ASAP7_75t_L g7409 ( 
.A(n_6894),
.B(n_4007),
.Y(n_7409)
);

AO22x2_ASAP7_75t_L g7410 ( 
.A1(n_7301),
.A2(n_4009),
.B1(n_4023),
.B2(n_4021),
.Y(n_7410)
);

AO22x2_ASAP7_75t_L g7411 ( 
.A1(n_6822),
.A2(n_4024),
.B1(n_4041),
.B2(n_4026),
.Y(n_7411)
);

INVx1_ASAP7_75t_L g7412 ( 
.A(n_7039),
.Y(n_7412)
);

CKINVDCx16_ASAP7_75t_R g7413 ( 
.A(n_7240),
.Y(n_7413)
);

AND2x2_ASAP7_75t_L g7414 ( 
.A(n_7076),
.B(n_4153),
.Y(n_7414)
);

BUFx8_ASAP7_75t_L g7415 ( 
.A(n_7258),
.Y(n_7415)
);

NAND2xp5_ASAP7_75t_L g7416 ( 
.A(n_7161),
.B(n_4042),
.Y(n_7416)
);

INVx1_ASAP7_75t_L g7417 ( 
.A(n_7041),
.Y(n_7417)
);

NAND2xp5_ASAP7_75t_L g7418 ( 
.A(n_7162),
.B(n_4055),
.Y(n_7418)
);

OAI221xp5_ASAP7_75t_L g7419 ( 
.A1(n_6920),
.A2(n_4082),
.B1(n_4105),
.B2(n_4098),
.C(n_4069),
.Y(n_7419)
);

INVx2_ASAP7_75t_SL g7420 ( 
.A(n_7028),
.Y(n_7420)
);

INVx2_ASAP7_75t_L g7421 ( 
.A(n_6815),
.Y(n_7421)
);

OR2x6_ASAP7_75t_L g7422 ( 
.A(n_7188),
.B(n_4109),
.Y(n_7422)
);

INVx1_ASAP7_75t_L g7423 ( 
.A(n_7060),
.Y(n_7423)
);

NOR2xp67_ASAP7_75t_L g7424 ( 
.A(n_6857),
.B(n_5),
.Y(n_7424)
);

INVx1_ASAP7_75t_L g7425 ( 
.A(n_7062),
.Y(n_7425)
);

INVx2_ASAP7_75t_L g7426 ( 
.A(n_6854),
.Y(n_7426)
);

NAND2x1p5_ASAP7_75t_L g7427 ( 
.A(n_6909),
.B(n_4116),
.Y(n_7427)
);

AO22x2_ASAP7_75t_L g7428 ( 
.A1(n_6838),
.A2(n_4125),
.B1(n_4139),
.B2(n_4131),
.Y(n_7428)
);

INVx2_ASAP7_75t_L g7429 ( 
.A(n_6860),
.Y(n_7429)
);

AND2x4_ASAP7_75t_L g7430 ( 
.A(n_6902),
.B(n_4141),
.Y(n_7430)
);

AND2x4_ASAP7_75t_L g7431 ( 
.A(n_6971),
.B(n_4146),
.Y(n_7431)
);

INVx1_ASAP7_75t_L g7432 ( 
.A(n_6868),
.Y(n_7432)
);

NAND2xp33_ASAP7_75t_L g7433 ( 
.A(n_7258),
.B(n_4156),
.Y(n_7433)
);

INVx2_ASAP7_75t_L g7434 ( 
.A(n_6869),
.Y(n_7434)
);

INVx1_ASAP7_75t_L g7435 ( 
.A(n_6873),
.Y(n_7435)
);

CKINVDCx5p33_ASAP7_75t_R g7436 ( 
.A(n_7229),
.Y(n_7436)
);

HAxp5_ASAP7_75t_SL g7437 ( 
.A(n_6983),
.B(n_4148),
.CON(n_7437),
.SN(n_7437)
);

INVx2_ASAP7_75t_L g7438 ( 
.A(n_6882),
.Y(n_7438)
);

INVx2_ASAP7_75t_L g7439 ( 
.A(n_6897),
.Y(n_7439)
);

NOR2xp33_ASAP7_75t_L g7440 ( 
.A(n_6817),
.B(n_4157),
.Y(n_7440)
);

INVxp67_ASAP7_75t_L g7441 ( 
.A(n_7139),
.Y(n_7441)
);

INVxp67_ASAP7_75t_L g7442 ( 
.A(n_7181),
.Y(n_7442)
);

OA22x2_ASAP7_75t_L g7443 ( 
.A1(n_6921),
.A2(n_4160),
.B1(n_4165),
.B2(n_4159),
.Y(n_7443)
);

INVx1_ASAP7_75t_L g7444 ( 
.A(n_6898),
.Y(n_7444)
);

INVx1_ASAP7_75t_L g7445 ( 
.A(n_6913),
.Y(n_7445)
);

NOR2xp33_ASAP7_75t_L g7446 ( 
.A(n_6938),
.B(n_6952),
.Y(n_7446)
);

NOR2xp33_ASAP7_75t_L g7447 ( 
.A(n_6835),
.B(n_4169),
.Y(n_7447)
);

INVx1_ASAP7_75t_L g7448 ( 
.A(n_6925),
.Y(n_7448)
);

OAI221xp5_ASAP7_75t_L g7449 ( 
.A1(n_7064),
.A2(n_4152),
.B1(n_4158),
.B2(n_4154),
.C(n_4151),
.Y(n_7449)
);

AND2x2_ASAP7_75t_L g7450 ( 
.A(n_6958),
.B(n_4170),
.Y(n_7450)
);

OAI221xp5_ASAP7_75t_L g7451 ( 
.A1(n_7066),
.A2(n_4163),
.B1(n_4166),
.B2(n_4164),
.C(n_4162),
.Y(n_7451)
);

AND2x4_ASAP7_75t_L g7452 ( 
.A(n_6971),
.B(n_4167),
.Y(n_7452)
);

INVx1_ASAP7_75t_L g7453 ( 
.A(n_6940),
.Y(n_7453)
);

NAND2xp5_ASAP7_75t_L g7454 ( 
.A(n_6956),
.B(n_4172),
.Y(n_7454)
);

OAI22xp5_ASAP7_75t_L g7455 ( 
.A1(n_6961),
.A2(n_6833),
.B1(n_6841),
.B2(n_6831),
.Y(n_7455)
);

NAND2xp5_ASAP7_75t_L g7456 ( 
.A(n_7166),
.B(n_4173),
.Y(n_7456)
);

INVx1_ASAP7_75t_L g7457 ( 
.A(n_7138),
.Y(n_7457)
);

NAND2xp5_ASAP7_75t_L g7458 ( 
.A(n_7068),
.B(n_4175),
.Y(n_7458)
);

AO22x2_ASAP7_75t_L g7459 ( 
.A1(n_7202),
.A2(n_3729),
.B1(n_8),
.B2(n_6),
.Y(n_7459)
);

BUFx8_ASAP7_75t_L g7460 ( 
.A(n_7258),
.Y(n_7460)
);

NAND2xp5_ASAP7_75t_L g7461 ( 
.A(n_6821),
.B(n_4176),
.Y(n_7461)
);

INVx1_ASAP7_75t_L g7462 ( 
.A(n_7063),
.Y(n_7462)
);

INVxp67_ASAP7_75t_L g7463 ( 
.A(n_7292),
.Y(n_7463)
);

OAI221xp5_ASAP7_75t_L g7464 ( 
.A1(n_7168),
.A2(n_6997),
.B1(n_7208),
.B2(n_7210),
.C(n_7207),
.Y(n_7464)
);

INVx1_ASAP7_75t_L g7465 ( 
.A(n_6948),
.Y(n_7465)
);

NAND2xp5_ASAP7_75t_L g7466 ( 
.A(n_6826),
.B(n_4177),
.Y(n_7466)
);

AO22x2_ASAP7_75t_L g7467 ( 
.A1(n_7137),
.A2(n_8),
.B1(n_6),
.B2(n_7),
.Y(n_7467)
);

INVx1_ASAP7_75t_L g7468 ( 
.A(n_6951),
.Y(n_7468)
);

AO22x2_ASAP7_75t_L g7469 ( 
.A1(n_6874),
.A2(n_8),
.B1(n_6),
.B2(n_7),
.Y(n_7469)
);

HB1xp67_ASAP7_75t_L g7470 ( 
.A(n_6879),
.Y(n_7470)
);

NOR2xp33_ASAP7_75t_L g7471 ( 
.A(n_6834),
.B(n_4181),
.Y(n_7471)
);

AO22x2_ASAP7_75t_L g7472 ( 
.A1(n_6904),
.A2(n_10),
.B1(n_7),
.B2(n_9),
.Y(n_7472)
);

OAI221xp5_ASAP7_75t_L g7473 ( 
.A1(n_7251),
.A2(n_4186),
.B1(n_4189),
.B2(n_4184),
.C(n_4182),
.Y(n_7473)
);

INVx1_ASAP7_75t_L g7474 ( 
.A(n_6955),
.Y(n_7474)
);

AO22x2_ASAP7_75t_L g7475 ( 
.A1(n_7252),
.A2(n_11),
.B1(n_9),
.B2(n_10),
.Y(n_7475)
);

INVx4_ASAP7_75t_SL g7476 ( 
.A(n_6911),
.Y(n_7476)
);

INVx1_ASAP7_75t_L g7477 ( 
.A(n_6972),
.Y(n_7477)
);

INVx1_ASAP7_75t_L g7478 ( 
.A(n_7021),
.Y(n_7478)
);

BUFx6f_ASAP7_75t_L g7479 ( 
.A(n_7188),
.Y(n_7479)
);

INVx1_ASAP7_75t_L g7480 ( 
.A(n_7026),
.Y(n_7480)
);

INVx2_ASAP7_75t_L g7481 ( 
.A(n_7048),
.Y(n_7481)
);

INVx1_ASAP7_75t_L g7482 ( 
.A(n_7070),
.Y(n_7482)
);

INVx2_ASAP7_75t_L g7483 ( 
.A(n_7078),
.Y(n_7483)
);

NAND2xp5_ASAP7_75t_L g7484 ( 
.A(n_6832),
.B(n_4194),
.Y(n_7484)
);

NAND2xp5_ASAP7_75t_L g7485 ( 
.A(n_7106),
.B(n_9),
.Y(n_7485)
);

OAI22xp5_ASAP7_75t_L g7486 ( 
.A1(n_7029),
.A2(n_568),
.B1(n_569),
.B2(n_567),
.Y(n_7486)
);

INVx2_ASAP7_75t_L g7487 ( 
.A(n_7080),
.Y(n_7487)
);

INVx1_ASAP7_75t_L g7488 ( 
.A(n_7114),
.Y(n_7488)
);

INVx1_ASAP7_75t_L g7489 ( 
.A(n_7117),
.Y(n_7489)
);

NOR2xp33_ASAP7_75t_L g7490 ( 
.A(n_6842),
.B(n_567),
.Y(n_7490)
);

AO22x2_ASAP7_75t_L g7491 ( 
.A1(n_7183),
.A2(n_12),
.B1(n_10),
.B2(n_11),
.Y(n_7491)
);

AND2x4_ASAP7_75t_L g7492 ( 
.A(n_7241),
.B(n_568),
.Y(n_7492)
);

HB1xp67_ASAP7_75t_L g7493 ( 
.A(n_7270),
.Y(n_7493)
);

INVx1_ASAP7_75t_L g7494 ( 
.A(n_7129),
.Y(n_7494)
);

AOI22xp5_ASAP7_75t_L g7495 ( 
.A1(n_6987),
.A2(n_572),
.B1(n_573),
.B2(n_570),
.Y(n_7495)
);

NAND2x1p5_ASAP7_75t_L g7496 ( 
.A(n_6911),
.B(n_572),
.Y(n_7496)
);

NAND2xp5_ASAP7_75t_L g7497 ( 
.A(n_6876),
.B(n_11),
.Y(n_7497)
);

NOR2xp33_ASAP7_75t_SL g7498 ( 
.A(n_6959),
.B(n_12),
.Y(n_7498)
);

BUFx3_ASAP7_75t_L g7499 ( 
.A(n_6950),
.Y(n_7499)
);

INVx1_ASAP7_75t_L g7500 ( 
.A(n_7133),
.Y(n_7500)
);

NAND2x1p5_ASAP7_75t_L g7501 ( 
.A(n_6950),
.B(n_573),
.Y(n_7501)
);

AO22x2_ASAP7_75t_L g7502 ( 
.A1(n_7190),
.A2(n_15),
.B1(n_13),
.B2(n_14),
.Y(n_7502)
);

INVx1_ASAP7_75t_L g7503 ( 
.A(n_7083),
.Y(n_7503)
);

NAND2xp5_ASAP7_75t_L g7504 ( 
.A(n_6828),
.B(n_13),
.Y(n_7504)
);

INVx1_ASAP7_75t_L g7505 ( 
.A(n_7092),
.Y(n_7505)
);

INVx1_ASAP7_75t_L g7506 ( 
.A(n_7093),
.Y(n_7506)
);

NAND2xp5_ASAP7_75t_L g7507 ( 
.A(n_7081),
.B(n_13),
.Y(n_7507)
);

NAND2x1p5_ASAP7_75t_L g7508 ( 
.A(n_7010),
.B(n_574),
.Y(n_7508)
);

AO22x2_ASAP7_75t_L g7509 ( 
.A1(n_7099),
.A2(n_16),
.B1(n_14),
.B2(n_15),
.Y(n_7509)
);

NAND2xp5_ASAP7_75t_L g7510 ( 
.A(n_6859),
.B(n_15),
.Y(n_7510)
);

OAI221xp5_ASAP7_75t_L g7511 ( 
.A1(n_7253),
.A2(n_18),
.B1(n_16),
.B2(n_17),
.C(n_19),
.Y(n_7511)
);

INVx1_ASAP7_75t_L g7512 ( 
.A(n_7096),
.Y(n_7512)
);

INVx1_ASAP7_75t_L g7513 ( 
.A(n_7120),
.Y(n_7513)
);

NAND2xp5_ASAP7_75t_L g7514 ( 
.A(n_6865),
.B(n_16),
.Y(n_7514)
);

AOI22xp33_ASAP7_75t_L g7515 ( 
.A1(n_6864),
.A2(n_19),
.B1(n_17),
.B2(n_18),
.Y(n_7515)
);

BUFx3_ASAP7_75t_L g7516 ( 
.A(n_7010),
.Y(n_7516)
);

BUFx6f_ASAP7_75t_SL g7517 ( 
.A(n_7274),
.Y(n_7517)
);

BUFx6f_ASAP7_75t_L g7518 ( 
.A(n_7113),
.Y(n_7518)
);

INVx1_ASAP7_75t_L g7519 ( 
.A(n_7123),
.Y(n_7519)
);

INVx1_ASAP7_75t_L g7520 ( 
.A(n_7154),
.Y(n_7520)
);

INVx1_ASAP7_75t_L g7521 ( 
.A(n_7159),
.Y(n_7521)
);

INVx2_ASAP7_75t_L g7522 ( 
.A(n_7179),
.Y(n_7522)
);

INVx1_ASAP7_75t_L g7523 ( 
.A(n_7182),
.Y(n_7523)
);

OAI22xp5_ASAP7_75t_L g7524 ( 
.A1(n_6990),
.A2(n_576),
.B1(n_577),
.B2(n_575),
.Y(n_7524)
);

NAND2x1p5_ASAP7_75t_L g7525 ( 
.A(n_7113),
.B(n_7170),
.Y(n_7525)
);

AND2x4_ASAP7_75t_L g7526 ( 
.A(n_7246),
.B(n_575),
.Y(n_7526)
);

AOI22xp5_ASAP7_75t_L g7527 ( 
.A1(n_7077),
.A2(n_577),
.B1(n_578),
.B2(n_576),
.Y(n_7527)
);

INVx1_ASAP7_75t_L g7528 ( 
.A(n_7196),
.Y(n_7528)
);

OAI22xp5_ASAP7_75t_SL g7529 ( 
.A1(n_6824),
.A2(n_19),
.B1(n_17),
.B2(n_18),
.Y(n_7529)
);

NAND2xp5_ASAP7_75t_SL g7530 ( 
.A(n_6954),
.B(n_579),
.Y(n_7530)
);

INVx1_ASAP7_75t_L g7531 ( 
.A(n_7215),
.Y(n_7531)
);

INVx1_ASAP7_75t_L g7532 ( 
.A(n_7216),
.Y(n_7532)
);

NAND2x1p5_ASAP7_75t_L g7533 ( 
.A(n_7170),
.B(n_580),
.Y(n_7533)
);

INVx1_ASAP7_75t_L g7534 ( 
.A(n_7220),
.Y(n_7534)
);

AO22x2_ASAP7_75t_L g7535 ( 
.A1(n_7124),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.Y(n_7535)
);

INVx1_ASAP7_75t_L g7536 ( 
.A(n_7231),
.Y(n_7536)
);

AOI22xp5_ASAP7_75t_L g7537 ( 
.A1(n_6819),
.A2(n_584),
.B1(n_585),
.B2(n_582),
.Y(n_7537)
);

INVx2_ASAP7_75t_L g7538 ( 
.A(n_7169),
.Y(n_7538)
);

NAND3xp33_ASAP7_75t_SL g7539 ( 
.A(n_6963),
.B(n_20),
.C(n_21),
.Y(n_7539)
);

OAI221xp5_ASAP7_75t_L g7540 ( 
.A1(n_7100),
.A2(n_23),
.B1(n_21),
.B2(n_22),
.C(n_24),
.Y(n_7540)
);

INVxp67_ASAP7_75t_L g7541 ( 
.A(n_7085),
.Y(n_7541)
);

INVx1_ASAP7_75t_L g7542 ( 
.A(n_7184),
.Y(n_7542)
);

AND2x2_ASAP7_75t_L g7543 ( 
.A(n_6999),
.B(n_584),
.Y(n_7543)
);

HB1xp67_ASAP7_75t_L g7544 ( 
.A(n_7239),
.Y(n_7544)
);

NAND2x1p5_ASAP7_75t_L g7545 ( 
.A(n_7239),
.B(n_585),
.Y(n_7545)
);

BUFx3_ASAP7_75t_L g7546 ( 
.A(n_7059),
.Y(n_7546)
);

NAND2x1p5_ASAP7_75t_L g7547 ( 
.A(n_7309),
.B(n_587),
.Y(n_7547)
);

OAI221xp5_ASAP7_75t_L g7548 ( 
.A1(n_7108),
.A2(n_24),
.B1(n_22),
.B2(n_23),
.C(n_25),
.Y(n_7548)
);

INVx1_ASAP7_75t_L g7549 ( 
.A(n_7195),
.Y(n_7549)
);

INVx1_ASAP7_75t_L g7550 ( 
.A(n_7200),
.Y(n_7550)
);

AND2x2_ASAP7_75t_L g7551 ( 
.A(n_7030),
.B(n_7037),
.Y(n_7551)
);

NOR2xp33_ASAP7_75t_L g7552 ( 
.A(n_7035),
.B(n_587),
.Y(n_7552)
);

HB1xp67_ASAP7_75t_L g7553 ( 
.A(n_7040),
.Y(n_7553)
);

NAND2xp5_ASAP7_75t_L g7554 ( 
.A(n_6939),
.B(n_24),
.Y(n_7554)
);

AND2x4_ASAP7_75t_L g7555 ( 
.A(n_7306),
.B(n_588),
.Y(n_7555)
);

AOI22xp5_ASAP7_75t_L g7556 ( 
.A1(n_6986),
.A2(n_589),
.B1(n_590),
.B2(n_588),
.Y(n_7556)
);

AOI22xp5_ASAP7_75t_L g7557 ( 
.A1(n_7214),
.A2(n_590),
.B1(n_591),
.B2(n_589),
.Y(n_7557)
);

BUFx8_ASAP7_75t_L g7558 ( 
.A(n_6849),
.Y(n_7558)
);

AO22x2_ASAP7_75t_L g7559 ( 
.A1(n_7101),
.A2(n_27),
.B1(n_25),
.B2(n_26),
.Y(n_7559)
);

CKINVDCx5p33_ASAP7_75t_R g7560 ( 
.A(n_7291),
.Y(n_7560)
);

AND2x4_ASAP7_75t_L g7561 ( 
.A(n_7172),
.B(n_593),
.Y(n_7561)
);

INVx1_ASAP7_75t_L g7562 ( 
.A(n_7206),
.Y(n_7562)
);

INVx1_ASAP7_75t_L g7563 ( 
.A(n_7212),
.Y(n_7563)
);

INVx1_ASAP7_75t_L g7564 ( 
.A(n_7230),
.Y(n_7564)
);

AO22x2_ASAP7_75t_L g7565 ( 
.A1(n_6980),
.A2(n_27),
.B1(n_25),
.B2(n_26),
.Y(n_7565)
);

AND2x2_ASAP7_75t_L g7566 ( 
.A(n_7102),
.B(n_593),
.Y(n_7566)
);

AO22x2_ASAP7_75t_L g7567 ( 
.A1(n_7178),
.A2(n_28),
.B1(n_26),
.B2(n_27),
.Y(n_7567)
);

NAND2xp5_ASAP7_75t_L g7568 ( 
.A(n_6877),
.B(n_28),
.Y(n_7568)
);

HB1xp67_ASAP7_75t_L g7569 ( 
.A(n_7044),
.Y(n_7569)
);

INVxp67_ASAP7_75t_L g7570 ( 
.A(n_7098),
.Y(n_7570)
);

OAI22xp5_ASAP7_75t_L g7571 ( 
.A1(n_7262),
.A2(n_595),
.B1(n_596),
.B2(n_594),
.Y(n_7571)
);

INVx1_ASAP7_75t_L g7572 ( 
.A(n_6998),
.Y(n_7572)
);

INVx1_ASAP7_75t_L g7573 ( 
.A(n_7004),
.Y(n_7573)
);

INVx1_ASAP7_75t_L g7574 ( 
.A(n_7006),
.Y(n_7574)
);

NAND2xp5_ASAP7_75t_SL g7575 ( 
.A(n_6895),
.B(n_594),
.Y(n_7575)
);

INVx1_ASAP7_75t_L g7576 ( 
.A(n_7012),
.Y(n_7576)
);

AO22x2_ASAP7_75t_L g7577 ( 
.A1(n_6840),
.A2(n_30),
.B1(n_28),
.B2(n_29),
.Y(n_7577)
);

AND2x4_ASAP7_75t_L g7578 ( 
.A(n_7171),
.B(n_595),
.Y(n_7578)
);

INVx1_ASAP7_75t_L g7579 ( 
.A(n_7013),
.Y(n_7579)
);

CKINVDCx5p33_ASAP7_75t_R g7580 ( 
.A(n_7176),
.Y(n_7580)
);

INVx1_ASAP7_75t_L g7581 ( 
.A(n_7017),
.Y(n_7581)
);

BUFx8_ASAP7_75t_L g7582 ( 
.A(n_7061),
.Y(n_7582)
);

INVx1_ASAP7_75t_L g7583 ( 
.A(n_7018),
.Y(n_7583)
);

INVx1_ASAP7_75t_L g7584 ( 
.A(n_7020),
.Y(n_7584)
);

INVx1_ASAP7_75t_L g7585 ( 
.A(n_7022),
.Y(n_7585)
);

AND2x4_ASAP7_75t_L g7586 ( 
.A(n_7280),
.B(n_597),
.Y(n_7586)
);

AND2x4_ASAP7_75t_L g7587 ( 
.A(n_7250),
.B(n_597),
.Y(n_7587)
);

INVx2_ASAP7_75t_L g7588 ( 
.A(n_7235),
.Y(n_7588)
);

BUFx8_ASAP7_75t_L g7589 ( 
.A(n_7136),
.Y(n_7589)
);

OAI221xp5_ASAP7_75t_L g7590 ( 
.A1(n_7128),
.A2(n_31),
.B1(n_29),
.B2(n_30),
.C(n_32),
.Y(n_7590)
);

BUFx8_ASAP7_75t_L g7591 ( 
.A(n_7173),
.Y(n_7591)
);

BUFx8_ASAP7_75t_L g7592 ( 
.A(n_7025),
.Y(n_7592)
);

BUFx8_ASAP7_75t_L g7593 ( 
.A(n_7145),
.Y(n_7593)
);

OR2x2_ASAP7_75t_L g7594 ( 
.A(n_7111),
.B(n_7185),
.Y(n_7594)
);

INVx1_ASAP7_75t_L g7595 ( 
.A(n_7024),
.Y(n_7595)
);

AND2x4_ASAP7_75t_L g7596 ( 
.A(n_7295),
.B(n_598),
.Y(n_7596)
);

AND2x4_ASAP7_75t_L g7597 ( 
.A(n_7309),
.B(n_599),
.Y(n_7597)
);

BUFx2_ASAP7_75t_L g7598 ( 
.A(n_7223),
.Y(n_7598)
);

NAND2x1p5_ASAP7_75t_L g7599 ( 
.A(n_7245),
.B(n_599),
.Y(n_7599)
);

INVx1_ASAP7_75t_L g7600 ( 
.A(n_7237),
.Y(n_7600)
);

AO22x2_ASAP7_75t_L g7601 ( 
.A1(n_6839),
.A2(n_31),
.B1(n_29),
.B2(n_30),
.Y(n_7601)
);

AND2x4_ASAP7_75t_L g7602 ( 
.A(n_7267),
.B(n_600),
.Y(n_7602)
);

NAND2x1p5_ASAP7_75t_L g7603 ( 
.A(n_6818),
.B(n_600),
.Y(n_7603)
);

INVxp67_ASAP7_75t_L g7604 ( 
.A(n_7087),
.Y(n_7604)
);

AO22x2_ASAP7_75t_L g7605 ( 
.A1(n_6989),
.A2(n_7121),
.B1(n_6837),
.B2(n_6941),
.Y(n_7605)
);

AO22x2_ASAP7_75t_L g7606 ( 
.A1(n_6861),
.A2(n_34),
.B1(n_32),
.B2(n_33),
.Y(n_7606)
);

CKINVDCx5p33_ASAP7_75t_R g7607 ( 
.A(n_6846),
.Y(n_7607)
);

A2O1A1Ixp33_ASAP7_75t_L g7608 ( 
.A1(n_7142),
.A2(n_35),
.B(n_32),
.C(n_33),
.Y(n_7608)
);

AO22x2_ASAP7_75t_L g7609 ( 
.A1(n_6995),
.A2(n_36),
.B1(n_33),
.B2(n_35),
.Y(n_7609)
);

INVxp67_ASAP7_75t_L g7610 ( 
.A(n_7090),
.Y(n_7610)
);

BUFx8_ASAP7_75t_L g7611 ( 
.A(n_7187),
.Y(n_7611)
);

BUFx2_ASAP7_75t_L g7612 ( 
.A(n_7204),
.Y(n_7612)
);

NAND2xp5_ASAP7_75t_L g7613 ( 
.A(n_6968),
.B(n_35),
.Y(n_7613)
);

INVx3_ASAP7_75t_L g7614 ( 
.A(n_7279),
.Y(n_7614)
);

INVx1_ASAP7_75t_L g7615 ( 
.A(n_7072),
.Y(n_7615)
);

NOR2xp67_ASAP7_75t_L g7616 ( 
.A(n_7289),
.B(n_36),
.Y(n_7616)
);

AOI22xp5_ASAP7_75t_L g7617 ( 
.A1(n_7228),
.A2(n_602),
.B1(n_604),
.B2(n_601),
.Y(n_7617)
);

BUFx6f_ASAP7_75t_L g7618 ( 
.A(n_7285),
.Y(n_7618)
);

AO22x2_ASAP7_75t_L g7619 ( 
.A1(n_7016),
.A2(n_39),
.B1(n_37),
.B2(n_38),
.Y(n_7619)
);

INVxp67_ASAP7_75t_L g7620 ( 
.A(n_7259),
.Y(n_7620)
);

INVx1_ASAP7_75t_L g7621 ( 
.A(n_7073),
.Y(n_7621)
);

AO22x2_ASAP7_75t_L g7622 ( 
.A1(n_6929),
.A2(n_40),
.B1(n_37),
.B2(n_38),
.Y(n_7622)
);

INVx1_ASAP7_75t_L g7623 ( 
.A(n_7032),
.Y(n_7623)
);

OR2x6_ASAP7_75t_L g7624 ( 
.A(n_6927),
.B(n_601),
.Y(n_7624)
);

BUFx3_ASAP7_75t_L g7625 ( 
.A(n_7256),
.Y(n_7625)
);

INVx1_ASAP7_75t_L g7626 ( 
.A(n_7034),
.Y(n_7626)
);

INVx1_ASAP7_75t_L g7627 ( 
.A(n_7036),
.Y(n_7627)
);

AO22x2_ASAP7_75t_L g7628 ( 
.A1(n_7307),
.A2(n_40),
.B1(n_37),
.B2(n_38),
.Y(n_7628)
);

AO22x2_ASAP7_75t_L g7629 ( 
.A1(n_6981),
.A2(n_42),
.B1(n_40),
.B2(n_41),
.Y(n_7629)
);

AO22x2_ASAP7_75t_L g7630 ( 
.A1(n_7053),
.A2(n_7058),
.B1(n_6887),
.B2(n_7009),
.Y(n_7630)
);

BUFx2_ASAP7_75t_L g7631 ( 
.A(n_7290),
.Y(n_7631)
);

NAND2xp5_ASAP7_75t_L g7632 ( 
.A(n_6962),
.B(n_41),
.Y(n_7632)
);

INVxp67_ASAP7_75t_L g7633 ( 
.A(n_7281),
.Y(n_7633)
);

INVx1_ASAP7_75t_L g7634 ( 
.A(n_7045),
.Y(n_7634)
);

INVx1_ASAP7_75t_L g7635 ( 
.A(n_7047),
.Y(n_7635)
);

AO22x2_ASAP7_75t_L g7636 ( 
.A1(n_7243),
.A2(n_43),
.B1(n_41),
.B2(n_42),
.Y(n_7636)
);

OAI221xp5_ASAP7_75t_L g7637 ( 
.A1(n_7300),
.A2(n_44),
.B1(n_42),
.B2(n_43),
.C(n_45),
.Y(n_7637)
);

INVx1_ASAP7_75t_L g7638 ( 
.A(n_7051),
.Y(n_7638)
);

OAI221xp5_ASAP7_75t_L g7639 ( 
.A1(n_7192),
.A2(n_45),
.B1(n_43),
.B2(n_44),
.C(n_46),
.Y(n_7639)
);

AND2x4_ASAP7_75t_L g7640 ( 
.A(n_7269),
.B(n_602),
.Y(n_7640)
);

NAND2xp5_ASAP7_75t_L g7641 ( 
.A(n_7097),
.B(n_44),
.Y(n_7641)
);

INVx2_ASAP7_75t_L g7642 ( 
.A(n_6883),
.Y(n_7642)
);

INVx1_ASAP7_75t_L g7643 ( 
.A(n_7052),
.Y(n_7643)
);

INVxp67_ASAP7_75t_L g7644 ( 
.A(n_7282),
.Y(n_7644)
);

BUFx2_ASAP7_75t_L g7645 ( 
.A(n_7278),
.Y(n_7645)
);

AO22x2_ASAP7_75t_L g7646 ( 
.A1(n_7191),
.A2(n_47),
.B1(n_45),
.B2(n_46),
.Y(n_7646)
);

AO22x2_ASAP7_75t_L g7647 ( 
.A1(n_7198),
.A2(n_48),
.B1(n_46),
.B2(n_47),
.Y(n_7647)
);

AND2x4_ASAP7_75t_L g7648 ( 
.A(n_7284),
.B(n_605),
.Y(n_7648)
);

HB1xp67_ASAP7_75t_L g7649 ( 
.A(n_6992),
.Y(n_7649)
);

INVx1_ASAP7_75t_L g7650 ( 
.A(n_7055),
.Y(n_7650)
);

INVx2_ASAP7_75t_L g7651 ( 
.A(n_6883),
.Y(n_7651)
);

AND2x4_ASAP7_75t_L g7652 ( 
.A(n_7287),
.B(n_605),
.Y(n_7652)
);

INVx1_ASAP7_75t_SL g7653 ( 
.A(n_7303),
.Y(n_7653)
);

INVx1_ASAP7_75t_L g7654 ( 
.A(n_6942),
.Y(n_7654)
);

AND2x2_ASAP7_75t_L g7655 ( 
.A(n_6907),
.B(n_606),
.Y(n_7655)
);

CKINVDCx5p33_ASAP7_75t_R g7656 ( 
.A(n_6936),
.Y(n_7656)
);

AO22x2_ASAP7_75t_L g7657 ( 
.A1(n_7091),
.A2(n_49),
.B1(n_47),
.B2(n_48),
.Y(n_7657)
);

NAND2x1p5_ASAP7_75t_L g7658 ( 
.A(n_7296),
.B(n_606),
.Y(n_7658)
);

AND2x2_ASAP7_75t_SL g7659 ( 
.A(n_7271),
.B(n_607),
.Y(n_7659)
);

NAND2xp5_ASAP7_75t_L g7660 ( 
.A(n_7110),
.B(n_48),
.Y(n_7660)
);

INVx1_ASAP7_75t_L g7661 ( 
.A(n_6943),
.Y(n_7661)
);

AO22x2_ASAP7_75t_L g7662 ( 
.A1(n_7103),
.A2(n_51),
.B1(n_49),
.B2(n_50),
.Y(n_7662)
);

INVx1_ASAP7_75t_L g7663 ( 
.A(n_6946),
.Y(n_7663)
);

AOI22xp33_ASAP7_75t_L g7664 ( 
.A1(n_7160),
.A2(n_7130),
.B1(n_7217),
.B2(n_7105),
.Y(n_7664)
);

CKINVDCx20_ASAP7_75t_R g7665 ( 
.A(n_6982),
.Y(n_7665)
);

AND2x4_ASAP7_75t_L g7666 ( 
.A(n_7297),
.B(n_607),
.Y(n_7666)
);

INVx1_ASAP7_75t_L g7667 ( 
.A(n_6878),
.Y(n_7667)
);

INVx1_ASAP7_75t_L g7668 ( 
.A(n_6881),
.Y(n_7668)
);

INVx1_ASAP7_75t_L g7669 ( 
.A(n_6884),
.Y(n_7669)
);

AO22x2_ASAP7_75t_L g7670 ( 
.A1(n_7156),
.A2(n_51),
.B1(n_49),
.B2(n_50),
.Y(n_7670)
);

INVx2_ASAP7_75t_L g7671 ( 
.A(n_6883),
.Y(n_7671)
);

INVx1_ASAP7_75t_L g7672 ( 
.A(n_6886),
.Y(n_7672)
);

AND2x2_ASAP7_75t_L g7673 ( 
.A(n_7272),
.B(n_608),
.Y(n_7673)
);

INVx1_ASAP7_75t_L g7674 ( 
.A(n_6891),
.Y(n_7674)
);

INVx2_ASAP7_75t_L g7675 ( 
.A(n_6883),
.Y(n_7675)
);

NOR2xp67_ASAP7_75t_L g7676 ( 
.A(n_7310),
.B(n_50),
.Y(n_7676)
);

INVxp67_ASAP7_75t_L g7677 ( 
.A(n_7286),
.Y(n_7677)
);

AND2x4_ASAP7_75t_L g7678 ( 
.A(n_7084),
.B(n_609),
.Y(n_7678)
);

NAND2xp5_ASAP7_75t_L g7679 ( 
.A(n_7116),
.B(n_51),
.Y(n_7679)
);

AO22x2_ASAP7_75t_L g7680 ( 
.A1(n_7180),
.A2(n_54),
.B1(n_52),
.B2(n_53),
.Y(n_7680)
);

INVxp67_ASAP7_75t_L g7681 ( 
.A(n_7115),
.Y(n_7681)
);

INVx1_ASAP7_75t_L g7682 ( 
.A(n_6893),
.Y(n_7682)
);

OAI221xp5_ASAP7_75t_L g7683 ( 
.A1(n_7193),
.A2(n_54),
.B1(n_52),
.B2(n_53),
.C(n_55),
.Y(n_7683)
);

INVx1_ASAP7_75t_L g7684 ( 
.A(n_6896),
.Y(n_7684)
);

AO22x2_ASAP7_75t_L g7685 ( 
.A1(n_7152),
.A2(n_54),
.B1(n_52),
.B2(n_53),
.Y(n_7685)
);

INVx2_ASAP7_75t_L g7686 ( 
.A(n_6923),
.Y(n_7686)
);

INVx2_ASAP7_75t_L g7687 ( 
.A(n_6923),
.Y(n_7687)
);

BUFx2_ASAP7_75t_L g7688 ( 
.A(n_7194),
.Y(n_7688)
);

INVx1_ASAP7_75t_L g7689 ( 
.A(n_6899),
.Y(n_7689)
);

INVx1_ASAP7_75t_SL g7690 ( 
.A(n_7288),
.Y(n_7690)
);

INVx2_ASAP7_75t_SL g7691 ( 
.A(n_7283),
.Y(n_7691)
);

OAI221xp5_ASAP7_75t_L g7692 ( 
.A1(n_6957),
.A2(n_58),
.B1(n_56),
.B2(n_57),
.C(n_59),
.Y(n_7692)
);

NAND2xp5_ASAP7_75t_L g7693 ( 
.A(n_7118),
.B(n_56),
.Y(n_7693)
);

NAND2xp5_ASAP7_75t_L g7694 ( 
.A(n_7119),
.B(n_56),
.Y(n_7694)
);

INVx1_ASAP7_75t_L g7695 ( 
.A(n_6900),
.Y(n_7695)
);

AO22x2_ASAP7_75t_L g7696 ( 
.A1(n_6970),
.A2(n_60),
.B1(n_57),
.B2(n_59),
.Y(n_7696)
);

NAND2xp33_ASAP7_75t_L g7697 ( 
.A(n_6923),
.B(n_57),
.Y(n_7697)
);

OAI221xp5_ASAP7_75t_L g7698 ( 
.A1(n_6977),
.A2(n_61),
.B1(n_59),
.B2(n_60),
.C(n_62),
.Y(n_7698)
);

NAND2x1p5_ASAP7_75t_L g7699 ( 
.A(n_7226),
.B(n_7174),
.Y(n_7699)
);

NAND2xp5_ASAP7_75t_L g7700 ( 
.A(n_7125),
.B(n_60),
.Y(n_7700)
);

NAND2xp5_ASAP7_75t_L g7701 ( 
.A(n_7126),
.B(n_61),
.Y(n_7701)
);

AND2x4_ASAP7_75t_L g7702 ( 
.A(n_7199),
.B(n_609),
.Y(n_7702)
);

INVx1_ASAP7_75t_L g7703 ( 
.A(n_6903),
.Y(n_7703)
);

INVxp67_ASAP7_75t_L g7704 ( 
.A(n_7260),
.Y(n_7704)
);

INVx1_ASAP7_75t_L g7705 ( 
.A(n_6908),
.Y(n_7705)
);

NOR2xp33_ASAP7_75t_L g7706 ( 
.A(n_7175),
.B(n_7146),
.Y(n_7706)
);

NAND2xp5_ASAP7_75t_L g7707 ( 
.A(n_7127),
.B(n_63),
.Y(n_7707)
);

NAND2x1p5_ASAP7_75t_L g7708 ( 
.A(n_7177),
.B(n_610),
.Y(n_7708)
);

NAND2x1p5_ASAP7_75t_L g7709 ( 
.A(n_7094),
.B(n_611),
.Y(n_7709)
);

NAND2xp5_ASAP7_75t_L g7710 ( 
.A(n_7131),
.B(n_63),
.Y(n_7710)
);

BUFx8_ASAP7_75t_L g7711 ( 
.A(n_7218),
.Y(n_7711)
);

INVx1_ASAP7_75t_L g7712 ( 
.A(n_6910),
.Y(n_7712)
);

OAI221xp5_ASAP7_75t_L g7713 ( 
.A1(n_6967),
.A2(n_65),
.B1(n_63),
.B2(n_64),
.C(n_66),
.Y(n_7713)
);

INVx1_ASAP7_75t_L g7714 ( 
.A(n_6914),
.Y(n_7714)
);

INVx1_ASAP7_75t_L g7715 ( 
.A(n_6918),
.Y(n_7715)
);

INVx1_ASAP7_75t_L g7716 ( 
.A(n_6919),
.Y(n_7716)
);

INVx1_ASAP7_75t_L g7717 ( 
.A(n_6928),
.Y(n_7717)
);

AO22x2_ASAP7_75t_L g7718 ( 
.A1(n_7201),
.A2(n_66),
.B1(n_64),
.B2(n_65),
.Y(n_7718)
);

INVx1_ASAP7_75t_L g7719 ( 
.A(n_6930),
.Y(n_7719)
);

INVx1_ASAP7_75t_L g7720 ( 
.A(n_6935),
.Y(n_7720)
);

AND2x6_ASAP7_75t_L g7721 ( 
.A(n_7203),
.B(n_7205),
.Y(n_7721)
);

AOI22xp5_ASAP7_75t_L g7722 ( 
.A1(n_7008),
.A2(n_612),
.B1(n_613),
.B2(n_611),
.Y(n_7722)
);

INVx1_ASAP7_75t_L g7723 ( 
.A(n_6937),
.Y(n_7723)
);

NAND2x1p5_ASAP7_75t_L g7724 ( 
.A(n_7095),
.B(n_612),
.Y(n_7724)
);

INVx1_ASAP7_75t_L g7725 ( 
.A(n_6862),
.Y(n_7725)
);

INVxp67_ASAP7_75t_L g7726 ( 
.A(n_7015),
.Y(n_7726)
);

AO22x2_ASAP7_75t_L g7727 ( 
.A1(n_7071),
.A2(n_67),
.B1(n_64),
.B2(n_66),
.Y(n_7727)
);

INVx1_ASAP7_75t_L g7728 ( 
.A(n_6969),
.Y(n_7728)
);

NAND2xp5_ASAP7_75t_L g7729 ( 
.A(n_7224),
.B(n_7150),
.Y(n_7729)
);

INVx1_ASAP7_75t_L g7730 ( 
.A(n_6966),
.Y(n_7730)
);

INVx1_ASAP7_75t_L g7731 ( 
.A(n_7232),
.Y(n_7731)
);

AND2x2_ASAP7_75t_L g7732 ( 
.A(n_6827),
.B(n_613),
.Y(n_7732)
);

INVxp67_ASAP7_75t_L g7733 ( 
.A(n_6870),
.Y(n_7733)
);

AO22x2_ASAP7_75t_L g7734 ( 
.A1(n_7244),
.A2(n_69),
.B1(n_67),
.B2(n_68),
.Y(n_7734)
);

AO22x2_ASAP7_75t_L g7735 ( 
.A1(n_6996),
.A2(n_72),
.B1(n_69),
.B2(n_71),
.Y(n_7735)
);

OR2x2_ASAP7_75t_SL g7736 ( 
.A(n_7268),
.B(n_71),
.Y(n_7736)
);

INVx2_ASAP7_75t_L g7737 ( 
.A(n_6923),
.Y(n_7737)
);

HB1xp67_ASAP7_75t_L g7738 ( 
.A(n_7273),
.Y(n_7738)
);

INVx1_ASAP7_75t_L g7739 ( 
.A(n_7109),
.Y(n_7739)
);

INVx1_ASAP7_75t_L g7740 ( 
.A(n_7109),
.Y(n_7740)
);

CKINVDCx5p33_ASAP7_75t_R g7741 ( 
.A(n_6936),
.Y(n_7741)
);

AND2x2_ASAP7_75t_L g7742 ( 
.A(n_7001),
.B(n_614),
.Y(n_7742)
);

INVx2_ASAP7_75t_L g7743 ( 
.A(n_6949),
.Y(n_7743)
);

NAND2xp5_ASAP7_75t_L g7744 ( 
.A(n_7155),
.B(n_71),
.Y(n_7744)
);

OR2x2_ASAP7_75t_L g7745 ( 
.A(n_7158),
.B(n_72),
.Y(n_7745)
);

AND2x4_ASAP7_75t_L g7746 ( 
.A(n_6931),
.B(n_614),
.Y(n_7746)
);

INVx2_ASAP7_75t_L g7747 ( 
.A(n_6949),
.Y(n_7747)
);

NAND2xp5_ASAP7_75t_SL g7748 ( 
.A(n_7132),
.B(n_615),
.Y(n_7748)
);

INVx1_ASAP7_75t_L g7749 ( 
.A(n_7109),
.Y(n_7749)
);

OR2x6_ASAP7_75t_SL g7750 ( 
.A(n_7276),
.B(n_7209),
.Y(n_7750)
);

AND2x4_ASAP7_75t_L g7751 ( 
.A(n_7069),
.B(n_615),
.Y(n_7751)
);

NAND2xp5_ASAP7_75t_L g7752 ( 
.A(n_7163),
.B(n_72),
.Y(n_7752)
);

BUFx8_ASAP7_75t_L g7753 ( 
.A(n_6974),
.Y(n_7753)
);

INVx1_ASAP7_75t_L g7754 ( 
.A(n_7079),
.Y(n_7754)
);

INVx1_ASAP7_75t_L g7755 ( 
.A(n_7086),
.Y(n_7755)
);

INVx2_ASAP7_75t_L g7756 ( 
.A(n_6949),
.Y(n_7756)
);

NAND2xp5_ASAP7_75t_L g7757 ( 
.A(n_7148),
.B(n_73),
.Y(n_7757)
);

INVx1_ASAP7_75t_L g7758 ( 
.A(n_7089),
.Y(n_7758)
);

INVx1_ASAP7_75t_L g7759 ( 
.A(n_7213),
.Y(n_7759)
);

INVx1_ASAP7_75t_L g7760 ( 
.A(n_6974),
.Y(n_7760)
);

INVx1_ASAP7_75t_L g7761 ( 
.A(n_6974),
.Y(n_7761)
);

BUFx6f_ASAP7_75t_L g7762 ( 
.A(n_6944),
.Y(n_7762)
);

OR2x2_ASAP7_75t_SL g7763 ( 
.A(n_7293),
.B(n_73),
.Y(n_7763)
);

INVx1_ASAP7_75t_L g7764 ( 
.A(n_7144),
.Y(n_7764)
);

BUFx3_ASAP7_75t_L g7765 ( 
.A(n_6944),
.Y(n_7765)
);

INVx1_ASAP7_75t_L g7766 ( 
.A(n_7225),
.Y(n_7766)
);

INVxp67_ASAP7_75t_L g7767 ( 
.A(n_7308),
.Y(n_7767)
);

AOI22xp5_ASAP7_75t_L g7768 ( 
.A1(n_6993),
.A2(n_617),
.B1(n_618),
.B2(n_616),
.Y(n_7768)
);

AO22x2_ASAP7_75t_L g7769 ( 
.A1(n_7088),
.A2(n_75),
.B1(n_73),
.B2(n_74),
.Y(n_7769)
);

INVx1_ASAP7_75t_L g7770 ( 
.A(n_7248),
.Y(n_7770)
);

NAND2xp5_ASAP7_75t_L g7771 ( 
.A(n_7255),
.B(n_74),
.Y(n_7771)
);

INVx1_ASAP7_75t_L g7772 ( 
.A(n_7263),
.Y(n_7772)
);

AO22x2_ASAP7_75t_L g7773 ( 
.A1(n_7027),
.A2(n_77),
.B1(n_75),
.B2(n_76),
.Y(n_7773)
);

INVx3_ASAP7_75t_L g7774 ( 
.A(n_6953),
.Y(n_7774)
);

NAND2xp5_ASAP7_75t_L g7775 ( 
.A(n_7264),
.B(n_75),
.Y(n_7775)
);

INVx1_ASAP7_75t_L g7776 ( 
.A(n_7277),
.Y(n_7776)
);

HB1xp67_ASAP7_75t_L g7777 ( 
.A(n_6953),
.Y(n_7777)
);

OAI221xp5_ASAP7_75t_L g7778 ( 
.A1(n_7249),
.A2(n_78),
.B1(n_76),
.B2(n_77),
.C(n_79),
.Y(n_7778)
);

AO22x2_ASAP7_75t_L g7779 ( 
.A1(n_7043),
.A2(n_6991),
.B1(n_7299),
.B2(n_7294),
.Y(n_7779)
);

AND2x4_ASAP7_75t_L g7780 ( 
.A(n_7236),
.B(n_616),
.Y(n_7780)
);

INVxp67_ASAP7_75t_L g7781 ( 
.A(n_7067),
.Y(n_7781)
);

INVx1_ASAP7_75t_L g7782 ( 
.A(n_7305),
.Y(n_7782)
);

OR2x2_ASAP7_75t_SL g7783 ( 
.A(n_6853),
.B(n_77),
.Y(n_7783)
);

INVx2_ASAP7_75t_L g7784 ( 
.A(n_6949),
.Y(n_7784)
);

NAND2x1p5_ASAP7_75t_L g7785 ( 
.A(n_6889),
.B(n_7189),
.Y(n_7785)
);

INVx2_ASAP7_75t_L g7786 ( 
.A(n_6945),
.Y(n_7786)
);

INVx2_ASAP7_75t_L g7787 ( 
.A(n_7122),
.Y(n_7787)
);

NAND2xp5_ASAP7_75t_L g7788 ( 
.A(n_6820),
.B(n_78),
.Y(n_7788)
);

NAND2xp5_ASAP7_75t_L g7789 ( 
.A(n_7135),
.B(n_78),
.Y(n_7789)
);

AO22x2_ASAP7_75t_L g7790 ( 
.A1(n_7247),
.A2(n_81),
.B1(n_79),
.B2(n_80),
.Y(n_7790)
);

BUFx3_ASAP7_75t_L g7791 ( 
.A(n_7266),
.Y(n_7791)
);

INVx1_ASAP7_75t_L g7792 ( 
.A(n_7238),
.Y(n_7792)
);

INVx1_ASAP7_75t_L g7793 ( 
.A(n_7003),
.Y(n_7793)
);

AO22x2_ASAP7_75t_L g7794 ( 
.A1(n_7254),
.A2(n_82),
.B1(n_79),
.B2(n_80),
.Y(n_7794)
);

INVx1_ASAP7_75t_L g7795 ( 
.A(n_7074),
.Y(n_7795)
);

AO22x2_ASAP7_75t_L g7796 ( 
.A1(n_7257),
.A2(n_84),
.B1(n_82),
.B2(n_83),
.Y(n_7796)
);

A2O1A1Ixp33_ASAP7_75t_L g7797 ( 
.A1(n_7219),
.A2(n_85),
.B(n_83),
.C(n_84),
.Y(n_7797)
);

CKINVDCx20_ASAP7_75t_R g7798 ( 
.A(n_7157),
.Y(n_7798)
);

NAND2xp5_ASAP7_75t_L g7799 ( 
.A(n_7023),
.B(n_83),
.Y(n_7799)
);

NAND2xp5_ASAP7_75t_L g7800 ( 
.A(n_7014),
.B(n_84),
.Y(n_7800)
);

INVx4_ASAP7_75t_L g7801 ( 
.A(n_7266),
.Y(n_7801)
);

NAND2xp5_ASAP7_75t_L g7802 ( 
.A(n_7197),
.B(n_85),
.Y(n_7802)
);

OAI221xp5_ASAP7_75t_L g7803 ( 
.A1(n_7054),
.A2(n_87),
.B1(n_85),
.B2(n_86),
.C(n_88),
.Y(n_7803)
);

INVxp67_ASAP7_75t_L g7804 ( 
.A(n_7234),
.Y(n_7804)
);

NAND2x1p5_ASAP7_75t_L g7805 ( 
.A(n_7304),
.B(n_617),
.Y(n_7805)
);

AOI22xp5_ASAP7_75t_L g7806 ( 
.A1(n_7134),
.A2(n_619),
.B1(n_620),
.B2(n_618),
.Y(n_7806)
);

INVx1_ASAP7_75t_L g7807 ( 
.A(n_7042),
.Y(n_7807)
);

INVx2_ASAP7_75t_L g7808 ( 
.A(n_7164),
.Y(n_7808)
);

O2A1O1Ixp5_ASAP7_75t_L g7809 ( 
.A1(n_7446),
.A2(n_7261),
.B(n_7141),
.C(n_7275),
.Y(n_7809)
);

OAI22xp5_ASAP7_75t_L g7810 ( 
.A1(n_7464),
.A2(n_7186),
.B1(n_7298),
.B2(n_7104),
.Y(n_7810)
);

OAI21xp5_ASAP7_75t_L g7811 ( 
.A1(n_7458),
.A2(n_7265),
.B(n_7298),
.Y(n_7811)
);

NAND2xp5_ASAP7_75t_L g7812 ( 
.A(n_7349),
.B(n_86),
.Y(n_7812)
);

INVx2_ASAP7_75t_L g7813 ( 
.A(n_7320),
.Y(n_7813)
);

BUFx6f_ASAP7_75t_L g7814 ( 
.A(n_7312),
.Y(n_7814)
);

AND2x4_ASAP7_75t_L g7815 ( 
.A(n_7329),
.B(n_619),
.Y(n_7815)
);

NOR2xp33_ASAP7_75t_L g7816 ( 
.A(n_7726),
.B(n_620),
.Y(n_7816)
);

BUFx6f_ASAP7_75t_L g7817 ( 
.A(n_7518),
.Y(n_7817)
);

AND2x2_ASAP7_75t_L g7818 ( 
.A(n_7551),
.B(n_86),
.Y(n_7818)
);

NAND2xp5_ASAP7_75t_SL g7819 ( 
.A(n_7607),
.B(n_621),
.Y(n_7819)
);

AOI21xp5_ASAP7_75t_L g7820 ( 
.A1(n_7729),
.A2(n_622),
.B(n_621),
.Y(n_7820)
);

AND2x2_ASAP7_75t_L g7821 ( 
.A(n_7414),
.B(n_87),
.Y(n_7821)
);

AOI21xp5_ASAP7_75t_L g7822 ( 
.A1(n_7455),
.A2(n_623),
.B(n_622),
.Y(n_7822)
);

NAND2xp5_ASAP7_75t_L g7823 ( 
.A(n_7351),
.B(n_87),
.Y(n_7823)
);

AOI21xp5_ASAP7_75t_L g7824 ( 
.A1(n_7697),
.A2(n_626),
.B(n_624),
.Y(n_7824)
);

AOI21xp5_ASAP7_75t_L g7825 ( 
.A1(n_7706),
.A2(n_626),
.B(n_624),
.Y(n_7825)
);

NAND2xp5_ASAP7_75t_L g7826 ( 
.A(n_7353),
.B(n_88),
.Y(n_7826)
);

NAND2xp5_ASAP7_75t_L g7827 ( 
.A(n_7357),
.B(n_88),
.Y(n_7827)
);

OAI21xp5_ASAP7_75t_L g7828 ( 
.A1(n_7454),
.A2(n_89),
.B(n_90),
.Y(n_7828)
);

NOR2xp33_ASAP7_75t_SL g7829 ( 
.A(n_7344),
.B(n_89),
.Y(n_7829)
);

OAI21xp5_ASAP7_75t_L g7830 ( 
.A1(n_7440),
.A2(n_90),
.B(n_91),
.Y(n_7830)
);

O2A1O1Ixp33_ASAP7_75t_L g7831 ( 
.A1(n_7807),
.A2(n_92),
.B(n_90),
.C(n_91),
.Y(n_7831)
);

NAND2xp5_ASAP7_75t_L g7832 ( 
.A(n_7388),
.B(n_92),
.Y(n_7832)
);

NAND3xp33_ASAP7_75t_SL g7833 ( 
.A(n_7471),
.B(n_92),
.C(n_93),
.Y(n_7833)
);

OAI21x1_ASAP7_75t_L g7834 ( 
.A1(n_7642),
.A2(n_93),
.B(n_94),
.Y(n_7834)
);

INVx1_ASAP7_75t_L g7835 ( 
.A(n_7322),
.Y(n_7835)
);

NAND2xp5_ASAP7_75t_SL g7836 ( 
.A(n_7604),
.B(n_627),
.Y(n_7836)
);

AOI21xp5_ASAP7_75t_L g7837 ( 
.A1(n_7433),
.A2(n_629),
.B(n_628),
.Y(n_7837)
);

AOI21xp5_ASAP7_75t_L g7838 ( 
.A1(n_7360),
.A2(n_631),
.B(n_630),
.Y(n_7838)
);

NOR2xp33_ASAP7_75t_L g7839 ( 
.A(n_7620),
.B(n_630),
.Y(n_7839)
);

INVx1_ASAP7_75t_L g7840 ( 
.A(n_7328),
.Y(n_7840)
);

INVx1_ASAP7_75t_L g7841 ( 
.A(n_7339),
.Y(n_7841)
);

AOI21xp5_ASAP7_75t_L g7842 ( 
.A1(n_7764),
.A2(n_633),
.B(n_632),
.Y(n_7842)
);

AOI22x1_ASAP7_75t_L g7843 ( 
.A1(n_7400),
.A2(n_95),
.B1(n_93),
.B2(n_94),
.Y(n_7843)
);

AOI22xp33_ASAP7_75t_L g7844 ( 
.A1(n_7539),
.A2(n_97),
.B1(n_95),
.B2(n_96),
.Y(n_7844)
);

AOI21xp5_ASAP7_75t_L g7845 ( 
.A1(n_7728),
.A2(n_633),
.B(n_632),
.Y(n_7845)
);

NOR2xp33_ASAP7_75t_L g7846 ( 
.A(n_7633),
.B(n_634),
.Y(n_7846)
);

NAND2xp5_ASAP7_75t_L g7847 ( 
.A(n_7730),
.B(n_96),
.Y(n_7847)
);

AOI21xp5_ASAP7_75t_L g7848 ( 
.A1(n_7381),
.A2(n_635),
.B(n_634),
.Y(n_7848)
);

BUFx3_ASAP7_75t_L g7849 ( 
.A(n_7313),
.Y(n_7849)
);

INVx1_ASAP7_75t_L g7850 ( 
.A(n_7348),
.Y(n_7850)
);

BUFx6f_ASAP7_75t_L g7851 ( 
.A(n_7518),
.Y(n_7851)
);

NAND2xp5_ASAP7_75t_SL g7852 ( 
.A(n_7610),
.B(n_635),
.Y(n_7852)
);

OAI21xp5_ASAP7_75t_L g7853 ( 
.A1(n_7447),
.A2(n_96),
.B(n_97),
.Y(n_7853)
);

AOI21xp5_ASAP7_75t_L g7854 ( 
.A1(n_7759),
.A2(n_7626),
.B(n_7623),
.Y(n_7854)
);

NAND2xp5_ASAP7_75t_L g7855 ( 
.A(n_7667),
.B(n_98),
.Y(n_7855)
);

INVx2_ASAP7_75t_L g7856 ( 
.A(n_7368),
.Y(n_7856)
);

BUFx2_ASAP7_75t_SL g7857 ( 
.A(n_7326),
.Y(n_7857)
);

NAND2xp5_ASAP7_75t_L g7858 ( 
.A(n_7668),
.B(n_98),
.Y(n_7858)
);

AOI21xp5_ASAP7_75t_L g7859 ( 
.A1(n_7627),
.A2(n_637),
.B(n_636),
.Y(n_7859)
);

INVx2_ASAP7_75t_L g7860 ( 
.A(n_7377),
.Y(n_7860)
);

AOI21xp5_ASAP7_75t_L g7861 ( 
.A1(n_7634),
.A2(n_640),
.B(n_639),
.Y(n_7861)
);

NOR2xp67_ASAP7_75t_L g7862 ( 
.A(n_7346),
.B(n_98),
.Y(n_7862)
);

NOR2xp33_ASAP7_75t_L g7863 ( 
.A(n_7644),
.B(n_7330),
.Y(n_7863)
);

INVx5_ASAP7_75t_L g7864 ( 
.A(n_7479),
.Y(n_7864)
);

AOI21xp5_ASAP7_75t_L g7865 ( 
.A1(n_7635),
.A2(n_641),
.B(n_639),
.Y(n_7865)
);

AOI21xp5_ASAP7_75t_L g7866 ( 
.A1(n_7638),
.A2(n_7650),
.B(n_7643),
.Y(n_7866)
);

OAI21xp5_ASAP7_75t_L g7867 ( 
.A1(n_7461),
.A2(n_99),
.B(n_100),
.Y(n_7867)
);

INVx2_ASAP7_75t_L g7868 ( 
.A(n_7404),
.Y(n_7868)
);

OAI21xp5_ASAP7_75t_L g7869 ( 
.A1(n_7466),
.A2(n_7484),
.B(n_7669),
.Y(n_7869)
);

NAND2xp5_ASAP7_75t_L g7870 ( 
.A(n_7672),
.B(n_99),
.Y(n_7870)
);

INVx1_ASAP7_75t_L g7871 ( 
.A(n_7315),
.Y(n_7871)
);

HB1xp67_ASAP7_75t_L g7872 ( 
.A(n_7493),
.Y(n_7872)
);

NOR2xp33_ASAP7_75t_L g7873 ( 
.A(n_7560),
.B(n_642),
.Y(n_7873)
);

NOR2xp33_ASAP7_75t_L g7874 ( 
.A(n_7690),
.B(n_642),
.Y(n_7874)
);

INVxp67_ASAP7_75t_L g7875 ( 
.A(n_7325),
.Y(n_7875)
);

OAI22xp5_ASAP7_75t_L g7876 ( 
.A1(n_7327),
.A2(n_101),
.B1(n_99),
.B2(n_100),
.Y(n_7876)
);

AND2x2_ASAP7_75t_L g7877 ( 
.A(n_7673),
.B(n_7543),
.Y(n_7877)
);

NAND2xp5_ASAP7_75t_L g7878 ( 
.A(n_7674),
.B(n_100),
.Y(n_7878)
);

NOR2x1_ASAP7_75t_L g7879 ( 
.A(n_7345),
.B(n_643),
.Y(n_7879)
);

NAND2xp5_ASAP7_75t_L g7880 ( 
.A(n_7682),
.B(n_101),
.Y(n_7880)
);

NAND2xp33_ASAP7_75t_L g7881 ( 
.A(n_7664),
.B(n_101),
.Y(n_7881)
);

HB1xp67_ASAP7_75t_L g7882 ( 
.A(n_7553),
.Y(n_7882)
);

INVx11_ASAP7_75t_L g7883 ( 
.A(n_7332),
.Y(n_7883)
);

AOI21xp5_ASAP7_75t_L g7884 ( 
.A1(n_7572),
.A2(n_645),
.B(n_644),
.Y(n_7884)
);

OAI22xp5_ASAP7_75t_L g7885 ( 
.A1(n_7314),
.A2(n_104),
.B1(n_102),
.B2(n_103),
.Y(n_7885)
);

OAI22xp5_ASAP7_75t_L g7886 ( 
.A1(n_7677),
.A2(n_7394),
.B1(n_7441),
.B2(n_7442),
.Y(n_7886)
);

AOI21xp5_ASAP7_75t_L g7887 ( 
.A1(n_7573),
.A2(n_645),
.B(n_644),
.Y(n_7887)
);

INVx2_ASAP7_75t_SL g7888 ( 
.A(n_7369),
.Y(n_7888)
);

NAND2xp5_ASAP7_75t_L g7889 ( 
.A(n_7684),
.B(n_102),
.Y(n_7889)
);

O2A1O1Ixp33_ASAP7_75t_L g7890 ( 
.A1(n_7490),
.A2(n_105),
.B(n_103),
.C(n_104),
.Y(n_7890)
);

NAND2xp5_ASAP7_75t_L g7891 ( 
.A(n_7689),
.B(n_103),
.Y(n_7891)
);

NAND2xp5_ASAP7_75t_L g7892 ( 
.A(n_7695),
.B(n_104),
.Y(n_7892)
);

NOR2x1_ASAP7_75t_L g7893 ( 
.A(n_7384),
.B(n_646),
.Y(n_7893)
);

NOR2xp33_ASAP7_75t_L g7894 ( 
.A(n_7703),
.B(n_647),
.Y(n_7894)
);

AOI21xp5_ASAP7_75t_L g7895 ( 
.A1(n_7574),
.A2(n_649),
.B(n_648),
.Y(n_7895)
);

AOI21xp5_ASAP7_75t_L g7896 ( 
.A1(n_7576),
.A2(n_649),
.B(n_648),
.Y(n_7896)
);

AOI21xp5_ASAP7_75t_L g7897 ( 
.A1(n_7579),
.A2(n_7583),
.B(n_7581),
.Y(n_7897)
);

AOI21xp5_ASAP7_75t_L g7898 ( 
.A1(n_7584),
.A2(n_7595),
.B(n_7585),
.Y(n_7898)
);

OAI21xp5_ASAP7_75t_L g7899 ( 
.A1(n_7705),
.A2(n_105),
.B(n_106),
.Y(n_7899)
);

AOI21xp5_ASAP7_75t_L g7900 ( 
.A1(n_7654),
.A2(n_651),
.B(n_650),
.Y(n_7900)
);

NOR2xp33_ASAP7_75t_L g7901 ( 
.A(n_7712),
.B(n_650),
.Y(n_7901)
);

AOI21xp5_ASAP7_75t_L g7902 ( 
.A1(n_7661),
.A2(n_7663),
.B(n_7621),
.Y(n_7902)
);

AOI21xp5_ASAP7_75t_L g7903 ( 
.A1(n_7615),
.A2(n_654),
.B(n_652),
.Y(n_7903)
);

AOI21xp5_ASAP7_75t_L g7904 ( 
.A1(n_7714),
.A2(n_654),
.B(n_652),
.Y(n_7904)
);

AOI21xp5_ASAP7_75t_L g7905 ( 
.A1(n_7715),
.A2(n_656),
.B(n_655),
.Y(n_7905)
);

INVxp67_ASAP7_75t_L g7906 ( 
.A(n_7399),
.Y(n_7906)
);

NAND2xp5_ASAP7_75t_L g7907 ( 
.A(n_7716),
.B(n_7717),
.Y(n_7907)
);

NAND2xp5_ASAP7_75t_SL g7908 ( 
.A(n_7364),
.B(n_655),
.Y(n_7908)
);

AND2x4_ASAP7_75t_L g7909 ( 
.A(n_7397),
.B(n_657),
.Y(n_7909)
);

NOR2xp33_ASAP7_75t_L g7910 ( 
.A(n_7719),
.B(n_657),
.Y(n_7910)
);

AOI21xp5_ASAP7_75t_L g7911 ( 
.A1(n_7720),
.A2(n_659),
.B(n_658),
.Y(n_7911)
);

INVx3_ASAP7_75t_L g7912 ( 
.A(n_7331),
.Y(n_7912)
);

AO32x2_ASAP7_75t_L g7913 ( 
.A1(n_7529),
.A2(n_107),
.A3(n_105),
.B1(n_106),
.B2(n_108),
.Y(n_7913)
);

AOI22xp5_ASAP7_75t_L g7914 ( 
.A1(n_7798),
.A2(n_109),
.B1(n_107),
.B2(n_108),
.Y(n_7914)
);

INVx3_ASAP7_75t_L g7915 ( 
.A(n_7403),
.Y(n_7915)
);

OAI22xp5_ASAP7_75t_L g7916 ( 
.A1(n_7541),
.A2(n_7570),
.B1(n_7767),
.B2(n_7361),
.Y(n_7916)
);

NAND2xp5_ASAP7_75t_L g7917 ( 
.A(n_7723),
.B(n_107),
.Y(n_7917)
);

AOI21xp5_ASAP7_75t_L g7918 ( 
.A1(n_7754),
.A2(n_659),
.B(n_658),
.Y(n_7918)
);

NAND2xp5_ASAP7_75t_L g7919 ( 
.A(n_7792),
.B(n_109),
.Y(n_7919)
);

NAND2xp5_ASAP7_75t_L g7920 ( 
.A(n_7352),
.B(n_110),
.Y(n_7920)
);

CKINVDCx10_ASAP7_75t_R g7921 ( 
.A(n_7517),
.Y(n_7921)
);

HB1xp67_ASAP7_75t_L g7922 ( 
.A(n_7470),
.Y(n_7922)
);

AOI21xp5_ASAP7_75t_L g7923 ( 
.A1(n_7755),
.A2(n_662),
.B(n_661),
.Y(n_7923)
);

NOR2xp33_ASAP7_75t_L g7924 ( 
.A(n_7580),
.B(n_662),
.Y(n_7924)
);

AOI21xp5_ASAP7_75t_L g7925 ( 
.A1(n_7758),
.A2(n_664),
.B(n_663),
.Y(n_7925)
);

NAND2xp5_ASAP7_75t_L g7926 ( 
.A(n_7770),
.B(n_110),
.Y(n_7926)
);

NAND2xp5_ASAP7_75t_L g7927 ( 
.A(n_7772),
.B(n_110),
.Y(n_7927)
);

AND2x6_ASAP7_75t_L g7928 ( 
.A(n_7651),
.B(n_111),
.Y(n_7928)
);

INVx1_ASAP7_75t_L g7929 ( 
.A(n_7317),
.Y(n_7929)
);

NAND2xp5_ASAP7_75t_L g7930 ( 
.A(n_7776),
.B(n_7782),
.Y(n_7930)
);

AOI21xp5_ASAP7_75t_L g7931 ( 
.A1(n_7795),
.A2(n_665),
.B(n_664),
.Y(n_7931)
);

AOI21xp5_ASAP7_75t_L g7932 ( 
.A1(n_7779),
.A2(n_666),
.B(n_665),
.Y(n_7932)
);

INVx2_ASAP7_75t_L g7933 ( 
.A(n_7421),
.Y(n_7933)
);

OAI22xp5_ASAP7_75t_L g7934 ( 
.A1(n_7336),
.A2(n_113),
.B1(n_111),
.B2(n_112),
.Y(n_7934)
);

AOI21xp5_ASAP7_75t_L g7935 ( 
.A1(n_7731),
.A2(n_668),
.B(n_667),
.Y(n_7935)
);

O2A1O1Ixp33_ASAP7_75t_L g7936 ( 
.A1(n_7504),
.A2(n_7608),
.B(n_7575),
.C(n_7789),
.Y(n_7936)
);

AND2x2_ASAP7_75t_L g7937 ( 
.A(n_7655),
.B(n_111),
.Y(n_7937)
);

AOI21xp5_ASAP7_75t_L g7938 ( 
.A1(n_7725),
.A2(n_670),
.B(n_669),
.Y(n_7938)
);

AO21x1_ASAP7_75t_L g7939 ( 
.A1(n_7486),
.A2(n_670),
.B(n_669),
.Y(n_7939)
);

CKINVDCx11_ASAP7_75t_R g7940 ( 
.A(n_7367),
.Y(n_7940)
);

AND3x2_ASAP7_75t_L g7941 ( 
.A(n_7804),
.B(n_112),
.C(n_113),
.Y(n_7941)
);

AOI21xp5_ASAP7_75t_L g7942 ( 
.A1(n_7605),
.A2(n_673),
.B(n_672),
.Y(n_7942)
);

A2O1A1Ixp33_ASAP7_75t_L g7943 ( 
.A1(n_7485),
.A2(n_116),
.B(n_114),
.C(n_115),
.Y(n_7943)
);

AOI21xp5_ASAP7_75t_L g7944 ( 
.A1(n_7630),
.A2(n_673),
.B(n_672),
.Y(n_7944)
);

A2O1A1Ixp33_ASAP7_75t_L g7945 ( 
.A1(n_7507),
.A2(n_116),
.B(n_114),
.C(n_115),
.Y(n_7945)
);

BUFx6f_ASAP7_75t_L g7946 ( 
.A(n_7479),
.Y(n_7946)
);

OAI21xp5_ASAP7_75t_L g7947 ( 
.A1(n_7510),
.A2(n_114),
.B(n_117),
.Y(n_7947)
);

OAI22xp5_ASAP7_75t_L g7948 ( 
.A1(n_7787),
.A2(n_119),
.B1(n_117),
.B2(n_118),
.Y(n_7948)
);

NOR2xp33_ASAP7_75t_L g7949 ( 
.A(n_7378),
.B(n_674),
.Y(n_7949)
);

INVx2_ASAP7_75t_L g7950 ( 
.A(n_7426),
.Y(n_7950)
);

NAND2xp5_ASAP7_75t_L g7951 ( 
.A(n_7450),
.B(n_117),
.Y(n_7951)
);

AOI21xp5_ASAP7_75t_L g7952 ( 
.A1(n_7641),
.A2(n_678),
.B(n_676),
.Y(n_7952)
);

NAND2xp5_ASAP7_75t_L g7953 ( 
.A(n_7497),
.B(n_7398),
.Y(n_7953)
);

NAND2xp5_ASAP7_75t_L g7954 ( 
.A(n_7401),
.B(n_118),
.Y(n_7954)
);

OAI22xp5_ASAP7_75t_L g7955 ( 
.A1(n_7681),
.A2(n_120),
.B1(n_118),
.B2(n_119),
.Y(n_7955)
);

INVx1_ASAP7_75t_L g7956 ( 
.A(n_7318),
.Y(n_7956)
);

AOI21xp5_ASAP7_75t_L g7957 ( 
.A1(n_7744),
.A2(n_679),
.B(n_678),
.Y(n_7957)
);

INVx2_ASAP7_75t_L g7958 ( 
.A(n_7429),
.Y(n_7958)
);

INVx3_ASAP7_75t_L g7959 ( 
.A(n_7415),
.Y(n_7959)
);

NAND2xp5_ASAP7_75t_L g7960 ( 
.A(n_7416),
.B(n_120),
.Y(n_7960)
);

NOR2xp33_ASAP7_75t_SL g7961 ( 
.A(n_7395),
.B(n_120),
.Y(n_7961)
);

A2O1A1Ixp33_ASAP7_75t_L g7962 ( 
.A1(n_7514),
.A2(n_123),
.B(n_121),
.C(n_122),
.Y(n_7962)
);

OAI21xp5_ASAP7_75t_L g7963 ( 
.A1(n_7554),
.A2(n_121),
.B(n_122),
.Y(n_7963)
);

AO22x1_ASAP7_75t_L g7964 ( 
.A1(n_7437),
.A2(n_123),
.B1(n_121),
.B2(n_122),
.Y(n_7964)
);

NAND2xp5_ASAP7_75t_L g7965 ( 
.A(n_7418),
.B(n_123),
.Y(n_7965)
);

NAND2xp5_ASAP7_75t_SL g7966 ( 
.A(n_7365),
.B(n_679),
.Y(n_7966)
);

NAND2xp5_ASAP7_75t_L g7967 ( 
.A(n_7568),
.B(n_124),
.Y(n_7967)
);

AOI21xp5_ASAP7_75t_L g7968 ( 
.A1(n_7752),
.A2(n_681),
.B(n_680),
.Y(n_7968)
);

OAI21xp5_ASAP7_75t_L g7969 ( 
.A1(n_7632),
.A2(n_124),
.B(n_125),
.Y(n_7969)
);

AND2x4_ASAP7_75t_L g7970 ( 
.A(n_7476),
.B(n_7369),
.Y(n_7970)
);

A2O1A1Ixp33_ASAP7_75t_L g7971 ( 
.A1(n_7660),
.A2(n_126),
.B(n_124),
.C(n_125),
.Y(n_7971)
);

INVx2_ASAP7_75t_L g7972 ( 
.A(n_7434),
.Y(n_7972)
);

CKINVDCx10_ASAP7_75t_R g7973 ( 
.A(n_7413),
.Y(n_7973)
);

NOR2xp33_ASAP7_75t_L g7974 ( 
.A(n_7704),
.B(n_681),
.Y(n_7974)
);

INVx1_ASAP7_75t_L g7975 ( 
.A(n_7319),
.Y(n_7975)
);

O2A1O1Ixp33_ASAP7_75t_L g7976 ( 
.A1(n_7639),
.A2(n_7373),
.B(n_7540),
.C(n_7511),
.Y(n_7976)
);

A2O1A1Ixp33_ASAP7_75t_L g7977 ( 
.A1(n_7679),
.A2(n_127),
.B(n_125),
.C(n_126),
.Y(n_7977)
);

NAND2xp5_ASAP7_75t_L g7978 ( 
.A(n_7693),
.B(n_126),
.Y(n_7978)
);

OAI21xp5_ASAP7_75t_L g7979 ( 
.A1(n_7694),
.A2(n_127),
.B(n_128),
.Y(n_7979)
);

OAI22xp5_ASAP7_75t_L g7980 ( 
.A1(n_7733),
.A2(n_129),
.B1(n_127),
.B2(n_128),
.Y(n_7980)
);

AOI21xp5_ASAP7_75t_L g7981 ( 
.A1(n_7757),
.A2(n_7701),
.B(n_7700),
.Y(n_7981)
);

NAND2xp5_ASAP7_75t_SL g7982 ( 
.A(n_7808),
.B(n_682),
.Y(n_7982)
);

AOI21xp5_ASAP7_75t_L g7983 ( 
.A1(n_7707),
.A2(n_683),
.B(n_682),
.Y(n_7983)
);

NOR2x1p5_ASAP7_75t_SL g7984 ( 
.A(n_7671),
.B(n_683),
.Y(n_7984)
);

AOI21xp5_ASAP7_75t_L g7985 ( 
.A1(n_7710),
.A2(n_685),
.B(n_684),
.Y(n_7985)
);

OAI21xp5_ASAP7_75t_L g7986 ( 
.A1(n_7613),
.A2(n_129),
.B(n_130),
.Y(n_7986)
);

AOI22x1_ASAP7_75t_L g7987 ( 
.A1(n_7385),
.A2(n_131),
.B1(n_129),
.B2(n_130),
.Y(n_7987)
);

AOI21xp5_ASAP7_75t_L g7988 ( 
.A1(n_7766),
.A2(n_686),
.B(n_685),
.Y(n_7988)
);

BUFx4f_ASAP7_75t_L g7989 ( 
.A(n_7347),
.Y(n_7989)
);

AOI21xp5_ASAP7_75t_L g7990 ( 
.A1(n_7675),
.A2(n_687),
.B(n_686),
.Y(n_7990)
);

NOR2xp67_ASAP7_75t_SL g7991 ( 
.A(n_7713),
.B(n_130),
.Y(n_7991)
);

NAND2xp5_ASAP7_75t_L g7992 ( 
.A(n_7334),
.B(n_131),
.Y(n_7992)
);

AOI21xp5_ASAP7_75t_L g7993 ( 
.A1(n_7686),
.A2(n_688),
.B(n_687),
.Y(n_7993)
);

INVx1_ASAP7_75t_L g7994 ( 
.A(n_7321),
.Y(n_7994)
);

INVx2_ASAP7_75t_L g7995 ( 
.A(n_7438),
.Y(n_7995)
);

OAI21xp5_ASAP7_75t_L g7996 ( 
.A1(n_7456),
.A2(n_132),
.B(n_133),
.Y(n_7996)
);

INVx4_ASAP7_75t_L g7997 ( 
.A(n_7402),
.Y(n_7997)
);

NAND2xp5_ASAP7_75t_L g7998 ( 
.A(n_7786),
.B(n_7649),
.Y(n_7998)
);

O2A1O1Ixp33_ASAP7_75t_SL g7999 ( 
.A1(n_7797),
.A2(n_690),
.B(n_691),
.C(n_689),
.Y(n_7999)
);

OAI21xp5_ASAP7_75t_L g8000 ( 
.A1(n_7771),
.A2(n_132),
.B(n_133),
.Y(n_8000)
);

AOI21xp5_ASAP7_75t_L g8001 ( 
.A1(n_7687),
.A2(n_690),
.B(n_689),
.Y(n_8001)
);

INVx1_ASAP7_75t_L g8002 ( 
.A(n_7324),
.Y(n_8002)
);

INVx2_ASAP7_75t_L g8003 ( 
.A(n_7439),
.Y(n_8003)
);

AOI21xp5_ASAP7_75t_L g8004 ( 
.A1(n_7737),
.A2(n_692),
.B(n_691),
.Y(n_8004)
);

AOI21xp5_ASAP7_75t_L g8005 ( 
.A1(n_7743),
.A2(n_693),
.B(n_692),
.Y(n_8005)
);

HB1xp67_ASAP7_75t_L g8006 ( 
.A(n_7316),
.Y(n_8006)
);

INVx1_ASAP7_75t_L g8007 ( 
.A(n_7333),
.Y(n_8007)
);

O2A1O1Ixp33_ASAP7_75t_L g8008 ( 
.A1(n_7548),
.A2(n_7590),
.B(n_7637),
.C(n_7530),
.Y(n_8008)
);

OAI21x1_ASAP7_75t_L g8009 ( 
.A1(n_7747),
.A2(n_132),
.B(n_133),
.Y(n_8009)
);

AND2x2_ASAP7_75t_L g8010 ( 
.A(n_7566),
.B(n_134),
.Y(n_8010)
);

AOI21xp5_ASAP7_75t_L g8011 ( 
.A1(n_7756),
.A2(n_694),
.B(n_693),
.Y(n_8011)
);

INVx2_ASAP7_75t_L g8012 ( 
.A(n_7481),
.Y(n_8012)
);

INVx2_ASAP7_75t_L g8013 ( 
.A(n_7483),
.Y(n_8013)
);

INVx1_ASAP7_75t_L g8014 ( 
.A(n_7335),
.Y(n_8014)
);

OR2x2_ASAP7_75t_L g8015 ( 
.A(n_7745),
.B(n_694),
.Y(n_8015)
);

NAND2xp5_ASAP7_75t_L g8016 ( 
.A(n_7343),
.B(n_7775),
.Y(n_8016)
);

AOI22xp5_ASAP7_75t_L g8017 ( 
.A1(n_7355),
.A2(n_137),
.B1(n_134),
.B2(n_136),
.Y(n_8017)
);

INVx2_ASAP7_75t_L g8018 ( 
.A(n_7487),
.Y(n_8018)
);

O2A1O1Ixp33_ASAP7_75t_L g8019 ( 
.A1(n_7748),
.A2(n_138),
.B(n_136),
.C(n_137),
.Y(n_8019)
);

AOI21xp5_ASAP7_75t_L g8020 ( 
.A1(n_7784),
.A2(n_696),
.B(n_695),
.Y(n_8020)
);

O2A1O1Ixp5_ASAP7_75t_L g8021 ( 
.A1(n_7524),
.A2(n_138),
.B(n_136),
.C(n_137),
.Y(n_8021)
);

NAND2xp5_ASAP7_75t_L g8022 ( 
.A(n_7390),
.B(n_138),
.Y(n_8022)
);

NOR2xp33_ASAP7_75t_L g8023 ( 
.A(n_7598),
.B(n_695),
.Y(n_8023)
);

NAND2xp5_ASAP7_75t_L g8024 ( 
.A(n_7799),
.B(n_139),
.Y(n_8024)
);

AOI21xp5_ASAP7_75t_L g8025 ( 
.A1(n_7793),
.A2(n_698),
.B(n_696),
.Y(n_8025)
);

BUFx3_ASAP7_75t_L g8026 ( 
.A(n_7499),
.Y(n_8026)
);

INVx1_ASAP7_75t_L g8027 ( 
.A(n_7338),
.Y(n_8027)
);

AOI221xp5_ASAP7_75t_SL g8028 ( 
.A1(n_7778),
.A2(n_141),
.B1(n_139),
.B2(n_140),
.C(n_143),
.Y(n_8028)
);

OAI21xp5_ASAP7_75t_L g8029 ( 
.A1(n_7802),
.A2(n_140),
.B(n_141),
.Y(n_8029)
);

AOI33xp33_ASAP7_75t_L g8030 ( 
.A1(n_7515),
.A2(n_143),
.A3(n_145),
.B1(n_140),
.B2(n_141),
.B3(n_144),
.Y(n_8030)
);

AOI21xp5_ASAP7_75t_L g8031 ( 
.A1(n_7382),
.A2(n_699),
.B(n_698),
.Y(n_8031)
);

NAND2xp5_ASAP7_75t_SL g8032 ( 
.A(n_7659),
.B(n_700),
.Y(n_8032)
);

AOI21x1_ASAP7_75t_L g8033 ( 
.A1(n_7363),
.A2(n_7761),
.B(n_7760),
.Y(n_8033)
);

NAND2xp5_ASAP7_75t_L g8034 ( 
.A(n_7742),
.B(n_144),
.Y(n_8034)
);

AOI21x1_ASAP7_75t_L g8035 ( 
.A1(n_7739),
.A2(n_146),
.B(n_147),
.Y(n_8035)
);

NAND2xp5_ASAP7_75t_L g8036 ( 
.A(n_7354),
.B(n_146),
.Y(n_8036)
);

HB1xp67_ASAP7_75t_L g8037 ( 
.A(n_7569),
.Y(n_8037)
);

AOI22x1_ASAP7_75t_L g8038 ( 
.A1(n_7380),
.A2(n_148),
.B1(n_146),
.B2(n_147),
.Y(n_8038)
);

NAND2xp5_ASAP7_75t_L g8039 ( 
.A(n_7371),
.B(n_148),
.Y(n_8039)
);

AOI21xp5_ASAP7_75t_L g8040 ( 
.A1(n_7457),
.A2(n_701),
.B(n_700),
.Y(n_8040)
);

CKINVDCx10_ASAP7_75t_R g8041 ( 
.A(n_7422),
.Y(n_8041)
);

INVx1_ASAP7_75t_L g8042 ( 
.A(n_7340),
.Y(n_8042)
);

NAND2xp5_ASAP7_75t_L g8043 ( 
.A(n_7391),
.B(n_148),
.Y(n_8043)
);

AOI22xp5_ASAP7_75t_L g8044 ( 
.A1(n_7376),
.A2(n_151),
.B1(n_149),
.B2(n_150),
.Y(n_8044)
);

INVx1_ASAP7_75t_SL g8045 ( 
.A(n_7594),
.Y(n_8045)
);

INVx2_ASAP7_75t_L g8046 ( 
.A(n_7341),
.Y(n_8046)
);

INVx3_ASAP7_75t_L g8047 ( 
.A(n_7460),
.Y(n_8047)
);

NAND2xp5_ASAP7_75t_L g8048 ( 
.A(n_7738),
.B(n_149),
.Y(n_8048)
);

A2O1A1Ixp33_ASAP7_75t_L g8049 ( 
.A1(n_7800),
.A2(n_152),
.B(n_150),
.C(n_151),
.Y(n_8049)
);

NOR2xp33_ASAP7_75t_L g8050 ( 
.A(n_7436),
.B(n_702),
.Y(n_8050)
);

AOI21xp5_ASAP7_75t_L g8051 ( 
.A1(n_7699),
.A2(n_703),
.B(n_702),
.Y(n_8051)
);

A2O1A1Ixp33_ASAP7_75t_L g8052 ( 
.A1(n_7803),
.A2(n_154),
.B(n_152),
.C(n_153),
.Y(n_8052)
);

AOI21x1_ASAP7_75t_L g8053 ( 
.A1(n_7740),
.A2(n_152),
.B(n_153),
.Y(n_8053)
);

NAND2xp5_ASAP7_75t_L g8054 ( 
.A(n_7732),
.B(n_153),
.Y(n_8054)
);

AND2x4_ASAP7_75t_L g8055 ( 
.A(n_7383),
.B(n_703),
.Y(n_8055)
);

OAI21xp5_ASAP7_75t_L g8056 ( 
.A1(n_7473),
.A2(n_154),
.B(n_155),
.Y(n_8056)
);

OAI22xp5_ASAP7_75t_L g8057 ( 
.A1(n_7781),
.A2(n_157),
.B1(n_155),
.B2(n_156),
.Y(n_8057)
);

OAI21xp5_ASAP7_75t_L g8058 ( 
.A1(n_7788),
.A2(n_155),
.B(n_157),
.Y(n_8058)
);

A2O1A1Ixp33_ASAP7_75t_L g8059 ( 
.A1(n_7676),
.A2(n_159),
.B(n_157),
.C(n_158),
.Y(n_8059)
);

OAI21xp5_ASAP7_75t_L g8060 ( 
.A1(n_7683),
.A2(n_158),
.B(n_159),
.Y(n_8060)
);

NAND2xp5_ASAP7_75t_L g8061 ( 
.A(n_7428),
.B(n_158),
.Y(n_8061)
);

NAND2xp5_ASAP7_75t_SL g8062 ( 
.A(n_7552),
.B(n_704),
.Y(n_8062)
);

OAI21xp5_ASAP7_75t_L g8063 ( 
.A1(n_7692),
.A2(n_159),
.B(n_160),
.Y(n_8063)
);

AO32x1_ASAP7_75t_L g8064 ( 
.A1(n_7571),
.A2(n_162),
.A3(n_160),
.B1(n_161),
.B2(n_163),
.Y(n_8064)
);

NOR2xp67_ASAP7_75t_SL g8065 ( 
.A(n_7698),
.B(n_160),
.Y(n_8065)
);

AOI21xp5_ASAP7_75t_L g8066 ( 
.A1(n_7342),
.A2(n_7359),
.B(n_7358),
.Y(n_8066)
);

NOR2xp33_ASAP7_75t_L g8067 ( 
.A(n_7356),
.B(n_705),
.Y(n_8067)
);

AND2x4_ASAP7_75t_L g8068 ( 
.A(n_7386),
.B(n_705),
.Y(n_8068)
);

AOI21xp5_ASAP7_75t_L g8069 ( 
.A1(n_7362),
.A2(n_708),
.B(n_707),
.Y(n_8069)
);

AOI21xp5_ASAP7_75t_L g8070 ( 
.A1(n_7370),
.A2(n_709),
.B(n_708),
.Y(n_8070)
);

NAND2xp5_ASAP7_75t_L g8071 ( 
.A(n_7432),
.B(n_161),
.Y(n_8071)
);

AOI21xp5_ASAP7_75t_L g8072 ( 
.A1(n_7372),
.A2(n_711),
.B(n_710),
.Y(n_8072)
);

NAND2xp5_ASAP7_75t_L g8073 ( 
.A(n_7435),
.B(n_161),
.Y(n_8073)
);

NAND2xp5_ASAP7_75t_L g8074 ( 
.A(n_7444),
.B(n_162),
.Y(n_8074)
);

BUFx3_ASAP7_75t_L g8075 ( 
.A(n_7516),
.Y(n_8075)
);

INVx1_ASAP7_75t_L g8076 ( 
.A(n_7375),
.Y(n_8076)
);

O2A1O1Ixp33_ASAP7_75t_SL g8077 ( 
.A1(n_7749),
.A2(n_711),
.B(n_712),
.C(n_710),
.Y(n_8077)
);

NAND2xp5_ASAP7_75t_L g8078 ( 
.A(n_7445),
.B(n_162),
.Y(n_8078)
);

AOI21xp5_ASAP7_75t_L g8079 ( 
.A1(n_7389),
.A2(n_715),
.B(n_714),
.Y(n_8079)
);

NAND2xp5_ASAP7_75t_L g8080 ( 
.A(n_7448),
.B(n_163),
.Y(n_8080)
);

NAND2xp5_ASAP7_75t_L g8081 ( 
.A(n_7453),
.B(n_163),
.Y(n_8081)
);

NAND2xp5_ASAP7_75t_L g8082 ( 
.A(n_7465),
.B(n_164),
.Y(n_8082)
);

A2O1A1Ixp33_ASAP7_75t_L g8083 ( 
.A1(n_7616),
.A2(n_166),
.B(n_164),
.C(n_165),
.Y(n_8083)
);

CKINVDCx10_ASAP7_75t_R g8084 ( 
.A(n_7337),
.Y(n_8084)
);

NAND2xp5_ASAP7_75t_SL g8085 ( 
.A(n_7785),
.B(n_714),
.Y(n_8085)
);

INVx1_ASAP7_75t_L g8086 ( 
.A(n_7393),
.Y(n_8086)
);

AND2x4_ASAP7_75t_L g8087 ( 
.A(n_7691),
.B(n_716),
.Y(n_8087)
);

BUFx4f_ASAP7_75t_L g8088 ( 
.A(n_7350),
.Y(n_8088)
);

NAND2xp5_ASAP7_75t_L g8089 ( 
.A(n_7468),
.B(n_7474),
.Y(n_8089)
);

AOI21xp5_ASAP7_75t_L g8090 ( 
.A1(n_7405),
.A2(n_717),
.B(n_716),
.Y(n_8090)
);

AND2x2_ASAP7_75t_SL g8091 ( 
.A(n_7557),
.B(n_717),
.Y(n_8091)
);

INVx1_ASAP7_75t_L g8092 ( 
.A(n_7406),
.Y(n_8092)
);

OAI22xp5_ASAP7_75t_L g8093 ( 
.A1(n_7750),
.A2(n_166),
.B1(n_164),
.B2(n_165),
.Y(n_8093)
);

AOI21xp5_ASAP7_75t_L g8094 ( 
.A1(n_7407),
.A2(n_719),
.B(n_718),
.Y(n_8094)
);

AND2x4_ASAP7_75t_L g8095 ( 
.A(n_7420),
.B(n_718),
.Y(n_8095)
);

INVxp67_ASAP7_75t_SL g8096 ( 
.A(n_7588),
.Y(n_8096)
);

AND2x2_ASAP7_75t_L g8097 ( 
.A(n_7467),
.B(n_165),
.Y(n_8097)
);

NAND2x1p5_ASAP7_75t_L g8098 ( 
.A(n_7631),
.B(n_7625),
.Y(n_8098)
);

NOR2xp33_ASAP7_75t_L g8099 ( 
.A(n_7688),
.B(n_7379),
.Y(n_8099)
);

OAI21xp33_ASAP7_75t_L g8100 ( 
.A1(n_7556),
.A2(n_7527),
.B(n_7495),
.Y(n_8100)
);

NAND2xp5_ASAP7_75t_L g8101 ( 
.A(n_7477),
.B(n_166),
.Y(n_8101)
);

BUFx2_ASAP7_75t_L g8102 ( 
.A(n_7544),
.Y(n_8102)
);

AOI21xp5_ASAP7_75t_L g8103 ( 
.A1(n_7412),
.A2(n_721),
.B(n_720),
.Y(n_8103)
);

O2A1O1Ixp33_ASAP7_75t_L g8104 ( 
.A1(n_7449),
.A2(n_169),
.B(n_167),
.C(n_168),
.Y(n_8104)
);

O2A1O1Ixp5_ASAP7_75t_L g8105 ( 
.A1(n_7417),
.A2(n_169),
.B(n_167),
.C(n_168),
.Y(n_8105)
);

NAND2xp5_ASAP7_75t_L g8106 ( 
.A(n_7478),
.B(n_167),
.Y(n_8106)
);

OAI22xp5_ASAP7_75t_L g8107 ( 
.A1(n_7783),
.A2(n_171),
.B1(n_168),
.B2(n_170),
.Y(n_8107)
);

NAND2xp5_ASAP7_75t_L g8108 ( 
.A(n_7480),
.B(n_7482),
.Y(n_8108)
);

NOR2xp33_ASAP7_75t_L g8109 ( 
.A(n_7463),
.B(n_720),
.Y(n_8109)
);

NAND2xp5_ASAP7_75t_L g8110 ( 
.A(n_7411),
.B(n_170),
.Y(n_8110)
);

NOR2xp33_ASAP7_75t_L g8111 ( 
.A(n_7665),
.B(n_7801),
.Y(n_8111)
);

AOI21xp5_ASAP7_75t_L g8112 ( 
.A1(n_7423),
.A2(n_722),
.B(n_721),
.Y(n_8112)
);

CKINVDCx14_ASAP7_75t_R g8113 ( 
.A(n_7656),
.Y(n_8113)
);

NAND2xp5_ASAP7_75t_L g8114 ( 
.A(n_7425),
.B(n_170),
.Y(n_8114)
);

AOI21xp5_ASAP7_75t_L g8115 ( 
.A1(n_7462),
.A2(n_723),
.B(n_722),
.Y(n_8115)
);

INVx2_ASAP7_75t_L g8116 ( 
.A(n_7494),
.Y(n_8116)
);

NOR2xp33_ASAP7_75t_L g8117 ( 
.A(n_7751),
.B(n_723),
.Y(n_8117)
);

INVx1_ASAP7_75t_L g8118 ( 
.A(n_7488),
.Y(n_8118)
);

OAI21xp5_ASAP7_75t_L g8119 ( 
.A1(n_7419),
.A2(n_172),
.B(n_173),
.Y(n_8119)
);

AOI21xp5_ASAP7_75t_L g8120 ( 
.A1(n_7489),
.A2(n_725),
.B(n_724),
.Y(n_8120)
);

INVx1_ASAP7_75t_L g8121 ( 
.A(n_7500),
.Y(n_8121)
);

NAND2xp5_ASAP7_75t_L g8122 ( 
.A(n_7503),
.B(n_172),
.Y(n_8122)
);

NOR2xp33_ASAP7_75t_L g8123 ( 
.A(n_7780),
.B(n_724),
.Y(n_8123)
);

NAND2xp5_ASAP7_75t_SL g8124 ( 
.A(n_7774),
.B(n_726),
.Y(n_8124)
);

INVx1_ASAP7_75t_L g8125 ( 
.A(n_7505),
.Y(n_8125)
);

NAND2xp5_ASAP7_75t_SL g8126 ( 
.A(n_7603),
.B(n_726),
.Y(n_8126)
);

NOR2xp33_ASAP7_75t_L g8127 ( 
.A(n_7724),
.B(n_727),
.Y(n_8127)
);

A2O1A1Ixp33_ASAP7_75t_L g8128 ( 
.A1(n_7722),
.A2(n_7806),
.B(n_7537),
.C(n_7617),
.Y(n_8128)
);

AOI21xp5_ASAP7_75t_L g8129 ( 
.A1(n_7323),
.A2(n_728),
.B(n_727),
.Y(n_8129)
);

INVx2_ASAP7_75t_L g8130 ( 
.A(n_7506),
.Y(n_8130)
);

AOI21xp5_ASAP7_75t_L g8131 ( 
.A1(n_7512),
.A2(n_729),
.B(n_728),
.Y(n_8131)
);

AND2x4_ASAP7_75t_L g8132 ( 
.A(n_7546),
.B(n_729),
.Y(n_8132)
);

NAND2xp5_ASAP7_75t_L g8133 ( 
.A(n_7513),
.B(n_172),
.Y(n_8133)
);

INVx1_ASAP7_75t_L g8134 ( 
.A(n_7519),
.Y(n_8134)
);

INVx2_ASAP7_75t_L g8135 ( 
.A(n_7522),
.Y(n_8135)
);

INVx1_ASAP7_75t_SL g8136 ( 
.A(n_7612),
.Y(n_8136)
);

AND2x2_ASAP7_75t_L g8137 ( 
.A(n_7509),
.B(n_173),
.Y(n_8137)
);

AOI21x1_ASAP7_75t_L g8138 ( 
.A1(n_7392),
.A2(n_173),
.B(n_174),
.Y(n_8138)
);

A2O1A1Ixp33_ASAP7_75t_L g8139 ( 
.A1(n_7768),
.A2(n_176),
.B(n_174),
.C(n_175),
.Y(n_8139)
);

NOR2xp33_ASAP7_75t_L g8140 ( 
.A(n_7777),
.B(n_730),
.Y(n_8140)
);

AOI21xp5_ASAP7_75t_L g8141 ( 
.A1(n_7559),
.A2(n_732),
.B(n_730),
.Y(n_8141)
);

AOI21xp5_ASAP7_75t_L g8142 ( 
.A1(n_7475),
.A2(n_733),
.B(n_732),
.Y(n_8142)
);

NAND2xp5_ASAP7_75t_L g8143 ( 
.A(n_7374),
.B(n_174),
.Y(n_8143)
);

NAND2xp5_ASAP7_75t_SL g8144 ( 
.A(n_7762),
.B(n_733),
.Y(n_8144)
);

BUFx2_ASAP7_75t_L g8145 ( 
.A(n_7387),
.Y(n_8145)
);

NAND2xp5_ASAP7_75t_L g8146 ( 
.A(n_7586),
.B(n_7492),
.Y(n_8146)
);

OAI21xp5_ASAP7_75t_L g8147 ( 
.A1(n_7451),
.A2(n_175),
.B(n_176),
.Y(n_8147)
);

NAND2xp5_ASAP7_75t_L g8148 ( 
.A(n_7526),
.B(n_175),
.Y(n_8148)
);

AOI22xp33_ASAP7_75t_L g8149 ( 
.A1(n_7606),
.A2(n_178),
.B1(n_176),
.B2(n_177),
.Y(n_8149)
);

AOI21xp5_ASAP7_75t_L g8150 ( 
.A1(n_7670),
.A2(n_735),
.B(n_734),
.Y(n_8150)
);

INVx1_ASAP7_75t_L g8151 ( 
.A(n_7542),
.Y(n_8151)
);

NAND2xp5_ASAP7_75t_L g8152 ( 
.A(n_7555),
.B(n_177),
.Y(n_8152)
);

AOI21x1_ASAP7_75t_L g8153 ( 
.A1(n_7549),
.A2(n_177),
.B(n_178),
.Y(n_8153)
);

BUFx4f_ASAP7_75t_L g8154 ( 
.A(n_7366),
.Y(n_8154)
);

OAI21xp5_ASAP7_75t_L g8155 ( 
.A1(n_7721),
.A2(n_179),
.B(n_180),
.Y(n_8155)
);

NAND2xp5_ASAP7_75t_L g8156 ( 
.A(n_7561),
.B(n_179),
.Y(n_8156)
);

NAND2xp5_ASAP7_75t_L g8157 ( 
.A(n_7721),
.B(n_179),
.Y(n_8157)
);

AOI22xp5_ASAP7_75t_L g8158 ( 
.A1(n_7702),
.A2(n_182),
.B1(n_180),
.B2(n_181),
.Y(n_8158)
);

NAND2xp5_ASAP7_75t_SL g8159 ( 
.A(n_7762),
.B(n_735),
.Y(n_8159)
);

AOI21xp5_ASAP7_75t_L g8160 ( 
.A1(n_7636),
.A2(n_737),
.B(n_736),
.Y(n_8160)
);

AO21x1_ASAP7_75t_L g8161 ( 
.A1(n_7805),
.A2(n_737),
.B(n_736),
.Y(n_8161)
);

AOI21xp5_ASAP7_75t_L g8162 ( 
.A1(n_7565),
.A2(n_739),
.B(n_738),
.Y(n_8162)
);

INVx2_ASAP7_75t_L g8163 ( 
.A(n_7538),
.Y(n_8163)
);

AOI21xp5_ASAP7_75t_L g8164 ( 
.A1(n_7721),
.A2(n_740),
.B(n_738),
.Y(n_8164)
);

INVx1_ASAP7_75t_L g8165 ( 
.A(n_7550),
.Y(n_8165)
);

NAND2xp5_ASAP7_75t_L g8166 ( 
.A(n_7578),
.B(n_180),
.Y(n_8166)
);

NOR2x1_ASAP7_75t_R g8167 ( 
.A(n_7741),
.B(n_740),
.Y(n_8167)
);

INVx3_ASAP7_75t_L g8168 ( 
.A(n_7618),
.Y(n_8168)
);

OAI21xp5_ASAP7_75t_L g8169 ( 
.A1(n_7424),
.A2(n_181),
.B(n_182),
.Y(n_8169)
);

NAND3xp33_ASAP7_75t_L g8170 ( 
.A(n_7498),
.B(n_182),
.C(n_183),
.Y(n_8170)
);

AOI21x1_ASAP7_75t_L g8171 ( 
.A1(n_7562),
.A2(n_183),
.B(n_184),
.Y(n_8171)
);

AOI21xp33_ASAP7_75t_L g8172 ( 
.A1(n_7535),
.A2(n_184),
.B(n_185),
.Y(n_8172)
);

AOI21xp5_ASAP7_75t_L g8173 ( 
.A1(n_7520),
.A2(n_742),
.B(n_741),
.Y(n_8173)
);

NAND2x1p5_ASAP7_75t_L g8174 ( 
.A(n_7618),
.B(n_741),
.Y(n_8174)
);

NAND2x1p5_ASAP7_75t_L g8175 ( 
.A(n_7653),
.B(n_743),
.Y(n_8175)
);

BUFx4f_ASAP7_75t_L g8176 ( 
.A(n_7525),
.Y(n_8176)
);

OAI21xp5_ASAP7_75t_L g8177 ( 
.A1(n_7443),
.A2(n_185),
.B(n_186),
.Y(n_8177)
);

INVx1_ASAP7_75t_L g8178 ( 
.A(n_7563),
.Y(n_8178)
);

AOI22xp33_ASAP7_75t_L g8179 ( 
.A1(n_7469),
.A2(n_187),
.B1(n_185),
.B2(n_186),
.Y(n_8179)
);

NAND2xp33_ASAP7_75t_L g8180 ( 
.A(n_7708),
.B(n_186),
.Y(n_8180)
);

OAI21xp5_ASAP7_75t_L g8181 ( 
.A1(n_7521),
.A2(n_187),
.B(n_188),
.Y(n_8181)
);

AND2x2_ASAP7_75t_L g8182 ( 
.A(n_7685),
.B(n_187),
.Y(n_8182)
);

NAND2xp5_ASAP7_75t_SL g8183 ( 
.A(n_7709),
.B(n_743),
.Y(n_8183)
);

NOR3xp33_ASAP7_75t_L g8184 ( 
.A(n_7678),
.B(n_188),
.C(n_189),
.Y(n_8184)
);

INVx1_ASAP7_75t_L g8185 ( 
.A(n_7564),
.Y(n_8185)
);

NAND2xp5_ASAP7_75t_L g8186 ( 
.A(n_7600),
.B(n_188),
.Y(n_8186)
);

NAND2xp5_ASAP7_75t_L g8187 ( 
.A(n_7410),
.B(n_189),
.Y(n_8187)
);

INVx2_ASAP7_75t_L g8188 ( 
.A(n_7523),
.Y(n_8188)
);

A2O1A1Ixp33_ASAP7_75t_L g8189 ( 
.A1(n_7528),
.A2(n_191),
.B(n_189),
.C(n_190),
.Y(n_8189)
);

NOR2xp33_ASAP7_75t_L g8190 ( 
.A(n_7599),
.B(n_745),
.Y(n_8190)
);

NAND2xp5_ASAP7_75t_SL g8191 ( 
.A(n_7746),
.B(n_745),
.Y(n_8191)
);

NAND2xp5_ASAP7_75t_L g8192 ( 
.A(n_7531),
.B(n_190),
.Y(n_8192)
);

AOI21xp5_ASAP7_75t_L g8193 ( 
.A1(n_7532),
.A2(n_747),
.B(n_746),
.Y(n_8193)
);

NAND2xp5_ASAP7_75t_L g8194 ( 
.A(n_7534),
.B(n_190),
.Y(n_8194)
);

NAND2xp5_ASAP7_75t_L g8195 ( 
.A(n_7536),
.B(n_191),
.Y(n_8195)
);

NAND2xp5_ASAP7_75t_L g8196 ( 
.A(n_7602),
.B(n_191),
.Y(n_8196)
);

OAI21xp5_ASAP7_75t_L g8197 ( 
.A1(n_7431),
.A2(n_192),
.B(n_193),
.Y(n_8197)
);

INVx1_ASAP7_75t_L g8198 ( 
.A(n_7645),
.Y(n_8198)
);

AOI21xp33_ASAP7_75t_L g8199 ( 
.A1(n_7472),
.A2(n_7680),
.B(n_7662),
.Y(n_8199)
);

AOI33xp33_ASAP7_75t_L g8200 ( 
.A1(n_7430),
.A2(n_194),
.A3(n_196),
.B1(n_192),
.B2(n_193),
.B3(n_195),
.Y(n_8200)
);

OAI321xp33_ASAP7_75t_L g8201 ( 
.A1(n_7624),
.A2(n_7547),
.A3(n_7496),
.B1(n_7508),
.B2(n_7545),
.C(n_7533),
.Y(n_8201)
);

XNOR2xp5_ASAP7_75t_L g8202 ( 
.A(n_7763),
.B(n_192),
.Y(n_8202)
);

NAND2xp5_ASAP7_75t_L g8203 ( 
.A(n_7614),
.B(n_193),
.Y(n_8203)
);

NOR2xp67_ASAP7_75t_L g8204 ( 
.A(n_7409),
.B(n_194),
.Y(n_8204)
);

OAI21xp5_ASAP7_75t_L g8205 ( 
.A1(n_7452),
.A2(n_194),
.B(n_195),
.Y(n_8205)
);

A2O1A1Ixp33_ASAP7_75t_L g8206 ( 
.A1(n_7765),
.A2(n_7791),
.B(n_7648),
.C(n_7652),
.Y(n_8206)
);

NAND2xp5_ASAP7_75t_L g8207 ( 
.A(n_7459),
.B(n_195),
.Y(n_8207)
);

INVx1_ASAP7_75t_L g8208 ( 
.A(n_7718),
.Y(n_8208)
);

NOR2xp33_ASAP7_75t_L g8209 ( 
.A(n_7408),
.B(n_748),
.Y(n_8209)
);

AND2x2_ASAP7_75t_L g8210 ( 
.A(n_7609),
.B(n_196),
.Y(n_8210)
);

AND2x2_ASAP7_75t_L g8211 ( 
.A(n_7619),
.B(n_197),
.Y(n_8211)
);

CKINVDCx14_ASAP7_75t_R g8212 ( 
.A(n_7597),
.Y(n_8212)
);

NAND2xp5_ASAP7_75t_L g8213 ( 
.A(n_7567),
.B(n_197),
.Y(n_8213)
);

AOI21xp5_ASAP7_75t_L g8214 ( 
.A1(n_7628),
.A2(n_750),
.B(n_748),
.Y(n_8214)
);

OAI22x1_ASAP7_75t_L g8215 ( 
.A1(n_7501),
.A2(n_199),
.B1(n_197),
.B2(n_198),
.Y(n_8215)
);

NOR2xp67_ASAP7_75t_L g8216 ( 
.A(n_7640),
.B(n_198),
.Y(n_8216)
);

INVx1_ASAP7_75t_L g8217 ( 
.A(n_7696),
.Y(n_8217)
);

NAND2xp5_ASAP7_75t_L g8218 ( 
.A(n_7396),
.B(n_198),
.Y(n_8218)
);

O2A1O1Ixp5_ASAP7_75t_L g8219 ( 
.A1(n_7666),
.A2(n_201),
.B(n_199),
.C(n_200),
.Y(n_8219)
);

NAND2xp5_ASAP7_75t_L g8220 ( 
.A(n_7734),
.B(n_199),
.Y(n_8220)
);

BUFx2_ASAP7_75t_L g8221 ( 
.A(n_7582),
.Y(n_8221)
);

NAND2xp5_ASAP7_75t_SL g8222 ( 
.A(n_7427),
.B(n_751),
.Y(n_8222)
);

NAND2xp5_ASAP7_75t_L g8223 ( 
.A(n_7735),
.B(n_200),
.Y(n_8223)
);

INVx4_ASAP7_75t_L g8224 ( 
.A(n_7587),
.Y(n_8224)
);

INVx3_ASAP7_75t_L g8225 ( 
.A(n_7589),
.Y(n_8225)
);

O2A1O1Ixp33_ASAP7_75t_SL g8226 ( 
.A1(n_7601),
.A2(n_752),
.B(n_753),
.C(n_751),
.Y(n_8226)
);

NAND2xp5_ASAP7_75t_SL g8227 ( 
.A(n_7658),
.B(n_752),
.Y(n_8227)
);

AOI21xp5_ASAP7_75t_L g8228 ( 
.A1(n_7577),
.A2(n_754),
.B(n_753),
.Y(n_8228)
);

NAND2xp5_ASAP7_75t_SL g8229 ( 
.A(n_7753),
.B(n_754),
.Y(n_8229)
);

AOI21xp5_ASAP7_75t_L g8230 ( 
.A1(n_7727),
.A2(n_756),
.B(n_755),
.Y(n_8230)
);

AOI21xp5_ASAP7_75t_L g8231 ( 
.A1(n_7769),
.A2(n_756),
.B(n_755),
.Y(n_8231)
);

NOR2xp33_ASAP7_75t_L g8232 ( 
.A(n_7736),
.B(n_757),
.Y(n_8232)
);

O2A1O1Ixp33_ASAP7_75t_L g8233 ( 
.A1(n_7596),
.A2(n_203),
.B(n_201),
.C(n_202),
.Y(n_8233)
);

INVx3_ASAP7_75t_L g8234 ( 
.A(n_7591),
.Y(n_8234)
);

NAND2xp5_ASAP7_75t_L g8235 ( 
.A(n_7622),
.B(n_201),
.Y(n_8235)
);

NAND2xp5_ASAP7_75t_L g8236 ( 
.A(n_7629),
.B(n_202),
.Y(n_8236)
);

OAI21xp5_ASAP7_75t_L g8237 ( 
.A1(n_7773),
.A2(n_202),
.B(n_203),
.Y(n_8237)
);

NAND2xp5_ASAP7_75t_L g8238 ( 
.A(n_7657),
.B(n_7790),
.Y(n_8238)
);

AO32x2_ASAP7_75t_L g8239 ( 
.A1(n_7491),
.A2(n_206),
.A3(n_204),
.B1(n_205),
.B2(n_207),
.Y(n_8239)
);

BUFx2_ASAP7_75t_L g8240 ( 
.A(n_7558),
.Y(n_8240)
);

NAND2xp5_ASAP7_75t_SL g8241 ( 
.A(n_7711),
.B(n_757),
.Y(n_8241)
);

AOI22xp5_ASAP7_75t_L g8242 ( 
.A1(n_7794),
.A2(n_206),
.B1(n_204),
.B2(n_205),
.Y(n_8242)
);

NOR2xp33_ASAP7_75t_L g8243 ( 
.A(n_7592),
.B(n_758),
.Y(n_8243)
);

AOI21xp5_ASAP7_75t_L g8244 ( 
.A1(n_7646),
.A2(n_7647),
.B(n_7502),
.Y(n_8244)
);

NAND2xp5_ASAP7_75t_L g8245 ( 
.A(n_7796),
.B(n_204),
.Y(n_8245)
);

INVx2_ASAP7_75t_L g8246 ( 
.A(n_7593),
.Y(n_8246)
);

NAND2xp5_ASAP7_75t_L g8247 ( 
.A(n_7611),
.B(n_207),
.Y(n_8247)
);

INVx3_ASAP7_75t_L g8248 ( 
.A(n_7312),
.Y(n_8248)
);

INVx2_ASAP7_75t_L g8249 ( 
.A(n_7320),
.Y(n_8249)
);

BUFx6f_ASAP7_75t_L g8250 ( 
.A(n_7518),
.Y(n_8250)
);

AOI21xp5_ASAP7_75t_L g8251 ( 
.A1(n_7446),
.A2(n_760),
.B(n_759),
.Y(n_8251)
);

AOI21xp5_ASAP7_75t_L g8252 ( 
.A1(n_7446),
.A2(n_760),
.B(n_759),
.Y(n_8252)
);

NOR2xp33_ASAP7_75t_L g8253 ( 
.A(n_7446),
.B(n_761),
.Y(n_8253)
);

AOI21xp5_ASAP7_75t_L g8254 ( 
.A1(n_7446),
.A2(n_762),
.B(n_761),
.Y(n_8254)
);

NOR2xp33_ASAP7_75t_L g8255 ( 
.A(n_7446),
.B(n_763),
.Y(n_8255)
);

NOR2x1_ASAP7_75t_L g8256 ( 
.A(n_7330),
.B(n_763),
.Y(n_8256)
);

NAND2xp5_ASAP7_75t_L g8257 ( 
.A(n_7446),
.B(n_208),
.Y(n_8257)
);

NOR2xp33_ASAP7_75t_L g8258 ( 
.A(n_7446),
.B(n_764),
.Y(n_8258)
);

INVx1_ASAP7_75t_SL g8259 ( 
.A(n_7316),
.Y(n_8259)
);

AOI21xp5_ASAP7_75t_L g8260 ( 
.A1(n_7446),
.A2(n_766),
.B(n_765),
.Y(n_8260)
);

OAI21xp33_ASAP7_75t_L g8261 ( 
.A1(n_7446),
.A2(n_208),
.B(n_209),
.Y(n_8261)
);

NAND2xp5_ASAP7_75t_L g8262 ( 
.A(n_7446),
.B(n_209),
.Y(n_8262)
);

OAI22xp5_ASAP7_75t_L g8263 ( 
.A1(n_7446),
.A2(n_211),
.B1(n_209),
.B2(n_210),
.Y(n_8263)
);

AOI21xp5_ASAP7_75t_L g8264 ( 
.A1(n_7446),
.A2(n_767),
.B(n_766),
.Y(n_8264)
);

NAND2xp5_ASAP7_75t_L g8265 ( 
.A(n_7446),
.B(n_210),
.Y(n_8265)
);

INVx1_ASAP7_75t_L g8266 ( 
.A(n_7320),
.Y(n_8266)
);

INVx2_ASAP7_75t_L g8267 ( 
.A(n_7320),
.Y(n_8267)
);

NAND2xp5_ASAP7_75t_L g8268 ( 
.A(n_7446),
.B(n_210),
.Y(n_8268)
);

AOI21xp5_ASAP7_75t_L g8269 ( 
.A1(n_7446),
.A2(n_769),
.B(n_768),
.Y(n_8269)
);

AOI21xp5_ASAP7_75t_L g8270 ( 
.A1(n_7446),
.A2(n_770),
.B(n_769),
.Y(n_8270)
);

INVx3_ASAP7_75t_L g8271 ( 
.A(n_7312),
.Y(n_8271)
);

INVx1_ASAP7_75t_L g8272 ( 
.A(n_7320),
.Y(n_8272)
);

BUFx3_ASAP7_75t_L g8273 ( 
.A(n_7312),
.Y(n_8273)
);

NAND2xp5_ASAP7_75t_SL g8274 ( 
.A(n_7446),
.B(n_770),
.Y(n_8274)
);

AOI21xp5_ASAP7_75t_L g8275 ( 
.A1(n_7446),
.A2(n_772),
.B(n_771),
.Y(n_8275)
);

NOR2xp33_ASAP7_75t_L g8276 ( 
.A(n_7446),
.B(n_772),
.Y(n_8276)
);

AOI21xp5_ASAP7_75t_L g8277 ( 
.A1(n_7446),
.A2(n_774),
.B(n_773),
.Y(n_8277)
);

NAND2xp5_ASAP7_75t_L g8278 ( 
.A(n_7446),
.B(n_211),
.Y(n_8278)
);

AOI21xp5_ASAP7_75t_L g8279 ( 
.A1(n_7446),
.A2(n_774),
.B(n_773),
.Y(n_8279)
);

AOI21x1_ASAP7_75t_L g8280 ( 
.A1(n_7605),
.A2(n_212),
.B(n_213),
.Y(n_8280)
);

NAND2xp5_ASAP7_75t_L g8281 ( 
.A(n_7446),
.B(n_212),
.Y(n_8281)
);

O2A1O1Ixp33_ASAP7_75t_L g8282 ( 
.A1(n_7446),
.A2(n_215),
.B(n_212),
.C(n_213),
.Y(n_8282)
);

AOI21xp5_ASAP7_75t_L g8283 ( 
.A1(n_7446),
.A2(n_776),
.B(n_775),
.Y(n_8283)
);

AOI21xp5_ASAP7_75t_L g8284 ( 
.A1(n_7446),
.A2(n_776),
.B(n_775),
.Y(n_8284)
);

AOI21xp5_ASAP7_75t_L g8285 ( 
.A1(n_7446),
.A2(n_778),
.B(n_777),
.Y(n_8285)
);

AOI21xp5_ASAP7_75t_L g8286 ( 
.A1(n_7446),
.A2(n_779),
.B(n_778),
.Y(n_8286)
);

NOR2xp33_ASAP7_75t_L g8287 ( 
.A(n_7446),
.B(n_779),
.Y(n_8287)
);

AOI21xp5_ASAP7_75t_L g8288 ( 
.A1(n_7446),
.A2(n_781),
.B(n_780),
.Y(n_8288)
);

O2A1O1Ixp33_ASAP7_75t_L g8289 ( 
.A1(n_7446),
.A2(n_216),
.B(n_213),
.C(n_215),
.Y(n_8289)
);

NOR2xp33_ASAP7_75t_L g8290 ( 
.A(n_7446),
.B(n_780),
.Y(n_8290)
);

NOR3xp33_ASAP7_75t_L g8291 ( 
.A(n_7446),
.B(n_216),
.C(n_217),
.Y(n_8291)
);

INVx2_ASAP7_75t_L g8292 ( 
.A(n_7320),
.Y(n_8292)
);

AOI21xp5_ASAP7_75t_L g8293 ( 
.A1(n_7446),
.A2(n_782),
.B(n_781),
.Y(n_8293)
);

BUFx2_ASAP7_75t_L g8294 ( 
.A(n_7553),
.Y(n_8294)
);

AOI21x1_ASAP7_75t_L g8295 ( 
.A1(n_7605),
.A2(n_217),
.B(n_218),
.Y(n_8295)
);

AOI22xp5_ASAP7_75t_L g8296 ( 
.A1(n_7446),
.A2(n_219),
.B1(n_217),
.B2(n_218),
.Y(n_8296)
);

BUFx6f_ASAP7_75t_L g8297 ( 
.A(n_7518),
.Y(n_8297)
);

AOI21xp5_ASAP7_75t_L g8298 ( 
.A1(n_7446),
.A2(n_783),
.B(n_782),
.Y(n_8298)
);

NAND2xp5_ASAP7_75t_L g8299 ( 
.A(n_7446),
.B(n_218),
.Y(n_8299)
);

O2A1O1Ixp33_ASAP7_75t_L g8300 ( 
.A1(n_7446),
.A2(n_221),
.B(n_219),
.C(n_220),
.Y(n_8300)
);

O2A1O1Ixp33_ASAP7_75t_L g8301 ( 
.A1(n_7446),
.A2(n_222),
.B(n_220),
.C(n_221),
.Y(n_8301)
);

CKINVDCx8_ASAP7_75t_R g8302 ( 
.A(n_7344),
.Y(n_8302)
);

BUFx2_ASAP7_75t_L g8303 ( 
.A(n_7553),
.Y(n_8303)
);

AOI21x1_ASAP7_75t_L g8304 ( 
.A1(n_7605),
.A2(n_220),
.B(n_221),
.Y(n_8304)
);

A2O1A1Ixp33_ASAP7_75t_L g8305 ( 
.A1(n_7446),
.A2(n_224),
.B(n_222),
.C(n_223),
.Y(n_8305)
);

BUFx8_ASAP7_75t_L g8306 ( 
.A(n_7326),
.Y(n_8306)
);

AOI21xp5_ASAP7_75t_L g8307 ( 
.A1(n_7446),
.A2(n_784),
.B(n_783),
.Y(n_8307)
);

INVx1_ASAP7_75t_SL g8308 ( 
.A(n_7316),
.Y(n_8308)
);

INVx2_ASAP7_75t_L g8309 ( 
.A(n_7320),
.Y(n_8309)
);

INVx1_ASAP7_75t_L g8310 ( 
.A(n_7320),
.Y(n_8310)
);

INVx1_ASAP7_75t_L g8311 ( 
.A(n_7320),
.Y(n_8311)
);

AOI21xp5_ASAP7_75t_L g8312 ( 
.A1(n_7446),
.A2(n_785),
.B(n_784),
.Y(n_8312)
);

AOI21xp5_ASAP7_75t_L g8313 ( 
.A1(n_7446),
.A2(n_786),
.B(n_785),
.Y(n_8313)
);

INVx2_ASAP7_75t_L g8314 ( 
.A(n_7320),
.Y(n_8314)
);

CKINVDCx10_ASAP7_75t_R g8315 ( 
.A(n_7517),
.Y(n_8315)
);

INVx1_ASAP7_75t_L g8316 ( 
.A(n_7320),
.Y(n_8316)
);

AOI22xp5_ASAP7_75t_L g8317 ( 
.A1(n_7446),
.A2(n_225),
.B1(n_223),
.B2(n_224),
.Y(n_8317)
);

NAND2xp5_ASAP7_75t_L g8318 ( 
.A(n_7446),
.B(n_223),
.Y(n_8318)
);

NAND2xp5_ASAP7_75t_L g8319 ( 
.A(n_7446),
.B(n_224),
.Y(n_8319)
);

NAND2xp5_ASAP7_75t_L g8320 ( 
.A(n_7446),
.B(n_225),
.Y(n_8320)
);

INVx1_ASAP7_75t_L g8321 ( 
.A(n_7320),
.Y(n_8321)
);

NAND2xp5_ASAP7_75t_L g8322 ( 
.A(n_7446),
.B(n_225),
.Y(n_8322)
);

INVx1_ASAP7_75t_L g8323 ( 
.A(n_7320),
.Y(n_8323)
);

OAI21xp33_ASAP7_75t_L g8324 ( 
.A1(n_7446),
.A2(n_226),
.B(n_227),
.Y(n_8324)
);

INVx2_ASAP7_75t_L g8325 ( 
.A(n_7320),
.Y(n_8325)
);

OAI21xp5_ASAP7_75t_L g8326 ( 
.A1(n_7446),
.A2(n_226),
.B(n_227),
.Y(n_8326)
);

INVx2_ASAP7_75t_L g8327 ( 
.A(n_7320),
.Y(n_8327)
);

AOI21xp5_ASAP7_75t_L g8328 ( 
.A1(n_7446),
.A2(n_788),
.B(n_787),
.Y(n_8328)
);

AOI21xp5_ASAP7_75t_L g8329 ( 
.A1(n_7446),
.A2(n_789),
.B(n_788),
.Y(n_8329)
);

AOI21xp5_ASAP7_75t_L g8330 ( 
.A1(n_7446),
.A2(n_790),
.B(n_789),
.Y(n_8330)
);

NOR2xp33_ASAP7_75t_L g8331 ( 
.A(n_7446),
.B(n_790),
.Y(n_8331)
);

INVx1_ASAP7_75t_L g8332 ( 
.A(n_7320),
.Y(n_8332)
);

NAND2xp5_ASAP7_75t_L g8333 ( 
.A(n_7446),
.B(n_226),
.Y(n_8333)
);

INVx3_ASAP7_75t_L g8334 ( 
.A(n_7312),
.Y(n_8334)
);

AOI21xp5_ASAP7_75t_L g8335 ( 
.A1(n_7446),
.A2(n_792),
.B(n_791),
.Y(n_8335)
);

INVx2_ASAP7_75t_L g8336 ( 
.A(n_7320),
.Y(n_8336)
);

INVx3_ASAP7_75t_L g8337 ( 
.A(n_7312),
.Y(n_8337)
);

A2O1A1Ixp33_ASAP7_75t_L g8338 ( 
.A1(n_7976),
.A2(n_792),
.B(n_793),
.C(n_791),
.Y(n_8338)
);

INVx2_ASAP7_75t_SL g8339 ( 
.A(n_7864),
.Y(n_8339)
);

CKINVDCx20_ASAP7_75t_R g8340 ( 
.A(n_7940),
.Y(n_8340)
);

OAI21xp5_ASAP7_75t_L g8341 ( 
.A1(n_7981),
.A2(n_227),
.B(n_228),
.Y(n_8341)
);

OR2x6_ASAP7_75t_SL g8342 ( 
.A(n_8238),
.B(n_8093),
.Y(n_8342)
);

NAND2xp5_ASAP7_75t_L g8343 ( 
.A(n_7907),
.B(n_7953),
.Y(n_8343)
);

AND2x2_ASAP7_75t_L g8344 ( 
.A(n_7877),
.B(n_793),
.Y(n_8344)
);

INVx2_ASAP7_75t_L g8345 ( 
.A(n_7813),
.Y(n_8345)
);

NAND2xp5_ASAP7_75t_L g8346 ( 
.A(n_7930),
.B(n_794),
.Y(n_8346)
);

AOI21xp5_ASAP7_75t_L g8347 ( 
.A1(n_7881),
.A2(n_796),
.B(n_795),
.Y(n_8347)
);

NOR2xp33_ASAP7_75t_L g8348 ( 
.A(n_7863),
.B(n_795),
.Y(n_8348)
);

AOI21xp5_ASAP7_75t_L g8349 ( 
.A1(n_7869),
.A2(n_797),
.B(n_796),
.Y(n_8349)
);

NOR2xp33_ASAP7_75t_L g8350 ( 
.A(n_8045),
.B(n_797),
.Y(n_8350)
);

INVx1_ASAP7_75t_L g8351 ( 
.A(n_7871),
.Y(n_8351)
);

NOR2xp33_ASAP7_75t_L g8352 ( 
.A(n_8259),
.B(n_798),
.Y(n_8352)
);

AOI21xp5_ASAP7_75t_L g8353 ( 
.A1(n_7824),
.A2(n_799),
.B(n_798),
.Y(n_8353)
);

NAND3xp33_ASAP7_75t_L g8354 ( 
.A(n_7830),
.B(n_228),
.C(n_229),
.Y(n_8354)
);

HB1xp67_ASAP7_75t_L g8355 ( 
.A(n_8037),
.Y(n_8355)
);

NAND2xp5_ASAP7_75t_SL g8356 ( 
.A(n_7866),
.B(n_799),
.Y(n_8356)
);

NOR2xp33_ASAP7_75t_R g8357 ( 
.A(n_8302),
.B(n_229),
.Y(n_8357)
);

OAI21x1_ASAP7_75t_L g8358 ( 
.A1(n_8066),
.A2(n_229),
.B(n_230),
.Y(n_8358)
);

OAI22x1_ASAP7_75t_L g8359 ( 
.A1(n_7843),
.A2(n_232),
.B1(n_230),
.B2(n_231),
.Y(n_8359)
);

BUFx3_ASAP7_75t_L g8360 ( 
.A(n_8026),
.Y(n_8360)
);

A2O1A1Ixp33_ASAP7_75t_L g8361 ( 
.A1(n_7936),
.A2(n_801),
.B(n_802),
.C(n_800),
.Y(n_8361)
);

BUFx6f_ASAP7_75t_L g8362 ( 
.A(n_7817),
.Y(n_8362)
);

AOI21xp5_ASAP7_75t_L g8363 ( 
.A1(n_7810),
.A2(n_801),
.B(n_800),
.Y(n_8363)
);

CKINVDCx20_ASAP7_75t_R g8364 ( 
.A(n_8306),
.Y(n_8364)
);

OAI22xp5_ASAP7_75t_L g8365 ( 
.A1(n_8253),
.A2(n_233),
.B1(n_231),
.B2(n_232),
.Y(n_8365)
);

AOI21xp5_ASAP7_75t_L g8366 ( 
.A1(n_7854),
.A2(n_804),
.B(n_803),
.Y(n_8366)
);

INVx1_ASAP7_75t_L g8367 ( 
.A(n_7929),
.Y(n_8367)
);

AOI22xp33_ASAP7_75t_L g8368 ( 
.A1(n_8100),
.A2(n_233),
.B1(n_231),
.B2(n_232),
.Y(n_8368)
);

NAND2xp5_ASAP7_75t_SL g8369 ( 
.A(n_7897),
.B(n_804),
.Y(n_8369)
);

BUFx2_ASAP7_75t_L g8370 ( 
.A(n_8294),
.Y(n_8370)
);

AOI22xp33_ASAP7_75t_L g8371 ( 
.A1(n_8091),
.A2(n_236),
.B1(n_234),
.B2(n_235),
.Y(n_8371)
);

NOR2xp33_ASAP7_75t_L g8372 ( 
.A(n_8308),
.B(n_805),
.Y(n_8372)
);

NAND2xp5_ASAP7_75t_L g8373 ( 
.A(n_7898),
.B(n_805),
.Y(n_8373)
);

O2A1O1Ixp33_ASAP7_75t_L g8374 ( 
.A1(n_8128),
.A2(n_236),
.B(n_234),
.C(n_235),
.Y(n_8374)
);

INVx1_ASAP7_75t_L g8375 ( 
.A(n_7956),
.Y(n_8375)
);

AOI22xp5_ASAP7_75t_L g8376 ( 
.A1(n_8255),
.A2(n_237),
.B1(n_235),
.B2(n_236),
.Y(n_8376)
);

INVx1_ASAP7_75t_L g8377 ( 
.A(n_7975),
.Y(n_8377)
);

CKINVDCx5p33_ASAP7_75t_R g8378 ( 
.A(n_8084),
.Y(n_8378)
);

NAND3xp33_ASAP7_75t_SL g8379 ( 
.A(n_7853),
.B(n_237),
.C(n_238),
.Y(n_8379)
);

INVx1_ASAP7_75t_L g8380 ( 
.A(n_7994),
.Y(n_8380)
);

O2A1O1Ixp5_ASAP7_75t_L g8381 ( 
.A1(n_7822),
.A2(n_8056),
.B(n_8065),
.C(n_7939),
.Y(n_8381)
);

NOR2xp33_ASAP7_75t_SL g8382 ( 
.A(n_7997),
.B(n_238),
.Y(n_8382)
);

NAND2xp5_ASAP7_75t_SL g8383 ( 
.A(n_7902),
.B(n_806),
.Y(n_8383)
);

AOI22x1_ASAP7_75t_SL g8384 ( 
.A1(n_8208),
.A2(n_241),
.B1(n_239),
.B2(n_240),
.Y(n_8384)
);

NAND2xp5_ASAP7_75t_SL g8385 ( 
.A(n_7811),
.B(n_7809),
.Y(n_8385)
);

INVx4_ASAP7_75t_L g8386 ( 
.A(n_7864),
.Y(n_8386)
);

HB1xp67_ASAP7_75t_L g8387 ( 
.A(n_7872),
.Y(n_8387)
);

BUFx3_ASAP7_75t_L g8388 ( 
.A(n_8075),
.Y(n_8388)
);

O2A1O1Ixp33_ASAP7_75t_L g8389 ( 
.A1(n_8258),
.A2(n_241),
.B(n_239),
.C(n_240),
.Y(n_8389)
);

NAND2xp5_ASAP7_75t_L g8390 ( 
.A(n_7882),
.B(n_807),
.Y(n_8390)
);

INVx4_ASAP7_75t_L g8391 ( 
.A(n_7864),
.Y(n_8391)
);

NOR2xp33_ASAP7_75t_L g8392 ( 
.A(n_8146),
.B(n_808),
.Y(n_8392)
);

OAI22xp5_ASAP7_75t_L g8393 ( 
.A1(n_8276),
.A2(n_243),
.B1(n_240),
.B2(n_242),
.Y(n_8393)
);

BUFx6f_ASAP7_75t_L g8394 ( 
.A(n_7817),
.Y(n_8394)
);

AOI21xp5_ASAP7_75t_L g8395 ( 
.A1(n_7837),
.A2(n_809),
.B(n_808),
.Y(n_8395)
);

INVx2_ASAP7_75t_L g8396 ( 
.A(n_7856),
.Y(n_8396)
);

NAND2xp5_ASAP7_75t_SL g8397 ( 
.A(n_8201),
.B(n_809),
.Y(n_8397)
);

NOR2xp67_ASAP7_75t_SL g8398 ( 
.A(n_7857),
.B(n_242),
.Y(n_8398)
);

A2O1A1Ixp33_ASAP7_75t_L g8399 ( 
.A1(n_8008),
.A2(n_811),
.B(n_812),
.C(n_810),
.Y(n_8399)
);

BUFx6f_ASAP7_75t_L g8400 ( 
.A(n_7817),
.Y(n_8400)
);

INVx1_ASAP7_75t_L g8401 ( 
.A(n_8002),
.Y(n_8401)
);

AND2x4_ASAP7_75t_L g8402 ( 
.A(n_7849),
.B(n_810),
.Y(n_8402)
);

AOI22xp5_ASAP7_75t_L g8403 ( 
.A1(n_8287),
.A2(n_244),
.B1(n_242),
.B2(n_243),
.Y(n_8403)
);

INVx1_ASAP7_75t_L g8404 ( 
.A(n_8007),
.Y(n_8404)
);

NOR2xp33_ASAP7_75t_L g8405 ( 
.A(n_8016),
.B(n_812),
.Y(n_8405)
);

NAND2xp5_ASAP7_75t_L g8406 ( 
.A(n_7922),
.B(n_8096),
.Y(n_8406)
);

NOR2xp33_ASAP7_75t_L g8407 ( 
.A(n_8067),
.B(n_813),
.Y(n_8407)
);

OAI22xp5_ASAP7_75t_L g8408 ( 
.A1(n_8290),
.A2(n_245),
.B1(n_243),
.B2(n_244),
.Y(n_8408)
);

BUFx2_ASAP7_75t_L g8409 ( 
.A(n_8303),
.Y(n_8409)
);

INVx2_ASAP7_75t_L g8410 ( 
.A(n_7860),
.Y(n_8410)
);

OAI21x1_ASAP7_75t_L g8411 ( 
.A1(n_7834),
.A2(n_245),
.B(n_246),
.Y(n_8411)
);

NAND2xp5_ASAP7_75t_SL g8412 ( 
.A(n_8256),
.B(n_813),
.Y(n_8412)
);

NOR2xp33_ASAP7_75t_L g8413 ( 
.A(n_8224),
.B(n_814),
.Y(n_8413)
);

NAND2xp5_ASAP7_75t_L g8414 ( 
.A(n_7998),
.B(n_814),
.Y(n_8414)
);

NAND2xp5_ASAP7_75t_L g8415 ( 
.A(n_7920),
.B(n_815),
.Y(n_8415)
);

AOI21x1_ASAP7_75t_L g8416 ( 
.A1(n_8033),
.A2(n_245),
.B(n_246),
.Y(n_8416)
);

INVx1_ASAP7_75t_SL g8417 ( 
.A(n_8136),
.Y(n_8417)
);

INVx3_ASAP7_75t_L g8418 ( 
.A(n_7814),
.Y(n_8418)
);

HB1xp67_ASAP7_75t_L g8419 ( 
.A(n_8198),
.Y(n_8419)
);

INVx1_ASAP7_75t_L g8420 ( 
.A(n_8014),
.Y(n_8420)
);

INVx1_ASAP7_75t_L g8421 ( 
.A(n_8027),
.Y(n_8421)
);

AOI21xp5_ASAP7_75t_L g8422 ( 
.A1(n_7828),
.A2(n_817),
.B(n_816),
.Y(n_8422)
);

AOI22xp5_ASAP7_75t_L g8423 ( 
.A1(n_8331),
.A2(n_8180),
.B1(n_7966),
.B2(n_8291),
.Y(n_8423)
);

AOI21xp5_ASAP7_75t_L g8424 ( 
.A1(n_7848),
.A2(n_817),
.B(n_816),
.Y(n_8424)
);

AOI22xp5_ASAP7_75t_L g8425 ( 
.A1(n_7833),
.A2(n_248),
.B1(n_246),
.B2(n_247),
.Y(n_8425)
);

INVx1_ASAP7_75t_SL g8426 ( 
.A(n_8006),
.Y(n_8426)
);

AOI21xp5_ASAP7_75t_L g8427 ( 
.A1(n_7867),
.A2(n_819),
.B(n_818),
.Y(n_8427)
);

AOI33xp33_ASAP7_75t_L g8428 ( 
.A1(n_8149),
.A2(n_249),
.A3(n_251),
.B1(n_247),
.B2(n_248),
.B3(n_250),
.Y(n_8428)
);

BUFx2_ASAP7_75t_L g8429 ( 
.A(n_8098),
.Y(n_8429)
);

AND2x2_ASAP7_75t_L g8430 ( 
.A(n_8010),
.B(n_7937),
.Y(n_8430)
);

AOI21xp5_ASAP7_75t_L g8431 ( 
.A1(n_8119),
.A2(n_820),
.B(n_819),
.Y(n_8431)
);

INVx2_ASAP7_75t_L g8432 ( 
.A(n_8249),
.Y(n_8432)
);

BUFx2_ASAP7_75t_L g8433 ( 
.A(n_8102),
.Y(n_8433)
);

INVx4_ASAP7_75t_L g8434 ( 
.A(n_7970),
.Y(n_8434)
);

OAI22xp5_ASAP7_75t_L g8435 ( 
.A1(n_8257),
.A2(n_8265),
.B1(n_8268),
.B2(n_8262),
.Y(n_8435)
);

OR2x6_ASAP7_75t_L g8436 ( 
.A(n_7959),
.B(n_821),
.Y(n_8436)
);

INVx1_ASAP7_75t_L g8437 ( 
.A(n_8042),
.Y(n_8437)
);

AOI21xp5_ASAP7_75t_L g8438 ( 
.A1(n_8147),
.A2(n_822),
.B(n_821),
.Y(n_8438)
);

O2A1O1Ixp33_ASAP7_75t_L g8439 ( 
.A1(n_7890),
.A2(n_250),
.B(n_248),
.C(n_249),
.Y(n_8439)
);

O2A1O1Ixp33_ASAP7_75t_L g8440 ( 
.A1(n_8274),
.A2(n_252),
.B(n_249),
.C(n_251),
.Y(n_8440)
);

NAND2xp5_ASAP7_75t_L g8441 ( 
.A(n_8029),
.B(n_822),
.Y(n_8441)
);

INVx1_ASAP7_75t_L g8442 ( 
.A(n_8076),
.Y(n_8442)
);

OR2x6_ASAP7_75t_SL g8443 ( 
.A(n_8157),
.B(n_252),
.Y(n_8443)
);

NAND2xp5_ASAP7_75t_L g8444 ( 
.A(n_8000),
.B(n_823),
.Y(n_8444)
);

NAND2xp5_ASAP7_75t_L g8445 ( 
.A(n_7947),
.B(n_7963),
.Y(n_8445)
);

INVx1_ASAP7_75t_L g8446 ( 
.A(n_8086),
.Y(n_8446)
);

INVx1_ASAP7_75t_L g8447 ( 
.A(n_8092),
.Y(n_8447)
);

NAND2xp5_ASAP7_75t_L g8448 ( 
.A(n_7969),
.B(n_823),
.Y(n_8448)
);

INVx1_ASAP7_75t_L g8449 ( 
.A(n_8118),
.Y(n_8449)
);

BUFx6f_ASAP7_75t_L g8450 ( 
.A(n_7851),
.Y(n_8450)
);

NOR3xp33_ASAP7_75t_SL g8451 ( 
.A(n_8172),
.B(n_252),
.C(n_253),
.Y(n_8451)
);

NAND2xp5_ASAP7_75t_SL g8452 ( 
.A(n_7916),
.B(n_824),
.Y(n_8452)
);

O2A1O1Ixp33_ASAP7_75t_L g8453 ( 
.A1(n_8052),
.A2(n_8326),
.B(n_7934),
.C(n_8032),
.Y(n_8453)
);

OAI22xp5_ASAP7_75t_L g8454 ( 
.A1(n_8278),
.A2(n_255),
.B1(n_253),
.B2(n_254),
.Y(n_8454)
);

NAND2xp5_ASAP7_75t_SL g8455 ( 
.A(n_7879),
.B(n_825),
.Y(n_8455)
);

NAND2xp5_ASAP7_75t_L g8456 ( 
.A(n_7979),
.B(n_7986),
.Y(n_8456)
);

AOI21xp5_ASAP7_75t_L g8457 ( 
.A1(n_8060),
.A2(n_826),
.B(n_825),
.Y(n_8457)
);

OAI21xp33_ASAP7_75t_L g8458 ( 
.A1(n_7996),
.A2(n_253),
.B(n_254),
.Y(n_8458)
);

CKINVDCx5p33_ASAP7_75t_R g8459 ( 
.A(n_7973),
.Y(n_8459)
);

BUFx6f_ASAP7_75t_L g8460 ( 
.A(n_7851),
.Y(n_8460)
);

AOI21xp5_ASAP7_75t_L g8461 ( 
.A1(n_7999),
.A2(n_828),
.B(n_827),
.Y(n_8461)
);

NAND2xp5_ASAP7_75t_SL g8462 ( 
.A(n_8281),
.B(n_8299),
.Y(n_8462)
);

A2O1A1Ixp33_ASAP7_75t_L g8463 ( 
.A1(n_8104),
.A2(n_828),
.B(n_829),
.C(n_827),
.Y(n_8463)
);

AOI33xp33_ASAP7_75t_L g8464 ( 
.A1(n_8179),
.A2(n_256),
.A3(n_258),
.B1(n_254),
.B2(n_255),
.B3(n_257),
.Y(n_8464)
);

AO21x1_ASAP7_75t_L g8465 ( 
.A1(n_8162),
.A2(n_255),
.B(n_256),
.Y(n_8465)
);

NAND2xp5_ASAP7_75t_SL g8466 ( 
.A(n_8318),
.B(n_829),
.Y(n_8466)
);

BUFx8_ASAP7_75t_L g8467 ( 
.A(n_8240),
.Y(n_8467)
);

AOI21x1_ASAP7_75t_L g8468 ( 
.A1(n_8280),
.A2(n_257),
.B(n_258),
.Y(n_8468)
);

AOI21xp5_ASAP7_75t_L g8469 ( 
.A1(n_8155),
.A2(n_832),
.B(n_831),
.Y(n_8469)
);

INVx4_ASAP7_75t_L g8470 ( 
.A(n_7851),
.Y(n_8470)
);

NOR2xp67_ASAP7_75t_L g8471 ( 
.A(n_7906),
.B(n_257),
.Y(n_8471)
);

OR2x6_ASAP7_75t_L g8472 ( 
.A(n_8047),
.B(n_831),
.Y(n_8472)
);

O2A1O1Ixp33_ASAP7_75t_L g8473 ( 
.A1(n_8139),
.A2(n_260),
.B(n_258),
.C(n_259),
.Y(n_8473)
);

NAND2xp5_ASAP7_75t_L g8474 ( 
.A(n_8054),
.B(n_833),
.Y(n_8474)
);

NAND2xp5_ASAP7_75t_L g8475 ( 
.A(n_8200),
.B(n_833),
.Y(n_8475)
);

AOI22xp5_ASAP7_75t_L g8476 ( 
.A1(n_7991),
.A2(n_261),
.B1(n_259),
.B2(n_260),
.Y(n_8476)
);

BUFx6f_ASAP7_75t_L g8477 ( 
.A(n_8250),
.Y(n_8477)
);

NOR2xp33_ASAP7_75t_L g8478 ( 
.A(n_8099),
.B(n_835),
.Y(n_8478)
);

AOI21xp5_ASAP7_75t_L g8479 ( 
.A1(n_8063),
.A2(n_836),
.B(n_835),
.Y(n_8479)
);

NAND2xp5_ASAP7_75t_SL g8480 ( 
.A(n_8319),
.B(n_836),
.Y(n_8480)
);

INVx2_ASAP7_75t_L g8481 ( 
.A(n_8267),
.Y(n_8481)
);

AOI21xp5_ASAP7_75t_L g8482 ( 
.A1(n_7988),
.A2(n_838),
.B(n_837),
.Y(n_8482)
);

BUFx6f_ASAP7_75t_L g8483 ( 
.A(n_8250),
.Y(n_8483)
);

O2A1O1Ixp33_ASAP7_75t_L g8484 ( 
.A1(n_8305),
.A2(n_262),
.B(n_260),
.C(n_261),
.Y(n_8484)
);

AOI21xp5_ASAP7_75t_L g8485 ( 
.A1(n_7899),
.A2(n_8181),
.B(n_8058),
.Y(n_8485)
);

AOI21xp5_ASAP7_75t_L g8486 ( 
.A1(n_7825),
.A2(n_839),
.B(n_837),
.Y(n_8486)
);

AOI21xp5_ASAP7_75t_L g8487 ( 
.A1(n_8025),
.A2(n_841),
.B(n_840),
.Y(n_8487)
);

NOR2xp33_ASAP7_75t_L g8488 ( 
.A(n_7875),
.B(n_840),
.Y(n_8488)
);

NAND2xp5_ASAP7_75t_SL g8489 ( 
.A(n_8320),
.B(n_842),
.Y(n_8489)
);

INVx2_ASAP7_75t_L g8490 ( 
.A(n_8292),
.Y(n_8490)
);

INVx2_ASAP7_75t_L g8491 ( 
.A(n_8309),
.Y(n_8491)
);

AND2x2_ASAP7_75t_L g8492 ( 
.A(n_7818),
.B(n_842),
.Y(n_8492)
);

AOI21xp5_ASAP7_75t_L g8493 ( 
.A1(n_8064),
.A2(n_844),
.B(n_843),
.Y(n_8493)
);

AOI21xp5_ASAP7_75t_L g8494 ( 
.A1(n_8064),
.A2(n_844),
.B(n_843),
.Y(n_8494)
);

AND2x2_ASAP7_75t_SL g8495 ( 
.A(n_8030),
.B(n_845),
.Y(n_8495)
);

AND2x4_ASAP7_75t_L g8496 ( 
.A(n_8273),
.B(n_845),
.Y(n_8496)
);

O2A1O1Ixp33_ASAP7_75t_L g8497 ( 
.A1(n_8062),
.A2(n_263),
.B(n_261),
.C(n_262),
.Y(n_8497)
);

NAND2xp5_ASAP7_75t_L g8498 ( 
.A(n_8314),
.B(n_846),
.Y(n_8498)
);

AND2x2_ASAP7_75t_L g8499 ( 
.A(n_8097),
.B(n_846),
.Y(n_8499)
);

NAND2xp5_ASAP7_75t_L g8500 ( 
.A(n_8325),
.B(n_847),
.Y(n_8500)
);

NOR2xp33_ASAP7_75t_L g8501 ( 
.A(n_8322),
.B(n_847),
.Y(n_8501)
);

NAND2xp5_ASAP7_75t_L g8502 ( 
.A(n_8327),
.B(n_848),
.Y(n_8502)
);

O2A1O1Ixp33_ASAP7_75t_L g8503 ( 
.A1(n_8282),
.A2(n_264),
.B(n_262),
.C(n_263),
.Y(n_8503)
);

NOR2xp33_ASAP7_75t_L g8504 ( 
.A(n_8333),
.B(n_848),
.Y(n_8504)
);

AOI22xp5_ASAP7_75t_L g8505 ( 
.A1(n_8017),
.A2(n_265),
.B1(n_263),
.B2(n_264),
.Y(n_8505)
);

INVx4_ASAP7_75t_L g8506 ( 
.A(n_8250),
.Y(n_8506)
);

AOI22xp5_ASAP7_75t_L g8507 ( 
.A1(n_7949),
.A2(n_266),
.B1(n_264),
.B2(n_265),
.Y(n_8507)
);

BUFx2_ASAP7_75t_L g8508 ( 
.A(n_8145),
.Y(n_8508)
);

NOR2xp33_ASAP7_75t_R g8509 ( 
.A(n_8113),
.B(n_265),
.Y(n_8509)
);

NOR2xp33_ASAP7_75t_L g8510 ( 
.A(n_7912),
.B(n_7886),
.Y(n_8510)
);

AOI21xp5_ASAP7_75t_L g8511 ( 
.A1(n_7938),
.A2(n_851),
.B(n_850),
.Y(n_8511)
);

HB1xp67_ASAP7_75t_L g8512 ( 
.A(n_8046),
.Y(n_8512)
);

OAI21xp5_ASAP7_75t_L g8513 ( 
.A1(n_8021),
.A2(n_266),
.B(n_267),
.Y(n_8513)
);

AOI21xp5_ASAP7_75t_L g8514 ( 
.A1(n_8261),
.A2(n_852),
.B(n_851),
.Y(n_8514)
);

NOR2xp67_ASAP7_75t_L g8515 ( 
.A(n_7915),
.B(n_266),
.Y(n_8515)
);

NAND2xp5_ASAP7_75t_L g8516 ( 
.A(n_8336),
.B(n_853),
.Y(n_8516)
);

OA21x2_ASAP7_75t_L g8517 ( 
.A1(n_7932),
.A2(n_7942),
.B(n_7944),
.Y(n_8517)
);

NOR2xp33_ASAP7_75t_L g8518 ( 
.A(n_8191),
.B(n_853),
.Y(n_8518)
);

NAND2xp5_ASAP7_75t_L g8519 ( 
.A(n_8163),
.B(n_854),
.Y(n_8519)
);

INVx4_ASAP7_75t_L g8520 ( 
.A(n_8297),
.Y(n_8520)
);

AOI21xp5_ASAP7_75t_L g8521 ( 
.A1(n_8324),
.A2(n_856),
.B(n_855),
.Y(n_8521)
);

NAND2xp5_ASAP7_75t_L g8522 ( 
.A(n_7835),
.B(n_855),
.Y(n_8522)
);

O2A1O1Ixp33_ASAP7_75t_L g8523 ( 
.A1(n_8289),
.A2(n_269),
.B(n_267),
.C(n_268),
.Y(n_8523)
);

INVx2_ASAP7_75t_L g8524 ( 
.A(n_8135),
.Y(n_8524)
);

OR2x2_ASAP7_75t_L g8525 ( 
.A(n_8217),
.B(n_856),
.Y(n_8525)
);

INVx1_ASAP7_75t_L g8526 ( 
.A(n_8151),
.Y(n_8526)
);

OAI22xp5_ASAP7_75t_L g8527 ( 
.A1(n_7844),
.A2(n_270),
.B1(n_267),
.B2(n_268),
.Y(n_8527)
);

AOI21xp5_ASAP7_75t_L g8528 ( 
.A1(n_8089),
.A2(n_858),
.B(n_857),
.Y(n_8528)
);

AOI21xp5_ASAP7_75t_L g8529 ( 
.A1(n_8108),
.A2(n_858),
.B(n_857),
.Y(n_8529)
);

CKINVDCx20_ASAP7_75t_R g8530 ( 
.A(n_8212),
.Y(n_8530)
);

OAI22x1_ASAP7_75t_L g8531 ( 
.A1(n_8242),
.A2(n_272),
.B1(n_270),
.B2(n_271),
.Y(n_8531)
);

AND2x2_ASAP7_75t_L g8532 ( 
.A(n_8137),
.B(n_859),
.Y(n_8532)
);

NAND2xp5_ASAP7_75t_L g8533 ( 
.A(n_7840),
.B(n_859),
.Y(n_8533)
);

NAND2xp5_ASAP7_75t_L g8534 ( 
.A(n_7841),
.B(n_860),
.Y(n_8534)
);

BUFx6f_ASAP7_75t_L g8535 ( 
.A(n_8297),
.Y(n_8535)
);

AND2x4_ASAP7_75t_SL g8536 ( 
.A(n_7814),
.B(n_8248),
.Y(n_8536)
);

INVx1_ASAP7_75t_L g8537 ( 
.A(n_8165),
.Y(n_8537)
);

INVx2_ASAP7_75t_L g8538 ( 
.A(n_8116),
.Y(n_8538)
);

O2A1O1Ixp33_ASAP7_75t_L g8539 ( 
.A1(n_8300),
.A2(n_8301),
.B(n_8049),
.C(n_7943),
.Y(n_8539)
);

NOR2xp67_ASAP7_75t_L g8540 ( 
.A(n_8271),
.B(n_271),
.Y(n_8540)
);

A2O1A1Ixp33_ASAP7_75t_L g8541 ( 
.A1(n_8251),
.A2(n_862),
.B(n_863),
.C(n_861),
.Y(n_8541)
);

OAI22xp5_ASAP7_75t_L g8542 ( 
.A1(n_8206),
.A2(n_274),
.B1(n_272),
.B2(n_273),
.Y(n_8542)
);

O2A1O1Ixp33_ASAP7_75t_SL g8543 ( 
.A1(n_7945),
.A2(n_7971),
.B(n_7977),
.C(n_7962),
.Y(n_8543)
);

INVx1_ASAP7_75t_L g8544 ( 
.A(n_8178),
.Y(n_8544)
);

NAND2xp5_ASAP7_75t_L g8545 ( 
.A(n_7850),
.B(n_8266),
.Y(n_8545)
);

NOR2xp33_ASAP7_75t_L g8546 ( 
.A(n_8022),
.B(n_862),
.Y(n_8546)
);

AOI21x1_ASAP7_75t_L g8547 ( 
.A1(n_8295),
.A2(n_272),
.B(n_273),
.Y(n_8547)
);

OAI22xp5_ASAP7_75t_L g8548 ( 
.A1(n_8170),
.A2(n_275),
.B1(n_273),
.B2(n_274),
.Y(n_8548)
);

BUFx2_ASAP7_75t_L g8549 ( 
.A(n_8168),
.Y(n_8549)
);

BUFx2_ASAP7_75t_R g8550 ( 
.A(n_8221),
.Y(n_8550)
);

NOR2xp33_ASAP7_75t_L g8551 ( 
.A(n_8085),
.B(n_863),
.Y(n_8551)
);

INVx2_ASAP7_75t_L g8552 ( 
.A(n_8188),
.Y(n_8552)
);

OAI22x1_ASAP7_75t_L g8553 ( 
.A1(n_8038),
.A2(n_276),
.B1(n_274),
.B2(n_275),
.Y(n_8553)
);

NOR2xp33_ASAP7_75t_L g8554 ( 
.A(n_8334),
.B(n_864),
.Y(n_8554)
);

CKINVDCx20_ASAP7_75t_R g8555 ( 
.A(n_7989),
.Y(n_8555)
);

INVx1_ASAP7_75t_SL g8556 ( 
.A(n_8337),
.Y(n_8556)
);

INVx1_ASAP7_75t_L g8557 ( 
.A(n_8185),
.Y(n_8557)
);

INVx4_ASAP7_75t_L g8558 ( 
.A(n_8297),
.Y(n_8558)
);

INVx2_ASAP7_75t_L g8559 ( 
.A(n_7868),
.Y(n_8559)
);

NOR2xp33_ASAP7_75t_SL g8560 ( 
.A(n_8088),
.B(n_275),
.Y(n_8560)
);

NAND2xp5_ASAP7_75t_L g8561 ( 
.A(n_8272),
.B(n_865),
.Y(n_8561)
);

BUFx6f_ASAP7_75t_L g8562 ( 
.A(n_7946),
.Y(n_8562)
);

INVx2_ASAP7_75t_SL g8563 ( 
.A(n_7946),
.Y(n_8563)
);

INVx1_ASAP7_75t_L g8564 ( 
.A(n_8121),
.Y(n_8564)
);

INVx3_ASAP7_75t_L g8565 ( 
.A(n_8176),
.Y(n_8565)
);

OAI21xp33_ASAP7_75t_SL g8566 ( 
.A1(n_8237),
.A2(n_867),
.B(n_866),
.Y(n_8566)
);

NOR2xp33_ASAP7_75t_L g8567 ( 
.A(n_7873),
.B(n_866),
.Y(n_8567)
);

OAI22xp5_ASAP7_75t_L g8568 ( 
.A1(n_8154),
.A2(n_278),
.B1(n_276),
.B2(n_277),
.Y(n_8568)
);

OR2x6_ASAP7_75t_L g8569 ( 
.A(n_7964),
.B(n_867),
.Y(n_8569)
);

HB1xp67_ASAP7_75t_L g8570 ( 
.A(n_8310),
.Y(n_8570)
);

NOR2xp33_ASAP7_75t_L g8571 ( 
.A(n_7908),
.B(n_868),
.Y(n_8571)
);

AOI21xp5_ASAP7_75t_L g8572 ( 
.A1(n_7838),
.A2(n_869),
.B(n_868),
.Y(n_8572)
);

A2O1A1Ixp33_ASAP7_75t_L g8573 ( 
.A1(n_8252),
.A2(n_871),
.B(n_872),
.C(n_870),
.Y(n_8573)
);

BUFx6f_ASAP7_75t_L g8574 ( 
.A(n_7946),
.Y(n_8574)
);

O2A1O1Ixp33_ASAP7_75t_L g8575 ( 
.A1(n_7819),
.A2(n_279),
.B(n_277),
.C(n_278),
.Y(n_8575)
);

OAI21x1_ASAP7_75t_L g8576 ( 
.A1(n_8009),
.A2(n_278),
.B(n_279),
.Y(n_8576)
);

INVx4_ASAP7_75t_L g8577 ( 
.A(n_7883),
.Y(n_8577)
);

NOR3xp33_ASAP7_75t_SL g8578 ( 
.A(n_8107),
.B(n_279),
.C(n_280),
.Y(n_8578)
);

OA22x2_ASAP7_75t_L g8579 ( 
.A1(n_7941),
.A2(n_282),
.B1(n_280),
.B2(n_281),
.Y(n_8579)
);

INVx2_ASAP7_75t_L g8580 ( 
.A(n_7933),
.Y(n_8580)
);

A2O1A1Ixp33_ASAP7_75t_L g8581 ( 
.A1(n_8254),
.A2(n_871),
.B(n_872),
.C(n_870),
.Y(n_8581)
);

O2A1O1Ixp33_ASAP7_75t_L g8582 ( 
.A1(n_7836),
.A2(n_282),
.B(n_280),
.C(n_281),
.Y(n_8582)
);

INVx1_ASAP7_75t_L g8583 ( 
.A(n_8125),
.Y(n_8583)
);

NAND2xp5_ASAP7_75t_SL g8584 ( 
.A(n_7992),
.B(n_873),
.Y(n_8584)
);

INVx2_ASAP7_75t_L g8585 ( 
.A(n_7950),
.Y(n_8585)
);

NAND2xp5_ASAP7_75t_L g8586 ( 
.A(n_8311),
.B(n_873),
.Y(n_8586)
);

AND2x4_ASAP7_75t_L g8587 ( 
.A(n_7888),
.B(n_874),
.Y(n_8587)
);

NAND2xp5_ASAP7_75t_SL g8588 ( 
.A(n_7893),
.B(n_874),
.Y(n_8588)
);

INVx3_ASAP7_75t_L g8589 ( 
.A(n_7909),
.Y(n_8589)
);

NAND2xp5_ASAP7_75t_L g8590 ( 
.A(n_8316),
.B(n_875),
.Y(n_8590)
);

BUFx6f_ASAP7_75t_L g8591 ( 
.A(n_7815),
.Y(n_8591)
);

OAI22xp5_ASAP7_75t_L g8592 ( 
.A1(n_7914),
.A2(n_284),
.B1(n_282),
.B2(n_283),
.Y(n_8592)
);

NOR2xp33_ASAP7_75t_L g8593 ( 
.A(n_8111),
.B(n_8034),
.Y(n_8593)
);

NOR2xp33_ASAP7_75t_L g8594 ( 
.A(n_8050),
.B(n_875),
.Y(n_8594)
);

HB1xp67_ASAP7_75t_L g8595 ( 
.A(n_8321),
.Y(n_8595)
);

NOR2xp33_ASAP7_75t_L g8596 ( 
.A(n_7894),
.B(n_876),
.Y(n_8596)
);

NAND2xp5_ASAP7_75t_L g8597 ( 
.A(n_8323),
.B(n_877),
.Y(n_8597)
);

AOI21xp5_ASAP7_75t_L g8598 ( 
.A1(n_7820),
.A2(n_879),
.B(n_877),
.Y(n_8598)
);

AO21x1_ASAP7_75t_L g8599 ( 
.A1(n_8228),
.A2(n_283),
.B(n_284),
.Y(n_8599)
);

BUFx6f_ASAP7_75t_L g8600 ( 
.A(n_8246),
.Y(n_8600)
);

AOI21xp5_ASAP7_75t_L g8601 ( 
.A1(n_8164),
.A2(n_881),
.B(n_880),
.Y(n_8601)
);

INVx1_ASAP7_75t_SL g8602 ( 
.A(n_7921),
.Y(n_8602)
);

NAND2xp5_ASAP7_75t_SL g8603 ( 
.A(n_8169),
.B(n_8051),
.Y(n_8603)
);

OAI21xp33_ASAP7_75t_SL g8604 ( 
.A1(n_8296),
.A2(n_881),
.B(n_880),
.Y(n_8604)
);

OAI22xp5_ASAP7_75t_L g8605 ( 
.A1(n_8317),
.A2(n_285),
.B1(n_283),
.B2(n_284),
.Y(n_8605)
);

NAND2xp5_ASAP7_75t_L g8606 ( 
.A(n_8332),
.B(n_882),
.Y(n_8606)
);

O2A1O1Ixp5_ASAP7_75t_L g8607 ( 
.A1(n_8304),
.A2(n_287),
.B(n_285),
.C(n_286),
.Y(n_8607)
);

OAI22x1_ASAP7_75t_L g8608 ( 
.A1(n_7987),
.A2(n_287),
.B1(n_285),
.B2(n_286),
.Y(n_8608)
);

O2A1O1Ixp33_ASAP7_75t_L g8609 ( 
.A1(n_7852),
.A2(n_288),
.B(n_286),
.C(n_287),
.Y(n_8609)
);

O2A1O1Ixp33_ASAP7_75t_L g8610 ( 
.A1(n_7876),
.A2(n_291),
.B(n_289),
.C(n_290),
.Y(n_8610)
);

A2O1A1Ixp33_ASAP7_75t_L g8611 ( 
.A1(n_8260),
.A2(n_8269),
.B(n_8270),
.C(n_8264),
.Y(n_8611)
);

NAND2xp5_ASAP7_75t_SL g8612 ( 
.A(n_7901),
.B(n_7910),
.Y(n_8612)
);

NAND2xp5_ASAP7_75t_SL g8613 ( 
.A(n_7954),
.B(n_883),
.Y(n_8613)
);

AND2x2_ASAP7_75t_L g8614 ( 
.A(n_7821),
.B(n_883),
.Y(n_8614)
);

NOR2xp33_ASAP7_75t_L g8615 ( 
.A(n_7951),
.B(n_884),
.Y(n_8615)
);

BUFx6f_ASAP7_75t_L g8616 ( 
.A(n_8225),
.Y(n_8616)
);

NAND2xp5_ASAP7_75t_L g8617 ( 
.A(n_8130),
.B(n_884),
.Y(n_8617)
);

INVx1_ASAP7_75t_L g8618 ( 
.A(n_8134),
.Y(n_8618)
);

INVx3_ASAP7_75t_L g8619 ( 
.A(n_8234),
.Y(n_8619)
);

BUFx6f_ASAP7_75t_L g8620 ( 
.A(n_8055),
.Y(n_8620)
);

CKINVDCx20_ASAP7_75t_R g8621 ( 
.A(n_8241),
.Y(n_8621)
);

AOI22xp33_ASAP7_75t_L g8622 ( 
.A1(n_8199),
.A2(n_291),
.B1(n_289),
.B2(n_290),
.Y(n_8622)
);

AND2x2_ASAP7_75t_L g8623 ( 
.A(n_8210),
.B(n_885),
.Y(n_8623)
);

AND2x2_ASAP7_75t_L g8624 ( 
.A(n_8211),
.B(n_885),
.Y(n_8624)
);

NAND3xp33_ASAP7_75t_SL g8625 ( 
.A(n_7829),
.B(n_290),
.C(n_292),
.Y(n_8625)
);

INVx1_ASAP7_75t_L g8626 ( 
.A(n_7958),
.Y(n_8626)
);

A2O1A1Ixp33_ASAP7_75t_L g8627 ( 
.A1(n_8275),
.A2(n_887),
.B(n_889),
.C(n_886),
.Y(n_8627)
);

NAND2xp5_ASAP7_75t_L g8628 ( 
.A(n_7972),
.B(n_886),
.Y(n_8628)
);

BUFx6f_ASAP7_75t_L g8629 ( 
.A(n_8068),
.Y(n_8629)
);

INVx1_ASAP7_75t_L g8630 ( 
.A(n_7995),
.Y(n_8630)
);

AO21x1_ASAP7_75t_L g8631 ( 
.A1(n_8214),
.A2(n_292),
.B(n_293),
.Y(n_8631)
);

AOI22xp5_ASAP7_75t_L g8632 ( 
.A1(n_8127),
.A2(n_294),
.B1(n_292),
.B2(n_293),
.Y(n_8632)
);

BUFx2_ASAP7_75t_L g8633 ( 
.A(n_8003),
.Y(n_8633)
);

OAI22xp5_ASAP7_75t_L g8634 ( 
.A1(n_8044),
.A2(n_295),
.B1(n_293),
.B2(n_294),
.Y(n_8634)
);

NAND2xp5_ASAP7_75t_SL g8635 ( 
.A(n_7960),
.B(n_889),
.Y(n_8635)
);

AOI21xp5_ASAP7_75t_L g8636 ( 
.A1(n_8077),
.A2(n_891),
.B(n_890),
.Y(n_8636)
);

O2A1O1Ixp33_ASAP7_75t_SL g8637 ( 
.A1(n_8059),
.A2(n_296),
.B(n_294),
.C(n_295),
.Y(n_8637)
);

NAND2xp5_ASAP7_75t_SL g8638 ( 
.A(n_7965),
.B(n_890),
.Y(n_8638)
);

NAND2xp5_ASAP7_75t_SL g8639 ( 
.A(n_8197),
.B(n_891),
.Y(n_8639)
);

OAI22xp5_ASAP7_75t_SL g8640 ( 
.A1(n_8202),
.A2(n_297),
.B1(n_295),
.B2(n_296),
.Y(n_8640)
);

OR2x2_ASAP7_75t_L g8641 ( 
.A(n_8015),
.B(n_892),
.Y(n_8641)
);

AND2x2_ASAP7_75t_L g8642 ( 
.A(n_8182),
.B(n_892),
.Y(n_8642)
);

BUFx6f_ASAP7_75t_L g8643 ( 
.A(n_8132),
.Y(n_8643)
);

INVx2_ASAP7_75t_L g8644 ( 
.A(n_8012),
.Y(n_8644)
);

NAND2xp5_ASAP7_75t_L g8645 ( 
.A(n_8013),
.B(n_893),
.Y(n_8645)
);

NAND2xp5_ASAP7_75t_SL g8646 ( 
.A(n_8205),
.B(n_894),
.Y(n_8646)
);

INVx1_ASAP7_75t_L g8647 ( 
.A(n_8018),
.Y(n_8647)
);

CKINVDCx16_ASAP7_75t_R g8648 ( 
.A(n_7961),
.Y(n_8648)
);

AND2x2_ASAP7_75t_L g8649 ( 
.A(n_8232),
.B(n_894),
.Y(n_8649)
);

CKINVDCx5p33_ASAP7_75t_R g8650 ( 
.A(n_8315),
.Y(n_8650)
);

AOI21xp5_ASAP7_75t_L g8651 ( 
.A1(n_7931),
.A2(n_896),
.B(n_895),
.Y(n_8651)
);

NAND2xp5_ASAP7_75t_SL g8652 ( 
.A(n_8019),
.B(n_895),
.Y(n_8652)
);

AOI21xp5_ASAP7_75t_L g8653 ( 
.A1(n_8277),
.A2(n_897),
.B(n_896),
.Y(n_8653)
);

NAND2xp5_ASAP7_75t_L g8654 ( 
.A(n_7812),
.B(n_897),
.Y(n_8654)
);

INVx1_ASAP7_75t_L g8655 ( 
.A(n_8153),
.Y(n_8655)
);

OAI22xp5_ASAP7_75t_L g8656 ( 
.A1(n_8024),
.A2(n_298),
.B1(n_296),
.B2(n_297),
.Y(n_8656)
);

AOI22xp5_ASAP7_75t_L g8657 ( 
.A1(n_8190),
.A2(n_299),
.B1(n_297),
.B2(n_298),
.Y(n_8657)
);

OAI21x1_ASAP7_75t_L g8658 ( 
.A1(n_8171),
.A2(n_298),
.B(n_299),
.Y(n_8658)
);

BUFx6f_ASAP7_75t_L g8659 ( 
.A(n_8087),
.Y(n_8659)
);

NOR2xp33_ASAP7_75t_R g8660 ( 
.A(n_8041),
.B(n_299),
.Y(n_8660)
);

AO21x1_ASAP7_75t_L g8661 ( 
.A1(n_8230),
.A2(n_300),
.B(n_301),
.Y(n_8661)
);

O2A1O1Ixp33_ASAP7_75t_L g8662 ( 
.A1(n_8126),
.A2(n_302),
.B(n_300),
.C(n_301),
.Y(n_8662)
);

INVx1_ASAP7_75t_L g8663 ( 
.A(n_8071),
.Y(n_8663)
);

NOR2xp33_ASAP7_75t_L g8664 ( 
.A(n_8227),
.B(n_898),
.Y(n_8664)
);

O2A1O1Ixp5_ASAP7_75t_L g8665 ( 
.A1(n_8279),
.A2(n_302),
.B(n_300),
.C(n_301),
.Y(n_8665)
);

AND2x2_ASAP7_75t_L g8666 ( 
.A(n_8177),
.B(n_898),
.Y(n_8666)
);

OR2x6_ASAP7_75t_L g8667 ( 
.A(n_8174),
.B(n_899),
.Y(n_8667)
);

INVx3_ASAP7_75t_L g8668 ( 
.A(n_8095),
.Y(n_8668)
);

BUFx6f_ASAP7_75t_L g8669 ( 
.A(n_8203),
.Y(n_8669)
);

INVx3_ASAP7_75t_L g8670 ( 
.A(n_7928),
.Y(n_8670)
);

HB1xp67_ASAP7_75t_L g8671 ( 
.A(n_8073),
.Y(n_8671)
);

NAND2xp5_ASAP7_75t_L g8672 ( 
.A(n_7823),
.B(n_899),
.Y(n_8672)
);

O2A1O1Ixp33_ASAP7_75t_L g8673 ( 
.A1(n_8183),
.A2(n_8083),
.B(n_7831),
.C(n_8220),
.Y(n_8673)
);

OAI21x1_ASAP7_75t_L g8674 ( 
.A1(n_8035),
.A2(n_8053),
.B(n_8105),
.Y(n_8674)
);

NAND2xp5_ASAP7_75t_SL g8675 ( 
.A(n_8028),
.B(n_900),
.Y(n_8675)
);

OAI22xp5_ASAP7_75t_L g8676 ( 
.A1(n_8244),
.A2(n_304),
.B1(n_302),
.B2(n_303),
.Y(n_8676)
);

O2A1O1Ixp33_ASAP7_75t_L g8677 ( 
.A1(n_8223),
.A2(n_305),
.B(n_303),
.C(n_304),
.Y(n_8677)
);

INVx1_ASAP7_75t_L g8678 ( 
.A(n_8074),
.Y(n_8678)
);

NOR3xp33_ASAP7_75t_SL g8679 ( 
.A(n_8150),
.B(n_305),
.C(n_306),
.Y(n_8679)
);

INVx2_ASAP7_75t_SL g8680 ( 
.A(n_8048),
.Y(n_8680)
);

INVx3_ASAP7_75t_L g8681 ( 
.A(n_7928),
.Y(n_8681)
);

NAND3xp33_ASAP7_75t_SL g8682 ( 
.A(n_8184),
.B(n_306),
.C(n_307),
.Y(n_8682)
);

INVx2_ASAP7_75t_L g8683 ( 
.A(n_8078),
.Y(n_8683)
);

INVxp67_ASAP7_75t_L g8684 ( 
.A(n_7974),
.Y(n_8684)
);

CKINVDCx5p33_ASAP7_75t_R g8685 ( 
.A(n_8243),
.Y(n_8685)
);

NAND2xp5_ASAP7_75t_SL g8686 ( 
.A(n_7982),
.B(n_900),
.Y(n_8686)
);

O2A1O1Ixp33_ASAP7_75t_L g8687 ( 
.A1(n_8207),
.A2(n_309),
.B(n_306),
.C(n_308),
.Y(n_8687)
);

NOR2xp33_ASAP7_75t_L g8688 ( 
.A(n_8222),
.B(n_902),
.Y(n_8688)
);

INVx2_ASAP7_75t_L g8689 ( 
.A(n_8080),
.Y(n_8689)
);

INVx2_ASAP7_75t_L g8690 ( 
.A(n_8081),
.Y(n_8690)
);

OAI21x1_ASAP7_75t_L g8691 ( 
.A1(n_8129),
.A2(n_308),
.B(n_309),
.Y(n_8691)
);

HB1xp67_ASAP7_75t_L g8692 ( 
.A(n_8082),
.Y(n_8692)
);

NOR2xp33_ASAP7_75t_L g8693 ( 
.A(n_8124),
.B(n_902),
.Y(n_8693)
);

O2A1O1Ixp5_ASAP7_75t_L g8694 ( 
.A1(n_8283),
.A2(n_310),
.B(n_308),
.C(n_309),
.Y(n_8694)
);

HB1xp67_ASAP7_75t_L g8695 ( 
.A(n_8101),
.Y(n_8695)
);

OAI21xp5_ASAP7_75t_L g8696 ( 
.A1(n_8284),
.A2(n_310),
.B(n_311),
.Y(n_8696)
);

AOI21xp5_ASAP7_75t_L g8697 ( 
.A1(n_8285),
.A2(n_904),
.B(n_903),
.Y(n_8697)
);

O2A1O1Ixp33_ASAP7_75t_L g8698 ( 
.A1(n_8036),
.A2(n_312),
.B(n_310),
.C(n_311),
.Y(n_8698)
);

NAND2xp5_ASAP7_75t_L g8699 ( 
.A(n_7826),
.B(n_905),
.Y(n_8699)
);

NOR2xp33_ASAP7_75t_SL g8700 ( 
.A(n_8167),
.B(n_312),
.Y(n_8700)
);

NAND2xp5_ASAP7_75t_L g8701 ( 
.A(n_7827),
.B(n_906),
.Y(n_8701)
);

AND2x4_ASAP7_75t_SL g8702 ( 
.A(n_8023),
.B(n_906),
.Y(n_8702)
);

OAI22x1_ASAP7_75t_L g8703 ( 
.A1(n_8158),
.A2(n_314),
.B1(n_312),
.B2(n_313),
.Y(n_8703)
);

NAND3xp33_ASAP7_75t_SL g8704 ( 
.A(n_8161),
.B(n_313),
.C(n_314),
.Y(n_8704)
);

AND2x2_ASAP7_75t_L g8705 ( 
.A(n_7967),
.B(n_907),
.Y(n_8705)
);

NOR3xp33_ASAP7_75t_L g8706 ( 
.A(n_8286),
.B(n_314),
.C(n_315),
.Y(n_8706)
);

OAI21x1_ASAP7_75t_L g8707 ( 
.A1(n_7990),
.A2(n_8001),
.B(n_7993),
.Y(n_8707)
);

A2O1A1Ixp33_ASAP7_75t_L g8708 ( 
.A1(n_8288),
.A2(n_908),
.B(n_909),
.C(n_907),
.Y(n_8708)
);

AOI21xp5_ASAP7_75t_L g8709 ( 
.A1(n_8293),
.A2(n_909),
.B(n_908),
.Y(n_8709)
);

AOI21xp5_ASAP7_75t_L g8710 ( 
.A1(n_8298),
.A2(n_8312),
.B(n_8307),
.Y(n_8710)
);

AOI21xp5_ASAP7_75t_L g8711 ( 
.A1(n_8313),
.A2(n_911),
.B(n_910),
.Y(n_8711)
);

NAND2xp5_ASAP7_75t_SL g8712 ( 
.A(n_7847),
.B(n_910),
.Y(n_8712)
);

AOI21xp5_ASAP7_75t_L g8713 ( 
.A1(n_8328),
.A2(n_912),
.B(n_911),
.Y(n_8713)
);

AOI22xp5_ASAP7_75t_L g8714 ( 
.A1(n_8209),
.A2(n_317),
.B1(n_315),
.B2(n_316),
.Y(n_8714)
);

NAND2xp5_ASAP7_75t_SL g8715 ( 
.A(n_7855),
.B(n_912),
.Y(n_8715)
);

NAND3xp33_ASAP7_75t_SL g8716 ( 
.A(n_8329),
.B(n_315),
.C(n_316),
.Y(n_8716)
);

BUFx8_ASAP7_75t_SL g8717 ( 
.A(n_8247),
.Y(n_8717)
);

NAND2xp5_ASAP7_75t_L g8718 ( 
.A(n_7832),
.B(n_7858),
.Y(n_8718)
);

NOR2xp33_ASAP7_75t_L g8719 ( 
.A(n_7870),
.B(n_913),
.Y(n_8719)
);

INVx1_ASAP7_75t_L g8720 ( 
.A(n_8106),
.Y(n_8720)
);

A2O1A1Ixp33_ASAP7_75t_L g8721 ( 
.A1(n_8330),
.A2(n_914),
.B(n_915),
.C(n_913),
.Y(n_8721)
);

A2O1A1Ixp33_ASAP7_75t_L g8722 ( 
.A1(n_8335),
.A2(n_916),
.B(n_917),
.C(n_915),
.Y(n_8722)
);

NAND2xp5_ASAP7_75t_L g8723 ( 
.A(n_7878),
.B(n_917),
.Y(n_8723)
);

INVx1_ASAP7_75t_L g8724 ( 
.A(n_8122),
.Y(n_8724)
);

NOR2x1_ASAP7_75t_L g8725 ( 
.A(n_7919),
.B(n_918),
.Y(n_8725)
);

INVx2_ASAP7_75t_L g8726 ( 
.A(n_8133),
.Y(n_8726)
);

NAND2xp5_ASAP7_75t_L g8727 ( 
.A(n_7880),
.B(n_919),
.Y(n_8727)
);

O2A1O1Ixp33_ASAP7_75t_L g8728 ( 
.A1(n_8235),
.A2(n_318),
.B(n_316),
.C(n_317),
.Y(n_8728)
);

OAI22xp5_ASAP7_75t_L g8729 ( 
.A1(n_7978),
.A2(n_319),
.B1(n_317),
.B2(n_318),
.Y(n_8729)
);

O2A1O1Ixp33_ASAP7_75t_L g8730 ( 
.A1(n_8236),
.A2(n_320),
.B(n_318),
.C(n_319),
.Y(n_8730)
);

NAND2xp5_ASAP7_75t_SL g8731 ( 
.A(n_7889),
.B(n_919),
.Y(n_8731)
);

NOR2xp33_ASAP7_75t_L g8732 ( 
.A(n_7891),
.B(n_920),
.Y(n_8732)
);

O2A1O1Ixp33_ASAP7_75t_L g8733 ( 
.A1(n_8226),
.A2(n_321),
.B(n_319),
.C(n_320),
.Y(n_8733)
);

INVx3_ASAP7_75t_L g8734 ( 
.A(n_7928),
.Y(n_8734)
);

BUFx2_ASAP7_75t_L g8735 ( 
.A(n_7928),
.Y(n_8735)
);

NAND2xp5_ASAP7_75t_L g8736 ( 
.A(n_7892),
.B(n_920),
.Y(n_8736)
);

INVx2_ASAP7_75t_SL g8737 ( 
.A(n_8166),
.Y(n_8737)
);

OAI21x1_ASAP7_75t_L g8738 ( 
.A1(n_8004),
.A2(n_320),
.B(n_321),
.Y(n_8738)
);

NAND2xp5_ASAP7_75t_SL g8739 ( 
.A(n_7917),
.B(n_921),
.Y(n_8739)
);

O2A1O1Ixp33_ASAP7_75t_L g8740 ( 
.A1(n_8213),
.A2(n_8245),
.B(n_8061),
.C(n_8110),
.Y(n_8740)
);

NAND2xp5_ASAP7_75t_SL g8741 ( 
.A(n_7926),
.B(n_922),
.Y(n_8741)
);

O2A1O1Ixp33_ASAP7_75t_L g8742 ( 
.A1(n_8043),
.A2(n_8039),
.B(n_8159),
.C(n_8144),
.Y(n_8742)
);

OAI22xp5_ASAP7_75t_SL g8743 ( 
.A1(n_8218),
.A2(n_323),
.B1(n_321),
.B2(n_322),
.Y(n_8743)
);

O2A1O1Ixp5_ASAP7_75t_L g8744 ( 
.A1(n_8141),
.A2(n_324),
.B(n_322),
.C(n_323),
.Y(n_8744)
);

INVx1_ASAP7_75t_L g8745 ( 
.A(n_8192),
.Y(n_8745)
);

NOR2xp33_ASAP7_75t_R g8746 ( 
.A(n_8138),
.B(n_322),
.Y(n_8746)
);

INVx1_ASAP7_75t_L g8747 ( 
.A(n_8194),
.Y(n_8747)
);

INVx1_ASAP7_75t_L g8748 ( 
.A(n_8195),
.Y(n_8748)
);

NAND2xp5_ASAP7_75t_L g8749 ( 
.A(n_7927),
.B(n_922),
.Y(n_8749)
);

AND2x2_ASAP7_75t_L g8750 ( 
.A(n_8114),
.B(n_923),
.Y(n_8750)
);

AOI21xp5_ASAP7_75t_L g8751 ( 
.A1(n_7918),
.A2(n_924),
.B(n_923),
.Y(n_8751)
);

NOR2xp33_ASAP7_75t_SL g8752 ( 
.A(n_7816),
.B(n_323),
.Y(n_8752)
);

INVx3_ASAP7_75t_L g8753 ( 
.A(n_8175),
.Y(n_8753)
);

NOR2xp33_ASAP7_75t_R g8754 ( 
.A(n_8148),
.B(n_8152),
.Y(n_8754)
);

INVx2_ASAP7_75t_L g8755 ( 
.A(n_8186),
.Y(n_8755)
);

NAND2xp5_ASAP7_75t_L g8756 ( 
.A(n_7952),
.B(n_924),
.Y(n_8756)
);

O2A1O1Ixp5_ASAP7_75t_L g8757 ( 
.A1(n_7957),
.A2(n_7983),
.B(n_7985),
.C(n_7968),
.Y(n_8757)
);

NAND2xp5_ASAP7_75t_SL g8758 ( 
.A(n_8031),
.B(n_8142),
.Y(n_8758)
);

NAND2xp5_ASAP7_75t_L g8759 ( 
.A(n_8160),
.B(n_925),
.Y(n_8759)
);

NAND2xp5_ASAP7_75t_SL g8760 ( 
.A(n_8233),
.B(n_925),
.Y(n_8760)
);

O2A1O1Ixp33_ASAP7_75t_L g8761 ( 
.A1(n_8143),
.A2(n_326),
.B(n_324),
.C(n_325),
.Y(n_8761)
);

AOI21xp5_ASAP7_75t_L g8762 ( 
.A1(n_7923),
.A2(n_7925),
.B(n_7845),
.Y(n_8762)
);

NAND2xp5_ASAP7_75t_L g8763 ( 
.A(n_8231),
.B(n_926),
.Y(n_8763)
);

INVx3_ASAP7_75t_L g8764 ( 
.A(n_8156),
.Y(n_8764)
);

NOR2xp33_ASAP7_75t_L g8765 ( 
.A(n_8117),
.B(n_926),
.Y(n_8765)
);

O2A1O1Ixp33_ASAP7_75t_L g8766 ( 
.A1(n_8189),
.A2(n_327),
.B(n_325),
.C(n_326),
.Y(n_8766)
);

NOR2xp33_ASAP7_75t_SL g8767 ( 
.A(n_7839),
.B(n_326),
.Y(n_8767)
);

OAI21xp33_ASAP7_75t_SL g8768 ( 
.A1(n_7842),
.A2(n_928),
.B(n_927),
.Y(n_8768)
);

NAND2xp5_ASAP7_75t_SL g8769 ( 
.A(n_8219),
.B(n_8216),
.Y(n_8769)
);

OAI22xp5_ASAP7_75t_L g8770 ( 
.A1(n_7846),
.A2(n_329),
.B1(n_327),
.B2(n_328),
.Y(n_8770)
);

NAND3xp33_ASAP7_75t_L g8771 ( 
.A(n_7859),
.B(n_327),
.C(n_328),
.Y(n_8771)
);

INVxp67_ASAP7_75t_SL g8772 ( 
.A(n_8196),
.Y(n_8772)
);

AOI21xp5_ASAP7_75t_L g8773 ( 
.A1(n_7861),
.A2(n_7904),
.B(n_7865),
.Y(n_8773)
);

OAI22x1_ASAP7_75t_L g8774 ( 
.A1(n_8229),
.A2(n_330),
.B1(n_328),
.B2(n_329),
.Y(n_8774)
);

AOI21xp5_ASAP7_75t_L g8775 ( 
.A1(n_7905),
.A2(n_929),
.B(n_927),
.Y(n_8775)
);

NAND2xp5_ASAP7_75t_L g8776 ( 
.A(n_8187),
.B(n_929),
.Y(n_8776)
);

NAND2xp5_ASAP7_75t_L g8777 ( 
.A(n_7935),
.B(n_930),
.Y(n_8777)
);

OAI21xp33_ASAP7_75t_L g8778 ( 
.A1(n_7911),
.A2(n_329),
.B(n_330),
.Y(n_8778)
);

INVx6_ASAP7_75t_L g8779 ( 
.A(n_8204),
.Y(n_8779)
);

NAND2xp5_ASAP7_75t_L g8780 ( 
.A(n_7884),
.B(n_930),
.Y(n_8780)
);

INVx1_ASAP7_75t_L g8781 ( 
.A(n_7984),
.Y(n_8781)
);

AOI21xp5_ASAP7_75t_L g8782 ( 
.A1(n_7887),
.A2(n_7896),
.B(n_7895),
.Y(n_8782)
);

NAND2xp5_ASAP7_75t_L g8783 ( 
.A(n_7900),
.B(n_931),
.Y(n_8783)
);

BUFx6f_ASAP7_75t_L g8784 ( 
.A(n_8109),
.Y(n_8784)
);

BUFx6f_ASAP7_75t_L g8785 ( 
.A(n_8123),
.Y(n_8785)
);

AOI22xp33_ASAP7_75t_L g8786 ( 
.A1(n_7885),
.A2(n_332),
.B1(n_330),
.B2(n_331),
.Y(n_8786)
);

BUFx2_ASAP7_75t_L g8787 ( 
.A(n_8239),
.Y(n_8787)
);

INVx6_ASAP7_75t_L g8788 ( 
.A(n_7862),
.Y(n_8788)
);

AND2x2_ASAP7_75t_L g8789 ( 
.A(n_8215),
.B(n_931),
.Y(n_8789)
);

O2A1O1Ixp33_ASAP7_75t_L g8790 ( 
.A1(n_8263),
.A2(n_333),
.B(n_331),
.C(n_332),
.Y(n_8790)
);

OAI22xp5_ASAP7_75t_L g8791 ( 
.A1(n_7924),
.A2(n_333),
.B1(n_331),
.B2(n_332),
.Y(n_8791)
);

NAND2xp5_ASAP7_75t_L g8792 ( 
.A(n_7903),
.B(n_932),
.Y(n_8792)
);

CKINVDCx5p33_ASAP7_75t_R g8793 ( 
.A(n_7874),
.Y(n_8793)
);

A2O1A1Ixp33_ASAP7_75t_L g8794 ( 
.A1(n_8069),
.A2(n_934),
.B(n_935),
.C(n_933),
.Y(n_8794)
);

INVx1_ASAP7_75t_SL g8795 ( 
.A(n_8140),
.Y(n_8795)
);

A2O1A1Ixp33_ASAP7_75t_L g8796 ( 
.A1(n_8070),
.A2(n_935),
.B(n_936),
.C(n_933),
.Y(n_8796)
);

NOR2xp67_ASAP7_75t_SL g8797 ( 
.A(n_8072),
.B(n_334),
.Y(n_8797)
);

NAND2xp5_ASAP7_75t_L g8798 ( 
.A(n_8115),
.B(n_937),
.Y(n_8798)
);

NAND2x1p5_ASAP7_75t_L g8799 ( 
.A(n_8005),
.B(n_938),
.Y(n_8799)
);

A2O1A1Ixp33_ASAP7_75t_SL g8800 ( 
.A1(n_8040),
.A2(n_336),
.B(n_334),
.C(n_335),
.Y(n_8800)
);

BUFx2_ASAP7_75t_L g8801 ( 
.A(n_8239),
.Y(n_8801)
);

NOR2xp33_ASAP7_75t_L g8802 ( 
.A(n_7980),
.B(n_939),
.Y(n_8802)
);

BUFx12f_ASAP7_75t_L g8803 ( 
.A(n_8173),
.Y(n_8803)
);

BUFx6f_ASAP7_75t_L g8804 ( 
.A(n_8239),
.Y(n_8804)
);

OAI21xp5_ASAP7_75t_L g8805 ( 
.A1(n_8079),
.A2(n_334),
.B(n_335),
.Y(n_8805)
);

AND2x2_ASAP7_75t_L g8806 ( 
.A(n_7913),
.B(n_940),
.Y(n_8806)
);

NAND2xp5_ASAP7_75t_L g8807 ( 
.A(n_7948),
.B(n_940),
.Y(n_8807)
);

INVx1_ASAP7_75t_L g8808 ( 
.A(n_7913),
.Y(n_8808)
);

A2O1A1Ixp33_ASAP7_75t_SL g8809 ( 
.A1(n_8131),
.A2(n_338),
.B(n_336),
.C(n_337),
.Y(n_8809)
);

NAND2xp5_ASAP7_75t_SL g8810 ( 
.A(n_8011),
.B(n_942),
.Y(n_8810)
);

HB1xp67_ASAP7_75t_L g8811 ( 
.A(n_8020),
.Y(n_8811)
);

INVx1_ASAP7_75t_SL g8812 ( 
.A(n_7955),
.Y(n_8812)
);

AOI21xp5_ASAP7_75t_L g8813 ( 
.A1(n_8090),
.A2(n_8103),
.B(n_8094),
.Y(n_8813)
);

INVx3_ASAP7_75t_L g8814 ( 
.A(n_8193),
.Y(n_8814)
);

AND2x2_ASAP7_75t_L g8815 ( 
.A(n_7913),
.B(n_8112),
.Y(n_8815)
);

INVx3_ASAP7_75t_L g8816 ( 
.A(n_8057),
.Y(n_8816)
);

HB1xp67_ASAP7_75t_L g8817 ( 
.A(n_8120),
.Y(n_8817)
);

INVx2_ASAP7_75t_L g8818 ( 
.A(n_7813),
.Y(n_8818)
);

O2A1O1Ixp33_ASAP7_75t_L g8819 ( 
.A1(n_7881),
.A2(n_338),
.B(n_336),
.C(n_337),
.Y(n_8819)
);

BUFx10_ASAP7_75t_L g8820 ( 
.A(n_7970),
.Y(n_8820)
);

BUFx6f_ASAP7_75t_L g8821 ( 
.A(n_7817),
.Y(n_8821)
);

INVx2_ASAP7_75t_L g8822 ( 
.A(n_7813),
.Y(n_8822)
);

AOI22xp5_ASAP7_75t_L g8823 ( 
.A1(n_7881),
.A2(n_340),
.B1(n_337),
.B2(n_339),
.Y(n_8823)
);

BUFx6f_ASAP7_75t_L g8824 ( 
.A(n_7817),
.Y(n_8824)
);

O2A1O1Ixp33_ASAP7_75t_L g8825 ( 
.A1(n_7881),
.A2(n_341),
.B(n_339),
.C(n_340),
.Y(n_8825)
);

AOI22xp5_ASAP7_75t_L g8826 ( 
.A1(n_7881),
.A2(n_342),
.B1(n_340),
.B2(n_341),
.Y(n_8826)
);

AND2x2_ASAP7_75t_L g8827 ( 
.A(n_7877),
.B(n_942),
.Y(n_8827)
);

O2A1O1Ixp33_ASAP7_75t_L g8828 ( 
.A1(n_7881),
.A2(n_344),
.B(n_342),
.C(n_343),
.Y(n_8828)
);

INVx4_ASAP7_75t_L g8829 ( 
.A(n_7864),
.Y(n_8829)
);

BUFx3_ASAP7_75t_L g8830 ( 
.A(n_8026),
.Y(n_8830)
);

AOI21xp5_ASAP7_75t_L g8831 ( 
.A1(n_7881),
.A2(n_944),
.B(n_943),
.Y(n_8831)
);

AO21x1_ASAP7_75t_L g8832 ( 
.A1(n_7822),
.A2(n_342),
.B(n_343),
.Y(n_8832)
);

NOR2xp33_ASAP7_75t_L g8833 ( 
.A(n_7863),
.B(n_943),
.Y(n_8833)
);

INVx2_ASAP7_75t_SL g8834 ( 
.A(n_7864),
.Y(n_8834)
);

NAND2xp5_ASAP7_75t_SL g8835 ( 
.A(n_7869),
.B(n_944),
.Y(n_8835)
);

HB1xp67_ASAP7_75t_L g8836 ( 
.A(n_8037),
.Y(n_8836)
);

O2A1O1Ixp33_ASAP7_75t_L g8837 ( 
.A1(n_7881),
.A2(n_346),
.B(n_344),
.C(n_345),
.Y(n_8837)
);

NOR2x1_ASAP7_75t_R g8838 ( 
.A(n_7940),
.B(n_344),
.Y(n_8838)
);

AOI33xp33_ASAP7_75t_L g8839 ( 
.A1(n_8149),
.A2(n_349),
.A3(n_351),
.B1(n_347),
.B2(n_348),
.B3(n_350),
.Y(n_8839)
);

NAND2xp5_ASAP7_75t_SL g8840 ( 
.A(n_7869),
.B(n_945),
.Y(n_8840)
);

INVx2_ASAP7_75t_L g8841 ( 
.A(n_7813),
.Y(n_8841)
);

AOI21xp5_ASAP7_75t_L g8842 ( 
.A1(n_7881),
.A2(n_946),
.B(n_945),
.Y(n_8842)
);

AND2x4_ASAP7_75t_L g8843 ( 
.A(n_7849),
.B(n_946),
.Y(n_8843)
);

AOI21xp5_ASAP7_75t_L g8844 ( 
.A1(n_7881),
.A2(n_948),
.B(n_947),
.Y(n_8844)
);

NAND2xp5_ASAP7_75t_L g8845 ( 
.A(n_7907),
.B(n_948),
.Y(n_8845)
);

INVx2_ASAP7_75t_L g8846 ( 
.A(n_7813),
.Y(n_8846)
);

NAND2xp5_ASAP7_75t_L g8847 ( 
.A(n_7907),
.B(n_949),
.Y(n_8847)
);

NOR2xp33_ASAP7_75t_L g8848 ( 
.A(n_7863),
.B(n_949),
.Y(n_8848)
);

NAND2xp5_ASAP7_75t_L g8849 ( 
.A(n_7907),
.B(n_950),
.Y(n_8849)
);

NAND2xp5_ASAP7_75t_L g8850 ( 
.A(n_7907),
.B(n_950),
.Y(n_8850)
);

NOR2xp33_ASAP7_75t_L g8851 ( 
.A(n_7863),
.B(n_951),
.Y(n_8851)
);

AOI21xp5_ASAP7_75t_L g8852 ( 
.A1(n_7881),
.A2(n_952),
.B(n_951),
.Y(n_8852)
);

OR2x6_ASAP7_75t_L g8853 ( 
.A(n_7857),
.B(n_952),
.Y(n_8853)
);

INVx3_ASAP7_75t_L g8854 ( 
.A(n_8302),
.Y(n_8854)
);

NAND2xp5_ASAP7_75t_L g8855 ( 
.A(n_7907),
.B(n_953),
.Y(n_8855)
);

A2O1A1Ixp33_ASAP7_75t_L g8856 ( 
.A1(n_7976),
.A2(n_954),
.B(n_955),
.C(n_953),
.Y(n_8856)
);

NOR2xp33_ASAP7_75t_L g8857 ( 
.A(n_7863),
.B(n_954),
.Y(n_8857)
);

INVx2_ASAP7_75t_SL g8858 ( 
.A(n_7864),
.Y(n_8858)
);

NAND2xp5_ASAP7_75t_L g8859 ( 
.A(n_7907),
.B(n_955),
.Y(n_8859)
);

INVx1_ASAP7_75t_L g8860 ( 
.A(n_7871),
.Y(n_8860)
);

INVx2_ASAP7_75t_SL g8861 ( 
.A(n_7864),
.Y(n_8861)
);

AOI21xp5_ASAP7_75t_L g8862 ( 
.A1(n_7881),
.A2(n_957),
.B(n_956),
.Y(n_8862)
);

INVx4_ASAP7_75t_L g8863 ( 
.A(n_7864),
.Y(n_8863)
);

NOR2xp33_ASAP7_75t_L g8864 ( 
.A(n_7863),
.B(n_956),
.Y(n_8864)
);

INVx1_ASAP7_75t_L g8865 ( 
.A(n_7871),
.Y(n_8865)
);

OR2x6_ASAP7_75t_L g8866 ( 
.A(n_7857),
.B(n_957),
.Y(n_8866)
);

INVx2_ASAP7_75t_SL g8867 ( 
.A(n_7864),
.Y(n_8867)
);

INVx2_ASAP7_75t_L g8868 ( 
.A(n_7813),
.Y(n_8868)
);

NAND2xp5_ASAP7_75t_L g8869 ( 
.A(n_7907),
.B(n_958),
.Y(n_8869)
);

O2A1O1Ixp33_ASAP7_75t_L g8870 ( 
.A1(n_7881),
.A2(n_349),
.B(n_347),
.C(n_348),
.Y(n_8870)
);

BUFx12f_ASAP7_75t_L g8871 ( 
.A(n_8378),
.Y(n_8871)
);

AOI22xp5_ASAP7_75t_L g8872 ( 
.A1(n_8423),
.A2(n_8456),
.B1(n_8445),
.B2(n_8612),
.Y(n_8872)
);

INVx2_ASAP7_75t_L g8873 ( 
.A(n_8538),
.Y(n_8873)
);

INVx1_ASAP7_75t_SL g8874 ( 
.A(n_8417),
.Y(n_8874)
);

HB1xp67_ASAP7_75t_L g8875 ( 
.A(n_8387),
.Y(n_8875)
);

INVx2_ASAP7_75t_L g8876 ( 
.A(n_8552),
.Y(n_8876)
);

OAI22xp5_ASAP7_75t_L g8877 ( 
.A1(n_8569),
.A2(n_351),
.B1(n_348),
.B2(n_350),
.Y(n_8877)
);

CKINVDCx5p33_ASAP7_75t_R g8878 ( 
.A(n_8459),
.Y(n_8878)
);

CKINVDCx5p33_ASAP7_75t_R g8879 ( 
.A(n_8650),
.Y(n_8879)
);

OAI22xp5_ASAP7_75t_L g8880 ( 
.A1(n_8569),
.A2(n_352),
.B1(n_350),
.B2(n_351),
.Y(n_8880)
);

A2O1A1Ixp33_ASAP7_75t_L g8881 ( 
.A1(n_8485),
.A2(n_960),
.B(n_961),
.C(n_959),
.Y(n_8881)
);

INVxp67_ASAP7_75t_L g8882 ( 
.A(n_8355),
.Y(n_8882)
);

OR2x6_ASAP7_75t_L g8883 ( 
.A(n_8434),
.B(n_8577),
.Y(n_8883)
);

INVx1_ASAP7_75t_L g8884 ( 
.A(n_8351),
.Y(n_8884)
);

INVx2_ASAP7_75t_L g8885 ( 
.A(n_8367),
.Y(n_8885)
);

INVx2_ASAP7_75t_L g8886 ( 
.A(n_8375),
.Y(n_8886)
);

AND2x2_ASAP7_75t_L g8887 ( 
.A(n_8512),
.B(n_959),
.Y(n_8887)
);

INVx1_ASAP7_75t_L g8888 ( 
.A(n_8377),
.Y(n_8888)
);

AOI22xp5_ASAP7_75t_L g8889 ( 
.A1(n_8379),
.A2(n_354),
.B1(n_352),
.B2(n_353),
.Y(n_8889)
);

OR2x2_ASAP7_75t_L g8890 ( 
.A(n_8406),
.B(n_960),
.Y(n_8890)
);

INVx1_ASAP7_75t_L g8891 ( 
.A(n_8380),
.Y(n_8891)
);

AND2x2_ASAP7_75t_L g8892 ( 
.A(n_8419),
.B(n_961),
.Y(n_8892)
);

INVx2_ASAP7_75t_L g8893 ( 
.A(n_8401),
.Y(n_8893)
);

OAI22xp33_ASAP7_75t_L g8894 ( 
.A1(n_8752),
.A2(n_354),
.B1(n_352),
.B2(n_353),
.Y(n_8894)
);

INVx1_ASAP7_75t_SL g8895 ( 
.A(n_8426),
.Y(n_8895)
);

BUFx3_ASAP7_75t_L g8896 ( 
.A(n_8360),
.Y(n_8896)
);

OAI21xp5_ASAP7_75t_L g8897 ( 
.A1(n_8611),
.A2(n_353),
.B(n_355),
.Y(n_8897)
);

AOI22xp33_ASAP7_75t_SL g8898 ( 
.A1(n_8354),
.A2(n_357),
.B1(n_355),
.B2(n_356),
.Y(n_8898)
);

INVx1_ASAP7_75t_L g8899 ( 
.A(n_8404),
.Y(n_8899)
);

INVx2_ASAP7_75t_SL g8900 ( 
.A(n_8388),
.Y(n_8900)
);

INVx1_ASAP7_75t_L g8901 ( 
.A(n_8420),
.Y(n_8901)
);

OR2x2_ASAP7_75t_L g8902 ( 
.A(n_8836),
.B(n_962),
.Y(n_8902)
);

BUFx2_ASAP7_75t_L g8903 ( 
.A(n_8370),
.Y(n_8903)
);

OAI22xp33_ASAP7_75t_L g8904 ( 
.A1(n_8767),
.A2(n_357),
.B1(n_355),
.B2(n_356),
.Y(n_8904)
);

NAND2xp5_ASAP7_75t_L g8905 ( 
.A(n_8343),
.B(n_8671),
.Y(n_8905)
);

NAND2xp5_ASAP7_75t_L g8906 ( 
.A(n_8692),
.B(n_962),
.Y(n_8906)
);

INVx1_ASAP7_75t_L g8907 ( 
.A(n_8421),
.Y(n_8907)
);

AOI22xp5_ASAP7_75t_L g8908 ( 
.A1(n_8452),
.A2(n_359),
.B1(n_357),
.B2(n_358),
.Y(n_8908)
);

INVx1_ASAP7_75t_L g8909 ( 
.A(n_8437),
.Y(n_8909)
);

INVx3_ASAP7_75t_L g8910 ( 
.A(n_8830),
.Y(n_8910)
);

BUFx3_ASAP7_75t_L g8911 ( 
.A(n_8643),
.Y(n_8911)
);

AOI22xp33_ASAP7_75t_L g8912 ( 
.A1(n_8458),
.A2(n_360),
.B1(n_358),
.B2(n_359),
.Y(n_8912)
);

INVx2_ASAP7_75t_L g8913 ( 
.A(n_8442),
.Y(n_8913)
);

BUFx6f_ASAP7_75t_L g8914 ( 
.A(n_8362),
.Y(n_8914)
);

NAND2xp5_ASAP7_75t_L g8915 ( 
.A(n_8695),
.B(n_963),
.Y(n_8915)
);

INVx1_ASAP7_75t_L g8916 ( 
.A(n_8446),
.Y(n_8916)
);

BUFx2_ASAP7_75t_SL g8917 ( 
.A(n_8555),
.Y(n_8917)
);

BUFx3_ASAP7_75t_L g8918 ( 
.A(n_8643),
.Y(n_8918)
);

BUFx3_ASAP7_75t_L g8919 ( 
.A(n_8433),
.Y(n_8919)
);

BUFx2_ASAP7_75t_L g8920 ( 
.A(n_8409),
.Y(n_8920)
);

NAND2xp5_ASAP7_75t_L g8921 ( 
.A(n_8570),
.B(n_963),
.Y(n_8921)
);

BUFx10_ASAP7_75t_L g8922 ( 
.A(n_8536),
.Y(n_8922)
);

INVx2_ASAP7_75t_L g8923 ( 
.A(n_8447),
.Y(n_8923)
);

AOI22xp33_ASAP7_75t_L g8924 ( 
.A1(n_8803),
.A2(n_362),
.B1(n_360),
.B2(n_361),
.Y(n_8924)
);

AND2x2_ASAP7_75t_L g8925 ( 
.A(n_8430),
.B(n_964),
.Y(n_8925)
);

OAI21xp33_ASAP7_75t_SL g8926 ( 
.A1(n_8341),
.A2(n_965),
.B(n_964),
.Y(n_8926)
);

INVx1_ASAP7_75t_L g8927 ( 
.A(n_8449),
.Y(n_8927)
);

INVx3_ASAP7_75t_L g8928 ( 
.A(n_8362),
.Y(n_8928)
);

NAND2xp5_ASAP7_75t_L g8929 ( 
.A(n_8595),
.B(n_966),
.Y(n_8929)
);

INVx1_ASAP7_75t_L g8930 ( 
.A(n_8526),
.Y(n_8930)
);

AOI21xp5_ASAP7_75t_L g8931 ( 
.A1(n_8710),
.A2(n_361),
.B(n_362),
.Y(n_8931)
);

INVxp67_ASAP7_75t_L g8932 ( 
.A(n_8680),
.Y(n_8932)
);

NAND2xp5_ASAP7_75t_L g8933 ( 
.A(n_8755),
.B(n_966),
.Y(n_8933)
);

BUFx2_ASAP7_75t_SL g8934 ( 
.A(n_8530),
.Y(n_8934)
);

AND2x4_ASAP7_75t_L g8935 ( 
.A(n_8429),
.B(n_8508),
.Y(n_8935)
);

INVx1_ASAP7_75t_SL g8936 ( 
.A(n_8556),
.Y(n_8936)
);

INVx2_ASAP7_75t_L g8937 ( 
.A(n_8537),
.Y(n_8937)
);

HB1xp67_ASAP7_75t_L g8938 ( 
.A(n_8633),
.Y(n_8938)
);

BUFx3_ASAP7_75t_L g8939 ( 
.A(n_8467),
.Y(n_8939)
);

A2O1A1Ixp33_ASAP7_75t_L g8940 ( 
.A1(n_8453),
.A2(n_8374),
.B(n_8479),
.C(n_8457),
.Y(n_8940)
);

O2A1O1Ixp33_ASAP7_75t_L g8941 ( 
.A1(n_8338),
.A2(n_363),
.B(n_361),
.C(n_362),
.Y(n_8941)
);

A2O1A1Ixp33_ASAP7_75t_L g8942 ( 
.A1(n_8381),
.A2(n_968),
.B(n_969),
.C(n_967),
.Y(n_8942)
);

BUFx3_ASAP7_75t_L g8943 ( 
.A(n_8820),
.Y(n_8943)
);

INVx2_ASAP7_75t_SL g8944 ( 
.A(n_8562),
.Y(n_8944)
);

NAND2xp5_ASAP7_75t_L g8945 ( 
.A(n_8683),
.B(n_967),
.Y(n_8945)
);

INVx1_ASAP7_75t_L g8946 ( 
.A(n_8544),
.Y(n_8946)
);

AOI22xp33_ASAP7_75t_L g8947 ( 
.A1(n_8706),
.A2(n_366),
.B1(n_363),
.B2(n_364),
.Y(n_8947)
);

NOR2xp33_ASAP7_75t_L g8948 ( 
.A(n_8793),
.B(n_969),
.Y(n_8948)
);

AOI21xp5_ASAP7_75t_L g8949 ( 
.A1(n_8813),
.A2(n_363),
.B(n_364),
.Y(n_8949)
);

BUFx2_ASAP7_75t_L g8950 ( 
.A(n_8735),
.Y(n_8950)
);

NAND2xp5_ASAP7_75t_SL g8951 ( 
.A(n_8385),
.B(n_8435),
.Y(n_8951)
);

INVx1_ASAP7_75t_SL g8952 ( 
.A(n_8550),
.Y(n_8952)
);

INVx1_ASAP7_75t_L g8953 ( 
.A(n_8557),
.Y(n_8953)
);

NOR2xp33_ASAP7_75t_SL g8954 ( 
.A(n_8340),
.B(n_364),
.Y(n_8954)
);

CKINVDCx5p33_ASAP7_75t_R g8955 ( 
.A(n_8364),
.Y(n_8955)
);

INVx1_ASAP7_75t_SL g8956 ( 
.A(n_8549),
.Y(n_8956)
);

OR2x6_ASAP7_75t_L g8957 ( 
.A(n_8854),
.B(n_970),
.Y(n_8957)
);

INVx2_ASAP7_75t_L g8958 ( 
.A(n_8860),
.Y(n_8958)
);

INVx1_ASAP7_75t_L g8959 ( 
.A(n_8865),
.Y(n_8959)
);

BUFx2_ASAP7_75t_L g8960 ( 
.A(n_8669),
.Y(n_8960)
);

NAND3xp33_ASAP7_75t_L g8961 ( 
.A(n_8349),
.B(n_366),
.C(n_367),
.Y(n_8961)
);

NOR2xp33_ASAP7_75t_L g8962 ( 
.A(n_8593),
.B(n_970),
.Y(n_8962)
);

BUFx2_ASAP7_75t_L g8963 ( 
.A(n_8669),
.Y(n_8963)
);

INVx4_ASAP7_75t_L g8964 ( 
.A(n_8394),
.Y(n_8964)
);

HB1xp67_ASAP7_75t_L g8965 ( 
.A(n_8564),
.Y(n_8965)
);

AOI22xp33_ASAP7_75t_SL g8966 ( 
.A1(n_8696),
.A2(n_368),
.B1(n_366),
.B2(n_367),
.Y(n_8966)
);

BUFx6f_ASAP7_75t_L g8967 ( 
.A(n_8394),
.Y(n_8967)
);

BUFx6f_ASAP7_75t_L g8968 ( 
.A(n_8400),
.Y(n_8968)
);

INVx3_ASAP7_75t_L g8969 ( 
.A(n_8400),
.Y(n_8969)
);

INVxp67_ASAP7_75t_SL g8970 ( 
.A(n_8817),
.Y(n_8970)
);

BUFx2_ASAP7_75t_L g8971 ( 
.A(n_8670),
.Y(n_8971)
);

HB1xp67_ASAP7_75t_L g8972 ( 
.A(n_8583),
.Y(n_8972)
);

INVx1_ASAP7_75t_L g8973 ( 
.A(n_8618),
.Y(n_8973)
);

INVx1_ASAP7_75t_L g8974 ( 
.A(n_8545),
.Y(n_8974)
);

OAI33xp33_ASAP7_75t_L g8975 ( 
.A1(n_8743),
.A2(n_369),
.A3(n_371),
.B1(n_367),
.B2(n_368),
.B3(n_370),
.Y(n_8975)
);

INVx2_ASAP7_75t_SL g8976 ( 
.A(n_8562),
.Y(n_8976)
);

O2A1O1Ixp33_ASAP7_75t_L g8977 ( 
.A1(n_8856),
.A2(n_371),
.B(n_368),
.C(n_369),
.Y(n_8977)
);

AO22x1_ASAP7_75t_L g8978 ( 
.A1(n_8806),
.A2(n_372),
.B1(n_369),
.B2(n_371),
.Y(n_8978)
);

CKINVDCx5p33_ASAP7_75t_R g8979 ( 
.A(n_8602),
.Y(n_8979)
);

AND2x4_ASAP7_75t_L g8980 ( 
.A(n_8681),
.B(n_971),
.Y(n_8980)
);

AND2x2_ASAP7_75t_L g8981 ( 
.A(n_8772),
.B(n_972),
.Y(n_8981)
);

INVx1_ASAP7_75t_SL g8982 ( 
.A(n_8754),
.Y(n_8982)
);

CKINVDCx11_ASAP7_75t_R g8983 ( 
.A(n_8443),
.Y(n_8983)
);

OR2x2_ASAP7_75t_L g8984 ( 
.A(n_8689),
.B(n_972),
.Y(n_8984)
);

INVx3_ASAP7_75t_L g8985 ( 
.A(n_8450),
.Y(n_8985)
);

NAND2xp5_ASAP7_75t_L g8986 ( 
.A(n_8690),
.B(n_973),
.Y(n_8986)
);

OAI22xp5_ASAP7_75t_L g8987 ( 
.A1(n_8371),
.A2(n_375),
.B1(n_373),
.B2(n_374),
.Y(n_8987)
);

O2A1O1Ixp5_ASAP7_75t_L g8988 ( 
.A1(n_8363),
.A2(n_8438),
.B(n_8431),
.C(n_8427),
.Y(n_8988)
);

BUFx6f_ASAP7_75t_L g8989 ( 
.A(n_8450),
.Y(n_8989)
);

NAND2xp5_ASAP7_75t_L g8990 ( 
.A(n_8726),
.B(n_973),
.Y(n_8990)
);

O2A1O1Ixp33_ASAP7_75t_SL g8991 ( 
.A1(n_8399),
.A2(n_375),
.B(n_373),
.C(n_374),
.Y(n_8991)
);

NAND2xp5_ASAP7_75t_L g8992 ( 
.A(n_8718),
.B(n_975),
.Y(n_8992)
);

BUFx6f_ASAP7_75t_L g8993 ( 
.A(n_8460),
.Y(n_8993)
);

BUFx2_ASAP7_75t_L g8994 ( 
.A(n_8734),
.Y(n_8994)
);

NAND2xp5_ASAP7_75t_L g8995 ( 
.A(n_8663),
.B(n_975),
.Y(n_8995)
);

NAND2xp5_ASAP7_75t_L g8996 ( 
.A(n_8678),
.B(n_976),
.Y(n_8996)
);

INVx3_ASAP7_75t_L g8997 ( 
.A(n_8460),
.Y(n_8997)
);

NAND2xp5_ASAP7_75t_L g8998 ( 
.A(n_8720),
.B(n_976),
.Y(n_8998)
);

AND2x4_ASAP7_75t_L g8999 ( 
.A(n_8345),
.B(n_978),
.Y(n_8999)
);

AND2x4_ASAP7_75t_L g9000 ( 
.A(n_8396),
.B(n_979),
.Y(n_9000)
);

OR2x2_ASAP7_75t_L g9001 ( 
.A(n_8724),
.B(n_980),
.Y(n_9001)
);

INVx2_ASAP7_75t_L g9002 ( 
.A(n_8410),
.Y(n_9002)
);

O2A1O1Ixp5_ASAP7_75t_L g9003 ( 
.A1(n_8422),
.A2(n_376),
.B(n_373),
.C(n_375),
.Y(n_9003)
);

AND2x4_ASAP7_75t_L g9004 ( 
.A(n_8432),
.B(n_981),
.Y(n_9004)
);

BUFx6f_ASAP7_75t_L g9005 ( 
.A(n_8477),
.Y(n_9005)
);

A2O1A1Ixp33_ASAP7_75t_L g9006 ( 
.A1(n_8819),
.A2(n_983),
.B(n_984),
.C(n_982),
.Y(n_9006)
);

NAND2xp5_ASAP7_75t_L g9007 ( 
.A(n_8745),
.B(n_982),
.Y(n_9007)
);

AND2x2_ASAP7_75t_L g9008 ( 
.A(n_8510),
.B(n_985),
.Y(n_9008)
);

INVx4_ASAP7_75t_L g9009 ( 
.A(n_8477),
.Y(n_9009)
);

AOI22xp5_ASAP7_75t_L g9010 ( 
.A1(n_8478),
.A2(n_378),
.B1(n_376),
.B2(n_377),
.Y(n_9010)
);

O2A1O1Ixp33_ASAP7_75t_SL g9011 ( 
.A1(n_8397),
.A2(n_379),
.B(n_377),
.C(n_378),
.Y(n_9011)
);

CKINVDCx8_ASAP7_75t_R g9012 ( 
.A(n_8648),
.Y(n_9012)
);

BUFx6f_ASAP7_75t_L g9013 ( 
.A(n_8483),
.Y(n_9013)
);

NAND2xp5_ASAP7_75t_L g9014 ( 
.A(n_8747),
.B(n_985),
.Y(n_9014)
);

HB1xp67_ASAP7_75t_L g9015 ( 
.A(n_8781),
.Y(n_9015)
);

BUFx2_ASAP7_75t_L g9016 ( 
.A(n_8386),
.Y(n_9016)
);

NAND2xp5_ASAP7_75t_L g9017 ( 
.A(n_8748),
.B(n_986),
.Y(n_9017)
);

INVx2_ASAP7_75t_SL g9018 ( 
.A(n_8574),
.Y(n_9018)
);

INVx1_ASAP7_75t_L g9019 ( 
.A(n_8626),
.Y(n_9019)
);

OAI22xp5_ASAP7_75t_L g9020 ( 
.A1(n_8823),
.A2(n_381),
.B1(n_379),
.B2(n_380),
.Y(n_9020)
);

BUFx12f_ASAP7_75t_L g9021 ( 
.A(n_8616),
.Y(n_9021)
);

AOI221xp5_ASAP7_75t_L g9022 ( 
.A1(n_8389),
.A2(n_381),
.B1(n_379),
.B2(n_380),
.C(n_382),
.Y(n_9022)
);

NAND3xp33_ASAP7_75t_L g9023 ( 
.A(n_8757),
.B(n_382),
.C(n_383),
.Y(n_9023)
);

BUFx2_ASAP7_75t_L g9024 ( 
.A(n_8391),
.Y(n_9024)
);

CKINVDCx20_ASAP7_75t_R g9025 ( 
.A(n_8717),
.Y(n_9025)
);

INVx2_ASAP7_75t_SL g9026 ( 
.A(n_8574),
.Y(n_9026)
);

OR2x6_ASAP7_75t_L g9027 ( 
.A(n_8565),
.B(n_987),
.Y(n_9027)
);

HAxp5_ASAP7_75t_L g9028 ( 
.A(n_8640),
.B(n_383),
.CON(n_9028),
.SN(n_9028)
);

INVx3_ASAP7_75t_L g9029 ( 
.A(n_8483),
.Y(n_9029)
);

INVx1_ASAP7_75t_L g9030 ( 
.A(n_8630),
.Y(n_9030)
);

OA21x2_ASAP7_75t_L g9031 ( 
.A1(n_8607),
.A2(n_383),
.B(n_384),
.Y(n_9031)
);

INVx1_ASAP7_75t_L g9032 ( 
.A(n_8647),
.Y(n_9032)
);

BUFx6f_ASAP7_75t_L g9033 ( 
.A(n_8535),
.Y(n_9033)
);

CKINVDCx11_ASAP7_75t_R g9034 ( 
.A(n_8621),
.Y(n_9034)
);

BUFx3_ASAP7_75t_L g9035 ( 
.A(n_8418),
.Y(n_9035)
);

NAND2xp5_ASAP7_75t_L g9036 ( 
.A(n_8740),
.B(n_987),
.Y(n_9036)
);

BUFx2_ASAP7_75t_L g9037 ( 
.A(n_8829),
.Y(n_9037)
);

OR2x6_ASAP7_75t_L g9038 ( 
.A(n_8620),
.B(n_988),
.Y(n_9038)
);

INVx1_ASAP7_75t_SL g9039 ( 
.A(n_8785),
.Y(n_9039)
);

BUFx6f_ASAP7_75t_L g9040 ( 
.A(n_8535),
.Y(n_9040)
);

CKINVDCx20_ASAP7_75t_R g9041 ( 
.A(n_8685),
.Y(n_9041)
);

AO221x1_ASAP7_75t_L g9042 ( 
.A1(n_8804),
.A2(n_386),
.B1(n_384),
.B2(n_385),
.C(n_387),
.Y(n_9042)
);

NOR2xp67_ASAP7_75t_L g9043 ( 
.A(n_8619),
.B(n_386),
.Y(n_9043)
);

OAI22xp5_ASAP7_75t_L g9044 ( 
.A1(n_8826),
.A2(n_388),
.B1(n_386),
.B2(n_387),
.Y(n_9044)
);

INVx3_ASAP7_75t_L g9045 ( 
.A(n_8821),
.Y(n_9045)
);

AND2x4_ASAP7_75t_L g9046 ( 
.A(n_8481),
.B(n_989),
.Y(n_9046)
);

BUFx6f_ASAP7_75t_L g9047 ( 
.A(n_8821),
.Y(n_9047)
);

INVx2_ASAP7_75t_L g9048 ( 
.A(n_8490),
.Y(n_9048)
);

INVx1_ASAP7_75t_L g9049 ( 
.A(n_8655),
.Y(n_9049)
);

NAND2xp5_ASAP7_75t_L g9050 ( 
.A(n_8462),
.B(n_8491),
.Y(n_9050)
);

INVx1_ASAP7_75t_L g9051 ( 
.A(n_8804),
.Y(n_9051)
);

A2O1A1Ixp33_ASAP7_75t_L g9052 ( 
.A1(n_8825),
.A2(n_991),
.B(n_992),
.C(n_990),
.Y(n_9052)
);

NAND2xp5_ASAP7_75t_L g9053 ( 
.A(n_8818),
.B(n_990),
.Y(n_9053)
);

CKINVDCx20_ASAP7_75t_R g9054 ( 
.A(n_8660),
.Y(n_9054)
);

INVx2_ASAP7_75t_L g9055 ( 
.A(n_8822),
.Y(n_9055)
);

OR2x6_ASAP7_75t_L g9056 ( 
.A(n_8620),
.B(n_992),
.Y(n_9056)
);

INVx1_ASAP7_75t_L g9057 ( 
.A(n_8841),
.Y(n_9057)
);

CKINVDCx5p33_ASAP7_75t_R g9058 ( 
.A(n_8357),
.Y(n_9058)
);

AND2x4_ASAP7_75t_L g9059 ( 
.A(n_8846),
.B(n_993),
.Y(n_9059)
);

INVx3_ASAP7_75t_L g9060 ( 
.A(n_8824),
.Y(n_9060)
);

BUFx6f_ASAP7_75t_L g9061 ( 
.A(n_8824),
.Y(n_9061)
);

INVx2_ASAP7_75t_L g9062 ( 
.A(n_8868),
.Y(n_9062)
);

INVx3_ASAP7_75t_L g9063 ( 
.A(n_8470),
.Y(n_9063)
);

BUFx12f_ASAP7_75t_L g9064 ( 
.A(n_8616),
.Y(n_9064)
);

AOI22xp5_ASAP7_75t_L g9065 ( 
.A1(n_8639),
.A2(n_390),
.B1(n_388),
.B2(n_389),
.Y(n_9065)
);

BUFx6f_ASAP7_75t_L g9066 ( 
.A(n_8629),
.Y(n_9066)
);

XOR2xp5_ASAP7_75t_L g9067 ( 
.A(n_8785),
.B(n_8591),
.Y(n_9067)
);

BUFx8_ASAP7_75t_SL g9068 ( 
.A(n_8600),
.Y(n_9068)
);

NAND2xp5_ASAP7_75t_L g9069 ( 
.A(n_8405),
.B(n_995),
.Y(n_9069)
);

BUFx6f_ASAP7_75t_L g9070 ( 
.A(n_8629),
.Y(n_9070)
);

INVx1_ASAP7_75t_L g9071 ( 
.A(n_8787),
.Y(n_9071)
);

OAI22xp5_ASAP7_75t_L g9072 ( 
.A1(n_8505),
.A2(n_391),
.B1(n_388),
.B2(n_389),
.Y(n_9072)
);

NAND2xp5_ASAP7_75t_L g9073 ( 
.A(n_8524),
.B(n_995),
.Y(n_9073)
);

BUFx2_ASAP7_75t_L g9074 ( 
.A(n_8863),
.Y(n_9074)
);

INVx2_ASAP7_75t_L g9075 ( 
.A(n_8559),
.Y(n_9075)
);

NAND2xp5_ASAP7_75t_SL g9076 ( 
.A(n_8673),
.B(n_996),
.Y(n_9076)
);

BUFx6f_ASAP7_75t_L g9077 ( 
.A(n_8591),
.Y(n_9077)
);

BUFx3_ASAP7_75t_L g9078 ( 
.A(n_8600),
.Y(n_9078)
);

AOI21xp5_ASAP7_75t_L g9079 ( 
.A1(n_8762),
.A2(n_8782),
.B(n_8773),
.Y(n_9079)
);

BUFx6f_ASAP7_75t_L g9080 ( 
.A(n_8659),
.Y(n_9080)
);

AOI22xp33_ASAP7_75t_SL g9081 ( 
.A1(n_8382),
.A2(n_393),
.B1(n_391),
.B2(n_392),
.Y(n_9081)
);

HB1xp67_ASAP7_75t_L g9082 ( 
.A(n_8811),
.Y(n_9082)
);

AOI22xp5_ASAP7_75t_L g9083 ( 
.A1(n_8646),
.A2(n_393),
.B1(n_391),
.B2(n_392),
.Y(n_9083)
);

NAND2x2_ASAP7_75t_L g9084 ( 
.A(n_8759),
.B(n_392),
.Y(n_9084)
);

BUFx3_ASAP7_75t_L g9085 ( 
.A(n_8589),
.Y(n_9085)
);

AOI21xp5_ASAP7_75t_L g9086 ( 
.A1(n_8603),
.A2(n_393),
.B(n_394),
.Y(n_9086)
);

INVx1_ASAP7_75t_L g9087 ( 
.A(n_8801),
.Y(n_9087)
);

AOI22xp33_ASAP7_75t_L g9088 ( 
.A1(n_8407),
.A2(n_396),
.B1(n_394),
.B2(n_395),
.Y(n_9088)
);

BUFx3_ASAP7_75t_L g9089 ( 
.A(n_8659),
.Y(n_9089)
);

AOI21xp5_ASAP7_75t_SL g9090 ( 
.A1(n_8828),
.A2(n_998),
.B(n_997),
.Y(n_9090)
);

CKINVDCx8_ASAP7_75t_R g9091 ( 
.A(n_8784),
.Y(n_9091)
);

INVx4_ASAP7_75t_L g9092 ( 
.A(n_8506),
.Y(n_9092)
);

NOR2xp33_ASAP7_75t_R g9093 ( 
.A(n_8560),
.B(n_394),
.Y(n_9093)
);

INVx2_ASAP7_75t_L g9094 ( 
.A(n_8580),
.Y(n_9094)
);

BUFx5_ASAP7_75t_L g9095 ( 
.A(n_8495),
.Y(n_9095)
);

BUFx3_ASAP7_75t_L g9096 ( 
.A(n_8563),
.Y(n_9096)
);

CKINVDCx20_ASAP7_75t_R g9097 ( 
.A(n_8509),
.Y(n_9097)
);

BUFx6f_ASAP7_75t_L g9098 ( 
.A(n_8520),
.Y(n_9098)
);

AND2x2_ASAP7_75t_L g9099 ( 
.A(n_8764),
.B(n_999),
.Y(n_9099)
);

AND2x4_ASAP7_75t_L g9100 ( 
.A(n_8585),
.B(n_8644),
.Y(n_9100)
);

INVx2_ASAP7_75t_L g9101 ( 
.A(n_8617),
.Y(n_9101)
);

BUFx6f_ASAP7_75t_L g9102 ( 
.A(n_8558),
.Y(n_9102)
);

INVx3_ASAP7_75t_L g9103 ( 
.A(n_8668),
.Y(n_9103)
);

NOR2xp33_ASAP7_75t_L g9104 ( 
.A(n_8795),
.B(n_999),
.Y(n_9104)
);

AND2x4_ASAP7_75t_L g9105 ( 
.A(n_8339),
.B(n_1000),
.Y(n_9105)
);

INVx1_ASAP7_75t_L g9106 ( 
.A(n_8808),
.Y(n_9106)
);

NOR2xp67_ASAP7_75t_L g9107 ( 
.A(n_8684),
.B(n_395),
.Y(n_9107)
);

BUFx2_ASAP7_75t_L g9108 ( 
.A(n_8834),
.Y(n_9108)
);

BUFx4_ASAP7_75t_SL g9109 ( 
.A(n_8853),
.Y(n_9109)
);

INVx2_ASAP7_75t_L g9110 ( 
.A(n_8522),
.Y(n_9110)
);

INVx2_ASAP7_75t_L g9111 ( 
.A(n_8533),
.Y(n_9111)
);

INVx2_ASAP7_75t_L g9112 ( 
.A(n_8534),
.Y(n_9112)
);

CKINVDCx5p33_ASAP7_75t_R g9113 ( 
.A(n_8784),
.Y(n_9113)
);

INVx3_ASAP7_75t_L g9114 ( 
.A(n_8858),
.Y(n_9114)
);

INVx2_ASAP7_75t_L g9115 ( 
.A(n_8561),
.Y(n_9115)
);

INVx2_ASAP7_75t_L g9116 ( 
.A(n_8586),
.Y(n_9116)
);

BUFx2_ASAP7_75t_L g9117 ( 
.A(n_8861),
.Y(n_9117)
);

O2A1O1Ixp33_ASAP7_75t_SL g9118 ( 
.A1(n_8361),
.A2(n_397),
.B(n_395),
.C(n_396),
.Y(n_9118)
);

AND2x4_ASAP7_75t_L g9119 ( 
.A(n_8867),
.B(n_1000),
.Y(n_9119)
);

AOI21xp33_ASAP7_75t_L g9120 ( 
.A1(n_8758),
.A2(n_396),
.B(n_397),
.Y(n_9120)
);

OR2x6_ASAP7_75t_L g9121 ( 
.A(n_8853),
.B(n_1001),
.Y(n_9121)
);

AOI22xp33_ASAP7_75t_SL g9122 ( 
.A1(n_8805),
.A2(n_400),
.B1(n_398),
.B2(n_399),
.Y(n_9122)
);

NOR2x1_ASAP7_75t_SL g9123 ( 
.A(n_8704),
.B(n_1002),
.Y(n_9123)
);

AOI21xp5_ASAP7_75t_L g9124 ( 
.A1(n_8469),
.A2(n_398),
.B(n_399),
.Y(n_9124)
);

BUFx3_ASAP7_75t_L g9125 ( 
.A(n_8788),
.Y(n_9125)
);

OR2x6_ASAP7_75t_L g9126 ( 
.A(n_8866),
.B(n_1002),
.Y(n_9126)
);

BUFx12f_ASAP7_75t_L g9127 ( 
.A(n_8866),
.Y(n_9127)
);

NAND2xp5_ASAP7_75t_L g9128 ( 
.A(n_8414),
.B(n_1003),
.Y(n_9128)
);

INVx2_ASAP7_75t_L g9129 ( 
.A(n_8590),
.Y(n_9129)
);

BUFx6f_ASAP7_75t_L g9130 ( 
.A(n_8496),
.Y(n_9130)
);

INVx2_ASAP7_75t_L g9131 ( 
.A(n_8597),
.Y(n_9131)
);

BUFx10_ASAP7_75t_L g9132 ( 
.A(n_8788),
.Y(n_9132)
);

INVx2_ASAP7_75t_L g9133 ( 
.A(n_8606),
.Y(n_9133)
);

AND2x4_ASAP7_75t_L g9134 ( 
.A(n_8737),
.B(n_8814),
.Y(n_9134)
);

BUFx6f_ASAP7_75t_L g9135 ( 
.A(n_8779),
.Y(n_9135)
);

AND2x4_ASAP7_75t_L g9136 ( 
.A(n_8402),
.B(n_1004),
.Y(n_9136)
);

INVx1_ASAP7_75t_L g9137 ( 
.A(n_8815),
.Y(n_9137)
);

BUFx2_ASAP7_75t_SL g9138 ( 
.A(n_8843),
.Y(n_9138)
);

AO21x2_ASAP7_75t_L g9139 ( 
.A1(n_8468),
.A2(n_398),
.B(n_400),
.Y(n_9139)
);

BUFx3_ASAP7_75t_L g9140 ( 
.A(n_8779),
.Y(n_9140)
);

INVx1_ASAP7_75t_L g9141 ( 
.A(n_8416),
.Y(n_9141)
);

INVx2_ASAP7_75t_L g9142 ( 
.A(n_8498),
.Y(n_9142)
);

AND2x4_ASAP7_75t_L g9143 ( 
.A(n_8691),
.B(n_1004),
.Y(n_9143)
);

INVx1_ASAP7_75t_L g9144 ( 
.A(n_8373),
.Y(n_9144)
);

INVx2_ASAP7_75t_L g9145 ( 
.A(n_8500),
.Y(n_9145)
);

OAI22xp5_ASAP7_75t_L g9146 ( 
.A1(n_8476),
.A2(n_403),
.B1(n_401),
.B2(n_402),
.Y(n_9146)
);

AOI22xp5_ASAP7_75t_L g9147 ( 
.A1(n_8760),
.A2(n_403),
.B1(n_401),
.B2(n_402),
.Y(n_9147)
);

INVx3_ASAP7_75t_L g9148 ( 
.A(n_8753),
.Y(n_9148)
);

NOR2xp33_ASAP7_75t_L g9149 ( 
.A(n_8838),
.B(n_1005),
.Y(n_9149)
);

AND2x2_ASAP7_75t_L g9150 ( 
.A(n_8344),
.B(n_8827),
.Y(n_9150)
);

NAND2xp5_ASAP7_75t_L g9151 ( 
.A(n_8346),
.B(n_1005),
.Y(n_9151)
);

AOI21xp5_ASAP7_75t_L g9152 ( 
.A1(n_8707),
.A2(n_401),
.B(n_403),
.Y(n_9152)
);

AND2x2_ASAP7_75t_SL g9153 ( 
.A(n_8441),
.B(n_404),
.Y(n_9153)
);

AND2x6_ASAP7_75t_L g9154 ( 
.A(n_8816),
.B(n_1006),
.Y(n_9154)
);

INVx3_ASAP7_75t_L g9155 ( 
.A(n_8436),
.Y(n_9155)
);

AND2x2_ASAP7_75t_L g9156 ( 
.A(n_8499),
.B(n_1006),
.Y(n_9156)
);

CKINVDCx5p33_ASAP7_75t_R g9157 ( 
.A(n_8702),
.Y(n_9157)
);

OAI22xp5_ASAP7_75t_L g9158 ( 
.A1(n_8425),
.A2(n_406),
.B1(n_404),
.B2(n_405),
.Y(n_9158)
);

BUFx3_ASAP7_75t_L g9159 ( 
.A(n_8587),
.Y(n_9159)
);

OR2x2_ASAP7_75t_L g9160 ( 
.A(n_8390),
.B(n_1007),
.Y(n_9160)
);

AOI22xp33_ASAP7_75t_L g9161 ( 
.A1(n_8716),
.A2(n_406),
.B1(n_404),
.B2(n_405),
.Y(n_9161)
);

BUFx8_ASAP7_75t_L g9162 ( 
.A(n_8492),
.Y(n_9162)
);

AOI22xp5_ASAP7_75t_L g9163 ( 
.A1(n_8551),
.A2(n_407),
.B1(n_405),
.B2(n_406),
.Y(n_9163)
);

CKINVDCx20_ASAP7_75t_R g9164 ( 
.A(n_8614),
.Y(n_9164)
);

BUFx12f_ASAP7_75t_L g9165 ( 
.A(n_8436),
.Y(n_9165)
);

AND2x2_ASAP7_75t_L g9166 ( 
.A(n_8532),
.B(n_1007),
.Y(n_9166)
);

INVx4_ASAP7_75t_L g9167 ( 
.A(n_8667),
.Y(n_9167)
);

NAND2xp5_ASAP7_75t_L g9168 ( 
.A(n_8845),
.B(n_1008),
.Y(n_9168)
);

BUFx6f_ASAP7_75t_L g9169 ( 
.A(n_8472),
.Y(n_9169)
);

AND2x2_ASAP7_75t_L g9170 ( 
.A(n_8623),
.B(n_1008),
.Y(n_9170)
);

NAND2xp5_ASAP7_75t_L g9171 ( 
.A(n_8847),
.B(n_1009),
.Y(n_9171)
);

BUFx2_ASAP7_75t_L g9172 ( 
.A(n_8517),
.Y(n_9172)
);

OAI22xp33_ASAP7_75t_L g9173 ( 
.A1(n_8376),
.A2(n_409),
.B1(n_407),
.B2(n_408),
.Y(n_9173)
);

INVx2_ASAP7_75t_L g9174 ( 
.A(n_8502),
.Y(n_9174)
);

INVx3_ASAP7_75t_L g9175 ( 
.A(n_8472),
.Y(n_9175)
);

NOR2x1_ASAP7_75t_SL g9176 ( 
.A(n_8356),
.B(n_1009),
.Y(n_9176)
);

BUFx2_ASAP7_75t_SL g9177 ( 
.A(n_8540),
.Y(n_9177)
);

NOR2xp33_ASAP7_75t_L g9178 ( 
.A(n_8700),
.B(n_1010),
.Y(n_9178)
);

NOR2xp67_ASAP7_75t_L g9179 ( 
.A(n_8849),
.B(n_407),
.Y(n_9179)
);

AND2x4_ASAP7_75t_L g9180 ( 
.A(n_8358),
.B(n_1010),
.Y(n_9180)
);

INVx3_ASAP7_75t_L g9181 ( 
.A(n_8667),
.Y(n_9181)
);

BUFx12f_ASAP7_75t_L g9182 ( 
.A(n_8641),
.Y(n_9182)
);

AOI222xp33_ASAP7_75t_L g9183 ( 
.A1(n_8682),
.A2(n_410),
.B1(n_412),
.B2(n_408),
.C1(n_409),
.C2(n_411),
.Y(n_9183)
);

INVx2_ASAP7_75t_L g9184 ( 
.A(n_8516),
.Y(n_9184)
);

INVx4_ASAP7_75t_L g9185 ( 
.A(n_8750),
.Y(n_9185)
);

INVx1_ASAP7_75t_L g9186 ( 
.A(n_8547),
.Y(n_9186)
);

INVx1_ASAP7_75t_L g9187 ( 
.A(n_8658),
.Y(n_9187)
);

INVx6_ASAP7_75t_SL g9188 ( 
.A(n_8413),
.Y(n_9188)
);

NOR2xp33_ASAP7_75t_L g9189 ( 
.A(n_8348),
.B(n_1011),
.Y(n_9189)
);

AOI22xp5_ASAP7_75t_L g9190 ( 
.A1(n_8652),
.A2(n_412),
.B1(n_409),
.B2(n_410),
.Y(n_9190)
);

AOI22xp5_ASAP7_75t_L g9191 ( 
.A1(n_8571),
.A2(n_413),
.B1(n_410),
.B2(n_412),
.Y(n_9191)
);

OR2x6_ASAP7_75t_L g9192 ( 
.A(n_8347),
.B(n_1011),
.Y(n_9192)
);

BUFx2_ASAP7_75t_L g9193 ( 
.A(n_8342),
.Y(n_9193)
);

BUFx3_ASAP7_75t_L g9194 ( 
.A(n_8705),
.Y(n_9194)
);

INVx8_ASAP7_75t_L g9195 ( 
.A(n_8624),
.Y(n_9195)
);

OR2x6_ASAP7_75t_L g9196 ( 
.A(n_8831),
.B(n_1012),
.Y(n_9196)
);

BUFx6f_ASAP7_75t_L g9197 ( 
.A(n_8519),
.Y(n_9197)
);

NAND2x1p5_ASAP7_75t_L g9198 ( 
.A(n_8369),
.B(n_1013),
.Y(n_9198)
);

OAI22xp5_ASAP7_75t_L g9199 ( 
.A1(n_8403),
.A2(n_415),
.B1(n_413),
.B2(n_414),
.Y(n_9199)
);

INVx3_ASAP7_75t_L g9200 ( 
.A(n_8525),
.Y(n_9200)
);

INVx2_ASAP7_75t_L g9201 ( 
.A(n_8628),
.Y(n_9201)
);

INVx1_ASAP7_75t_L g9202 ( 
.A(n_8645),
.Y(n_9202)
);

INVx3_ASAP7_75t_L g9203 ( 
.A(n_8579),
.Y(n_9203)
);

INVx2_ASAP7_75t_SL g9204 ( 
.A(n_8776),
.Y(n_9204)
);

BUFx6f_ASAP7_75t_L g9205 ( 
.A(n_8554),
.Y(n_9205)
);

AND2x4_ASAP7_75t_L g9206 ( 
.A(n_8411),
.B(n_1013),
.Y(n_9206)
);

INVx1_ASAP7_75t_L g9207 ( 
.A(n_8576),
.Y(n_9207)
);

INVx2_ASAP7_75t_L g9208 ( 
.A(n_8674),
.Y(n_9208)
);

AND2x2_ASAP7_75t_L g9209 ( 
.A(n_8642),
.B(n_1014),
.Y(n_9209)
);

BUFx4f_ASAP7_75t_L g9210 ( 
.A(n_8799),
.Y(n_9210)
);

INVx2_ASAP7_75t_L g9211 ( 
.A(n_8850),
.Y(n_9211)
);

AO21x2_ASAP7_75t_L g9212 ( 
.A1(n_8746),
.A2(n_413),
.B(n_414),
.Y(n_9212)
);

BUFx12f_ASAP7_75t_L g9213 ( 
.A(n_8789),
.Y(n_9213)
);

A2O1A1Ixp33_ASAP7_75t_L g9214 ( 
.A1(n_8837),
.A2(n_1015),
.B(n_1016),
.C(n_1014),
.Y(n_9214)
);

OAI22xp5_ASAP7_75t_L g9215 ( 
.A1(n_8368),
.A2(n_417),
.B1(n_415),
.B2(n_416),
.Y(n_9215)
);

BUFx5_ASAP7_75t_L g9216 ( 
.A(n_8666),
.Y(n_9216)
);

INVx2_ASAP7_75t_L g9217 ( 
.A(n_8855),
.Y(n_9217)
);

INVx1_ASAP7_75t_L g9218 ( 
.A(n_8763),
.Y(n_9218)
);

INVx1_ASAP7_75t_L g9219 ( 
.A(n_8465),
.Y(n_9219)
);

INVx1_ASAP7_75t_L g9220 ( 
.A(n_8599),
.Y(n_9220)
);

INVx3_ASAP7_75t_L g9221 ( 
.A(n_8738),
.Y(n_9221)
);

CKINVDCx8_ASAP7_75t_R g9222 ( 
.A(n_8833),
.Y(n_9222)
);

BUFx2_ASAP7_75t_L g9223 ( 
.A(n_8725),
.Y(n_9223)
);

OAI21x1_ASAP7_75t_SL g9224 ( 
.A1(n_8733),
.A2(n_416),
.B(n_417),
.Y(n_9224)
);

INVx2_ASAP7_75t_L g9225 ( 
.A(n_8859),
.Y(n_9225)
);

INVx8_ASAP7_75t_L g9226 ( 
.A(n_8649),
.Y(n_9226)
);

NAND2xp5_ASAP7_75t_L g9227 ( 
.A(n_8869),
.B(n_1015),
.Y(n_9227)
);

BUFx2_ASAP7_75t_SL g9228 ( 
.A(n_8515),
.Y(n_9228)
);

INVx1_ASAP7_75t_SL g9229 ( 
.A(n_8474),
.Y(n_9229)
);

BUFx3_ASAP7_75t_L g9230 ( 
.A(n_8350),
.Y(n_9230)
);

INVx1_ASAP7_75t_L g9231 ( 
.A(n_8631),
.Y(n_9231)
);

NOR2xp33_ASAP7_75t_SL g9232 ( 
.A(n_8848),
.B(n_418),
.Y(n_9232)
);

AND2x2_ASAP7_75t_L g9233 ( 
.A(n_8392),
.B(n_8488),
.Y(n_9233)
);

CKINVDCx6p67_ASAP7_75t_R g9234 ( 
.A(n_8774),
.Y(n_9234)
);

CKINVDCx14_ASAP7_75t_R g9235 ( 
.A(n_8765),
.Y(n_9235)
);

INVx1_ASAP7_75t_L g9236 ( 
.A(n_8661),
.Y(n_9236)
);

NAND2xp5_ASAP7_75t_SL g9237 ( 
.A(n_8835),
.B(n_1016),
.Y(n_9237)
);

CKINVDCx11_ASAP7_75t_R g9238 ( 
.A(n_8812),
.Y(n_9238)
);

INVx2_ASAP7_75t_L g9239 ( 
.A(n_8383),
.Y(n_9239)
);

OAI22xp5_ASAP7_75t_L g9240 ( 
.A1(n_8622),
.A2(n_8463),
.B1(n_8507),
.B2(n_8842),
.Y(n_9240)
);

BUFx2_ASAP7_75t_L g9241 ( 
.A(n_8566),
.Y(n_9241)
);

OAI22xp5_ASAP7_75t_L g9242 ( 
.A1(n_8844),
.A2(n_420),
.B1(n_418),
.B2(n_419),
.Y(n_9242)
);

BUFx4f_ASAP7_75t_L g9243 ( 
.A(n_8384),
.Y(n_9243)
);

BUFx3_ASAP7_75t_L g9244 ( 
.A(n_8352),
.Y(n_9244)
);

INVx1_ASAP7_75t_L g9245 ( 
.A(n_8756),
.Y(n_9245)
);

AND2x4_ASAP7_75t_L g9246 ( 
.A(n_8679),
.B(n_1017),
.Y(n_9246)
);

INVx1_ASAP7_75t_L g9247 ( 
.A(n_8777),
.Y(n_9247)
);

BUFx3_ASAP7_75t_L g9248 ( 
.A(n_8372),
.Y(n_9248)
);

BUFx3_ASAP7_75t_L g9249 ( 
.A(n_8415),
.Y(n_9249)
);

NOR2xp33_ASAP7_75t_L g9250 ( 
.A(n_8851),
.B(n_1017),
.Y(n_9250)
);

INVxp67_ASAP7_75t_L g9251 ( 
.A(n_8857),
.Y(n_9251)
);

OAI22xp5_ASAP7_75t_L g9252 ( 
.A1(n_8852),
.A2(n_420),
.B1(n_418),
.B2(n_419),
.Y(n_9252)
);

INVx1_ASAP7_75t_L g9253 ( 
.A(n_8780),
.Y(n_9253)
);

BUFx12f_ASAP7_75t_L g9254 ( 
.A(n_8398),
.Y(n_9254)
);

BUFx4f_ASAP7_75t_L g9255 ( 
.A(n_8742),
.Y(n_9255)
);

INVx1_ASAP7_75t_L g9256 ( 
.A(n_8783),
.Y(n_9256)
);

INVx1_ASAP7_75t_L g9257 ( 
.A(n_8792),
.Y(n_9257)
);

BUFx3_ASAP7_75t_L g9258 ( 
.A(n_8654),
.Y(n_9258)
);

INVx2_ASAP7_75t_L g9259 ( 
.A(n_8798),
.Y(n_9259)
);

NAND2xp5_ASAP7_75t_L g9260 ( 
.A(n_8501),
.B(n_1018),
.Y(n_9260)
);

AOI22xp33_ASAP7_75t_SL g9261 ( 
.A1(n_8444),
.A2(n_423),
.B1(n_421),
.B2(n_422),
.Y(n_9261)
);

BUFx6f_ASAP7_75t_L g9262 ( 
.A(n_8672),
.Y(n_9262)
);

AND2x4_ASAP7_75t_L g9263 ( 
.A(n_8584),
.B(n_1018),
.Y(n_9263)
);

INVx2_ASAP7_75t_L g9264 ( 
.A(n_8699),
.Y(n_9264)
);

INVx1_ASAP7_75t_L g9265 ( 
.A(n_8832),
.Y(n_9265)
);

AOI22xp33_ASAP7_75t_L g9266 ( 
.A1(n_8596),
.A2(n_424),
.B1(n_422),
.B2(n_423),
.Y(n_9266)
);

INVx1_ASAP7_75t_L g9267 ( 
.A(n_8840),
.Y(n_9267)
);

HB1xp67_ASAP7_75t_L g9268 ( 
.A(n_8769),
.Y(n_9268)
);

A2O1A1Ixp33_ASAP7_75t_SL g9269 ( 
.A1(n_8802),
.A2(n_427),
.B(n_423),
.C(n_426),
.Y(n_9269)
);

AND2x2_ASAP7_75t_L g9270 ( 
.A(n_8719),
.B(n_1019),
.Y(n_9270)
);

INVx1_ASAP7_75t_L g9271 ( 
.A(n_8744),
.Y(n_9271)
);

NAND2xp5_ASAP7_75t_L g9272 ( 
.A(n_8504),
.B(n_1020),
.Y(n_9272)
);

AND2x2_ASAP7_75t_L g9273 ( 
.A(n_8732),
.B(n_1021),
.Y(n_9273)
);

AOI21xp5_ASAP7_75t_L g9274 ( 
.A1(n_8461),
.A2(n_426),
.B(n_427),
.Y(n_9274)
);

INVx5_ASAP7_75t_L g9275 ( 
.A(n_8471),
.Y(n_9275)
);

BUFx6f_ASAP7_75t_L g9276 ( 
.A(n_8701),
.Y(n_9276)
);

BUFx6f_ASAP7_75t_L g9277 ( 
.A(n_8723),
.Y(n_9277)
);

A2O1A1Ixp33_ASAP7_75t_L g9278 ( 
.A1(n_8870),
.A2(n_1023),
.B(n_1024),
.C(n_1022),
.Y(n_9278)
);

INVx1_ASAP7_75t_L g9279 ( 
.A(n_8553),
.Y(n_9279)
);

AND2x4_ASAP7_75t_L g9280 ( 
.A(n_8686),
.B(n_1024),
.Y(n_9280)
);

INVx1_ASAP7_75t_L g9281 ( 
.A(n_8608),
.Y(n_9281)
);

OAI22xp5_ASAP7_75t_L g9282 ( 
.A1(n_8862),
.A2(n_429),
.B1(n_426),
.B2(n_428),
.Y(n_9282)
);

OAI22xp33_ASAP7_75t_L g9283 ( 
.A1(n_8632),
.A2(n_8657),
.B1(n_8714),
.B2(n_8448),
.Y(n_9283)
);

NAND2xp5_ASAP7_75t_L g9284 ( 
.A(n_8864),
.B(n_1026),
.Y(n_9284)
);

INVx2_ASAP7_75t_L g9285 ( 
.A(n_8727),
.Y(n_9285)
);

O2A1O1Ixp5_ASAP7_75t_SL g9286 ( 
.A1(n_8676),
.A2(n_431),
.B(n_429),
.C(n_430),
.Y(n_9286)
);

BUFx6f_ASAP7_75t_L g9287 ( 
.A(n_8736),
.Y(n_9287)
);

INVx2_ASAP7_75t_L g9288 ( 
.A(n_8749),
.Y(n_9288)
);

INVx2_ASAP7_75t_L g9289 ( 
.A(n_8359),
.Y(n_9289)
);

INVx1_ASAP7_75t_L g9290 ( 
.A(n_8771),
.Y(n_9290)
);

AOI21xp5_ASAP7_75t_SL g9291 ( 
.A1(n_8541),
.A2(n_1027),
.B(n_1026),
.Y(n_9291)
);

OAI22xp5_ASAP7_75t_L g9292 ( 
.A1(n_8578),
.A2(n_8475),
.B1(n_8786),
.B2(n_8592),
.Y(n_9292)
);

INVx1_ASAP7_75t_SL g9293 ( 
.A(n_8466),
.Y(n_9293)
);

BUFx2_ASAP7_75t_SL g9294 ( 
.A(n_8412),
.Y(n_9294)
);

INVx3_ASAP7_75t_L g9295 ( 
.A(n_8807),
.Y(n_9295)
);

NOR4xp25_ASAP7_75t_L g9296 ( 
.A(n_8728),
.B(n_431),
.C(n_429),
.D(n_430),
.Y(n_9296)
);

INVx2_ASAP7_75t_L g9297 ( 
.A(n_8665),
.Y(n_9297)
);

BUFx3_ASAP7_75t_L g9298 ( 
.A(n_8615),
.Y(n_9298)
);

BUFx2_ASAP7_75t_L g9299 ( 
.A(n_8604),
.Y(n_9299)
);

AO21x1_ASAP7_75t_L g9300 ( 
.A1(n_8636),
.A2(n_430),
.B(n_431),
.Y(n_9300)
);

NAND2xp5_ASAP7_75t_L g9301 ( 
.A(n_8480),
.B(n_1028),
.Y(n_9301)
);

AOI21xp33_ASAP7_75t_L g9302 ( 
.A1(n_8539),
.A2(n_432),
.B(n_433),
.Y(n_9302)
);

INVx4_ASAP7_75t_L g9303 ( 
.A(n_8588),
.Y(n_9303)
);

AND2x2_ASAP7_75t_L g9304 ( 
.A(n_8546),
.B(n_1028),
.Y(n_9304)
);

INVx1_ASAP7_75t_L g9305 ( 
.A(n_8712),
.Y(n_9305)
);

INVx5_ASAP7_75t_L g9306 ( 
.A(n_8797),
.Y(n_9306)
);

NAND2xp5_ASAP7_75t_L g9307 ( 
.A(n_8489),
.B(n_1029),
.Y(n_9307)
);

AOI21xp5_ASAP7_75t_L g9308 ( 
.A1(n_8543),
.A2(n_432),
.B(n_433),
.Y(n_9308)
);

INVx1_ASAP7_75t_L g9309 ( 
.A(n_8715),
.Y(n_9309)
);

HB1xp67_ASAP7_75t_L g9310 ( 
.A(n_8810),
.Y(n_9310)
);

INVx2_ASAP7_75t_SL g9311 ( 
.A(n_8455),
.Y(n_9311)
);

AND2x6_ASAP7_75t_L g9312 ( 
.A(n_8664),
.B(n_1029),
.Y(n_9312)
);

OR2x6_ASAP7_75t_L g9313 ( 
.A(n_8601),
.B(n_1030),
.Y(n_9313)
);

NAND2xp5_ASAP7_75t_L g9314 ( 
.A(n_8731),
.B(n_1030),
.Y(n_9314)
);

INVx1_ASAP7_75t_L g9315 ( 
.A(n_8739),
.Y(n_9315)
);

HB1xp67_ASAP7_75t_L g9316 ( 
.A(n_8741),
.Y(n_9316)
);

INVx1_ASAP7_75t_SL g9317 ( 
.A(n_8613),
.Y(n_9317)
);

INVx1_ASAP7_75t_L g9318 ( 
.A(n_8730),
.Y(n_9318)
);

NOR2xp33_ASAP7_75t_L g9319 ( 
.A(n_8567),
.B(n_1031),
.Y(n_9319)
);

INVx1_ASAP7_75t_L g9320 ( 
.A(n_8635),
.Y(n_9320)
);

INVx2_ASAP7_75t_L g9321 ( 
.A(n_8694),
.Y(n_9321)
);

CKINVDCx5p33_ASAP7_75t_R g9322 ( 
.A(n_8879),
.Y(n_9322)
);

AND2x4_ASAP7_75t_L g9323 ( 
.A(n_8919),
.B(n_8638),
.Y(n_9323)
);

AOI21xp5_ASAP7_75t_L g9324 ( 
.A1(n_9079),
.A2(n_8395),
.B(n_8778),
.Y(n_9324)
);

INVx8_ASAP7_75t_L g9325 ( 
.A(n_8871),
.Y(n_9325)
);

AND2x4_ASAP7_75t_L g9326 ( 
.A(n_8903),
.B(n_8528),
.Y(n_9326)
);

O2A1O1Ixp33_ASAP7_75t_L g9327 ( 
.A1(n_8940),
.A2(n_8439),
.B(n_8581),
.C(n_8573),
.Y(n_9327)
);

AOI21xp5_ASAP7_75t_L g9328 ( 
.A1(n_8897),
.A2(n_8424),
.B(n_8513),
.Y(n_9328)
);

AND2x2_ASAP7_75t_SL g9329 ( 
.A(n_9255),
.B(n_8464),
.Y(n_9329)
);

INVx2_ASAP7_75t_L g9330 ( 
.A(n_8885),
.Y(n_9330)
);

BUFx2_ASAP7_75t_L g9331 ( 
.A(n_8950),
.Y(n_9331)
);

AND2x2_ASAP7_75t_L g9332 ( 
.A(n_8875),
.B(n_8594),
.Y(n_9332)
);

INVxp67_ASAP7_75t_L g9333 ( 
.A(n_8938),
.Y(n_9333)
);

OR2x6_ASAP7_75t_L g9334 ( 
.A(n_8934),
.B(n_8366),
.Y(n_9334)
);

NOR2xp67_ASAP7_75t_SL g9335 ( 
.A(n_9090),
.B(n_8653),
.Y(n_9335)
);

OR2x2_ASAP7_75t_L g9336 ( 
.A(n_9137),
.B(n_8598),
.Y(n_9336)
);

BUFx4f_ASAP7_75t_L g9337 ( 
.A(n_9135),
.Y(n_9337)
);

INVx1_ASAP7_75t_L g9338 ( 
.A(n_8965),
.Y(n_9338)
);

NAND2xp5_ASAP7_75t_SL g9339 ( 
.A(n_9306),
.B(n_8687),
.Y(n_9339)
);

INVx1_ASAP7_75t_L g9340 ( 
.A(n_8972),
.Y(n_9340)
);

INVx1_ASAP7_75t_SL g9341 ( 
.A(n_8982),
.Y(n_9341)
);

AOI21xp5_ASAP7_75t_L g9342 ( 
.A1(n_8951),
.A2(n_8482),
.B(n_8487),
.Y(n_9342)
);

NAND3xp33_ASAP7_75t_L g9343 ( 
.A(n_8988),
.B(n_8709),
.C(n_8697),
.Y(n_9343)
);

AND2x4_ASAP7_75t_L g9344 ( 
.A(n_8920),
.B(n_8529),
.Y(n_9344)
);

XNOR2xp5_ASAP7_75t_L g9345 ( 
.A(n_8955),
.B(n_8791),
.Y(n_9345)
);

INVx3_ASAP7_75t_SL g9346 ( 
.A(n_8878),
.Y(n_9346)
);

NAND2xp5_ASAP7_75t_L g9347 ( 
.A(n_8905),
.B(n_8688),
.Y(n_9347)
);

AOI21xp5_ASAP7_75t_L g9348 ( 
.A1(n_9023),
.A2(n_8353),
.B(n_8514),
.Y(n_9348)
);

INVx2_ASAP7_75t_L g9349 ( 
.A(n_8886),
.Y(n_9349)
);

INVx1_ASAP7_75t_L g9350 ( 
.A(n_8884),
.Y(n_9350)
);

AND2x2_ASAP7_75t_L g9351 ( 
.A(n_8882),
.B(n_8693),
.Y(n_9351)
);

AND2x4_ASAP7_75t_L g9352 ( 
.A(n_8935),
.B(n_8572),
.Y(n_9352)
);

OAI22xp5_ASAP7_75t_L g9353 ( 
.A1(n_8872),
.A2(n_8708),
.B1(n_8721),
.B2(n_8627),
.Y(n_9353)
);

INVx3_ASAP7_75t_SL g9354 ( 
.A(n_8979),
.Y(n_9354)
);

NAND2x1p5_ASAP7_75t_L g9355 ( 
.A(n_8895),
.B(n_8675),
.Y(n_9355)
);

AOI21xp5_ASAP7_75t_L g9356 ( 
.A1(n_8931),
.A2(n_8521),
.B(n_8503),
.Y(n_9356)
);

INVx4_ASAP7_75t_L g9357 ( 
.A(n_9113),
.Y(n_9357)
);

BUFx2_ASAP7_75t_SL g9358 ( 
.A(n_8939),
.Y(n_9358)
);

AND2x2_ASAP7_75t_L g9359 ( 
.A(n_8960),
.B(n_8518),
.Y(n_9359)
);

INVx3_ASAP7_75t_L g9360 ( 
.A(n_8896),
.Y(n_9360)
);

OAI21xp33_ASAP7_75t_L g9361 ( 
.A1(n_9296),
.A2(n_8722),
.B(n_8428),
.Y(n_9361)
);

OR2x2_ASAP7_75t_L g9362 ( 
.A(n_9071),
.B(n_8486),
.Y(n_9362)
);

NAND2xp5_ASAP7_75t_L g9363 ( 
.A(n_8974),
.B(n_8677),
.Y(n_9363)
);

OR2x2_ASAP7_75t_L g9364 ( 
.A(n_9087),
.B(n_8711),
.Y(n_9364)
);

INVx3_ASAP7_75t_L g9365 ( 
.A(n_9091),
.Y(n_9365)
);

BUFx6f_ASAP7_75t_L g9366 ( 
.A(n_8914),
.Y(n_9366)
);

OR2x2_ASAP7_75t_L g9367 ( 
.A(n_9082),
.B(n_8713),
.Y(n_9367)
);

AOI22xp33_ASAP7_75t_L g9368 ( 
.A1(n_9095),
.A2(n_8625),
.B1(n_8605),
.B2(n_8527),
.Y(n_9368)
);

INVx2_ASAP7_75t_L g9369 ( 
.A(n_8893),
.Y(n_9369)
);

AND2x2_ASAP7_75t_L g9370 ( 
.A(n_8963),
.B(n_8531),
.Y(n_9370)
);

OAI22xp5_ASAP7_75t_L g9371 ( 
.A1(n_8966),
.A2(n_8542),
.B1(n_8796),
.B2(n_8794),
.Y(n_9371)
);

BUFx12f_ASAP7_75t_L g9372 ( 
.A(n_9058),
.Y(n_9372)
);

BUFx2_ASAP7_75t_L g9373 ( 
.A(n_8971),
.Y(n_9373)
);

AND2x6_ASAP7_75t_L g9374 ( 
.A(n_9290),
.B(n_8768),
.Y(n_9374)
);

AND2x2_ASAP7_75t_L g9375 ( 
.A(n_8956),
.B(n_8451),
.Y(n_9375)
);

AND2x2_ASAP7_75t_L g9376 ( 
.A(n_9200),
.B(n_8703),
.Y(n_9376)
);

INVx1_ASAP7_75t_L g9377 ( 
.A(n_8888),
.Y(n_9377)
);

AOI21xp5_ASAP7_75t_L g9378 ( 
.A1(n_8949),
.A2(n_8523),
.B(n_8511),
.Y(n_9378)
);

NAND2xp5_ASAP7_75t_L g9379 ( 
.A(n_9144),
.B(n_8698),
.Y(n_9379)
);

OR2x2_ASAP7_75t_L g9380 ( 
.A(n_8970),
.B(n_8751),
.Y(n_9380)
);

AND2x2_ASAP7_75t_L g9381 ( 
.A(n_9194),
.B(n_8568),
.Y(n_9381)
);

INVx3_ASAP7_75t_L g9382 ( 
.A(n_9096),
.Y(n_9382)
);

A2O1A1Ixp33_ASAP7_75t_L g9383 ( 
.A1(n_8941),
.A2(n_8761),
.B(n_8484),
.C(n_8473),
.Y(n_9383)
);

OAI22xp5_ASAP7_75t_L g9384 ( 
.A1(n_8889),
.A2(n_8610),
.B1(n_8634),
.B2(n_8393),
.Y(n_9384)
);

O2A1O1Ixp33_ASAP7_75t_SL g9385 ( 
.A1(n_9076),
.A2(n_8408),
.B(n_8365),
.C(n_8770),
.Y(n_9385)
);

INVx2_ASAP7_75t_L g9386 ( 
.A(n_8913),
.Y(n_9386)
);

AOI22xp33_ASAP7_75t_L g9387 ( 
.A1(n_9095),
.A2(n_8775),
.B1(n_8651),
.B2(n_8548),
.Y(n_9387)
);

NAND2xp5_ASAP7_75t_L g9388 ( 
.A(n_9245),
.B(n_8454),
.Y(n_9388)
);

INVx2_ASAP7_75t_L g9389 ( 
.A(n_8923),
.Y(n_9389)
);

AOI22xp5_ASAP7_75t_L g9390 ( 
.A1(n_9240),
.A2(n_8656),
.B1(n_8729),
.B2(n_8637),
.Y(n_9390)
);

BUFx10_ASAP7_75t_L g9391 ( 
.A(n_9135),
.Y(n_9391)
);

NAND2x1p5_ASAP7_75t_L g9392 ( 
.A(n_9134),
.B(n_8493),
.Y(n_9392)
);

AND2x2_ASAP7_75t_SL g9393 ( 
.A(n_9193),
.B(n_8839),
.Y(n_9393)
);

BUFx3_ASAP7_75t_L g9394 ( 
.A(n_9021),
.Y(n_9394)
);

NAND2xp5_ASAP7_75t_L g9395 ( 
.A(n_9247),
.B(n_8494),
.Y(n_9395)
);

BUFx3_ASAP7_75t_L g9396 ( 
.A(n_9064),
.Y(n_9396)
);

AND2x4_ASAP7_75t_L g9397 ( 
.A(n_8994),
.B(n_1031),
.Y(n_9397)
);

NAND2x1p5_ASAP7_75t_L g9398 ( 
.A(n_9306),
.B(n_8800),
.Y(n_9398)
);

INVx1_ASAP7_75t_L g9399 ( 
.A(n_8891),
.Y(n_9399)
);

OR2x6_ASAP7_75t_L g9400 ( 
.A(n_8917),
.B(n_8766),
.Y(n_9400)
);

AND2x4_ASAP7_75t_L g9401 ( 
.A(n_9108),
.B(n_1032),
.Y(n_9401)
);

AND2x4_ASAP7_75t_L g9402 ( 
.A(n_9117),
.B(n_1032),
.Y(n_9402)
);

CKINVDCx5p33_ASAP7_75t_R g9403 ( 
.A(n_9041),
.Y(n_9403)
);

INVx4_ASAP7_75t_L g9404 ( 
.A(n_8914),
.Y(n_9404)
);

HB1xp67_ASAP7_75t_L g9405 ( 
.A(n_9015),
.Y(n_9405)
);

BUFx2_ASAP7_75t_L g9406 ( 
.A(n_9016),
.Y(n_9406)
);

OR2x4_ASAP7_75t_L g9407 ( 
.A(n_9149),
.B(n_8575),
.Y(n_9407)
);

AND2x2_ASAP7_75t_L g9408 ( 
.A(n_8874),
.B(n_8582),
.Y(n_9408)
);

INVx1_ASAP7_75t_SL g9409 ( 
.A(n_9039),
.Y(n_9409)
);

OR2x2_ASAP7_75t_L g9410 ( 
.A(n_9049),
.B(n_8809),
.Y(n_9410)
);

INVx1_ASAP7_75t_L g9411 ( 
.A(n_8899),
.Y(n_9411)
);

NAND2xp5_ASAP7_75t_L g9412 ( 
.A(n_9253),
.B(n_9256),
.Y(n_9412)
);

AND2x4_ASAP7_75t_L g9413 ( 
.A(n_8873),
.B(n_1033),
.Y(n_9413)
);

INVx1_ASAP7_75t_L g9414 ( 
.A(n_8901),
.Y(n_9414)
);

INVx1_ASAP7_75t_L g9415 ( 
.A(n_8907),
.Y(n_9415)
);

AOI21xp5_ASAP7_75t_L g9416 ( 
.A1(n_8961),
.A2(n_8440),
.B(n_8790),
.Y(n_9416)
);

BUFx2_ASAP7_75t_L g9417 ( 
.A(n_9024),
.Y(n_9417)
);

OAI21xp33_ASAP7_75t_L g9418 ( 
.A1(n_9291),
.A2(n_8497),
.B(n_8609),
.Y(n_9418)
);

INVx1_ASAP7_75t_L g9419 ( 
.A(n_8909),
.Y(n_9419)
);

INVx2_ASAP7_75t_SL g9420 ( 
.A(n_8910),
.Y(n_9420)
);

BUFx2_ASAP7_75t_L g9421 ( 
.A(n_9037),
.Y(n_9421)
);

OR2x6_ASAP7_75t_L g9422 ( 
.A(n_9294),
.B(n_8662),
.Y(n_9422)
);

O2A1O1Ixp33_ASAP7_75t_L g9423 ( 
.A1(n_8942),
.A2(n_434),
.B(n_432),
.C(n_433),
.Y(n_9423)
);

OR2x2_ASAP7_75t_L g9424 ( 
.A(n_9106),
.B(n_1035),
.Y(n_9424)
);

INVx3_ASAP7_75t_SL g9425 ( 
.A(n_9157),
.Y(n_9425)
);

BUFx12f_ASAP7_75t_L g9426 ( 
.A(n_9132),
.Y(n_9426)
);

AO21x2_ASAP7_75t_L g9427 ( 
.A1(n_9141),
.A2(n_434),
.B(n_435),
.Y(n_9427)
);

OAI22xp5_ASAP7_75t_L g9428 ( 
.A1(n_9122),
.A2(n_437),
.B1(n_435),
.B2(n_436),
.Y(n_9428)
);

NOR2xp67_ASAP7_75t_L g9429 ( 
.A(n_8932),
.B(n_435),
.Y(n_9429)
);

BUFx2_ASAP7_75t_SL g9430 ( 
.A(n_9012),
.Y(n_9430)
);

BUFx6f_ASAP7_75t_L g9431 ( 
.A(n_8967),
.Y(n_9431)
);

INVx1_ASAP7_75t_L g9432 ( 
.A(n_8916),
.Y(n_9432)
);

INVx1_ASAP7_75t_L g9433 ( 
.A(n_8927),
.Y(n_9433)
);

OAI21x1_ASAP7_75t_L g9434 ( 
.A1(n_9152),
.A2(n_436),
.B(n_437),
.Y(n_9434)
);

NAND2xp5_ASAP7_75t_L g9435 ( 
.A(n_9257),
.B(n_1035),
.Y(n_9435)
);

INVx3_ASAP7_75t_L g9436 ( 
.A(n_8964),
.Y(n_9436)
);

NOR2xp33_ASAP7_75t_L g9437 ( 
.A(n_9251),
.B(n_1036),
.Y(n_9437)
);

INVx2_ASAP7_75t_L g9438 ( 
.A(n_8937),
.Y(n_9438)
);

BUFx4f_ASAP7_75t_L g9439 ( 
.A(n_9066),
.Y(n_9439)
);

BUFx4f_ASAP7_75t_SL g9440 ( 
.A(n_9025),
.Y(n_9440)
);

OAI22xp5_ASAP7_75t_L g9441 ( 
.A1(n_9147),
.A2(n_438),
.B1(n_436),
.B2(n_437),
.Y(n_9441)
);

INVx1_ASAP7_75t_L g9442 ( 
.A(n_8930),
.Y(n_9442)
);

NOR2x1_ASAP7_75t_L g9443 ( 
.A(n_9223),
.B(n_438),
.Y(n_9443)
);

AOI21xp5_ASAP7_75t_L g9444 ( 
.A1(n_9308),
.A2(n_438),
.B(n_439),
.Y(n_9444)
);

AND2x2_ASAP7_75t_L g9445 ( 
.A(n_9150),
.B(n_1036),
.Y(n_9445)
);

INVx1_ASAP7_75t_L g9446 ( 
.A(n_8946),
.Y(n_9446)
);

AOI21xp5_ASAP7_75t_L g9447 ( 
.A1(n_9274),
.A2(n_439),
.B(n_440),
.Y(n_9447)
);

A2O1A1Ixp33_ASAP7_75t_SL g9448 ( 
.A1(n_9124),
.A2(n_441),
.B(n_439),
.C(n_440),
.Y(n_9448)
);

INVx2_ASAP7_75t_L g9449 ( 
.A(n_8958),
.Y(n_9449)
);

NAND2xp5_ASAP7_75t_L g9450 ( 
.A(n_9259),
.B(n_9218),
.Y(n_9450)
);

INVx2_ASAP7_75t_SL g9451 ( 
.A(n_9078),
.Y(n_9451)
);

BUFx2_ASAP7_75t_L g9452 ( 
.A(n_9074),
.Y(n_9452)
);

INVx1_ASAP7_75t_L g9453 ( 
.A(n_8953),
.Y(n_9453)
);

CKINVDCx5p33_ASAP7_75t_R g9454 ( 
.A(n_9068),
.Y(n_9454)
);

NAND2xp5_ASAP7_75t_L g9455 ( 
.A(n_9211),
.B(n_9217),
.Y(n_9455)
);

BUFx3_ASAP7_75t_L g9456 ( 
.A(n_8911),
.Y(n_9456)
);

NAND2xp5_ASAP7_75t_L g9457 ( 
.A(n_9225),
.B(n_1037),
.Y(n_9457)
);

AND2x2_ASAP7_75t_L g9458 ( 
.A(n_9205),
.B(n_1037),
.Y(n_9458)
);

AOI21xp5_ASAP7_75t_L g9459 ( 
.A1(n_8977),
.A2(n_9210),
.B(n_9283),
.Y(n_9459)
);

NOR2xp33_ASAP7_75t_L g9460 ( 
.A(n_9222),
.B(n_1038),
.Y(n_9460)
);

AOI21xp5_ASAP7_75t_L g9461 ( 
.A1(n_9192),
.A2(n_9196),
.B(n_9118),
.Y(n_9461)
);

NAND2xp5_ASAP7_75t_L g9462 ( 
.A(n_9019),
.B(n_1038),
.Y(n_9462)
);

AOI21xp33_ASAP7_75t_L g9463 ( 
.A1(n_9318),
.A2(n_440),
.B(n_441),
.Y(n_9463)
);

INVx1_ASAP7_75t_L g9464 ( 
.A(n_8959),
.Y(n_9464)
);

OAI22xp5_ASAP7_75t_L g9465 ( 
.A1(n_9243),
.A2(n_444),
.B1(n_442),
.B2(n_443),
.Y(n_9465)
);

INVx1_ASAP7_75t_SL g9466 ( 
.A(n_9238),
.Y(n_9466)
);

AOI21xp5_ASAP7_75t_L g9467 ( 
.A1(n_9237),
.A2(n_9036),
.B(n_9006),
.Y(n_9467)
);

AOI21xp5_ASAP7_75t_L g9468 ( 
.A1(n_9052),
.A2(n_442),
.B(n_443),
.Y(n_9468)
);

CKINVDCx5p33_ASAP7_75t_R g9469 ( 
.A(n_9034),
.Y(n_9469)
);

OR2x6_ASAP7_75t_L g9470 ( 
.A(n_9138),
.B(n_9268),
.Y(n_9470)
);

INVx1_ASAP7_75t_L g9471 ( 
.A(n_8973),
.Y(n_9471)
);

BUFx2_ASAP7_75t_L g9472 ( 
.A(n_9051),
.Y(n_9472)
);

INVx5_ASAP7_75t_L g9473 ( 
.A(n_9154),
.Y(n_9473)
);

NAND2xp5_ASAP7_75t_L g9474 ( 
.A(n_9030),
.B(n_1039),
.Y(n_9474)
);

OAI22xp5_ASAP7_75t_L g9475 ( 
.A1(n_8912),
.A2(n_444),
.B1(n_442),
.B2(n_443),
.Y(n_9475)
);

AOI21xp5_ASAP7_75t_L g9476 ( 
.A1(n_9214),
.A2(n_444),
.B(n_445),
.Y(n_9476)
);

AOI211xp5_ASAP7_75t_L g9477 ( 
.A1(n_8894),
.A2(n_448),
.B(n_446),
.C(n_447),
.Y(n_9477)
);

AND2x2_ASAP7_75t_L g9478 ( 
.A(n_9205),
.B(n_9185),
.Y(n_9478)
);

AOI22xp33_ASAP7_75t_L g9479 ( 
.A1(n_9095),
.A2(n_1040),
.B1(n_1041),
.B2(n_1039),
.Y(n_9479)
);

OAI22xp5_ASAP7_75t_L g9480 ( 
.A1(n_8947),
.A2(n_448),
.B1(n_446),
.B2(n_447),
.Y(n_9480)
);

INVx2_ASAP7_75t_SL g9481 ( 
.A(n_8900),
.Y(n_9481)
);

OR2x2_ASAP7_75t_L g9482 ( 
.A(n_9172),
.B(n_1040),
.Y(n_9482)
);

BUFx3_ASAP7_75t_L g9483 ( 
.A(n_8918),
.Y(n_9483)
);

INVx4_ASAP7_75t_L g9484 ( 
.A(n_8967),
.Y(n_9484)
);

INVx2_ASAP7_75t_L g9485 ( 
.A(n_9032),
.Y(n_9485)
);

INVx2_ASAP7_75t_SL g9486 ( 
.A(n_9140),
.Y(n_9486)
);

INVx2_ASAP7_75t_SL g9487 ( 
.A(n_9125),
.Y(n_9487)
);

AND2x2_ASAP7_75t_L g9488 ( 
.A(n_9204),
.B(n_1041),
.Y(n_9488)
);

NAND2xp5_ASAP7_75t_SL g9489 ( 
.A(n_9303),
.B(n_9197),
.Y(n_9489)
);

AND2x4_ASAP7_75t_L g9490 ( 
.A(n_8876),
.B(n_1042),
.Y(n_9490)
);

INVx2_ASAP7_75t_L g9491 ( 
.A(n_9057),
.Y(n_9491)
);

AOI21xp5_ASAP7_75t_L g9492 ( 
.A1(n_9278),
.A2(n_446),
.B(n_447),
.Y(n_9492)
);

NAND2xp5_ASAP7_75t_L g9493 ( 
.A(n_9142),
.B(n_1042),
.Y(n_9493)
);

AOI222xp33_ASAP7_75t_L g9494 ( 
.A1(n_9022),
.A2(n_451),
.B1(n_453),
.B2(n_449),
.C1(n_450),
.C2(n_452),
.Y(n_9494)
);

OAI22xp33_ASAP7_75t_SL g9495 ( 
.A1(n_9232),
.A2(n_9219),
.B1(n_9231),
.B2(n_9220),
.Y(n_9495)
);

CKINVDCx5p33_ASAP7_75t_R g9496 ( 
.A(n_9054),
.Y(n_9496)
);

AND2x4_ASAP7_75t_L g9497 ( 
.A(n_9002),
.B(n_1044),
.Y(n_9497)
);

OAI21xp5_ASAP7_75t_L g9498 ( 
.A1(n_9003),
.A2(n_449),
.B(n_450),
.Y(n_9498)
);

AND2x6_ASAP7_75t_L g9499 ( 
.A(n_9267),
.B(n_449),
.Y(n_9499)
);

INVx1_ASAP7_75t_L g9500 ( 
.A(n_9048),
.Y(n_9500)
);

NAND2xp5_ASAP7_75t_L g9501 ( 
.A(n_9145),
.B(n_1044),
.Y(n_9501)
);

AND2x2_ASAP7_75t_L g9502 ( 
.A(n_8936),
.B(n_1045),
.Y(n_9502)
);

AND2x4_ASAP7_75t_L g9503 ( 
.A(n_9055),
.B(n_1045),
.Y(n_9503)
);

NAND2xp5_ASAP7_75t_L g9504 ( 
.A(n_9174),
.B(n_1046),
.Y(n_9504)
);

NAND2xp5_ASAP7_75t_SL g9505 ( 
.A(n_9197),
.B(n_1046),
.Y(n_9505)
);

BUFx6f_ASAP7_75t_L g9506 ( 
.A(n_8968),
.Y(n_9506)
);

OAI22xp5_ASAP7_75t_L g9507 ( 
.A1(n_9190),
.A2(n_452),
.B1(n_450),
.B2(n_451),
.Y(n_9507)
);

AND2x2_ASAP7_75t_L g9508 ( 
.A(n_9262),
.B(n_1047),
.Y(n_9508)
);

AOI22xp33_ASAP7_75t_L g9509 ( 
.A1(n_9312),
.A2(n_9241),
.B1(n_9302),
.B2(n_9250),
.Y(n_9509)
);

INVx1_ASAP7_75t_L g9510 ( 
.A(n_9062),
.Y(n_9510)
);

AOI21xp5_ASAP7_75t_L g9511 ( 
.A1(n_9120),
.A2(n_451),
.B(n_452),
.Y(n_9511)
);

CKINVDCx20_ASAP7_75t_R g9512 ( 
.A(n_9097),
.Y(n_9512)
);

INVx1_ASAP7_75t_SL g9513 ( 
.A(n_8952),
.Y(n_9513)
);

AOI21xp5_ASAP7_75t_L g9514 ( 
.A1(n_8991),
.A2(n_453),
.B(n_454),
.Y(n_9514)
);

INVx1_ASAP7_75t_L g9515 ( 
.A(n_9075),
.Y(n_9515)
);

AOI21xp5_ASAP7_75t_L g9516 ( 
.A1(n_9269),
.A2(n_454),
.B(n_455),
.Y(n_9516)
);

AND2x4_ASAP7_75t_L g9517 ( 
.A(n_9094),
.B(n_1048),
.Y(n_9517)
);

CKINVDCx6p67_ASAP7_75t_R g9518 ( 
.A(n_9127),
.Y(n_9518)
);

AOI22xp33_ASAP7_75t_L g9519 ( 
.A1(n_9312),
.A2(n_1050),
.B1(n_1051),
.B2(n_1049),
.Y(n_9519)
);

NOR2xp33_ASAP7_75t_L g9520 ( 
.A(n_9235),
.B(n_1049),
.Y(n_9520)
);

INVx1_ASAP7_75t_SL g9521 ( 
.A(n_9035),
.Y(n_9521)
);

OAI21x1_ASAP7_75t_L g9522 ( 
.A1(n_9208),
.A2(n_454),
.B(n_455),
.Y(n_9522)
);

CKINVDCx20_ASAP7_75t_R g9523 ( 
.A(n_9164),
.Y(n_9523)
);

OAI22xp5_ASAP7_75t_L g9524 ( 
.A1(n_8898),
.A2(n_457),
.B1(n_455),
.B2(n_456),
.Y(n_9524)
);

NAND2xp5_ASAP7_75t_L g9525 ( 
.A(n_9184),
.B(n_1051),
.Y(n_9525)
);

BUFx2_ASAP7_75t_L g9526 ( 
.A(n_9103),
.Y(n_9526)
);

AOI21xp5_ASAP7_75t_L g9527 ( 
.A1(n_8926),
.A2(n_456),
.B(n_457),
.Y(n_9527)
);

BUFx3_ASAP7_75t_L g9528 ( 
.A(n_9066),
.Y(n_9528)
);

AO21x2_ASAP7_75t_L g9529 ( 
.A1(n_9186),
.A2(n_456),
.B(n_457),
.Y(n_9529)
);

AOI21xp5_ASAP7_75t_L g9530 ( 
.A1(n_9313),
.A2(n_458),
.B(n_459),
.Y(n_9530)
);

AOI22xp5_ASAP7_75t_L g9531 ( 
.A1(n_9312),
.A2(n_461),
.B1(n_458),
.B2(n_460),
.Y(n_9531)
);

AND2x4_ASAP7_75t_L g9532 ( 
.A(n_9100),
.B(n_1052),
.Y(n_9532)
);

INVx2_ASAP7_75t_L g9533 ( 
.A(n_9050),
.Y(n_9533)
);

INVx1_ASAP7_75t_L g9534 ( 
.A(n_9187),
.Y(n_9534)
);

AND2x2_ASAP7_75t_L g9535 ( 
.A(n_9262),
.B(n_1052),
.Y(n_9535)
);

NAND2xp5_ASAP7_75t_L g9536 ( 
.A(n_9201),
.B(n_1053),
.Y(n_9536)
);

AOI21xp5_ASAP7_75t_L g9537 ( 
.A1(n_9297),
.A2(n_460),
.B(n_461),
.Y(n_9537)
);

NOR2x1_ASAP7_75t_L g9538 ( 
.A(n_9202),
.B(n_460),
.Y(n_9538)
);

NOR2xp33_ASAP7_75t_SL g9539 ( 
.A(n_9092),
.B(n_1053),
.Y(n_9539)
);

BUFx3_ASAP7_75t_L g9540 ( 
.A(n_9070),
.Y(n_9540)
);

AND2x4_ASAP7_75t_L g9541 ( 
.A(n_9114),
.B(n_9085),
.Y(n_9541)
);

AOI22xp5_ASAP7_75t_L g9542 ( 
.A1(n_9292),
.A2(n_463),
.B1(n_461),
.B2(n_462),
.Y(n_9542)
);

NAND2xp5_ASAP7_75t_L g9543 ( 
.A(n_9110),
.B(n_1054),
.Y(n_9543)
);

NAND2xp5_ASAP7_75t_L g9544 ( 
.A(n_9111),
.B(n_1055),
.Y(n_9544)
);

INVx2_ASAP7_75t_SL g9545 ( 
.A(n_9089),
.Y(n_9545)
);

INVx3_ASAP7_75t_L g9546 ( 
.A(n_9009),
.Y(n_9546)
);

OAI21x1_ASAP7_75t_L g9547 ( 
.A1(n_9221),
.A2(n_462),
.B(n_463),
.Y(n_9547)
);

AND2x2_ASAP7_75t_L g9548 ( 
.A(n_9276),
.B(n_1055),
.Y(n_9548)
);

INVxp67_ASAP7_75t_SL g9549 ( 
.A(n_9207),
.Y(n_9549)
);

NAND2xp5_ASAP7_75t_L g9550 ( 
.A(n_9112),
.B(n_1056),
.Y(n_9550)
);

INVx1_ASAP7_75t_SL g9551 ( 
.A(n_9067),
.Y(n_9551)
);

INVx1_ASAP7_75t_L g9552 ( 
.A(n_9289),
.Y(n_9552)
);

INVx2_ASAP7_75t_L g9553 ( 
.A(n_9115),
.Y(n_9553)
);

AND3x1_ASAP7_75t_SL g9554 ( 
.A(n_9028),
.B(n_462),
.C(n_464),
.Y(n_9554)
);

INVx3_ASAP7_75t_SL g9555 ( 
.A(n_9226),
.Y(n_9555)
);

AOI21xp5_ASAP7_75t_L g9556 ( 
.A1(n_9321),
.A2(n_464),
.B(n_465),
.Y(n_9556)
);

AOI21x1_ASAP7_75t_L g9557 ( 
.A1(n_8978),
.A2(n_465),
.B(n_466),
.Y(n_9557)
);

INVx2_ASAP7_75t_L g9558 ( 
.A(n_9116),
.Y(n_9558)
);

AO21x2_ASAP7_75t_L g9559 ( 
.A1(n_9042),
.A2(n_465),
.B(n_466),
.Y(n_9559)
);

NOR2xp33_ASAP7_75t_SL g9560 ( 
.A(n_9254),
.B(n_1057),
.Y(n_9560)
);

INVx1_ASAP7_75t_L g9561 ( 
.A(n_9279),
.Y(n_9561)
);

BUFx2_ASAP7_75t_L g9562 ( 
.A(n_9148),
.Y(n_9562)
);

AOI21xp5_ASAP7_75t_L g9563 ( 
.A1(n_9300),
.A2(n_467),
.B(n_468),
.Y(n_9563)
);

NAND2xp5_ASAP7_75t_L g9564 ( 
.A(n_9129),
.B(n_1057),
.Y(n_9564)
);

INVx2_ASAP7_75t_SL g9565 ( 
.A(n_9070),
.Y(n_9565)
);

OAI22xp5_ASAP7_75t_L g9566 ( 
.A1(n_8908),
.A2(n_470),
.B1(n_467),
.B2(n_469),
.Y(n_9566)
);

INVx3_ASAP7_75t_L g9567 ( 
.A(n_9098),
.Y(n_9567)
);

BUFx3_ASAP7_75t_L g9568 ( 
.A(n_9077),
.Y(n_9568)
);

NOR2xp67_ASAP7_75t_SL g9569 ( 
.A(n_9275),
.B(n_467),
.Y(n_9569)
);

CKINVDCx6p67_ASAP7_75t_R g9570 ( 
.A(n_8883),
.Y(n_9570)
);

BUFx3_ASAP7_75t_L g9571 ( 
.A(n_9077),
.Y(n_9571)
);

OR2x6_ASAP7_75t_L g9572 ( 
.A(n_9177),
.B(n_1058),
.Y(n_9572)
);

INVxp67_ASAP7_75t_L g9573 ( 
.A(n_9276),
.Y(n_9573)
);

AOI22xp5_ASAP7_75t_L g9574 ( 
.A1(n_9242),
.A2(n_471),
.B1(n_469),
.B2(n_470),
.Y(n_9574)
);

AOI22xp33_ASAP7_75t_L g9575 ( 
.A1(n_9189),
.A2(n_1060),
.B1(n_1061),
.B2(n_1059),
.Y(n_9575)
);

AND2x4_ASAP7_75t_L g9576 ( 
.A(n_9063),
.B(n_1059),
.Y(n_9576)
);

AND2x2_ASAP7_75t_L g9577 ( 
.A(n_9277),
.B(n_1061),
.Y(n_9577)
);

INVx3_ASAP7_75t_SL g9578 ( 
.A(n_9195),
.Y(n_9578)
);

AND2x2_ASAP7_75t_L g9579 ( 
.A(n_9277),
.B(n_1062),
.Y(n_9579)
);

AND2x4_ASAP7_75t_L g9580 ( 
.A(n_8943),
.B(n_1063),
.Y(n_9580)
);

A2O1A1Ixp33_ASAP7_75t_L g9581 ( 
.A1(n_8881),
.A2(n_1065),
.B(n_1066),
.C(n_1064),
.Y(n_9581)
);

INVx1_ASAP7_75t_L g9582 ( 
.A(n_9281),
.Y(n_9582)
);

AOI21xp5_ASAP7_75t_L g9583 ( 
.A1(n_9271),
.A2(n_469),
.B(n_470),
.Y(n_9583)
);

AND2x4_ASAP7_75t_L g9584 ( 
.A(n_8928),
.B(n_1064),
.Y(n_9584)
);

AND2x2_ASAP7_75t_L g9585 ( 
.A(n_9287),
.B(n_1065),
.Y(n_9585)
);

BUFx6f_ASAP7_75t_L g9586 ( 
.A(n_8968),
.Y(n_9586)
);

AND2x2_ASAP7_75t_L g9587 ( 
.A(n_9287),
.B(n_1066),
.Y(n_9587)
);

BUFx4_ASAP7_75t_SL g9588 ( 
.A(n_9121),
.Y(n_9588)
);

AND2x4_ASAP7_75t_L g9589 ( 
.A(n_8969),
.B(n_1067),
.Y(n_9589)
);

AND2x2_ASAP7_75t_L g9590 ( 
.A(n_9258),
.B(n_1067),
.Y(n_9590)
);

INVx1_ASAP7_75t_L g9591 ( 
.A(n_8921),
.Y(n_9591)
);

INVx2_ASAP7_75t_L g9592 ( 
.A(n_9131),
.Y(n_9592)
);

BUFx3_ASAP7_75t_L g9593 ( 
.A(n_9080),
.Y(n_9593)
);

CKINVDCx20_ASAP7_75t_R g9594 ( 
.A(n_8983),
.Y(n_9594)
);

NOR2xp33_ASAP7_75t_SL g9595 ( 
.A(n_9167),
.B(n_1068),
.Y(n_9595)
);

BUFx3_ASAP7_75t_L g9596 ( 
.A(n_9080),
.Y(n_9596)
);

INVx1_ASAP7_75t_L g9597 ( 
.A(n_8929),
.Y(n_9597)
);

CKINVDCx8_ASAP7_75t_R g9598 ( 
.A(n_9130),
.Y(n_9598)
);

BUFx6f_ASAP7_75t_L g9599 ( 
.A(n_8989),
.Y(n_9599)
);

CKINVDCx20_ASAP7_75t_R g9600 ( 
.A(n_9162),
.Y(n_9600)
);

AOI21xp5_ASAP7_75t_L g9601 ( 
.A1(n_9265),
.A2(n_471),
.B(n_472),
.Y(n_9601)
);

BUFx3_ASAP7_75t_L g9602 ( 
.A(n_9130),
.Y(n_9602)
);

INVx8_ASAP7_75t_L g9603 ( 
.A(n_9126),
.Y(n_9603)
);

NAND2xp5_ASAP7_75t_L g9604 ( 
.A(n_9133),
.B(n_1068),
.Y(n_9604)
);

CKINVDCx5p33_ASAP7_75t_R g9605 ( 
.A(n_9109),
.Y(n_9605)
);

NOR2xp33_ASAP7_75t_L g9606 ( 
.A(n_9244),
.B(n_1069),
.Y(n_9606)
);

INVx2_ASAP7_75t_L g9607 ( 
.A(n_9101),
.Y(n_9607)
);

NAND2xp5_ASAP7_75t_L g9608 ( 
.A(n_9295),
.B(n_1069),
.Y(n_9608)
);

BUFx12f_ASAP7_75t_L g9609 ( 
.A(n_8922),
.Y(n_9609)
);

O2A1O1Ixp5_ASAP7_75t_L g9610 ( 
.A1(n_8975),
.A2(n_473),
.B(n_471),
.C(n_472),
.Y(n_9610)
);

INVx1_ASAP7_75t_L g9611 ( 
.A(n_9236),
.Y(n_9611)
);

A2O1A1Ixp33_ASAP7_75t_L g9612 ( 
.A1(n_9086),
.A2(n_1071),
.B(n_1072),
.C(n_1070),
.Y(n_9612)
);

O2A1O1Ixp5_ASAP7_75t_L g9613 ( 
.A1(n_8877),
.A2(n_474),
.B(n_472),
.C(n_473),
.Y(n_9613)
);

BUFx6f_ASAP7_75t_L g9614 ( 
.A(n_8989),
.Y(n_9614)
);

BUFx2_ASAP7_75t_L g9615 ( 
.A(n_9316),
.Y(n_9615)
);

OAI22xp5_ASAP7_75t_L g9616 ( 
.A1(n_9065),
.A2(n_475),
.B1(n_473),
.B2(n_474),
.Y(n_9616)
);

INVx1_ASAP7_75t_SL g9617 ( 
.A(n_9229),
.Y(n_9617)
);

OAI22xp5_ASAP7_75t_L g9618 ( 
.A1(n_9083),
.A2(n_477),
.B1(n_475),
.B2(n_476),
.Y(n_9618)
);

INVx1_ASAP7_75t_L g9619 ( 
.A(n_9310),
.Y(n_9619)
);

OAI21xp33_ASAP7_75t_L g9620 ( 
.A1(n_9010),
.A2(n_475),
.B(n_476),
.Y(n_9620)
);

INVx2_ASAP7_75t_L g9621 ( 
.A(n_8890),
.Y(n_9621)
);

OR2x6_ASAP7_75t_L g9622 ( 
.A(n_9228),
.B(n_1070),
.Y(n_9622)
);

AOI21xp5_ASAP7_75t_L g9623 ( 
.A1(n_9239),
.A2(n_476),
.B(n_477),
.Y(n_9623)
);

OR2x2_ASAP7_75t_L g9624 ( 
.A(n_9264),
.B(n_1071),
.Y(n_9624)
);

OR2x6_ASAP7_75t_L g9625 ( 
.A(n_9299),
.B(n_1072),
.Y(n_9625)
);

INVx1_ASAP7_75t_L g9626 ( 
.A(n_8902),
.Y(n_9626)
);

INVx1_ASAP7_75t_SL g9627 ( 
.A(n_9249),
.Y(n_9627)
);

INVx5_ASAP7_75t_L g9628 ( 
.A(n_9154),
.Y(n_9628)
);

INVx3_ASAP7_75t_L g9629 ( 
.A(n_9098),
.Y(n_9629)
);

NAND2xp5_ASAP7_75t_L g9630 ( 
.A(n_9285),
.B(n_1073),
.Y(n_9630)
);

INVx2_ASAP7_75t_SL g9631 ( 
.A(n_8993),
.Y(n_9631)
);

INVx1_ASAP7_75t_L g9632 ( 
.A(n_9053),
.Y(n_9632)
);

AOI21xp5_ASAP7_75t_L g9633 ( 
.A1(n_9011),
.A2(n_477),
.B(n_478),
.Y(n_9633)
);

BUFx3_ASAP7_75t_L g9634 ( 
.A(n_8993),
.Y(n_9634)
);

AOI21xp5_ASAP7_75t_L g9635 ( 
.A1(n_9252),
.A2(n_478),
.B(n_479),
.Y(n_9635)
);

INVx1_ASAP7_75t_L g9636 ( 
.A(n_9073),
.Y(n_9636)
);

INVx2_ASAP7_75t_L g9637 ( 
.A(n_9216),
.Y(n_9637)
);

AOI21xp5_ASAP7_75t_L g9638 ( 
.A1(n_9282),
.A2(n_478),
.B(n_479),
.Y(n_9638)
);

O2A1O1Ixp5_ASAP7_75t_L g9639 ( 
.A1(n_8880),
.A2(n_482),
.B(n_480),
.C(n_481),
.Y(n_9639)
);

NAND3xp33_ASAP7_75t_L g9640 ( 
.A(n_9183),
.B(n_480),
.C(n_481),
.Y(n_9640)
);

AOI22xp33_ASAP7_75t_L g9641 ( 
.A1(n_9319),
.A2(n_1075),
.B1(n_1076),
.B2(n_1074),
.Y(n_9641)
);

OAI21xp5_ASAP7_75t_L g9642 ( 
.A1(n_9286),
.A2(n_480),
.B(n_481),
.Y(n_9642)
);

INVx2_ASAP7_75t_L g9643 ( 
.A(n_9216),
.Y(n_9643)
);

BUFx8_ASAP7_75t_SL g9644 ( 
.A(n_9165),
.Y(n_9644)
);

INVx2_ASAP7_75t_L g9645 ( 
.A(n_9216),
.Y(n_9645)
);

INVx1_ASAP7_75t_L g9646 ( 
.A(n_8984),
.Y(n_9646)
);

NAND2x1p5_ASAP7_75t_L g9647 ( 
.A(n_9275),
.B(n_1074),
.Y(n_9647)
);

INVxp67_ASAP7_75t_SL g9648 ( 
.A(n_9320),
.Y(n_9648)
);

BUFx6f_ASAP7_75t_L g9649 ( 
.A(n_9005),
.Y(n_9649)
);

INVx1_ASAP7_75t_L g9650 ( 
.A(n_9305),
.Y(n_9650)
);

INVx1_ASAP7_75t_L g9651 ( 
.A(n_9309),
.Y(n_9651)
);

INVx3_ASAP7_75t_L g9652 ( 
.A(n_9102),
.Y(n_9652)
);

INVx2_ASAP7_75t_L g9653 ( 
.A(n_9288),
.Y(n_9653)
);

NAND2xp5_ASAP7_75t_L g9654 ( 
.A(n_9315),
.B(n_1075),
.Y(n_9654)
);

NAND2xp5_ASAP7_75t_L g9655 ( 
.A(n_9293),
.B(n_1077),
.Y(n_9655)
);

INVx2_ASAP7_75t_L g9656 ( 
.A(n_8887),
.Y(n_9656)
);

NAND2xp5_ASAP7_75t_L g9657 ( 
.A(n_9317),
.B(n_1078),
.Y(n_9657)
);

INVx2_ASAP7_75t_SL g9658 ( 
.A(n_9005),
.Y(n_9658)
);

O2A1O1Ixp33_ASAP7_75t_L g9659 ( 
.A1(n_9158),
.A2(n_484),
.B(n_482),
.C(n_483),
.Y(n_9659)
);

O2A1O1Ixp33_ASAP7_75t_L g9660 ( 
.A1(n_9224),
.A2(n_485),
.B(n_483),
.C(n_484),
.Y(n_9660)
);

AOI21xp5_ASAP7_75t_L g9661 ( 
.A1(n_9198),
.A2(n_483),
.B(n_484),
.Y(n_9661)
);

INVx1_ASAP7_75t_L g9662 ( 
.A(n_9001),
.Y(n_9662)
);

AOI21xp5_ASAP7_75t_L g9663 ( 
.A1(n_9123),
.A2(n_485),
.B(n_486),
.Y(n_9663)
);

INVx1_ASAP7_75t_L g9664 ( 
.A(n_8906),
.Y(n_9664)
);

AND2x2_ASAP7_75t_L g9665 ( 
.A(n_9298),
.B(n_1078),
.Y(n_9665)
);

A2O1A1Ixp33_ASAP7_75t_L g9666 ( 
.A1(n_9163),
.A2(n_1080),
.B(n_1081),
.C(n_1079),
.Y(n_9666)
);

INVx2_ASAP7_75t_L g9667 ( 
.A(n_8892),
.Y(n_9667)
);

BUFx2_ASAP7_75t_L g9668 ( 
.A(n_9188),
.Y(n_9668)
);

HB1xp67_ASAP7_75t_L g9669 ( 
.A(n_9180),
.Y(n_9669)
);

AND2x4_ASAP7_75t_L g9670 ( 
.A(n_8985),
.B(n_1079),
.Y(n_9670)
);

OAI22xp5_ASAP7_75t_L g9671 ( 
.A1(n_9161),
.A2(n_487),
.B1(n_485),
.B2(n_486),
.Y(n_9671)
);

NAND2xp5_ASAP7_75t_L g9672 ( 
.A(n_8981),
.B(n_1080),
.Y(n_9672)
);

NOR2xp33_ASAP7_75t_SL g9673 ( 
.A(n_8954),
.B(n_1082),
.Y(n_9673)
);

AND2x4_ASAP7_75t_L g9674 ( 
.A(n_8997),
.B(n_1082),
.Y(n_9674)
);

INVx1_ASAP7_75t_L g9675 ( 
.A(n_8915),
.Y(n_9675)
);

AND2x2_ASAP7_75t_L g9676 ( 
.A(n_9248),
.B(n_1083),
.Y(n_9676)
);

AOI21xp5_ASAP7_75t_L g9677 ( 
.A1(n_9176),
.A2(n_9215),
.B(n_9173),
.Y(n_9677)
);

AND2x4_ASAP7_75t_L g9678 ( 
.A(n_9029),
.B(n_1084),
.Y(n_9678)
);

INVx1_ASAP7_75t_L g9679 ( 
.A(n_8933),
.Y(n_9679)
);

NAND2xp5_ASAP7_75t_L g9680 ( 
.A(n_9153),
.B(n_1084),
.Y(n_9680)
);

INVx4_ASAP7_75t_L g9681 ( 
.A(n_9013),
.Y(n_9681)
);

INVx3_ASAP7_75t_L g9682 ( 
.A(n_9102),
.Y(n_9682)
);

AND2x4_ASAP7_75t_L g9683 ( 
.A(n_9045),
.B(n_9060),
.Y(n_9683)
);

INVx2_ASAP7_75t_SL g9684 ( 
.A(n_9013),
.Y(n_9684)
);

INVx2_ASAP7_75t_L g9685 ( 
.A(n_9311),
.Y(n_9685)
);

AND2x4_ASAP7_75t_L g9686 ( 
.A(n_8944),
.B(n_1085),
.Y(n_9686)
);

INVx2_ASAP7_75t_L g9687 ( 
.A(n_8976),
.Y(n_9687)
);

INVx2_ASAP7_75t_L g9688 ( 
.A(n_9619),
.Y(n_9688)
);

AOI22xp33_ASAP7_75t_SL g9689 ( 
.A1(n_9329),
.A2(n_9093),
.B1(n_9154),
.B2(n_9212),
.Y(n_9689)
);

INVx1_ASAP7_75t_L g9690 ( 
.A(n_9350),
.Y(n_9690)
);

INVx1_ASAP7_75t_SL g9691 ( 
.A(n_9466),
.Y(n_9691)
);

OAI22xp33_ASAP7_75t_L g9692 ( 
.A1(n_9328),
.A2(n_9234),
.B1(n_9191),
.B2(n_9084),
.Y(n_9692)
);

AOI22xp33_ASAP7_75t_L g9693 ( 
.A1(n_9640),
.A2(n_9213),
.B1(n_8962),
.B2(n_9199),
.Y(n_9693)
);

INVx6_ASAP7_75t_L g9694 ( 
.A(n_9391),
.Y(n_9694)
);

BUFx4_ASAP7_75t_SL g9695 ( 
.A(n_9600),
.Y(n_9695)
);

AOI22xp33_ASAP7_75t_L g9696 ( 
.A1(n_9335),
.A2(n_9072),
.B1(n_9146),
.B2(n_9044),
.Y(n_9696)
);

AOI22xp5_ASAP7_75t_L g9697 ( 
.A1(n_9353),
.A2(n_9371),
.B1(n_9418),
.B2(n_9384),
.Y(n_9697)
);

OAI22xp33_ASAP7_75t_L g9698 ( 
.A1(n_9473),
.A2(n_9203),
.B1(n_9020),
.B2(n_9284),
.Y(n_9698)
);

BUFx6f_ASAP7_75t_L g9699 ( 
.A(n_9366),
.Y(n_9699)
);

INVx2_ASAP7_75t_L g9700 ( 
.A(n_9650),
.Y(n_9700)
);

AOI22xp33_ASAP7_75t_SL g9701 ( 
.A1(n_9393),
.A2(n_9495),
.B1(n_9459),
.B2(n_9473),
.Y(n_9701)
);

INVx2_ASAP7_75t_L g9702 ( 
.A(n_9651),
.Y(n_9702)
);

HB1xp67_ASAP7_75t_L g9703 ( 
.A(n_9405),
.Y(n_9703)
);

INVx1_ASAP7_75t_SL g9704 ( 
.A(n_9354),
.Y(n_9704)
);

CKINVDCx20_ASAP7_75t_R g9705 ( 
.A(n_9440),
.Y(n_9705)
);

AOI22xp33_ASAP7_75t_L g9706 ( 
.A1(n_9620),
.A2(n_9178),
.B1(n_8987),
.B2(n_9246),
.Y(n_9706)
);

BUFx4f_ASAP7_75t_L g9707 ( 
.A(n_9372),
.Y(n_9707)
);

INVx6_ASAP7_75t_L g9708 ( 
.A(n_9357),
.Y(n_9708)
);

INVx1_ASAP7_75t_SL g9709 ( 
.A(n_9617),
.Y(n_9709)
);

INVx3_ASAP7_75t_L g9710 ( 
.A(n_9541),
.Y(n_9710)
);

INVx2_ASAP7_75t_L g9711 ( 
.A(n_9552),
.Y(n_9711)
);

INVx1_ASAP7_75t_L g9712 ( 
.A(n_9377),
.Y(n_9712)
);

BUFx2_ASAP7_75t_L g9713 ( 
.A(n_9470),
.Y(n_9713)
);

AOI22xp5_ASAP7_75t_L g9714 ( 
.A1(n_9361),
.A2(n_8904),
.B1(n_9261),
.B2(n_9175),
.Y(n_9714)
);

NAND2x1p5_ASAP7_75t_L g9715 ( 
.A(n_9628),
.B(n_9155),
.Y(n_9715)
);

CKINVDCx20_ASAP7_75t_R g9716 ( 
.A(n_9512),
.Y(n_9716)
);

BUFx10_ASAP7_75t_L g9717 ( 
.A(n_9469),
.Y(n_9717)
);

INVxp67_ASAP7_75t_L g9718 ( 
.A(n_9615),
.Y(n_9718)
);

INVx1_ASAP7_75t_L g9719 ( 
.A(n_9399),
.Y(n_9719)
);

AOI22xp33_ASAP7_75t_L g9720 ( 
.A1(n_9494),
.A2(n_9182),
.B1(n_9230),
.B2(n_9081),
.Y(n_9720)
);

OAI22xp5_ASAP7_75t_L g9721 ( 
.A1(n_9383),
.A2(n_8924),
.B1(n_9266),
.B2(n_9088),
.Y(n_9721)
);

INVx6_ASAP7_75t_L g9722 ( 
.A(n_9426),
.Y(n_9722)
);

CKINVDCx11_ASAP7_75t_R g9723 ( 
.A(n_9594),
.Y(n_9723)
);

AOI22xp5_ASAP7_75t_L g9724 ( 
.A1(n_9390),
.A2(n_9181),
.B1(n_9008),
.B2(n_9143),
.Y(n_9724)
);

BUFx6f_ASAP7_75t_L g9725 ( 
.A(n_9366),
.Y(n_9725)
);

OAI22xp5_ASAP7_75t_L g9726 ( 
.A1(n_9509),
.A2(n_9368),
.B1(n_9628),
.B2(n_9581),
.Y(n_9726)
);

CKINVDCx5p33_ASAP7_75t_R g9727 ( 
.A(n_9403),
.Y(n_9727)
);

INVx2_ASAP7_75t_L g9728 ( 
.A(n_9331),
.Y(n_9728)
);

BUFx2_ASAP7_75t_L g9729 ( 
.A(n_9470),
.Y(n_9729)
);

NAND2xp5_ASAP7_75t_L g9730 ( 
.A(n_9533),
.B(n_9648),
.Y(n_9730)
);

INVx1_ASAP7_75t_L g9731 ( 
.A(n_9411),
.Y(n_9731)
);

AOI21xp5_ASAP7_75t_L g9732 ( 
.A1(n_9324),
.A2(n_9307),
.B(n_9301),
.Y(n_9732)
);

INVx5_ASAP7_75t_L g9733 ( 
.A(n_9572),
.Y(n_9733)
);

BUFx2_ASAP7_75t_L g9734 ( 
.A(n_9406),
.Y(n_9734)
);

OAI22xp5_ASAP7_75t_L g9735 ( 
.A1(n_9387),
.A2(n_9069),
.B1(n_9169),
.B2(n_9314),
.Y(n_9735)
);

INVx4_ASAP7_75t_L g9736 ( 
.A(n_9346),
.Y(n_9736)
);

CKINVDCx6p67_ASAP7_75t_R g9737 ( 
.A(n_9425),
.Y(n_9737)
);

INVx3_ASAP7_75t_L g9738 ( 
.A(n_9528),
.Y(n_9738)
);

INVx1_ASAP7_75t_L g9739 ( 
.A(n_9414),
.Y(n_9739)
);

AND2x2_ASAP7_75t_L g9740 ( 
.A(n_9373),
.B(n_9233),
.Y(n_9740)
);

BUFx8_ASAP7_75t_L g9741 ( 
.A(n_9676),
.Y(n_9741)
);

INVx3_ASAP7_75t_L g9742 ( 
.A(n_9540),
.Y(n_9742)
);

INVx6_ASAP7_75t_L g9743 ( 
.A(n_9325),
.Y(n_9743)
);

INVx1_ASAP7_75t_L g9744 ( 
.A(n_9415),
.Y(n_9744)
);

INVx2_ASAP7_75t_SL g9745 ( 
.A(n_9478),
.Y(n_9745)
);

INVx1_ASAP7_75t_L g9746 ( 
.A(n_9419),
.Y(n_9746)
);

INVx8_ASAP7_75t_L g9747 ( 
.A(n_9325),
.Y(n_9747)
);

INVx1_ASAP7_75t_L g9748 ( 
.A(n_9432),
.Y(n_9748)
);

INVx1_ASAP7_75t_L g9749 ( 
.A(n_9433),
.Y(n_9749)
);

INVx1_ASAP7_75t_L g9750 ( 
.A(n_9442),
.Y(n_9750)
);

CKINVDCx11_ASAP7_75t_R g9751 ( 
.A(n_9598),
.Y(n_9751)
);

AOI21xp5_ASAP7_75t_SL g9752 ( 
.A1(n_9327),
.A2(n_9206),
.B(n_9031),
.Y(n_9752)
);

INVxp67_ASAP7_75t_SL g9753 ( 
.A(n_9611),
.Y(n_9753)
);

NAND2xp5_ASAP7_75t_L g9754 ( 
.A(n_9561),
.B(n_9179),
.Y(n_9754)
);

BUFx6f_ASAP7_75t_L g9755 ( 
.A(n_9431),
.Y(n_9755)
);

OAI22xp5_ASAP7_75t_L g9756 ( 
.A1(n_9531),
.A2(n_9169),
.B1(n_9272),
.B2(n_9260),
.Y(n_9756)
);

INVx1_ASAP7_75t_SL g9757 ( 
.A(n_9627),
.Y(n_9757)
);

BUFx2_ASAP7_75t_L g9758 ( 
.A(n_9417),
.Y(n_9758)
);

INVx2_ASAP7_75t_L g9759 ( 
.A(n_9637),
.Y(n_9759)
);

HB1xp67_ASAP7_75t_L g9760 ( 
.A(n_9582),
.Y(n_9760)
);

CKINVDCx11_ASAP7_75t_R g9761 ( 
.A(n_9523),
.Y(n_9761)
);

INVx4_ASAP7_75t_L g9762 ( 
.A(n_9454),
.Y(n_9762)
);

AOI22xp33_ASAP7_75t_L g9763 ( 
.A1(n_9356),
.A2(n_8948),
.B1(n_9273),
.B2(n_9270),
.Y(n_9763)
);

OAI22xp5_ASAP7_75t_L g9764 ( 
.A1(n_9422),
.A2(n_9159),
.B1(n_9107),
.B2(n_9151),
.Y(n_9764)
);

AOI22xp33_ASAP7_75t_SL g9765 ( 
.A1(n_9343),
.A2(n_9673),
.B1(n_9595),
.B2(n_9498),
.Y(n_9765)
);

INVx1_ASAP7_75t_L g9766 ( 
.A(n_9446),
.Y(n_9766)
);

AOI22xp33_ASAP7_75t_L g9767 ( 
.A1(n_9378),
.A2(n_9304),
.B1(n_9263),
.B2(n_9280),
.Y(n_9767)
);

INVx1_ASAP7_75t_L g9768 ( 
.A(n_9453),
.Y(n_9768)
);

INVx2_ASAP7_75t_L g9769 ( 
.A(n_9643),
.Y(n_9769)
);

BUFx6f_ASAP7_75t_L g9770 ( 
.A(n_9431),
.Y(n_9770)
);

INVx2_ASAP7_75t_L g9771 ( 
.A(n_9645),
.Y(n_9771)
);

AOI22xp33_ASAP7_75t_L g9772 ( 
.A1(n_9342),
.A2(n_9139),
.B1(n_8957),
.B2(n_9104),
.Y(n_9772)
);

INVx1_ASAP7_75t_L g9773 ( 
.A(n_9464),
.Y(n_9773)
);

INVx3_ASAP7_75t_L g9774 ( 
.A(n_9568),
.Y(n_9774)
);

CKINVDCx14_ASAP7_75t_R g9775 ( 
.A(n_9605),
.Y(n_9775)
);

AOI22xp33_ASAP7_75t_L g9776 ( 
.A1(n_9348),
.A2(n_9038),
.B1(n_9056),
.B2(n_9027),
.Y(n_9776)
);

INVx2_ASAP7_75t_L g9777 ( 
.A(n_9471),
.Y(n_9777)
);

AOI22xp33_ASAP7_75t_L g9778 ( 
.A1(n_9334),
.A2(n_9156),
.B1(n_9170),
.B2(n_9166),
.Y(n_9778)
);

INVx6_ASAP7_75t_L g9779 ( 
.A(n_9609),
.Y(n_9779)
);

AOI22xp33_ASAP7_75t_SL g9780 ( 
.A1(n_9467),
.A2(n_9168),
.B1(n_9227),
.B2(n_9171),
.Y(n_9780)
);

INVx2_ASAP7_75t_SL g9781 ( 
.A(n_9456),
.Y(n_9781)
);

CKINVDCx5p33_ASAP7_75t_R g9782 ( 
.A(n_9322),
.Y(n_9782)
);

AOI22xp33_ASAP7_75t_L g9783 ( 
.A1(n_9334),
.A2(n_9339),
.B1(n_9416),
.B2(n_9352),
.Y(n_9783)
);

INVx1_ASAP7_75t_L g9784 ( 
.A(n_9485),
.Y(n_9784)
);

AOI22xp33_ASAP7_75t_L g9785 ( 
.A1(n_9465),
.A2(n_9476),
.B1(n_9492),
.B2(n_9468),
.Y(n_9785)
);

OAI22xp5_ASAP7_75t_L g9786 ( 
.A1(n_9422),
.A2(n_9128),
.B1(n_8996),
.B2(n_8998),
.Y(n_9786)
);

BUFx3_ASAP7_75t_L g9787 ( 
.A(n_9483),
.Y(n_9787)
);

AOI22xp33_ASAP7_75t_SL g9788 ( 
.A1(n_9560),
.A2(n_9000),
.B1(n_9004),
.B2(n_8999),
.Y(n_9788)
);

BUFx4_ASAP7_75t_SL g9789 ( 
.A(n_9496),
.Y(n_9789)
);

INVx3_ASAP7_75t_L g9790 ( 
.A(n_9571),
.Y(n_9790)
);

BUFx2_ASAP7_75t_L g9791 ( 
.A(n_9421),
.Y(n_9791)
);

OAI22xp5_ASAP7_75t_L g9792 ( 
.A1(n_9400),
.A2(n_9007),
.B1(n_9014),
.B2(n_8995),
.Y(n_9792)
);

INVx2_ASAP7_75t_L g9793 ( 
.A(n_9491),
.Y(n_9793)
);

CKINVDCx5p33_ASAP7_75t_R g9794 ( 
.A(n_9644),
.Y(n_9794)
);

BUFx8_ASAP7_75t_SL g9795 ( 
.A(n_9337),
.Y(n_9795)
);

OR2x2_ASAP7_75t_L g9796 ( 
.A(n_9338),
.B(n_9160),
.Y(n_9796)
);

CKINVDCx11_ASAP7_75t_R g9797 ( 
.A(n_9578),
.Y(n_9797)
);

AOI22xp33_ASAP7_75t_SL g9798 ( 
.A1(n_9539),
.A2(n_9059),
.B1(n_9046),
.B2(n_8980),
.Y(n_9798)
);

INVx1_ASAP7_75t_L g9799 ( 
.A(n_9340),
.Y(n_9799)
);

INVx1_ASAP7_75t_L g9800 ( 
.A(n_9534),
.Y(n_9800)
);

BUFx3_ASAP7_75t_L g9801 ( 
.A(n_9394),
.Y(n_9801)
);

INVx1_ASAP7_75t_L g9802 ( 
.A(n_9330),
.Y(n_9802)
);

NAND2xp5_ASAP7_75t_L g9803 ( 
.A(n_9333),
.B(n_8992),
.Y(n_9803)
);

BUFx12f_ASAP7_75t_L g9804 ( 
.A(n_9580),
.Y(n_9804)
);

AOI22xp5_ASAP7_75t_L g9805 ( 
.A1(n_9542),
.A2(n_9043),
.B1(n_8925),
.B2(n_9209),
.Y(n_9805)
);

INVx2_ASAP7_75t_L g9806 ( 
.A(n_9349),
.Y(n_9806)
);

BUFx12f_ASAP7_75t_L g9807 ( 
.A(n_9572),
.Y(n_9807)
);

BUFx3_ASAP7_75t_L g9808 ( 
.A(n_9396),
.Y(n_9808)
);

INVx1_ASAP7_75t_L g9809 ( 
.A(n_9369),
.Y(n_9809)
);

BUFx3_ASAP7_75t_L g9810 ( 
.A(n_9555),
.Y(n_9810)
);

INVx4_ASAP7_75t_L g9811 ( 
.A(n_9365),
.Y(n_9811)
);

INVx1_ASAP7_75t_L g9812 ( 
.A(n_9386),
.Y(n_9812)
);

OAI22xp33_ASAP7_75t_R g9813 ( 
.A1(n_9520),
.A2(n_489),
.B1(n_487),
.B2(n_488),
.Y(n_9813)
);

HB1xp67_ASAP7_75t_L g9814 ( 
.A(n_9336),
.Y(n_9814)
);

INVx2_ASAP7_75t_L g9815 ( 
.A(n_9389),
.Y(n_9815)
);

BUFx3_ASAP7_75t_L g9816 ( 
.A(n_9668),
.Y(n_9816)
);

INVx6_ASAP7_75t_L g9817 ( 
.A(n_9602),
.Y(n_9817)
);

INVx1_ASAP7_75t_L g9818 ( 
.A(n_9438),
.Y(n_9818)
);

OAI22xp5_ASAP7_75t_L g9819 ( 
.A1(n_9400),
.A2(n_9017),
.B1(n_8986),
.B2(n_8990),
.Y(n_9819)
);

INVx6_ASAP7_75t_L g9820 ( 
.A(n_9506),
.Y(n_9820)
);

INVx1_ASAP7_75t_L g9821 ( 
.A(n_9449),
.Y(n_9821)
);

AOI22xp33_ASAP7_75t_L g9822 ( 
.A1(n_9374),
.A2(n_9136),
.B1(n_9099),
.B2(n_9119),
.Y(n_9822)
);

INVx1_ASAP7_75t_L g9823 ( 
.A(n_9500),
.Y(n_9823)
);

BUFx6f_ASAP7_75t_L g9824 ( 
.A(n_9506),
.Y(n_9824)
);

OAI22xp5_ASAP7_75t_L g9825 ( 
.A1(n_9519),
.A2(n_8945),
.B1(n_9026),
.B2(n_9018),
.Y(n_9825)
);

AOI22xp33_ASAP7_75t_SL g9826 ( 
.A1(n_9461),
.A2(n_9105),
.B1(n_9040),
.B2(n_9047),
.Y(n_9826)
);

BUFx3_ASAP7_75t_L g9827 ( 
.A(n_9360),
.Y(n_9827)
);

INVx2_ASAP7_75t_L g9828 ( 
.A(n_9452),
.Y(n_9828)
);

INVx1_ASAP7_75t_L g9829 ( 
.A(n_9510),
.Y(n_9829)
);

INVx1_ASAP7_75t_SL g9830 ( 
.A(n_9341),
.Y(n_9830)
);

OAI22xp33_ASAP7_75t_L g9831 ( 
.A1(n_9625),
.A2(n_9040),
.B1(n_9047),
.B2(n_9033),
.Y(n_9831)
);

CKINVDCx11_ASAP7_75t_R g9832 ( 
.A(n_9518),
.Y(n_9832)
);

CKINVDCx11_ASAP7_75t_R g9833 ( 
.A(n_9551),
.Y(n_9833)
);

INVxp33_ASAP7_75t_SL g9834 ( 
.A(n_9430),
.Y(n_9834)
);

AND2x2_ASAP7_75t_L g9835 ( 
.A(n_9526),
.B(n_9033),
.Y(n_9835)
);

OAI22xp33_ASAP7_75t_L g9836 ( 
.A1(n_9625),
.A2(n_9061),
.B1(n_1087),
.B2(n_1088),
.Y(n_9836)
);

INVx6_ASAP7_75t_L g9837 ( 
.A(n_9586),
.Y(n_9837)
);

NAND2xp5_ASAP7_75t_L g9838 ( 
.A(n_9450),
.B(n_9061),
.Y(n_9838)
);

CKINVDCx11_ASAP7_75t_R g9839 ( 
.A(n_9513),
.Y(n_9839)
);

BUFx8_ASAP7_75t_SL g9840 ( 
.A(n_9439),
.Y(n_9840)
);

NAND2x1p5_ASAP7_75t_L g9841 ( 
.A(n_9562),
.B(n_1086),
.Y(n_9841)
);

CKINVDCx11_ASAP7_75t_R g9842 ( 
.A(n_9603),
.Y(n_9842)
);

AOI22xp33_ASAP7_75t_L g9843 ( 
.A1(n_9374),
.A2(n_1087),
.B1(n_1089),
.B2(n_1086),
.Y(n_9843)
);

INVx2_ASAP7_75t_SL g9844 ( 
.A(n_9382),
.Y(n_9844)
);

CKINVDCx14_ASAP7_75t_R g9845 ( 
.A(n_9570),
.Y(n_9845)
);

BUFx12f_ASAP7_75t_L g9846 ( 
.A(n_9622),
.Y(n_9846)
);

BUFx10_ASAP7_75t_L g9847 ( 
.A(n_9460),
.Y(n_9847)
);

INVx1_ASAP7_75t_L g9848 ( 
.A(n_9515),
.Y(n_9848)
);

INVx2_ASAP7_75t_SL g9849 ( 
.A(n_9420),
.Y(n_9849)
);

BUFx2_ASAP7_75t_SL g9850 ( 
.A(n_9429),
.Y(n_9850)
);

BUFx2_ASAP7_75t_L g9851 ( 
.A(n_9472),
.Y(n_9851)
);

OAI22xp5_ASAP7_75t_L g9852 ( 
.A1(n_9477),
.A2(n_489),
.B1(n_487),
.B2(n_488),
.Y(n_9852)
);

AOI22xp33_ASAP7_75t_SL g9853 ( 
.A1(n_9499),
.A2(n_1090),
.B1(n_1091),
.B2(n_1089),
.Y(n_9853)
);

OAI21xp5_ASAP7_75t_L g9854 ( 
.A1(n_9583),
.A2(n_1092),
.B(n_1091),
.Y(n_9854)
);

AOI22xp33_ASAP7_75t_L g9855 ( 
.A1(n_9374),
.A2(n_1093),
.B1(n_1094),
.B2(n_1092),
.Y(n_9855)
);

AOI22xp5_ASAP7_75t_L g9856 ( 
.A1(n_9499),
.A2(n_1094),
.B1(n_1095),
.B2(n_1093),
.Y(n_9856)
);

CKINVDCx20_ASAP7_75t_R g9857 ( 
.A(n_9358),
.Y(n_9857)
);

BUFx3_ASAP7_75t_L g9858 ( 
.A(n_9593),
.Y(n_9858)
);

BUFx12f_ASAP7_75t_L g9859 ( 
.A(n_9622),
.Y(n_9859)
);

AOI22xp33_ASAP7_75t_L g9860 ( 
.A1(n_9326),
.A2(n_1097),
.B1(n_1098),
.B2(n_1096),
.Y(n_9860)
);

AOI22xp33_ASAP7_75t_L g9861 ( 
.A1(n_9344),
.A2(n_1097),
.B1(n_1099),
.B2(n_1096),
.Y(n_9861)
);

INVx1_ASAP7_75t_L g9862 ( 
.A(n_9607),
.Y(n_9862)
);

BUFx2_ASAP7_75t_L g9863 ( 
.A(n_9669),
.Y(n_9863)
);

AOI22xp33_ASAP7_75t_L g9864 ( 
.A1(n_9677),
.A2(n_1100),
.B1(n_1101),
.B2(n_1099),
.Y(n_9864)
);

INVx1_ASAP7_75t_L g9865 ( 
.A(n_9553),
.Y(n_9865)
);

AOI22xp33_ASAP7_75t_L g9866 ( 
.A1(n_9527),
.A2(n_9428),
.B1(n_9444),
.B2(n_9447),
.Y(n_9866)
);

OAI22xp5_ASAP7_75t_L g9867 ( 
.A1(n_9666),
.A2(n_490),
.B1(n_488),
.B2(n_489),
.Y(n_9867)
);

BUFx3_ASAP7_75t_L g9868 ( 
.A(n_9596),
.Y(n_9868)
);

AND2x2_ASAP7_75t_L g9869 ( 
.A(n_9621),
.B(n_9332),
.Y(n_9869)
);

NAND2xp5_ASAP7_75t_L g9870 ( 
.A(n_9412),
.B(n_1100),
.Y(n_9870)
);

INVx1_ASAP7_75t_SL g9871 ( 
.A(n_9521),
.Y(n_9871)
);

INVx1_ASAP7_75t_L g9872 ( 
.A(n_9558),
.Y(n_9872)
);

INVx2_ASAP7_75t_L g9873 ( 
.A(n_9653),
.Y(n_9873)
);

OAI22xp5_ASAP7_75t_L g9874 ( 
.A1(n_9423),
.A2(n_9479),
.B1(n_9407),
.B2(n_9398),
.Y(n_9874)
);

BUFx4_ASAP7_75t_SL g9875 ( 
.A(n_9634),
.Y(n_9875)
);

INVx2_ASAP7_75t_L g9876 ( 
.A(n_9592),
.Y(n_9876)
);

INVx1_ASAP7_75t_L g9877 ( 
.A(n_9549),
.Y(n_9877)
);

INVx6_ASAP7_75t_L g9878 ( 
.A(n_9586),
.Y(n_9878)
);

INVx2_ASAP7_75t_SL g9879 ( 
.A(n_9481),
.Y(n_9879)
);

AOI22xp33_ASAP7_75t_L g9880 ( 
.A1(n_9441),
.A2(n_1102),
.B1(n_1103),
.B2(n_1101),
.Y(n_9880)
);

INVx1_ASAP7_75t_L g9881 ( 
.A(n_9455),
.Y(n_9881)
);

INVx1_ASAP7_75t_L g9882 ( 
.A(n_9646),
.Y(n_9882)
);

BUFx6f_ASAP7_75t_L g9883 ( 
.A(n_9599),
.Y(n_9883)
);

INVx4_ASAP7_75t_L g9884 ( 
.A(n_9599),
.Y(n_9884)
);

INVx6_ASAP7_75t_L g9885 ( 
.A(n_9614),
.Y(n_9885)
);

AOI21xp5_ASAP7_75t_L g9886 ( 
.A1(n_9563),
.A2(n_490),
.B(n_491),
.Y(n_9886)
);

BUFx12f_ASAP7_75t_L g9887 ( 
.A(n_9647),
.Y(n_9887)
);

HB1xp67_ASAP7_75t_L g9888 ( 
.A(n_9362),
.Y(n_9888)
);

AND2x2_ASAP7_75t_L g9889 ( 
.A(n_9359),
.B(n_490),
.Y(n_9889)
);

INVx1_ASAP7_75t_L g9890 ( 
.A(n_9626),
.Y(n_9890)
);

INVxp67_ASAP7_75t_SL g9891 ( 
.A(n_9395),
.Y(n_9891)
);

CKINVDCx11_ASAP7_75t_R g9892 ( 
.A(n_9603),
.Y(n_9892)
);

INVx1_ASAP7_75t_L g9893 ( 
.A(n_9662),
.Y(n_9893)
);

BUFx10_ASAP7_75t_L g9894 ( 
.A(n_9606),
.Y(n_9894)
);

AOI22xp5_ASAP7_75t_L g9895 ( 
.A1(n_9499),
.A2(n_1104),
.B1(n_1105),
.B2(n_1102),
.Y(n_9895)
);

BUFx5_ASAP7_75t_L g9896 ( 
.A(n_9632),
.Y(n_9896)
);

AOI22xp5_ASAP7_75t_L g9897 ( 
.A1(n_9507),
.A2(n_1106),
.B1(n_1107),
.B2(n_1104),
.Y(n_9897)
);

INVx1_ASAP7_75t_L g9898 ( 
.A(n_9364),
.Y(n_9898)
);

INVx1_ASAP7_75t_SL g9899 ( 
.A(n_9409),
.Y(n_9899)
);

CKINVDCx6p67_ASAP7_75t_R g9900 ( 
.A(n_9401),
.Y(n_9900)
);

INVx1_ASAP7_75t_L g9901 ( 
.A(n_9685),
.Y(n_9901)
);

CKINVDCx20_ASAP7_75t_R g9902 ( 
.A(n_9486),
.Y(n_9902)
);

OAI22xp33_ASAP7_75t_L g9903 ( 
.A1(n_9514),
.A2(n_1108),
.B1(n_1110),
.B2(n_1106),
.Y(n_9903)
);

INVx2_ASAP7_75t_SL g9904 ( 
.A(n_9451),
.Y(n_9904)
);

CKINVDCx11_ASAP7_75t_R g9905 ( 
.A(n_9614),
.Y(n_9905)
);

INVx2_ASAP7_75t_L g9906 ( 
.A(n_9687),
.Y(n_9906)
);

CKINVDCx20_ASAP7_75t_R g9907 ( 
.A(n_9487),
.Y(n_9907)
);

INVx1_ASAP7_75t_L g9908 ( 
.A(n_9636),
.Y(n_9908)
);

OAI21xp5_ASAP7_75t_L g9909 ( 
.A1(n_9537),
.A2(n_1110),
.B(n_1108),
.Y(n_9909)
);

INVxp67_ASAP7_75t_SL g9910 ( 
.A(n_9367),
.Y(n_9910)
);

INVx1_ASAP7_75t_L g9911 ( 
.A(n_9410),
.Y(n_9911)
);

INVx1_ASAP7_75t_SL g9912 ( 
.A(n_9351),
.Y(n_9912)
);

CKINVDCx5p33_ASAP7_75t_R g9913 ( 
.A(n_9649),
.Y(n_9913)
);

CKINVDCx6p67_ASAP7_75t_R g9914 ( 
.A(n_9402),
.Y(n_9914)
);

AOI22xp33_ASAP7_75t_SL g9915 ( 
.A1(n_9559),
.A2(n_1112),
.B1(n_1114),
.B2(n_1111),
.Y(n_9915)
);

AOI22xp33_ASAP7_75t_L g9916 ( 
.A1(n_9616),
.A2(n_1112),
.B1(n_1115),
.B2(n_1111),
.Y(n_9916)
);

INVx6_ASAP7_75t_L g9917 ( 
.A(n_9649),
.Y(n_9917)
);

AOI22xp33_ASAP7_75t_SL g9918 ( 
.A1(n_9379),
.A2(n_1117),
.B1(n_1118),
.B2(n_1116),
.Y(n_9918)
);

INVx2_ASAP7_75t_L g9919 ( 
.A(n_9656),
.Y(n_9919)
);

INVx6_ASAP7_75t_L g9920 ( 
.A(n_9683),
.Y(n_9920)
);

CKINVDCx6p67_ASAP7_75t_R g9921 ( 
.A(n_9397),
.Y(n_9921)
);

AOI22x1_ASAP7_75t_SL g9922 ( 
.A1(n_9567),
.A2(n_493),
.B1(n_491),
.B2(n_492),
.Y(n_9922)
);

BUFx3_ASAP7_75t_L g9923 ( 
.A(n_9629),
.Y(n_9923)
);

INVx4_ASAP7_75t_L g9924 ( 
.A(n_9404),
.Y(n_9924)
);

INVx2_ASAP7_75t_L g9925 ( 
.A(n_9667),
.Y(n_9925)
);

AOI22xp33_ASAP7_75t_L g9926 ( 
.A1(n_9618),
.A2(n_1117),
.B1(n_1118),
.B2(n_1116),
.Y(n_9926)
);

AOI22xp33_ASAP7_75t_L g9927 ( 
.A1(n_9566),
.A2(n_9524),
.B1(n_9463),
.B2(n_9671),
.Y(n_9927)
);

INVx2_ASAP7_75t_L g9928 ( 
.A(n_9591),
.Y(n_9928)
);

OAI21xp5_ASAP7_75t_SL g9929 ( 
.A1(n_9575),
.A2(n_491),
.B(n_492),
.Y(n_9929)
);

OAI22xp33_ASAP7_75t_L g9930 ( 
.A1(n_9355),
.A2(n_1120),
.B1(n_1121),
.B2(n_1119),
.Y(n_9930)
);

AOI22xp33_ASAP7_75t_L g9931 ( 
.A1(n_9480),
.A2(n_1121),
.B1(n_1122),
.B2(n_1120),
.Y(n_9931)
);

BUFx3_ASAP7_75t_L g9932 ( 
.A(n_9652),
.Y(n_9932)
);

AOI22xp33_ASAP7_75t_L g9933 ( 
.A1(n_9475),
.A2(n_1124),
.B1(n_1125),
.B2(n_1123),
.Y(n_9933)
);

AOI22xp33_ASAP7_75t_L g9934 ( 
.A1(n_9641),
.A2(n_1126),
.B1(n_1127),
.B2(n_1125),
.Y(n_9934)
);

INVx2_ASAP7_75t_SL g9935 ( 
.A(n_9545),
.Y(n_9935)
);

INVx6_ASAP7_75t_L g9936 ( 
.A(n_9484),
.Y(n_9936)
);

AOI22xp33_ASAP7_75t_L g9937 ( 
.A1(n_9556),
.A2(n_1127),
.B1(n_1128),
.B2(n_1126),
.Y(n_9937)
);

BUFx3_ASAP7_75t_L g9938 ( 
.A(n_9682),
.Y(n_9938)
);

OAI22xp5_ASAP7_75t_L g9939 ( 
.A1(n_9574),
.A2(n_494),
.B1(n_492),
.B2(n_493),
.Y(n_9939)
);

AOI22xp33_ASAP7_75t_SL g9940 ( 
.A1(n_9408),
.A2(n_1131),
.B1(n_1132),
.B2(n_1130),
.Y(n_9940)
);

AOI22xp33_ASAP7_75t_L g9941 ( 
.A1(n_9511),
.A2(n_1131),
.B1(n_1132),
.B2(n_1130),
.Y(n_9941)
);

AOI22xp33_ASAP7_75t_SL g9942 ( 
.A1(n_9680),
.A2(n_1134),
.B1(n_1135),
.B2(n_1133),
.Y(n_9942)
);

INVx2_ASAP7_75t_L g9943 ( 
.A(n_9597),
.Y(n_9943)
);

INVx1_ASAP7_75t_L g9944 ( 
.A(n_9664),
.Y(n_9944)
);

INVx2_ASAP7_75t_R g9945 ( 
.A(n_9675),
.Y(n_9945)
);

NAND2x1p5_ASAP7_75t_L g9946 ( 
.A(n_9489),
.B(n_1133),
.Y(n_9946)
);

AOI22xp33_ASAP7_75t_L g9947 ( 
.A1(n_9516),
.A2(n_1136),
.B1(n_1137),
.B2(n_1135),
.Y(n_9947)
);

BUFx12f_ASAP7_75t_L g9948 ( 
.A(n_9458),
.Y(n_9948)
);

AOI22xp33_ASAP7_75t_SL g9949 ( 
.A1(n_9363),
.A2(n_1137),
.B1(n_1138),
.B2(n_1136),
.Y(n_9949)
);

CKINVDCx6p67_ASAP7_75t_R g9950 ( 
.A(n_9681),
.Y(n_9950)
);

AOI22xp33_ASAP7_75t_L g9951 ( 
.A1(n_9635),
.A2(n_1140),
.B1(n_1141),
.B2(n_1139),
.Y(n_9951)
);

INVx1_ASAP7_75t_L g9952 ( 
.A(n_9679),
.Y(n_9952)
);

BUFx6f_ASAP7_75t_L g9953 ( 
.A(n_9631),
.Y(n_9953)
);

CKINVDCx11_ASAP7_75t_R g9954 ( 
.A(n_9576),
.Y(n_9954)
);

OAI22xp5_ASAP7_75t_L g9955 ( 
.A1(n_9612),
.A2(n_495),
.B1(n_493),
.B2(n_494),
.Y(n_9955)
);

BUFx2_ASAP7_75t_L g9956 ( 
.A(n_9573),
.Y(n_9956)
);

AOI21xp33_ASAP7_75t_L g9957 ( 
.A1(n_9380),
.A2(n_1141),
.B(n_1139),
.Y(n_9957)
);

BUFx2_ASAP7_75t_SL g9958 ( 
.A(n_9436),
.Y(n_9958)
);

INVx6_ASAP7_75t_L g9959 ( 
.A(n_9584),
.Y(n_9959)
);

OAI22xp5_ASAP7_75t_L g9960 ( 
.A1(n_9557),
.A2(n_496),
.B1(n_494),
.B2(n_495),
.Y(n_9960)
);

INVx1_ASAP7_75t_L g9961 ( 
.A(n_9424),
.Y(n_9961)
);

OAI21xp33_ASAP7_75t_L g9962 ( 
.A1(n_9601),
.A2(n_495),
.B(n_497),
.Y(n_9962)
);

BUFx2_ASAP7_75t_L g9963 ( 
.A(n_9323),
.Y(n_9963)
);

INVx6_ASAP7_75t_L g9964 ( 
.A(n_9589),
.Y(n_9964)
);

INVx2_ASAP7_75t_L g9965 ( 
.A(n_9482),
.Y(n_9965)
);

CKINVDCx20_ASAP7_75t_R g9966 ( 
.A(n_9554),
.Y(n_9966)
);

NAND2x1p5_ASAP7_75t_L g9967 ( 
.A(n_9546),
.B(n_1142),
.Y(n_9967)
);

AOI22xp33_ASAP7_75t_L g9968 ( 
.A1(n_9638),
.A2(n_1143),
.B1(n_1144),
.B2(n_1142),
.Y(n_9968)
);

AOI22xp33_ASAP7_75t_L g9969 ( 
.A1(n_9569),
.A2(n_1144),
.B1(n_1145),
.B2(n_1143),
.Y(n_9969)
);

INVx6_ASAP7_75t_L g9970 ( 
.A(n_9532),
.Y(n_9970)
);

OAI22xp5_ASAP7_75t_L g9971 ( 
.A1(n_9633),
.A2(n_499),
.B1(n_497),
.B2(n_498),
.Y(n_9971)
);

AOI22xp33_ASAP7_75t_SL g9972 ( 
.A1(n_9376),
.A2(n_1146),
.B1(n_1147),
.B2(n_1145),
.Y(n_9972)
);

INVx2_ASAP7_75t_L g9973 ( 
.A(n_9392),
.Y(n_9973)
);

BUFx10_ASAP7_75t_L g9974 ( 
.A(n_9670),
.Y(n_9974)
);

INVx1_ASAP7_75t_L g9975 ( 
.A(n_9462),
.Y(n_9975)
);

OAI22xp5_ASAP7_75t_L g9976 ( 
.A1(n_9660),
.A2(n_499),
.B1(n_497),
.B2(n_498),
.Y(n_9976)
);

INVx1_ASAP7_75t_L g9977 ( 
.A(n_9474),
.Y(n_9977)
);

AOI22xp33_ASAP7_75t_L g9978 ( 
.A1(n_9375),
.A2(n_1149),
.B1(n_1150),
.B2(n_1148),
.Y(n_9978)
);

OAI22xp33_ASAP7_75t_L g9979 ( 
.A1(n_9388),
.A2(n_1151),
.B1(n_1152),
.B2(n_1149),
.Y(n_9979)
);

AOI22xp33_ASAP7_75t_L g9980 ( 
.A1(n_9661),
.A2(n_1152),
.B1(n_1153),
.B2(n_1151),
.Y(n_9980)
);

BUFx2_ASAP7_75t_SL g9981 ( 
.A(n_9565),
.Y(n_9981)
);

INVx1_ASAP7_75t_L g9982 ( 
.A(n_9624),
.Y(n_9982)
);

INVx1_ASAP7_75t_SL g9983 ( 
.A(n_9665),
.Y(n_9983)
);

INVx1_ASAP7_75t_SL g9984 ( 
.A(n_9588),
.Y(n_9984)
);

BUFx3_ASAP7_75t_L g9985 ( 
.A(n_9658),
.Y(n_9985)
);

BUFx12f_ASAP7_75t_L g9986 ( 
.A(n_9674),
.Y(n_9986)
);

INVx2_ASAP7_75t_L g9987 ( 
.A(n_9896),
.Y(n_9987)
);

AO21x1_ASAP7_75t_L g9988 ( 
.A1(n_9911),
.A2(n_9663),
.B(n_9347),
.Y(n_9988)
);

INVx1_ASAP7_75t_L g9989 ( 
.A(n_9760),
.Y(n_9989)
);

INVx1_ASAP7_75t_L g9990 ( 
.A(n_9800),
.Y(n_9990)
);

AOI222xp33_ASAP7_75t_L g9991 ( 
.A1(n_9852),
.A2(n_9642),
.B1(n_9437),
.B2(n_9443),
.C1(n_9448),
.C2(n_9505),
.Y(n_9991)
);

HB1xp67_ASAP7_75t_L g9992 ( 
.A(n_9888),
.Y(n_9992)
);

INVx1_ASAP7_75t_L g9993 ( 
.A(n_9753),
.Y(n_9993)
);

INVx2_ASAP7_75t_L g9994 ( 
.A(n_9896),
.Y(n_9994)
);

INVx2_ASAP7_75t_L g9995 ( 
.A(n_9896),
.Y(n_9995)
);

INVx3_ASAP7_75t_L g9996 ( 
.A(n_9816),
.Y(n_9996)
);

INVx1_ASAP7_75t_L g9997 ( 
.A(n_9690),
.Y(n_9997)
);

BUFx3_ASAP7_75t_L g9998 ( 
.A(n_9857),
.Y(n_9998)
);

INVx1_ASAP7_75t_L g9999 ( 
.A(n_9712),
.Y(n_9999)
);

BUFx3_ASAP7_75t_L g10000 ( 
.A(n_9795),
.Y(n_10000)
);

BUFx2_ASAP7_75t_L g10001 ( 
.A(n_9734),
.Y(n_10001)
);

NAND2xp5_ASAP7_75t_L g10002 ( 
.A(n_9891),
.B(n_9370),
.Y(n_10002)
);

INVx1_ASAP7_75t_L g10003 ( 
.A(n_9719),
.Y(n_10003)
);

AOI22xp33_ASAP7_75t_L g10004 ( 
.A1(n_9701),
.A2(n_9530),
.B1(n_9623),
.B2(n_9381),
.Y(n_10004)
);

INVx1_ASAP7_75t_L g10005 ( 
.A(n_9731),
.Y(n_10005)
);

INVx2_ASAP7_75t_L g10006 ( 
.A(n_9896),
.Y(n_10006)
);

INVx2_ASAP7_75t_SL g10007 ( 
.A(n_9875),
.Y(n_10007)
);

AND2x2_ASAP7_75t_L g10008 ( 
.A(n_9713),
.B(n_9684),
.Y(n_10008)
);

CKINVDCx8_ASAP7_75t_R g10009 ( 
.A(n_9794),
.Y(n_10009)
);

INVx1_ASAP7_75t_L g10010 ( 
.A(n_9739),
.Y(n_10010)
);

INVx1_ASAP7_75t_L g10011 ( 
.A(n_9744),
.Y(n_10011)
);

INVx1_ASAP7_75t_L g10012 ( 
.A(n_9746),
.Y(n_10012)
);

INVx1_ASAP7_75t_L g10013 ( 
.A(n_9748),
.Y(n_10013)
);

OR2x6_ASAP7_75t_L g10014 ( 
.A(n_9958),
.B(n_9538),
.Y(n_10014)
);

AO21x1_ASAP7_75t_L g10015 ( 
.A1(n_9874),
.A2(n_9726),
.B(n_9697),
.Y(n_10015)
);

INVx3_ASAP7_75t_L g10016 ( 
.A(n_9950),
.Y(n_10016)
);

OAI21xp5_ASAP7_75t_L g10017 ( 
.A1(n_9732),
.A2(n_9610),
.B(n_9613),
.Y(n_10017)
);

INVx1_ASAP7_75t_L g10018 ( 
.A(n_9749),
.Y(n_10018)
);

INVx1_ASAP7_75t_SL g10019 ( 
.A(n_9839),
.Y(n_10019)
);

INVx1_ASAP7_75t_L g10020 ( 
.A(n_9750),
.Y(n_10020)
);

INVx1_ASAP7_75t_L g10021 ( 
.A(n_9766),
.Y(n_10021)
);

HB1xp67_ASAP7_75t_L g10022 ( 
.A(n_9814),
.Y(n_10022)
);

INVx2_ASAP7_75t_L g10023 ( 
.A(n_9711),
.Y(n_10023)
);

INVx1_ASAP7_75t_L g10024 ( 
.A(n_9768),
.Y(n_10024)
);

AOI22xp33_ASAP7_75t_SL g10025 ( 
.A1(n_9721),
.A2(n_9427),
.B1(n_9529),
.B2(n_9434),
.Y(n_10025)
);

BUFx2_ASAP7_75t_L g10026 ( 
.A(n_9758),
.Y(n_10026)
);

INVx1_ASAP7_75t_L g10027 ( 
.A(n_9773),
.Y(n_10027)
);

OAI21xp5_ASAP7_75t_L g10028 ( 
.A1(n_9752),
.A2(n_9639),
.B(n_9608),
.Y(n_10028)
);

INVx2_ASAP7_75t_L g10029 ( 
.A(n_9700),
.Y(n_10029)
);

INVx3_ASAP7_75t_L g10030 ( 
.A(n_9924),
.Y(n_10030)
);

HB1xp67_ASAP7_75t_L g10031 ( 
.A(n_9703),
.Y(n_10031)
);

INVx1_ASAP7_75t_L g10032 ( 
.A(n_9777),
.Y(n_10032)
);

INVxp33_ASAP7_75t_L g10033 ( 
.A(n_9723),
.Y(n_10033)
);

INVx2_ASAP7_75t_L g10034 ( 
.A(n_9702),
.Y(n_10034)
);

INVx2_ASAP7_75t_L g10035 ( 
.A(n_9759),
.Y(n_10035)
);

NAND2xp5_ASAP7_75t_L g10036 ( 
.A(n_9910),
.B(n_9488),
.Y(n_10036)
);

OR2x2_ASAP7_75t_L g10037 ( 
.A(n_9898),
.B(n_9672),
.Y(n_10037)
);

HB1xp67_ASAP7_75t_L g10038 ( 
.A(n_9877),
.Y(n_10038)
);

INVx2_ASAP7_75t_L g10039 ( 
.A(n_9769),
.Y(n_10039)
);

AO21x1_ASAP7_75t_L g10040 ( 
.A1(n_9764),
.A2(n_9657),
.B(n_9655),
.Y(n_10040)
);

INVx1_ASAP7_75t_L g10041 ( 
.A(n_9823),
.Y(n_10041)
);

AOI22xp33_ASAP7_75t_SL g10042 ( 
.A1(n_9922),
.A2(n_9590),
.B1(n_9535),
.B2(n_9548),
.Y(n_10042)
);

INVx1_ASAP7_75t_L g10043 ( 
.A(n_9829),
.Y(n_10043)
);

HB1xp67_ASAP7_75t_L g10044 ( 
.A(n_9851),
.Y(n_10044)
);

INVx1_ASAP7_75t_L g10045 ( 
.A(n_9848),
.Y(n_10045)
);

INVx1_ASAP7_75t_L g10046 ( 
.A(n_9784),
.Y(n_10046)
);

INVx1_ASAP7_75t_L g10047 ( 
.A(n_9908),
.Y(n_10047)
);

INVx2_ASAP7_75t_L g10048 ( 
.A(n_9771),
.Y(n_10048)
);

BUFx2_ASAP7_75t_SL g10049 ( 
.A(n_9902),
.Y(n_10049)
);

AOI21x1_ASAP7_75t_L g10050 ( 
.A1(n_9786),
.A2(n_9435),
.B(n_9654),
.Y(n_10050)
);

INVx2_ASAP7_75t_L g10051 ( 
.A(n_9973),
.Y(n_10051)
);

INVx2_ASAP7_75t_L g10052 ( 
.A(n_9863),
.Y(n_10052)
);

INVx1_ASAP7_75t_L g10053 ( 
.A(n_9952),
.Y(n_10053)
);

HB1xp67_ASAP7_75t_L g10054 ( 
.A(n_9791),
.Y(n_10054)
);

INVx3_ASAP7_75t_L g10055 ( 
.A(n_9810),
.Y(n_10055)
);

INVx1_ASAP7_75t_SL g10056 ( 
.A(n_9761),
.Y(n_10056)
);

BUFx6f_ASAP7_75t_L g10057 ( 
.A(n_9797),
.Y(n_10057)
);

INVx3_ASAP7_75t_L g10058 ( 
.A(n_9694),
.Y(n_10058)
);

AO21x2_ASAP7_75t_L g10059 ( 
.A1(n_9870),
.A2(n_9630),
.B(n_9457),
.Y(n_10059)
);

INVx1_ASAP7_75t_L g10060 ( 
.A(n_9944),
.Y(n_10060)
);

OAI21x1_ASAP7_75t_L g10061 ( 
.A1(n_9715),
.A2(n_9730),
.B(n_9928),
.Y(n_10061)
);

INVx2_ASAP7_75t_SL g10062 ( 
.A(n_9708),
.Y(n_10062)
);

BUFx4f_ASAP7_75t_SL g10063 ( 
.A(n_9705),
.Y(n_10063)
);

INVx1_ASAP7_75t_L g10064 ( 
.A(n_9799),
.Y(n_10064)
);

INVx2_ASAP7_75t_L g10065 ( 
.A(n_9963),
.Y(n_10065)
);

INVx1_ASAP7_75t_L g10066 ( 
.A(n_9943),
.Y(n_10066)
);

BUFx6f_ASAP7_75t_L g10067 ( 
.A(n_9905),
.Y(n_10067)
);

INVx1_ASAP7_75t_L g10068 ( 
.A(n_9890),
.Y(n_10068)
);

INVx1_ASAP7_75t_L g10069 ( 
.A(n_9881),
.Y(n_10069)
);

INVx1_ASAP7_75t_L g10070 ( 
.A(n_9802),
.Y(n_10070)
);

INVx1_ASAP7_75t_L g10071 ( 
.A(n_9809),
.Y(n_10071)
);

INVx1_ASAP7_75t_L g10072 ( 
.A(n_9812),
.Y(n_10072)
);

INVx1_ASAP7_75t_L g10073 ( 
.A(n_9818),
.Y(n_10073)
);

OAI222xp33_ASAP7_75t_L g10074 ( 
.A1(n_9689),
.A2(n_9659),
.B1(n_9345),
.B2(n_9579),
.C1(n_9585),
.C2(n_9577),
.Y(n_10074)
);

INVx2_ASAP7_75t_L g10075 ( 
.A(n_9793),
.Y(n_10075)
);

HB1xp67_ASAP7_75t_L g10076 ( 
.A(n_9688),
.Y(n_10076)
);

INVx2_ASAP7_75t_L g10077 ( 
.A(n_9806),
.Y(n_10077)
);

INVx1_ASAP7_75t_L g10078 ( 
.A(n_9821),
.Y(n_10078)
);

INVx1_ASAP7_75t_L g10079 ( 
.A(n_9893),
.Y(n_10079)
);

CKINVDCx5p33_ASAP7_75t_R g10080 ( 
.A(n_9789),
.Y(n_10080)
);

INVx2_ASAP7_75t_L g10081 ( 
.A(n_9815),
.Y(n_10081)
);

BUFx2_ASAP7_75t_SL g10082 ( 
.A(n_9907),
.Y(n_10082)
);

INVx3_ASAP7_75t_L g10083 ( 
.A(n_9694),
.Y(n_10083)
);

NAND2x1p5_ASAP7_75t_L g10084 ( 
.A(n_9709),
.B(n_9413),
.Y(n_10084)
);

AO31x2_ASAP7_75t_L g10085 ( 
.A1(n_9729),
.A2(n_9544),
.A3(n_9550),
.B(n_9543),
.Y(n_10085)
);

HB1xp67_ASAP7_75t_L g10086 ( 
.A(n_9718),
.Y(n_10086)
);

INVx2_ASAP7_75t_L g10087 ( 
.A(n_9873),
.Y(n_10087)
);

INVx2_ASAP7_75t_L g10088 ( 
.A(n_9876),
.Y(n_10088)
);

HB1xp67_ASAP7_75t_L g10089 ( 
.A(n_9862),
.Y(n_10089)
);

AO21x2_ASAP7_75t_L g10090 ( 
.A1(n_9975),
.A2(n_9604),
.B(n_9564),
.Y(n_10090)
);

NAND2x1p5_ASAP7_75t_L g10091 ( 
.A(n_9899),
.B(n_9490),
.Y(n_10091)
);

INVx2_ASAP7_75t_L g10092 ( 
.A(n_9906),
.Y(n_10092)
);

OAI221xp5_ASAP7_75t_SL g10093 ( 
.A1(n_9785),
.A2(n_9493),
.B1(n_9525),
.B2(n_9504),
.C(n_9501),
.Y(n_10093)
);

INVx2_ASAP7_75t_L g10094 ( 
.A(n_9865),
.Y(n_10094)
);

AND2x4_ASAP7_75t_L g10095 ( 
.A(n_9745),
.B(n_9497),
.Y(n_10095)
);

OR2x6_ASAP7_75t_L g10096 ( 
.A(n_9981),
.B(n_9547),
.Y(n_10096)
);

OA21x2_ASAP7_75t_L g10097 ( 
.A1(n_9754),
.A2(n_9522),
.B(n_9536),
.Y(n_10097)
);

AOI22xp33_ASAP7_75t_SL g10098 ( 
.A1(n_9966),
.A2(n_9508),
.B1(n_9587),
.B2(n_9517),
.Y(n_10098)
);

CKINVDCx5p33_ASAP7_75t_R g10099 ( 
.A(n_9716),
.Y(n_10099)
);

INVx2_ASAP7_75t_L g10100 ( 
.A(n_9872),
.Y(n_10100)
);

AOI22xp33_ASAP7_75t_L g10101 ( 
.A1(n_9765),
.A2(n_9813),
.B1(n_9696),
.B2(n_9854),
.Y(n_10101)
);

HB1xp67_ASAP7_75t_L g10102 ( 
.A(n_9912),
.Y(n_10102)
);

INVx2_ASAP7_75t_L g10103 ( 
.A(n_9828),
.Y(n_10103)
);

INVx2_ASAP7_75t_L g10104 ( 
.A(n_9901),
.Y(n_10104)
);

AND2x2_ASAP7_75t_L g10105 ( 
.A(n_9710),
.B(n_9445),
.Y(n_10105)
);

INVx2_ASAP7_75t_L g10106 ( 
.A(n_9882),
.Y(n_10106)
);

AND2x4_ASAP7_75t_L g10107 ( 
.A(n_9728),
.B(n_9503),
.Y(n_10107)
);

OAI21xp5_ASAP7_75t_L g10108 ( 
.A1(n_9886),
.A2(n_9502),
.B(n_9385),
.Y(n_10108)
);

INVx1_ASAP7_75t_L g10109 ( 
.A(n_9982),
.Y(n_10109)
);

INVx2_ASAP7_75t_SL g10110 ( 
.A(n_9708),
.Y(n_10110)
);

HB1xp67_ASAP7_75t_L g10111 ( 
.A(n_9965),
.Y(n_10111)
);

INVx1_ASAP7_75t_L g10112 ( 
.A(n_9961),
.Y(n_10112)
);

INVx2_ASAP7_75t_SL g10113 ( 
.A(n_9747),
.Y(n_10113)
);

OAI22xp5_ASAP7_75t_L g10114 ( 
.A1(n_9783),
.A2(n_9686),
.B1(n_9678),
.B2(n_500),
.Y(n_10114)
);

OAI21x1_ASAP7_75t_L g10115 ( 
.A1(n_9977),
.A2(n_498),
.B(n_499),
.Y(n_10115)
);

INVxp67_ASAP7_75t_L g10116 ( 
.A(n_9850),
.Y(n_10116)
);

NAND2xp5_ASAP7_75t_L g10117 ( 
.A(n_9803),
.B(n_9869),
.Y(n_10117)
);

INVx1_ASAP7_75t_L g10118 ( 
.A(n_9796),
.Y(n_10118)
);

HB1xp67_ASAP7_75t_L g10119 ( 
.A(n_9740),
.Y(n_10119)
);

NAND2xp5_ASAP7_75t_L g10120 ( 
.A(n_9919),
.B(n_1154),
.Y(n_10120)
);

CKINVDCx6p67_ASAP7_75t_R g10121 ( 
.A(n_9832),
.Y(n_10121)
);

INVx2_ASAP7_75t_L g10122 ( 
.A(n_9956),
.Y(n_10122)
);

INVx1_ASAP7_75t_L g10123 ( 
.A(n_9925),
.Y(n_10123)
);

AOI22xp33_ASAP7_75t_L g10124 ( 
.A1(n_9866),
.A2(n_1155),
.B1(n_1156),
.B2(n_1154),
.Y(n_10124)
);

INVx1_ASAP7_75t_L g10125 ( 
.A(n_9838),
.Y(n_10125)
);

INVx2_ASAP7_75t_L g10126 ( 
.A(n_9849),
.Y(n_10126)
);

OR2x2_ASAP7_75t_L g10127 ( 
.A(n_9945),
.B(n_500),
.Y(n_10127)
);

INVx1_ASAP7_75t_SL g10128 ( 
.A(n_9833),
.Y(n_10128)
);

INVx2_ASAP7_75t_SL g10129 ( 
.A(n_9747),
.Y(n_10129)
);

INVx5_ASAP7_75t_L g10130 ( 
.A(n_9722),
.Y(n_10130)
);

BUFx2_ASAP7_75t_L g10131 ( 
.A(n_9845),
.Y(n_10131)
);

INVx1_ASAP7_75t_L g10132 ( 
.A(n_9835),
.Y(n_10132)
);

HB1xp67_ASAP7_75t_L g10133 ( 
.A(n_9830),
.Y(n_10133)
);

AND2x2_ASAP7_75t_L g10134 ( 
.A(n_9844),
.B(n_501),
.Y(n_10134)
);

INVx2_ASAP7_75t_L g10135 ( 
.A(n_9879),
.Y(n_10135)
);

INVx2_ASAP7_75t_L g10136 ( 
.A(n_9904),
.Y(n_10136)
);

INVx1_ASAP7_75t_L g10137 ( 
.A(n_9757),
.Y(n_10137)
);

BUFx3_ASAP7_75t_L g10138 ( 
.A(n_9840),
.Y(n_10138)
);

HB1xp67_ASAP7_75t_L g10139 ( 
.A(n_9871),
.Y(n_10139)
);

INVx1_ASAP7_75t_L g10140 ( 
.A(n_9935),
.Y(n_10140)
);

AOI22xp33_ASAP7_75t_L g10141 ( 
.A1(n_9927),
.A2(n_1156),
.B1(n_1157),
.B2(n_1155),
.Y(n_10141)
);

INVx3_ASAP7_75t_L g10142 ( 
.A(n_9743),
.Y(n_10142)
);

INVx2_ASAP7_75t_L g10143 ( 
.A(n_9985),
.Y(n_10143)
);

INVx1_ASAP7_75t_L g10144 ( 
.A(n_9827),
.Y(n_10144)
);

OA21x2_ASAP7_75t_L g10145 ( 
.A1(n_9778),
.A2(n_501),
.B(n_502),
.Y(n_10145)
);

INVx1_ASAP7_75t_L g10146 ( 
.A(n_9738),
.Y(n_10146)
);

AND2x2_ASAP7_75t_L g10147 ( 
.A(n_9742),
.B(n_502),
.Y(n_10147)
);

INVx1_ASAP7_75t_L g10148 ( 
.A(n_9774),
.Y(n_10148)
);

INVx2_ASAP7_75t_L g10149 ( 
.A(n_9790),
.Y(n_10149)
);

INVx1_ASAP7_75t_L g10150 ( 
.A(n_9983),
.Y(n_10150)
);

BUFx3_ASAP7_75t_L g10151 ( 
.A(n_9842),
.Y(n_10151)
);

INVx1_ASAP7_75t_L g10152 ( 
.A(n_9819),
.Y(n_10152)
);

OAI22xp5_ASAP7_75t_L g10153 ( 
.A1(n_9826),
.A2(n_504),
.B1(n_502),
.B2(n_503),
.Y(n_10153)
);

INVx2_ASAP7_75t_L g10154 ( 
.A(n_9953),
.Y(n_10154)
);

INVx1_ASAP7_75t_L g10155 ( 
.A(n_9923),
.Y(n_10155)
);

OA21x2_ASAP7_75t_L g10156 ( 
.A1(n_9772),
.A2(n_503),
.B(n_504),
.Y(n_10156)
);

AOI22xp33_ASAP7_75t_L g10157 ( 
.A1(n_9867),
.A2(n_1158),
.B1(n_1159),
.B2(n_1157),
.Y(n_10157)
);

INVx1_ASAP7_75t_L g10158 ( 
.A(n_9932),
.Y(n_10158)
);

INVx1_ASAP7_75t_L g10159 ( 
.A(n_9938),
.Y(n_10159)
);

BUFx2_ASAP7_75t_L g10160 ( 
.A(n_9737),
.Y(n_10160)
);

AOI22xp33_ASAP7_75t_SL g10161 ( 
.A1(n_9733),
.A2(n_1161),
.B1(n_1162),
.B2(n_1160),
.Y(n_10161)
);

INVxp67_ASAP7_75t_L g10162 ( 
.A(n_9792),
.Y(n_10162)
);

INVx1_ASAP7_75t_L g10163 ( 
.A(n_9781),
.Y(n_10163)
);

AND2x4_ASAP7_75t_L g10164 ( 
.A(n_9811),
.B(n_1160),
.Y(n_10164)
);

INVx1_ASAP7_75t_L g10165 ( 
.A(n_9920),
.Y(n_10165)
);

INVx2_ASAP7_75t_L g10166 ( 
.A(n_9953),
.Y(n_10166)
);

OAI21x1_ASAP7_75t_L g10167 ( 
.A1(n_9735),
.A2(n_503),
.B(n_504),
.Y(n_10167)
);

HB1xp67_ASAP7_75t_L g10168 ( 
.A(n_9841),
.Y(n_10168)
);

NAND2xp5_ASAP7_75t_L g10169 ( 
.A(n_9780),
.B(n_1162),
.Y(n_10169)
);

HB1xp67_ASAP7_75t_L g10170 ( 
.A(n_9889),
.Y(n_10170)
);

INVx3_ASAP7_75t_L g10171 ( 
.A(n_9736),
.Y(n_10171)
);

INVx2_ASAP7_75t_L g10172 ( 
.A(n_9917),
.Y(n_10172)
);

BUFx2_ASAP7_75t_L g10173 ( 
.A(n_9787),
.Y(n_10173)
);

OAI21x1_ASAP7_75t_L g10174 ( 
.A1(n_9946),
.A2(n_506),
.B(n_507),
.Y(n_10174)
);

INVx1_ASAP7_75t_L g10175 ( 
.A(n_9858),
.Y(n_10175)
);

INVx1_ASAP7_75t_L g10176 ( 
.A(n_9868),
.Y(n_10176)
);

INVx2_ASAP7_75t_L g10177 ( 
.A(n_9917),
.Y(n_10177)
);

OAI21x1_ASAP7_75t_L g10178 ( 
.A1(n_9967),
.A2(n_506),
.B(n_507),
.Y(n_10178)
);

HB1xp67_ASAP7_75t_L g10179 ( 
.A(n_9691),
.Y(n_10179)
);

INVx2_ASAP7_75t_L g10180 ( 
.A(n_9817),
.Y(n_10180)
);

NAND2xp5_ASAP7_75t_L g10181 ( 
.A(n_9763),
.B(n_1163),
.Y(n_10181)
);

BUFx3_ASAP7_75t_L g10182 ( 
.A(n_9892),
.Y(n_10182)
);

INVx1_ASAP7_75t_L g10183 ( 
.A(n_9724),
.Y(n_10183)
);

AOI21x1_ASAP7_75t_L g10184 ( 
.A1(n_9756),
.A2(n_506),
.B(n_508),
.Y(n_10184)
);

BUFx2_ASAP7_75t_L g10185 ( 
.A(n_9807),
.Y(n_10185)
);

INVx2_ASAP7_75t_L g10186 ( 
.A(n_9884),
.Y(n_10186)
);

INVx2_ASAP7_75t_L g10187 ( 
.A(n_9699),
.Y(n_10187)
);

INVx2_ASAP7_75t_SL g10188 ( 
.A(n_9936),
.Y(n_10188)
);

OR2x2_ASAP7_75t_L g10189 ( 
.A(n_9767),
.B(n_508),
.Y(n_10189)
);

AND2x2_ASAP7_75t_L g10190 ( 
.A(n_9921),
.B(n_509),
.Y(n_10190)
);

BUFx2_ASAP7_75t_L g10191 ( 
.A(n_9846),
.Y(n_10191)
);

INVx2_ASAP7_75t_L g10192 ( 
.A(n_9699),
.Y(n_10192)
);

INVx1_ASAP7_75t_L g10193 ( 
.A(n_9970),
.Y(n_10193)
);

INVx1_ASAP7_75t_L g10194 ( 
.A(n_9970),
.Y(n_10194)
);

INVx2_ASAP7_75t_L g10195 ( 
.A(n_9725),
.Y(n_10195)
);

INVx1_ASAP7_75t_L g10196 ( 
.A(n_9725),
.Y(n_10196)
);

INVx2_ASAP7_75t_L g10197 ( 
.A(n_9755),
.Y(n_10197)
);

AOI22xp33_ASAP7_75t_SL g10198 ( 
.A1(n_9733),
.A2(n_1164),
.B1(n_1165),
.B2(n_1163),
.Y(n_10198)
);

INVx3_ASAP7_75t_L g10199 ( 
.A(n_9801),
.Y(n_10199)
);

INVx2_ASAP7_75t_L g10200 ( 
.A(n_9755),
.Y(n_10200)
);

HB1xp67_ASAP7_75t_L g10201 ( 
.A(n_9770),
.Y(n_10201)
);

BUFx2_ASAP7_75t_L g10202 ( 
.A(n_9859),
.Y(n_10202)
);

OAI21x1_ASAP7_75t_L g10203 ( 
.A1(n_9822),
.A2(n_509),
.B(n_510),
.Y(n_10203)
);

INVxp67_ASAP7_75t_L g10204 ( 
.A(n_9847),
.Y(n_10204)
);

INVx2_ASAP7_75t_L g10205 ( 
.A(n_9770),
.Y(n_10205)
);

INVx1_ASAP7_75t_L g10206 ( 
.A(n_9824),
.Y(n_10206)
);

OAI22xp5_ASAP7_75t_L g10207 ( 
.A1(n_9856),
.A2(n_511),
.B1(n_509),
.B2(n_510),
.Y(n_10207)
);

INVx8_ASAP7_75t_L g10208 ( 
.A(n_9887),
.Y(n_10208)
);

BUFx3_ASAP7_75t_L g10209 ( 
.A(n_9717),
.Y(n_10209)
);

OA21x2_ASAP7_75t_L g10210 ( 
.A1(n_9984),
.A2(n_510),
.B(n_511),
.Y(n_10210)
);

INVx3_ASAP7_75t_L g10211 ( 
.A(n_9808),
.Y(n_10211)
);

HB1xp67_ASAP7_75t_L g10212 ( 
.A(n_9824),
.Y(n_10212)
);

INVx1_ASAP7_75t_L g10213 ( 
.A(n_9883),
.Y(n_10213)
);

INVx2_ASAP7_75t_L g10214 ( 
.A(n_9883),
.Y(n_10214)
);

INVx1_ASAP7_75t_L g10215 ( 
.A(n_9820),
.Y(n_10215)
);

INVx1_ASAP7_75t_L g10216 ( 
.A(n_9837),
.Y(n_10216)
);

INVx1_ASAP7_75t_L g10217 ( 
.A(n_9878),
.Y(n_10217)
);

BUFx2_ASAP7_75t_L g10218 ( 
.A(n_9948),
.Y(n_10218)
);

INVx1_ASAP7_75t_L g10219 ( 
.A(n_9885),
.Y(n_10219)
);

HB1xp67_ASAP7_75t_L g10220 ( 
.A(n_9704),
.Y(n_10220)
);

BUFx3_ASAP7_75t_L g10221 ( 
.A(n_9707),
.Y(n_10221)
);

INVx3_ASAP7_75t_L g10222 ( 
.A(n_9722),
.Y(n_10222)
);

INVx1_ASAP7_75t_L g10223 ( 
.A(n_9831),
.Y(n_10223)
);

INVx2_ASAP7_75t_L g10224 ( 
.A(n_9974),
.Y(n_10224)
);

INVx8_ASAP7_75t_L g10225 ( 
.A(n_9804),
.Y(n_10225)
);

OAI21x1_ASAP7_75t_L g10226 ( 
.A1(n_9776),
.A2(n_511),
.B(n_512),
.Y(n_10226)
);

AOI22xp33_ASAP7_75t_SL g10227 ( 
.A1(n_9976),
.A2(n_1167),
.B1(n_1169),
.B2(n_1166),
.Y(n_10227)
);

BUFx2_ASAP7_75t_L g10228 ( 
.A(n_9741),
.Y(n_10228)
);

INVx2_ASAP7_75t_L g10229 ( 
.A(n_9959),
.Y(n_10229)
);

INVx3_ASAP7_75t_L g10230 ( 
.A(n_9779),
.Y(n_10230)
);

BUFx6f_ASAP7_75t_L g10231 ( 
.A(n_9751),
.Y(n_10231)
);

BUFx4f_ASAP7_75t_L g10232 ( 
.A(n_9986),
.Y(n_10232)
);

AND2x2_ASAP7_75t_L g10233 ( 
.A(n_9900),
.B(n_512),
.Y(n_10233)
);

INVx3_ASAP7_75t_L g10234 ( 
.A(n_9964),
.Y(n_10234)
);

INVx2_ASAP7_75t_SL g10235 ( 
.A(n_9913),
.Y(n_10235)
);

INVx2_ASAP7_75t_L g10236 ( 
.A(n_9894),
.Y(n_10236)
);

INVx1_ASAP7_75t_SL g10237 ( 
.A(n_9695),
.Y(n_10237)
);

INVx1_ASAP7_75t_L g10238 ( 
.A(n_9960),
.Y(n_10238)
);

INVx1_ASAP7_75t_L g10239 ( 
.A(n_9914),
.Y(n_10239)
);

AND2x2_ASAP7_75t_L g10240 ( 
.A(n_9775),
.B(n_512),
.Y(n_10240)
);

CKINVDCx11_ASAP7_75t_R g10241 ( 
.A(n_9954),
.Y(n_10241)
);

INVx3_ASAP7_75t_L g10242 ( 
.A(n_9762),
.Y(n_10242)
);

OR2x2_ASAP7_75t_L g10243 ( 
.A(n_9698),
.B(n_9714),
.Y(n_10243)
);

HB1xp67_ASAP7_75t_L g10244 ( 
.A(n_9834),
.Y(n_10244)
);

OR2x6_ASAP7_75t_L g10245 ( 
.A(n_9909),
.B(n_1167),
.Y(n_10245)
);

OAI22xp5_ASAP7_75t_L g10246 ( 
.A1(n_9895),
.A2(n_515),
.B1(n_513),
.B2(n_514),
.Y(n_10246)
);

INVx1_ASAP7_75t_L g10247 ( 
.A(n_9971),
.Y(n_10247)
);

HB1xp67_ASAP7_75t_L g10248 ( 
.A(n_9825),
.Y(n_10248)
);

INVx2_ASAP7_75t_L g10249 ( 
.A(n_9805),
.Y(n_10249)
);

INVx2_ASAP7_75t_L g10250 ( 
.A(n_9727),
.Y(n_10250)
);

INVx2_ASAP7_75t_L g10251 ( 
.A(n_9782),
.Y(n_10251)
);

AO21x2_ASAP7_75t_L g10252 ( 
.A1(n_9957),
.A2(n_513),
.B(n_514),
.Y(n_10252)
);

INVx1_ASAP7_75t_L g10253 ( 
.A(n_9692),
.Y(n_10253)
);

AOI221xp5_ASAP7_75t_L g10254 ( 
.A1(n_9979),
.A2(n_516),
.B1(n_513),
.B2(n_515),
.C(n_517),
.Y(n_10254)
);

INVxp67_ASAP7_75t_SL g10255 ( 
.A(n_9930),
.Y(n_10255)
);

INVx1_ASAP7_75t_L g10256 ( 
.A(n_9962),
.Y(n_10256)
);

INVx1_ASAP7_75t_L g10257 ( 
.A(n_9915),
.Y(n_10257)
);

AOI221xp5_ASAP7_75t_L g10258 ( 
.A1(n_9903),
.A2(n_517),
.B1(n_515),
.B2(n_516),
.C(n_518),
.Y(n_10258)
);

BUFx3_ASAP7_75t_L g10259 ( 
.A(n_9897),
.Y(n_10259)
);

BUFx2_ASAP7_75t_L g10260 ( 
.A(n_9836),
.Y(n_10260)
);

NAND2xp5_ASAP7_75t_L g10261 ( 
.A(n_9693),
.B(n_1169),
.Y(n_10261)
);

HB1xp67_ASAP7_75t_L g10262 ( 
.A(n_9955),
.Y(n_10262)
);

BUFx3_ASAP7_75t_L g10263 ( 
.A(n_9788),
.Y(n_10263)
);

NAND2xp5_ASAP7_75t_L g10264 ( 
.A(n_9972),
.B(n_1170),
.Y(n_10264)
);

HB1xp67_ASAP7_75t_L g10265 ( 
.A(n_9939),
.Y(n_10265)
);

INVx1_ASAP7_75t_L g10266 ( 
.A(n_9798),
.Y(n_10266)
);

INVx1_ASAP7_75t_L g10267 ( 
.A(n_9942),
.Y(n_10267)
);

INVx2_ASAP7_75t_L g10268 ( 
.A(n_9853),
.Y(n_10268)
);

AOI21x1_ASAP7_75t_L g10269 ( 
.A1(n_9940),
.A2(n_9720),
.B(n_9918),
.Y(n_10269)
);

AOI22xp33_ASAP7_75t_L g10270 ( 
.A1(n_9864),
.A2(n_1171),
.B1(n_1172),
.B2(n_1170),
.Y(n_10270)
);

OAI21x1_ASAP7_75t_L g10271 ( 
.A1(n_9843),
.A2(n_518),
.B(n_519),
.Y(n_10271)
);

BUFx3_ASAP7_75t_L g10272 ( 
.A(n_9706),
.Y(n_10272)
);

AND2x2_ASAP7_75t_L g10273 ( 
.A(n_9860),
.B(n_518),
.Y(n_10273)
);

OAI22xp5_ASAP7_75t_L g10274 ( 
.A1(n_9855),
.A2(n_521),
.B1(n_519),
.B2(n_520),
.Y(n_10274)
);

HB1xp67_ASAP7_75t_L g10275 ( 
.A(n_9929),
.Y(n_10275)
);

INVx1_ASAP7_75t_L g10276 ( 
.A(n_9941),
.Y(n_10276)
);

OAI21x1_ASAP7_75t_L g10277 ( 
.A1(n_9861),
.A2(n_519),
.B(n_520),
.Y(n_10277)
);

CKINVDCx20_ASAP7_75t_R g10278 ( 
.A(n_10063),
.Y(n_10278)
);

INVx1_ASAP7_75t_L g10279 ( 
.A(n_10041),
.Y(n_10279)
);

INVx2_ASAP7_75t_L g10280 ( 
.A(n_10001),
.Y(n_10280)
);

BUFx3_ASAP7_75t_L g10281 ( 
.A(n_10057),
.Y(n_10281)
);

INVx2_ASAP7_75t_L g10282 ( 
.A(n_10026),
.Y(n_10282)
);

INVx3_ASAP7_75t_L g10283 ( 
.A(n_10151),
.Y(n_10283)
);

OAI21xp5_ASAP7_75t_L g10284 ( 
.A1(n_10101),
.A2(n_9937),
.B(n_9949),
.Y(n_10284)
);

INVx2_ASAP7_75t_L g10285 ( 
.A(n_10116),
.Y(n_10285)
);

BUFx6f_ASAP7_75t_L g10286 ( 
.A(n_10057),
.Y(n_10286)
);

OAI21xp5_ASAP7_75t_L g10287 ( 
.A1(n_10028),
.A2(n_9947),
.B(n_9980),
.Y(n_10287)
);

OR2x2_ASAP7_75t_L g10288 ( 
.A(n_9992),
.B(n_10022),
.Y(n_10288)
);

NOR2x1_ASAP7_75t_SL g10289 ( 
.A(n_10127),
.B(n_9969),
.Y(n_10289)
);

INVx1_ASAP7_75t_L g10290 ( 
.A(n_10043),
.Y(n_10290)
);

INVx1_ASAP7_75t_L g10291 ( 
.A(n_10045),
.Y(n_10291)
);

INVx2_ASAP7_75t_L g10292 ( 
.A(n_10122),
.Y(n_10292)
);

INVx3_ASAP7_75t_L g10293 ( 
.A(n_10182),
.Y(n_10293)
);

NAND3xp33_ASAP7_75t_L g10294 ( 
.A(n_10025),
.B(n_9978),
.C(n_9968),
.Y(n_10294)
);

INVx1_ASAP7_75t_L g10295 ( 
.A(n_9990),
.Y(n_10295)
);

INVx1_ASAP7_75t_L g10296 ( 
.A(n_9997),
.Y(n_10296)
);

INVx1_ASAP7_75t_L g10297 ( 
.A(n_9999),
.Y(n_10297)
);

INVx2_ASAP7_75t_L g10298 ( 
.A(n_10051),
.Y(n_10298)
);

INVx1_ASAP7_75t_L g10299 ( 
.A(n_10003),
.Y(n_10299)
);

INVx2_ASAP7_75t_L g10300 ( 
.A(n_10061),
.Y(n_10300)
);

INVx2_ASAP7_75t_L g10301 ( 
.A(n_10236),
.Y(n_10301)
);

OA21x2_ASAP7_75t_L g10302 ( 
.A1(n_10162),
.A2(n_9951),
.B(n_9916),
.Y(n_10302)
);

BUFx6f_ASAP7_75t_L g10303 ( 
.A(n_10067),
.Y(n_10303)
);

INVx2_ASAP7_75t_SL g10304 ( 
.A(n_10130),
.Y(n_10304)
);

INVx2_ASAP7_75t_L g10305 ( 
.A(n_10065),
.Y(n_10305)
);

INVx2_ASAP7_75t_L g10306 ( 
.A(n_10035),
.Y(n_10306)
);

INVx1_ASAP7_75t_L g10307 ( 
.A(n_10005),
.Y(n_10307)
);

BUFx2_ASAP7_75t_L g10308 ( 
.A(n_10131),
.Y(n_10308)
);

AND2x2_ASAP7_75t_L g10309 ( 
.A(n_10223),
.B(n_9880),
.Y(n_10309)
);

INVx2_ASAP7_75t_L g10310 ( 
.A(n_10039),
.Y(n_10310)
);

OR2x6_ASAP7_75t_L g10311 ( 
.A(n_10208),
.B(n_10049),
.Y(n_10311)
);

CKINVDCx20_ASAP7_75t_R g10312 ( 
.A(n_10241),
.Y(n_10312)
);

BUFx4f_ASAP7_75t_L g10313 ( 
.A(n_10067),
.Y(n_10313)
);

INVx2_ASAP7_75t_SL g10314 ( 
.A(n_10130),
.Y(n_10314)
);

INVx2_ASAP7_75t_L g10315 ( 
.A(n_10048),
.Y(n_10315)
);

INVx1_ASAP7_75t_L g10316 ( 
.A(n_10010),
.Y(n_10316)
);

AND2x2_ASAP7_75t_L g10317 ( 
.A(n_10054),
.B(n_9926),
.Y(n_10317)
);

HB1xp67_ASAP7_75t_L g10318 ( 
.A(n_10031),
.Y(n_10318)
);

INVx1_ASAP7_75t_L g10319 ( 
.A(n_10011),
.Y(n_10319)
);

INVx2_ASAP7_75t_L g10320 ( 
.A(n_10092),
.Y(n_10320)
);

HB1xp67_ASAP7_75t_L g10321 ( 
.A(n_10044),
.Y(n_10321)
);

AND2x4_ASAP7_75t_L g10322 ( 
.A(n_10058),
.B(n_9933),
.Y(n_10322)
);

INVx1_ASAP7_75t_L g10323 ( 
.A(n_10012),
.Y(n_10323)
);

BUFx12f_ASAP7_75t_L g10324 ( 
.A(n_10231),
.Y(n_10324)
);

INVx1_ASAP7_75t_L g10325 ( 
.A(n_10013),
.Y(n_10325)
);

AND2x2_ASAP7_75t_L g10326 ( 
.A(n_10244),
.B(n_9931),
.Y(n_10326)
);

OAI21x1_ASAP7_75t_L g10327 ( 
.A1(n_9987),
.A2(n_9934),
.B(n_520),
.Y(n_10327)
);

AND2x2_ASAP7_75t_L g10328 ( 
.A(n_10119),
.B(n_521),
.Y(n_10328)
);

INVx1_ASAP7_75t_L g10329 ( 
.A(n_10018),
.Y(n_10329)
);

INVx1_ASAP7_75t_L g10330 ( 
.A(n_10020),
.Y(n_10330)
);

HB1xp67_ASAP7_75t_L g10331 ( 
.A(n_10102),
.Y(n_10331)
);

INVx1_ASAP7_75t_L g10332 ( 
.A(n_10021),
.Y(n_10332)
);

INVx1_ASAP7_75t_L g10333 ( 
.A(n_10024),
.Y(n_10333)
);

INVx2_ASAP7_75t_L g10334 ( 
.A(n_10077),
.Y(n_10334)
);

NAND2x1p5_ASAP7_75t_L g10335 ( 
.A(n_9996),
.B(n_521),
.Y(n_10335)
);

OR2x2_ASAP7_75t_L g10336 ( 
.A(n_10118),
.B(n_10002),
.Y(n_10336)
);

INVx2_ASAP7_75t_L g10337 ( 
.A(n_10081),
.Y(n_10337)
);

INVx1_ASAP7_75t_L g10338 ( 
.A(n_10027),
.Y(n_10338)
);

INVx1_ASAP7_75t_L g10339 ( 
.A(n_10047),
.Y(n_10339)
);

INVx1_ASAP7_75t_L g10340 ( 
.A(n_10053),
.Y(n_10340)
);

INVx2_ASAP7_75t_L g10341 ( 
.A(n_10087),
.Y(n_10341)
);

NAND2xp5_ASAP7_75t_L g10342 ( 
.A(n_10152),
.B(n_1171),
.Y(n_10342)
);

NAND2xp5_ASAP7_75t_L g10343 ( 
.A(n_10090),
.B(n_1173),
.Y(n_10343)
);

OAI21x1_ASAP7_75t_L g10344 ( 
.A1(n_9994),
.A2(n_522),
.B(n_523),
.Y(n_10344)
);

OR2x2_ASAP7_75t_L g10345 ( 
.A(n_10037),
.B(n_522),
.Y(n_10345)
);

INVx1_ASAP7_75t_L g10346 ( 
.A(n_10060),
.Y(n_10346)
);

AND2x2_ASAP7_75t_L g10347 ( 
.A(n_10052),
.B(n_522),
.Y(n_10347)
);

AND2x2_ASAP7_75t_L g10348 ( 
.A(n_10008),
.B(n_523),
.Y(n_10348)
);

INVx1_ASAP7_75t_L g10349 ( 
.A(n_10068),
.Y(n_10349)
);

HB1xp67_ASAP7_75t_L g10350 ( 
.A(n_10089),
.Y(n_10350)
);

AND2x2_ASAP7_75t_L g10351 ( 
.A(n_10224),
.B(n_524),
.Y(n_10351)
);

INVx1_ASAP7_75t_L g10352 ( 
.A(n_10079),
.Y(n_10352)
);

OR2x2_ASAP7_75t_L g10353 ( 
.A(n_10111),
.B(n_524),
.Y(n_10353)
);

INVx1_ASAP7_75t_L g10354 ( 
.A(n_10064),
.Y(n_10354)
);

AND2x4_ASAP7_75t_L g10355 ( 
.A(n_10083),
.B(n_524),
.Y(n_10355)
);

INVx1_ASAP7_75t_L g10356 ( 
.A(n_10038),
.Y(n_10356)
);

INVx2_ASAP7_75t_L g10357 ( 
.A(n_10088),
.Y(n_10357)
);

INVx2_ASAP7_75t_L g10358 ( 
.A(n_10075),
.Y(n_10358)
);

INVx2_ASAP7_75t_L g10359 ( 
.A(n_10104),
.Y(n_10359)
);

BUFx6f_ASAP7_75t_L g10360 ( 
.A(n_10231),
.Y(n_10360)
);

INVx1_ASAP7_75t_L g10361 ( 
.A(n_10046),
.Y(n_10361)
);

AND2x2_ASAP7_75t_L g10362 ( 
.A(n_10193),
.B(n_525),
.Y(n_10362)
);

AOI21x1_ASAP7_75t_L g10363 ( 
.A1(n_10160),
.A2(n_525),
.B(n_526),
.Y(n_10363)
);

INVx1_ASAP7_75t_L g10364 ( 
.A(n_10106),
.Y(n_10364)
);

INVx2_ASAP7_75t_L g10365 ( 
.A(n_10029),
.Y(n_10365)
);

INVx1_ASAP7_75t_L g10366 ( 
.A(n_10069),
.Y(n_10366)
);

INVx2_ASAP7_75t_L g10367 ( 
.A(n_10034),
.Y(n_10367)
);

INVx1_ASAP7_75t_L g10368 ( 
.A(n_10070),
.Y(n_10368)
);

INVx2_ASAP7_75t_L g10369 ( 
.A(n_10023),
.Y(n_10369)
);

INVx1_ASAP7_75t_L g10370 ( 
.A(n_10071),
.Y(n_10370)
);

INVx1_ASAP7_75t_L g10371 ( 
.A(n_10072),
.Y(n_10371)
);

NOR2xp33_ASAP7_75t_SL g10372 ( 
.A(n_10121),
.B(n_1173),
.Y(n_10372)
);

BUFx2_ASAP7_75t_L g10373 ( 
.A(n_10014),
.Y(n_10373)
);

AND2x2_ASAP7_75t_L g10374 ( 
.A(n_10194),
.B(n_525),
.Y(n_10374)
);

INVx3_ASAP7_75t_L g10375 ( 
.A(n_10222),
.Y(n_10375)
);

INVx1_ASAP7_75t_L g10376 ( 
.A(n_10073),
.Y(n_10376)
);

AND2x2_ASAP7_75t_L g10377 ( 
.A(n_10172),
.B(n_527),
.Y(n_10377)
);

AND2x2_ASAP7_75t_L g10378 ( 
.A(n_10177),
.B(n_527),
.Y(n_10378)
);

INVx2_ASAP7_75t_L g10379 ( 
.A(n_10094),
.Y(n_10379)
);

INVx2_ASAP7_75t_SL g10380 ( 
.A(n_10225),
.Y(n_10380)
);

INVx4_ASAP7_75t_SL g10381 ( 
.A(n_10221),
.Y(n_10381)
);

INVx3_ASAP7_75t_L g10382 ( 
.A(n_10016),
.Y(n_10382)
);

INVx2_ASAP7_75t_L g10383 ( 
.A(n_10100),
.Y(n_10383)
);

INVx1_ASAP7_75t_L g10384 ( 
.A(n_10078),
.Y(n_10384)
);

INVx2_ASAP7_75t_L g10385 ( 
.A(n_10103),
.Y(n_10385)
);

AND2x2_ASAP7_75t_L g10386 ( 
.A(n_10149),
.B(n_527),
.Y(n_10386)
);

INVx2_ASAP7_75t_L g10387 ( 
.A(n_9995),
.Y(n_10387)
);

INVx2_ASAP7_75t_L g10388 ( 
.A(n_10006),
.Y(n_10388)
);

INVx1_ASAP7_75t_L g10389 ( 
.A(n_9993),
.Y(n_10389)
);

AO21x2_ASAP7_75t_L g10390 ( 
.A1(n_10015),
.A2(n_528),
.B(n_529),
.Y(n_10390)
);

OR2x2_ASAP7_75t_L g10391 ( 
.A(n_10117),
.B(n_528),
.Y(n_10391)
);

INVx4_ASAP7_75t_L g10392 ( 
.A(n_10080),
.Y(n_10392)
);

HB1xp67_ASAP7_75t_L g10393 ( 
.A(n_10097),
.Y(n_10393)
);

INVx1_ASAP7_75t_L g10394 ( 
.A(n_9989),
.Y(n_10394)
);

INVx2_ASAP7_75t_L g10395 ( 
.A(n_10032),
.Y(n_10395)
);

AND2x2_ASAP7_75t_L g10396 ( 
.A(n_10179),
.B(n_529),
.Y(n_10396)
);

NOR2xp33_ASAP7_75t_SL g10397 ( 
.A(n_10128),
.B(n_1174),
.Y(n_10397)
);

INVx1_ASAP7_75t_L g10398 ( 
.A(n_10112),
.Y(n_10398)
);

HB1xp67_ASAP7_75t_L g10399 ( 
.A(n_10133),
.Y(n_10399)
);

INVx1_ASAP7_75t_L g10400 ( 
.A(n_10109),
.Y(n_10400)
);

INVx3_ASAP7_75t_L g10401 ( 
.A(n_10209),
.Y(n_10401)
);

INVxp67_ASAP7_75t_L g10402 ( 
.A(n_10210),
.Y(n_10402)
);

CKINVDCx20_ASAP7_75t_R g10403 ( 
.A(n_10099),
.Y(n_10403)
);

INVx1_ASAP7_75t_L g10404 ( 
.A(n_10076),
.Y(n_10404)
);

INVx3_ASAP7_75t_L g10405 ( 
.A(n_10225),
.Y(n_10405)
);

OAI21xp5_ASAP7_75t_L g10406 ( 
.A1(n_10017),
.A2(n_530),
.B(n_531),
.Y(n_10406)
);

INVx2_ASAP7_75t_L g10407 ( 
.A(n_10066),
.Y(n_10407)
);

INVx1_ASAP7_75t_L g10408 ( 
.A(n_10086),
.Y(n_10408)
);

INVx1_ASAP7_75t_L g10409 ( 
.A(n_10123),
.Y(n_10409)
);

INVx3_ASAP7_75t_L g10410 ( 
.A(n_10230),
.Y(n_10410)
);

INVx2_ASAP7_75t_SL g10411 ( 
.A(n_10208),
.Y(n_10411)
);

AO21x2_ASAP7_75t_L g10412 ( 
.A1(n_9988),
.A2(n_530),
.B(n_531),
.Y(n_10412)
);

AO21x2_ASAP7_75t_L g10413 ( 
.A1(n_10040),
.A2(n_530),
.B(n_531),
.Y(n_10413)
);

BUFx2_ASAP7_75t_L g10414 ( 
.A(n_10014),
.Y(n_10414)
);

INVx1_ASAP7_75t_L g10415 ( 
.A(n_10139),
.Y(n_10415)
);

INVx1_ASAP7_75t_L g10416 ( 
.A(n_10150),
.Y(n_10416)
);

INVx2_ASAP7_75t_L g10417 ( 
.A(n_10186),
.Y(n_10417)
);

INVx2_ASAP7_75t_L g10418 ( 
.A(n_10126),
.Y(n_10418)
);

AND2x2_ASAP7_75t_L g10419 ( 
.A(n_10201),
.B(n_532),
.Y(n_10419)
);

OR2x6_ASAP7_75t_L g10420 ( 
.A(n_10082),
.B(n_1174),
.Y(n_10420)
);

INVx2_ASAP7_75t_SL g10421 ( 
.A(n_10007),
.Y(n_10421)
);

INVx1_ASAP7_75t_SL g10422 ( 
.A(n_10019),
.Y(n_10422)
);

BUFx3_ASAP7_75t_L g10423 ( 
.A(n_10000),
.Y(n_10423)
);

INVx2_ASAP7_75t_L g10424 ( 
.A(n_10220),
.Y(n_10424)
);

INVx2_ASAP7_75t_L g10425 ( 
.A(n_10135),
.Y(n_10425)
);

INVx2_ASAP7_75t_L g10426 ( 
.A(n_10136),
.Y(n_10426)
);

INVx1_ASAP7_75t_L g10427 ( 
.A(n_10120),
.Y(n_10427)
);

BUFx6f_ASAP7_75t_L g10428 ( 
.A(n_10138),
.Y(n_10428)
);

AND2x2_ASAP7_75t_L g10429 ( 
.A(n_10212),
.B(n_532),
.Y(n_10429)
);

AND2x2_ASAP7_75t_L g10430 ( 
.A(n_10132),
.B(n_532),
.Y(n_10430)
);

INVx1_ASAP7_75t_L g10431 ( 
.A(n_10125),
.Y(n_10431)
);

INVx1_ASAP7_75t_L g10432 ( 
.A(n_10085),
.Y(n_10432)
);

INVx2_ASAP7_75t_L g10433 ( 
.A(n_10185),
.Y(n_10433)
);

AND2x2_ASAP7_75t_L g10434 ( 
.A(n_10170),
.B(n_533),
.Y(n_10434)
);

INVx3_ASAP7_75t_L g10435 ( 
.A(n_10055),
.Y(n_10435)
);

INVx1_ASAP7_75t_L g10436 ( 
.A(n_10085),
.Y(n_10436)
);

INVx1_ASAP7_75t_L g10437 ( 
.A(n_10036),
.Y(n_10437)
);

OAI21x1_ASAP7_75t_L g10438 ( 
.A1(n_10146),
.A2(n_533),
.B(n_534),
.Y(n_10438)
);

BUFx2_ASAP7_75t_L g10439 ( 
.A(n_10191),
.Y(n_10439)
);

HB1xp67_ASAP7_75t_L g10440 ( 
.A(n_10096),
.Y(n_10440)
);

HB1xp67_ASAP7_75t_L g10441 ( 
.A(n_10096),
.Y(n_10441)
);

INVx1_ASAP7_75t_L g10442 ( 
.A(n_10137),
.Y(n_10442)
);

OA21x2_ASAP7_75t_L g10443 ( 
.A1(n_10253),
.A2(n_534),
.B(n_535),
.Y(n_10443)
);

INVx1_ASAP7_75t_SL g10444 ( 
.A(n_10228),
.Y(n_10444)
);

INVx2_ASAP7_75t_L g10445 ( 
.A(n_10202),
.Y(n_10445)
);

OA21x2_ASAP7_75t_L g10446 ( 
.A1(n_10266),
.A2(n_534),
.B(n_535),
.Y(n_10446)
);

INVx1_ASAP7_75t_L g10447 ( 
.A(n_10238),
.Y(n_10447)
);

OAI21x1_ASAP7_75t_L g10448 ( 
.A1(n_10148),
.A2(n_536),
.B(n_537),
.Y(n_10448)
);

HB1xp67_ASAP7_75t_L g10449 ( 
.A(n_10059),
.Y(n_10449)
);

INVx2_ASAP7_75t_L g10450 ( 
.A(n_10173),
.Y(n_10450)
);

INVx1_ASAP7_75t_L g10451 ( 
.A(n_10115),
.Y(n_10451)
);

INVx2_ASAP7_75t_L g10452 ( 
.A(n_10187),
.Y(n_10452)
);

HB1xp67_ASAP7_75t_L g10453 ( 
.A(n_10248),
.Y(n_10453)
);

INVx2_ASAP7_75t_L g10454 ( 
.A(n_10192),
.Y(n_10454)
);

OR2x2_ASAP7_75t_L g10455 ( 
.A(n_10249),
.B(n_536),
.Y(n_10455)
);

INVx2_ASAP7_75t_L g10456 ( 
.A(n_10195),
.Y(n_10456)
);

BUFx3_ASAP7_75t_L g10457 ( 
.A(n_9998),
.Y(n_10457)
);

INVx1_ASAP7_75t_L g10458 ( 
.A(n_10050),
.Y(n_10458)
);

INVx1_ASAP7_75t_L g10459 ( 
.A(n_10247),
.Y(n_10459)
);

INVx2_ASAP7_75t_L g10460 ( 
.A(n_10197),
.Y(n_10460)
);

INVx1_ASAP7_75t_L g10461 ( 
.A(n_10140),
.Y(n_10461)
);

INVx1_ASAP7_75t_L g10462 ( 
.A(n_10262),
.Y(n_10462)
);

NAND2xp5_ASAP7_75t_L g10463 ( 
.A(n_10183),
.B(n_1175),
.Y(n_10463)
);

INVx2_ASAP7_75t_L g10464 ( 
.A(n_10200),
.Y(n_10464)
);

INVx1_ASAP7_75t_L g10465 ( 
.A(n_10134),
.Y(n_10465)
);

OA21x2_ASAP7_75t_L g10466 ( 
.A1(n_10204),
.A2(n_536),
.B(n_537),
.Y(n_10466)
);

BUFx3_ASAP7_75t_L g10467 ( 
.A(n_10232),
.Y(n_10467)
);

INVx1_ASAP7_75t_L g10468 ( 
.A(n_10265),
.Y(n_10468)
);

AO21x1_ASAP7_75t_SL g10469 ( 
.A1(n_10243),
.A2(n_537),
.B(n_538),
.Y(n_10469)
);

AO21x2_ASAP7_75t_L g10470 ( 
.A1(n_10169),
.A2(n_538),
.B(n_539),
.Y(n_10470)
);

INVxp67_ASAP7_75t_SL g10471 ( 
.A(n_10263),
.Y(n_10471)
);

OA21x2_ASAP7_75t_L g10472 ( 
.A1(n_10239),
.A2(n_538),
.B(n_539),
.Y(n_10472)
);

INVx2_ASAP7_75t_SL g10473 ( 
.A(n_10218),
.Y(n_10473)
);

HB1xp67_ASAP7_75t_L g10474 ( 
.A(n_10168),
.Y(n_10474)
);

HB1xp67_ASAP7_75t_L g10475 ( 
.A(n_10156),
.Y(n_10475)
);

INVx3_ASAP7_75t_L g10476 ( 
.A(n_10171),
.Y(n_10476)
);

INVx2_ASAP7_75t_L g10477 ( 
.A(n_10205),
.Y(n_10477)
);

AND2x2_ASAP7_75t_L g10478 ( 
.A(n_10154),
.B(n_540),
.Y(n_10478)
);

INVx2_ASAP7_75t_L g10479 ( 
.A(n_10214),
.Y(n_10479)
);

BUFx2_ASAP7_75t_L g10480 ( 
.A(n_10062),
.Y(n_10480)
);

AND2x2_ASAP7_75t_L g10481 ( 
.A(n_10166),
.B(n_540),
.Y(n_10481)
);

CKINVDCx16_ASAP7_75t_R g10482 ( 
.A(n_10240),
.Y(n_10482)
);

HB1xp67_ASAP7_75t_L g10483 ( 
.A(n_10145),
.Y(n_10483)
);

INVx2_ASAP7_75t_L g10484 ( 
.A(n_10196),
.Y(n_10484)
);

AND2x2_ASAP7_75t_L g10485 ( 
.A(n_10229),
.B(n_10206),
.Y(n_10485)
);

INVx1_ASAP7_75t_L g10486 ( 
.A(n_10213),
.Y(n_10486)
);

INVx1_ASAP7_75t_L g10487 ( 
.A(n_10163),
.Y(n_10487)
);

BUFx3_ASAP7_75t_L g10488 ( 
.A(n_10009),
.Y(n_10488)
);

INVx1_ASAP7_75t_L g10489 ( 
.A(n_10107),
.Y(n_10489)
);

INVx1_ASAP7_75t_L g10490 ( 
.A(n_10147),
.Y(n_10490)
);

OAI21xp5_ASAP7_75t_L g10491 ( 
.A1(n_10275),
.A2(n_540),
.B(n_541),
.Y(n_10491)
);

INVx2_ASAP7_75t_L g10492 ( 
.A(n_10110),
.Y(n_10492)
);

INVx1_ASAP7_75t_L g10493 ( 
.A(n_10084),
.Y(n_10493)
);

INVx1_ASAP7_75t_L g10494 ( 
.A(n_10091),
.Y(n_10494)
);

BUFx2_ASAP7_75t_L g10495 ( 
.A(n_10030),
.Y(n_10495)
);

AND2x2_ASAP7_75t_L g10496 ( 
.A(n_10105),
.B(n_10165),
.Y(n_10496)
);

INVx1_ASAP7_75t_L g10497 ( 
.A(n_10256),
.Y(n_10497)
);

INVx1_ASAP7_75t_L g10498 ( 
.A(n_10144),
.Y(n_10498)
);

AND2x2_ASAP7_75t_L g10499 ( 
.A(n_10143),
.B(n_10155),
.Y(n_10499)
);

OR2x2_ASAP7_75t_L g10500 ( 
.A(n_10158),
.B(n_541),
.Y(n_10500)
);

INVx2_ASAP7_75t_L g10501 ( 
.A(n_10159),
.Y(n_10501)
);

INVx2_ASAP7_75t_SL g10502 ( 
.A(n_10199),
.Y(n_10502)
);

INVxp67_ASAP7_75t_SL g10503 ( 
.A(n_10211),
.Y(n_10503)
);

INVx4_ASAP7_75t_L g10504 ( 
.A(n_10164),
.Y(n_10504)
);

BUFx2_ASAP7_75t_L g10505 ( 
.A(n_10242),
.Y(n_10505)
);

INVx2_ASAP7_75t_L g10506 ( 
.A(n_10095),
.Y(n_10506)
);

INVx1_ASAP7_75t_L g10507 ( 
.A(n_10184),
.Y(n_10507)
);

INVx2_ASAP7_75t_L g10508 ( 
.A(n_10175),
.Y(n_10508)
);

INVx1_ASAP7_75t_L g10509 ( 
.A(n_10176),
.Y(n_10509)
);

INVx2_ASAP7_75t_L g10510 ( 
.A(n_10215),
.Y(n_10510)
);

NOR2x1_ASAP7_75t_SL g10511 ( 
.A(n_10245),
.B(n_541),
.Y(n_10511)
);

INVx1_ASAP7_75t_L g10512 ( 
.A(n_10276),
.Y(n_10512)
);

OAI21x1_ASAP7_75t_L g10513 ( 
.A1(n_10234),
.A2(n_542),
.B(n_543),
.Y(n_10513)
);

BUFx3_ASAP7_75t_L g10514 ( 
.A(n_10237),
.Y(n_10514)
);

INVx2_ASAP7_75t_L g10515 ( 
.A(n_10216),
.Y(n_10515)
);

OR2x6_ASAP7_75t_L g10516 ( 
.A(n_10245),
.B(n_1175),
.Y(n_10516)
);

OR2x2_ASAP7_75t_L g10517 ( 
.A(n_10255),
.B(n_542),
.Y(n_10517)
);

INVx1_ASAP7_75t_L g10518 ( 
.A(n_10217),
.Y(n_10518)
);

AO21x2_ASAP7_75t_L g10519 ( 
.A1(n_10190),
.A2(n_542),
.B(n_543),
.Y(n_10519)
);

AO21x2_ASAP7_75t_L g10520 ( 
.A1(n_10233),
.A2(n_543),
.B(n_544),
.Y(n_10520)
);

AND2x2_ASAP7_75t_L g10521 ( 
.A(n_10219),
.B(n_544),
.Y(n_10521)
);

INVx3_ASAP7_75t_L g10522 ( 
.A(n_10142),
.Y(n_10522)
);

AND2x2_ASAP7_75t_L g10523 ( 
.A(n_10180),
.B(n_544),
.Y(n_10523)
);

INVx2_ASAP7_75t_SL g10524 ( 
.A(n_10235),
.Y(n_10524)
);

BUFx3_ASAP7_75t_L g10525 ( 
.A(n_10056),
.Y(n_10525)
);

INVx1_ASAP7_75t_L g10526 ( 
.A(n_10272),
.Y(n_10526)
);

AND2x4_ASAP7_75t_L g10527 ( 
.A(n_10188),
.B(n_545),
.Y(n_10527)
);

INVx3_ASAP7_75t_L g10528 ( 
.A(n_10113),
.Y(n_10528)
);

INVx1_ASAP7_75t_L g10529 ( 
.A(n_10257),
.Y(n_10529)
);

CKINVDCx20_ASAP7_75t_R g10530 ( 
.A(n_10129),
.Y(n_10530)
);

INVx2_ASAP7_75t_L g10531 ( 
.A(n_10260),
.Y(n_10531)
);

INVx1_ASAP7_75t_L g10532 ( 
.A(n_10252),
.Y(n_10532)
);

AND2x2_ASAP7_75t_L g10533 ( 
.A(n_10033),
.B(n_545),
.Y(n_10533)
);

INVx1_ASAP7_75t_L g10534 ( 
.A(n_10167),
.Y(n_10534)
);

INVx2_ASAP7_75t_L g10535 ( 
.A(n_10259),
.Y(n_10535)
);

INVx2_ASAP7_75t_L g10536 ( 
.A(n_10226),
.Y(n_10536)
);

BUFx2_ASAP7_75t_L g10537 ( 
.A(n_10251),
.Y(n_10537)
);

HB1xp67_ASAP7_75t_L g10538 ( 
.A(n_10203),
.Y(n_10538)
);

INVx1_ASAP7_75t_L g10539 ( 
.A(n_10189),
.Y(n_10539)
);

AND2x2_ASAP7_75t_L g10540 ( 
.A(n_10098),
.B(n_545),
.Y(n_10540)
);

INVx1_ASAP7_75t_L g10541 ( 
.A(n_10181),
.Y(n_10541)
);

INVx1_ASAP7_75t_L g10542 ( 
.A(n_10267),
.Y(n_10542)
);

HB1xp67_ASAP7_75t_L g10543 ( 
.A(n_10178),
.Y(n_10543)
);

INVx2_ASAP7_75t_L g10544 ( 
.A(n_10268),
.Y(n_10544)
);

BUFx3_ASAP7_75t_L g10545 ( 
.A(n_10250),
.Y(n_10545)
);

INVx2_ASAP7_75t_L g10546 ( 
.A(n_10174),
.Y(n_10546)
);

INVx1_ASAP7_75t_L g10547 ( 
.A(n_10093),
.Y(n_10547)
);

BUFx6f_ASAP7_75t_L g10548 ( 
.A(n_10261),
.Y(n_10548)
);

AO21x2_ASAP7_75t_L g10549 ( 
.A1(n_10269),
.A2(n_10108),
.B(n_10264),
.Y(n_10549)
);

NAND2xp5_ASAP7_75t_L g10550 ( 
.A(n_10004),
.B(n_1176),
.Y(n_10550)
);

INVx1_ASAP7_75t_L g10551 ( 
.A(n_9991),
.Y(n_10551)
);

AND2x2_ASAP7_75t_L g10552 ( 
.A(n_10042),
.B(n_10114),
.Y(n_10552)
);

INVx2_ASAP7_75t_L g10553 ( 
.A(n_10271),
.Y(n_10553)
);

INVx2_ASAP7_75t_L g10554 ( 
.A(n_10277),
.Y(n_10554)
);

AND2x2_ASAP7_75t_L g10555 ( 
.A(n_10153),
.B(n_10273),
.Y(n_10555)
);

AND2x2_ASAP7_75t_L g10556 ( 
.A(n_10161),
.B(n_546),
.Y(n_10556)
);

INVx2_ASAP7_75t_L g10557 ( 
.A(n_10207),
.Y(n_10557)
);

INVx2_ASAP7_75t_L g10558 ( 
.A(n_10246),
.Y(n_10558)
);

OAI21xp5_ASAP7_75t_SL g10559 ( 
.A1(n_10074),
.A2(n_10254),
.B(n_10141),
.Y(n_10559)
);

INVx1_ASAP7_75t_L g10560 ( 
.A(n_10274),
.Y(n_10560)
);

INVx2_ASAP7_75t_L g10561 ( 
.A(n_10198),
.Y(n_10561)
);

OR2x6_ASAP7_75t_L g10562 ( 
.A(n_10258),
.B(n_1176),
.Y(n_10562)
);

INVxp67_ASAP7_75t_L g10563 ( 
.A(n_10227),
.Y(n_10563)
);

INVx2_ASAP7_75t_L g10564 ( 
.A(n_10124),
.Y(n_10564)
);

INVx2_ASAP7_75t_L g10565 ( 
.A(n_10157),
.Y(n_10565)
);

AND2x2_ASAP7_75t_L g10566 ( 
.A(n_10270),
.B(n_546),
.Y(n_10566)
);

AND2x4_ASAP7_75t_L g10567 ( 
.A(n_10116),
.B(n_547),
.Y(n_10567)
);

INVx1_ASAP7_75t_L g10568 ( 
.A(n_10041),
.Y(n_10568)
);

INVx1_ASAP7_75t_L g10569 ( 
.A(n_10041),
.Y(n_10569)
);

INVx2_ASAP7_75t_SL g10570 ( 
.A(n_10130),
.Y(n_10570)
);

AND2x2_ASAP7_75t_L g10571 ( 
.A(n_10001),
.B(n_547),
.Y(n_10571)
);

INVx1_ASAP7_75t_L g10572 ( 
.A(n_10041),
.Y(n_10572)
);

INVx1_ASAP7_75t_L g10573 ( 
.A(n_10041),
.Y(n_10573)
);

AND2x2_ASAP7_75t_L g10574 ( 
.A(n_10001),
.B(n_547),
.Y(n_10574)
);

INVx1_ASAP7_75t_L g10575 ( 
.A(n_10041),
.Y(n_10575)
);

INVx1_ASAP7_75t_L g10576 ( 
.A(n_10041),
.Y(n_10576)
);

INVx3_ASAP7_75t_L g10577 ( 
.A(n_10151),
.Y(n_10577)
);

INVx2_ASAP7_75t_L g10578 ( 
.A(n_10001),
.Y(n_10578)
);

AO21x2_ASAP7_75t_L g10579 ( 
.A1(n_10015),
.A2(n_548),
.B(n_549),
.Y(n_10579)
);

AND2x4_ASAP7_75t_L g10580 ( 
.A(n_10116),
.B(n_548),
.Y(n_10580)
);

INVx1_ASAP7_75t_L g10581 ( 
.A(n_10041),
.Y(n_10581)
);

INVx1_ASAP7_75t_L g10582 ( 
.A(n_10041),
.Y(n_10582)
);

INVx1_ASAP7_75t_L g10583 ( 
.A(n_10041),
.Y(n_10583)
);

INVx2_ASAP7_75t_L g10584 ( 
.A(n_10001),
.Y(n_10584)
);

AND2x2_ASAP7_75t_L g10585 ( 
.A(n_10001),
.B(n_548),
.Y(n_10585)
);

INVx2_ASAP7_75t_SL g10586 ( 
.A(n_10130),
.Y(n_10586)
);

HB1xp67_ASAP7_75t_L g10587 ( 
.A(n_10031),
.Y(n_10587)
);

INVx2_ASAP7_75t_L g10588 ( 
.A(n_10001),
.Y(n_10588)
);

INVx2_ASAP7_75t_L g10589 ( 
.A(n_10001),
.Y(n_10589)
);

AO21x2_ASAP7_75t_L g10590 ( 
.A1(n_10015),
.A2(n_549),
.B(n_550),
.Y(n_10590)
);

INVx2_ASAP7_75t_L g10591 ( 
.A(n_10001),
.Y(n_10591)
);

BUFx5_ASAP7_75t_L g10592 ( 
.A(n_10151),
.Y(n_10592)
);

OAI21xp5_ASAP7_75t_L g10593 ( 
.A1(n_10559),
.A2(n_549),
.B(n_550),
.Y(n_10593)
);

AND2x2_ASAP7_75t_L g10594 ( 
.A(n_10308),
.B(n_550),
.Y(n_10594)
);

NOR2xp33_ASAP7_75t_L g10595 ( 
.A(n_10444),
.B(n_551),
.Y(n_10595)
);

OAI211xp5_ASAP7_75t_SL g10596 ( 
.A1(n_10551),
.A2(n_553),
.B(n_551),
.C(n_552),
.Y(n_10596)
);

AOI21xp5_ASAP7_75t_L g10597 ( 
.A1(n_10549),
.A2(n_552),
.B(n_553),
.Y(n_10597)
);

AND2x2_ASAP7_75t_L g10598 ( 
.A(n_10439),
.B(n_10433),
.Y(n_10598)
);

NOR2xp33_ASAP7_75t_L g10599 ( 
.A(n_10312),
.B(n_554),
.Y(n_10599)
);

BUFx2_ASAP7_75t_L g10600 ( 
.A(n_10311),
.Y(n_10600)
);

AND2x2_ASAP7_75t_L g10601 ( 
.A(n_10445),
.B(n_554),
.Y(n_10601)
);

O2A1O1Ixp33_ASAP7_75t_SL g10602 ( 
.A1(n_10402),
.A2(n_556),
.B(n_554),
.C(n_555),
.Y(n_10602)
);

A2O1A1Ixp33_ASAP7_75t_L g10603 ( 
.A1(n_10294),
.A2(n_558),
.B(n_556),
.C(n_557),
.Y(n_10603)
);

NOR2xp33_ASAP7_75t_L g10604 ( 
.A(n_10405),
.B(n_556),
.Y(n_10604)
);

AND2x2_ASAP7_75t_L g10605 ( 
.A(n_10473),
.B(n_557),
.Y(n_10605)
);

INVx1_ASAP7_75t_L g10606 ( 
.A(n_10399),
.Y(n_10606)
);

AO32x2_ASAP7_75t_L g10607 ( 
.A1(n_10502),
.A2(n_560),
.A3(n_558),
.B1(n_559),
.B2(n_561),
.Y(n_10607)
);

NOR2xp33_ASAP7_75t_L g10608 ( 
.A(n_10324),
.B(n_558),
.Y(n_10608)
);

BUFx3_ASAP7_75t_L g10609 ( 
.A(n_10313),
.Y(n_10609)
);

AND2x2_ASAP7_75t_L g10610 ( 
.A(n_10373),
.B(n_559),
.Y(n_10610)
);

AND2x2_ASAP7_75t_L g10611 ( 
.A(n_10414),
.B(n_559),
.Y(n_10611)
);

NAND2xp33_ASAP7_75t_L g10612 ( 
.A(n_10592),
.B(n_560),
.Y(n_10612)
);

INVx1_ASAP7_75t_L g10613 ( 
.A(n_10331),
.Y(n_10613)
);

AND2x2_ASAP7_75t_L g10614 ( 
.A(n_10480),
.B(n_560),
.Y(n_10614)
);

OR2x6_ASAP7_75t_L g10615 ( 
.A(n_10311),
.B(n_561),
.Y(n_10615)
);

CKINVDCx5p33_ASAP7_75t_R g10616 ( 
.A(n_10278),
.Y(n_10616)
);

OAI22xp5_ASAP7_75t_L g10617 ( 
.A1(n_10475),
.A2(n_563),
.B1(n_561),
.B2(n_562),
.Y(n_10617)
);

OAI21xp5_ASAP7_75t_L g10618 ( 
.A1(n_10287),
.A2(n_562),
.B(n_563),
.Y(n_10618)
);

AND2x2_ASAP7_75t_L g10619 ( 
.A(n_10495),
.B(n_10505),
.Y(n_10619)
);

OR2x6_ASAP7_75t_L g10620 ( 
.A(n_10304),
.B(n_562),
.Y(n_10620)
);

OR2x2_ASAP7_75t_L g10621 ( 
.A(n_10531),
.B(n_564),
.Y(n_10621)
);

INVx2_ASAP7_75t_L g10622 ( 
.A(n_10421),
.Y(n_10622)
);

NAND2xp5_ASAP7_75t_L g10623 ( 
.A(n_10526),
.B(n_564),
.Y(n_10623)
);

INVx1_ASAP7_75t_L g10624 ( 
.A(n_10279),
.Y(n_10624)
);

OAI21x1_ASAP7_75t_L g10625 ( 
.A1(n_10424),
.A2(n_564),
.B(n_565),
.Y(n_10625)
);

INVx1_ASAP7_75t_L g10626 ( 
.A(n_10290),
.Y(n_10626)
);

AO22x2_ASAP7_75t_L g10627 ( 
.A1(n_10468),
.A2(n_10462),
.B1(n_10450),
.B2(n_10408),
.Y(n_10627)
);

AND2x2_ASAP7_75t_L g10628 ( 
.A(n_10503),
.B(n_566),
.Y(n_10628)
);

OR2x6_ASAP7_75t_L g10629 ( 
.A(n_10314),
.B(n_566),
.Y(n_10629)
);

AND2x2_ASAP7_75t_L g10630 ( 
.A(n_10570),
.B(n_10586),
.Y(n_10630)
);

OA21x2_ASAP7_75t_L g10631 ( 
.A1(n_10471),
.A2(n_10458),
.B(n_10436),
.Y(n_10631)
);

AND2x2_ASAP7_75t_L g10632 ( 
.A(n_10375),
.B(n_566),
.Y(n_10632)
);

HB1xp67_ASAP7_75t_L g10633 ( 
.A(n_10321),
.Y(n_10633)
);

OR2x2_ASAP7_75t_L g10634 ( 
.A(n_10288),
.B(n_10415),
.Y(n_10634)
);

O2A1O1Ixp33_ASAP7_75t_L g10635 ( 
.A1(n_10483),
.A2(n_1179),
.B(n_1177),
.C(n_1178),
.Y(n_10635)
);

OAI21xp5_ASAP7_75t_L g10636 ( 
.A1(n_10406),
.A2(n_1178),
.B(n_1179),
.Y(n_10636)
);

A2O1A1Ixp33_ASAP7_75t_L g10637 ( 
.A1(n_10284),
.A2(n_1182),
.B(n_1180),
.C(n_1181),
.Y(n_10637)
);

OR2x6_ASAP7_75t_L g10638 ( 
.A(n_10516),
.B(n_1180),
.Y(n_10638)
);

INVx2_ASAP7_75t_L g10639 ( 
.A(n_10592),
.Y(n_10639)
);

NAND2xp5_ASAP7_75t_L g10640 ( 
.A(n_10390),
.B(n_1181),
.Y(n_10640)
);

INVx3_ASAP7_75t_L g10641 ( 
.A(n_10281),
.Y(n_10641)
);

BUFx3_ASAP7_75t_L g10642 ( 
.A(n_10303),
.Y(n_10642)
);

O2A1O1Ixp33_ASAP7_75t_SL g10643 ( 
.A1(n_10563),
.A2(n_1184),
.B(n_1182),
.C(n_1183),
.Y(n_10643)
);

OR2x6_ASAP7_75t_L g10644 ( 
.A(n_10516),
.B(n_1185),
.Y(n_10644)
);

AND2x2_ASAP7_75t_L g10645 ( 
.A(n_10382),
.B(n_1186),
.Y(n_10645)
);

O2A1O1Ixp33_ASAP7_75t_SL g10646 ( 
.A1(n_10343),
.A2(n_1188),
.B(n_1186),
.C(n_1187),
.Y(n_10646)
);

INVx1_ASAP7_75t_L g10647 ( 
.A(n_10291),
.Y(n_10647)
);

OA21x2_ASAP7_75t_L g10648 ( 
.A1(n_10432),
.A2(n_1188),
.B(n_1189),
.Y(n_10648)
);

AND2x4_ASAP7_75t_L g10649 ( 
.A(n_10410),
.B(n_1190),
.Y(n_10649)
);

AND2x2_ASAP7_75t_L g10650 ( 
.A(n_10476),
.B(n_1190),
.Y(n_10650)
);

AND2x2_ASAP7_75t_L g10651 ( 
.A(n_10285),
.B(n_1191),
.Y(n_10651)
);

AOI22xp5_ASAP7_75t_L g10652 ( 
.A1(n_10579),
.A2(n_1195),
.B1(n_1191),
.B2(n_1193),
.Y(n_10652)
);

AOI221xp5_ASAP7_75t_L g10653 ( 
.A1(n_10547),
.A2(n_1197),
.B1(n_1193),
.B2(n_1196),
.C(n_1198),
.Y(n_10653)
);

HB1xp67_ASAP7_75t_L g10654 ( 
.A(n_10318),
.Y(n_10654)
);

INVx1_ASAP7_75t_SL g10655 ( 
.A(n_10422),
.Y(n_10655)
);

NAND2xp5_ASAP7_75t_L g10656 ( 
.A(n_10590),
.B(n_1196),
.Y(n_10656)
);

INVx1_ASAP7_75t_L g10657 ( 
.A(n_10295),
.Y(n_10657)
);

AND2x2_ASAP7_75t_L g10658 ( 
.A(n_10435),
.B(n_1197),
.Y(n_10658)
);

AOI221xp5_ASAP7_75t_L g10659 ( 
.A1(n_10453),
.A2(n_10491),
.B1(n_10552),
.B2(n_10393),
.C(n_10532),
.Y(n_10659)
);

INVx2_ASAP7_75t_L g10660 ( 
.A(n_10592),
.Y(n_10660)
);

INVx1_ASAP7_75t_L g10661 ( 
.A(n_10296),
.Y(n_10661)
);

NOR2xp33_ASAP7_75t_L g10662 ( 
.A(n_10283),
.B(n_10293),
.Y(n_10662)
);

INVx2_ASAP7_75t_L g10663 ( 
.A(n_10514),
.Y(n_10663)
);

INVx1_ASAP7_75t_L g10664 ( 
.A(n_10297),
.Y(n_10664)
);

AND2x2_ASAP7_75t_L g10665 ( 
.A(n_10535),
.B(n_1198),
.Y(n_10665)
);

AND2x2_ASAP7_75t_L g10666 ( 
.A(n_10522),
.B(n_1199),
.Y(n_10666)
);

AND2x2_ASAP7_75t_L g10667 ( 
.A(n_10544),
.B(n_1199),
.Y(n_10667)
);

BUFx3_ASAP7_75t_L g10668 ( 
.A(n_10303),
.Y(n_10668)
);

NAND2xp5_ASAP7_75t_L g10669 ( 
.A(n_10451),
.B(n_1200),
.Y(n_10669)
);

AND2x2_ASAP7_75t_L g10670 ( 
.A(n_10280),
.B(n_1200),
.Y(n_10670)
);

AND2x2_ASAP7_75t_L g10671 ( 
.A(n_10282),
.B(n_1201),
.Y(n_10671)
);

OR2x6_ASAP7_75t_L g10672 ( 
.A(n_10380),
.B(n_1202),
.Y(n_10672)
);

INVx2_ASAP7_75t_L g10673 ( 
.A(n_10525),
.Y(n_10673)
);

OAI22xp5_ASAP7_75t_L g10674 ( 
.A1(n_10482),
.A2(n_1204),
.B1(n_1202),
.B2(n_1203),
.Y(n_10674)
);

A2O1A1Ixp33_ASAP7_75t_L g10675 ( 
.A1(n_10550),
.A2(n_1205),
.B(n_1203),
.C(n_1204),
.Y(n_10675)
);

AND2x2_ASAP7_75t_L g10676 ( 
.A(n_10578),
.B(n_1205),
.Y(n_10676)
);

NOR2xp33_ASAP7_75t_L g10677 ( 
.A(n_10577),
.B(n_1206),
.Y(n_10677)
);

INVx2_ASAP7_75t_L g10678 ( 
.A(n_10528),
.Y(n_10678)
);

OR2x2_ASAP7_75t_L g10679 ( 
.A(n_10336),
.B(n_1206),
.Y(n_10679)
);

A2O1A1Ixp33_ASAP7_75t_L g10680 ( 
.A1(n_10507),
.A2(n_1209),
.B(n_1207),
.C(n_1208),
.Y(n_10680)
);

BUFx3_ASAP7_75t_L g10681 ( 
.A(n_10360),
.Y(n_10681)
);

AND2x4_ASAP7_75t_SL g10682 ( 
.A(n_10286),
.B(n_1207),
.Y(n_10682)
);

BUFx6f_ASAP7_75t_L g10683 ( 
.A(n_10360),
.Y(n_10683)
);

NAND2xp5_ASAP7_75t_L g10684 ( 
.A(n_10543),
.B(n_1208),
.Y(n_10684)
);

AND2x4_ASAP7_75t_L g10685 ( 
.A(n_10401),
.B(n_1210),
.Y(n_10685)
);

INVx1_ASAP7_75t_L g10686 ( 
.A(n_10299),
.Y(n_10686)
);

O2A1O1Ixp33_ASAP7_75t_SL g10687 ( 
.A1(n_10561),
.A2(n_1213),
.B(n_1210),
.C(n_1212),
.Y(n_10687)
);

AO32x2_ASAP7_75t_L g10688 ( 
.A1(n_10524),
.A2(n_1214),
.A3(n_1212),
.B1(n_1213),
.B2(n_1215),
.Y(n_10688)
);

NAND2xp5_ASAP7_75t_L g10689 ( 
.A(n_10553),
.B(n_1215),
.Y(n_10689)
);

OA21x2_ASAP7_75t_L g10690 ( 
.A1(n_10300),
.A2(n_10588),
.B(n_10584),
.Y(n_10690)
);

AND2x2_ASAP7_75t_L g10691 ( 
.A(n_10589),
.B(n_1216),
.Y(n_10691)
);

NAND2xp5_ASAP7_75t_L g10692 ( 
.A(n_10554),
.B(n_1216),
.Y(n_10692)
);

INVx3_ASAP7_75t_L g10693 ( 
.A(n_10286),
.Y(n_10693)
);

AND2x4_ASAP7_75t_L g10694 ( 
.A(n_10411),
.B(n_1218),
.Y(n_10694)
);

AND2x2_ASAP7_75t_L g10695 ( 
.A(n_10591),
.B(n_1218),
.Y(n_10695)
);

INVxp67_ASAP7_75t_L g10696 ( 
.A(n_10469),
.Y(n_10696)
);

HB1xp67_ASAP7_75t_L g10697 ( 
.A(n_10587),
.Y(n_10697)
);

AO21x1_ASAP7_75t_L g10698 ( 
.A1(n_10449),
.A2(n_1219),
.B(n_1220),
.Y(n_10698)
);

OAI21xp5_ASAP7_75t_L g10699 ( 
.A1(n_10538),
.A2(n_1219),
.B(n_1220),
.Y(n_10699)
);

NAND4xp25_ASAP7_75t_L g10700 ( 
.A(n_10529),
.B(n_1223),
.C(n_1221),
.D(n_1222),
.Y(n_10700)
);

AND2x4_ASAP7_75t_L g10701 ( 
.A(n_10492),
.B(n_1221),
.Y(n_10701)
);

NAND2xp5_ASAP7_75t_L g10702 ( 
.A(n_10541),
.B(n_1224),
.Y(n_10702)
);

OAI21xp5_ASAP7_75t_L g10703 ( 
.A1(n_10562),
.A2(n_1224),
.B(n_1225),
.Y(n_10703)
);

INVx1_ASAP7_75t_L g10704 ( 
.A(n_10307),
.Y(n_10704)
);

INVx1_ASAP7_75t_L g10705 ( 
.A(n_10316),
.Y(n_10705)
);

INVx2_ASAP7_75t_L g10706 ( 
.A(n_10537),
.Y(n_10706)
);

AND2x2_ASAP7_75t_L g10707 ( 
.A(n_10417),
.B(n_1226),
.Y(n_10707)
);

HB1xp67_ASAP7_75t_L g10708 ( 
.A(n_10350),
.Y(n_10708)
);

AOI22xp5_ASAP7_75t_L g10709 ( 
.A1(n_10413),
.A2(n_1229),
.B1(n_1227),
.B2(n_1228),
.Y(n_10709)
);

INVx1_ASAP7_75t_L g10710 ( 
.A(n_10319),
.Y(n_10710)
);

OR2x2_ASAP7_75t_L g10711 ( 
.A(n_10512),
.B(n_1227),
.Y(n_10711)
);

OR2x2_ASAP7_75t_L g10712 ( 
.A(n_10542),
.B(n_1229),
.Y(n_10712)
);

AND2x2_ASAP7_75t_L g10713 ( 
.A(n_10301),
.B(n_1230),
.Y(n_10713)
);

AND2x2_ASAP7_75t_L g10714 ( 
.A(n_10447),
.B(n_1230),
.Y(n_10714)
);

OAI21x1_ASAP7_75t_L g10715 ( 
.A1(n_10305),
.A2(n_10425),
.B(n_10418),
.Y(n_10715)
);

INVx1_ASAP7_75t_L g10716 ( 
.A(n_10323),
.Y(n_10716)
);

INVx3_ASAP7_75t_L g10717 ( 
.A(n_10423),
.Y(n_10717)
);

AND2x2_ASAP7_75t_L g10718 ( 
.A(n_10485),
.B(n_1231),
.Y(n_10718)
);

AND2x2_ASAP7_75t_L g10719 ( 
.A(n_10510),
.B(n_1231),
.Y(n_10719)
);

NOR2x1_ASAP7_75t_SL g10720 ( 
.A(n_10412),
.B(n_10420),
.Y(n_10720)
);

AO21x1_ASAP7_75t_L g10721 ( 
.A1(n_10517),
.A2(n_1233),
.B(n_1234),
.Y(n_10721)
);

INVx2_ASAP7_75t_SL g10722 ( 
.A(n_10467),
.Y(n_10722)
);

O2A1O1Ixp33_ASAP7_75t_SL g10723 ( 
.A1(n_10534),
.A2(n_1236),
.B(n_1234),
.C(n_1235),
.Y(n_10723)
);

AND4x1_ASAP7_75t_L g10724 ( 
.A(n_10372),
.B(n_10397),
.C(n_10540),
.D(n_10556),
.Y(n_10724)
);

AND2x2_ASAP7_75t_L g10725 ( 
.A(n_10515),
.B(n_10459),
.Y(n_10725)
);

OR2x2_ASAP7_75t_L g10726 ( 
.A(n_10437),
.B(n_1236),
.Y(n_10726)
);

A2O1A1Ixp33_ASAP7_75t_L g10727 ( 
.A1(n_10536),
.A2(n_1239),
.B(n_1237),
.C(n_1238),
.Y(n_10727)
);

AO32x2_ASAP7_75t_L g10728 ( 
.A1(n_10504),
.A2(n_1239),
.A3(n_1237),
.B1(n_1238),
.B2(n_1240),
.Y(n_10728)
);

INVx3_ASAP7_75t_L g10729 ( 
.A(n_10428),
.Y(n_10729)
);

HB1xp67_ASAP7_75t_L g10730 ( 
.A(n_10474),
.Y(n_10730)
);

OR2x6_ASAP7_75t_L g10731 ( 
.A(n_10420),
.B(n_1240),
.Y(n_10731)
);

INVx1_ASAP7_75t_L g10732 ( 
.A(n_10325),
.Y(n_10732)
);

OR2x2_ASAP7_75t_L g10733 ( 
.A(n_10497),
.B(n_10539),
.Y(n_10733)
);

OR2x2_ASAP7_75t_L g10734 ( 
.A(n_10292),
.B(n_1241),
.Y(n_10734)
);

AND2x2_ASAP7_75t_L g10735 ( 
.A(n_10452),
.B(n_1242),
.Y(n_10735)
);

OAI21xp5_ASAP7_75t_L g10736 ( 
.A1(n_10562),
.A2(n_1242),
.B(n_1243),
.Y(n_10736)
);

AOI221xp5_ASAP7_75t_L g10737 ( 
.A1(n_10560),
.A2(n_10558),
.B1(n_10557),
.B2(n_10548),
.C(n_10564),
.Y(n_10737)
);

AOI221xp5_ASAP7_75t_L g10738 ( 
.A1(n_10548),
.A2(n_1247),
.B1(n_1243),
.B2(n_1246),
.C(n_1248),
.Y(n_10738)
);

HB1xp67_ASAP7_75t_L g10739 ( 
.A(n_10356),
.Y(n_10739)
);

AND2x4_ASAP7_75t_L g10740 ( 
.A(n_10496),
.B(n_1246),
.Y(n_10740)
);

AND2x2_ASAP7_75t_L g10741 ( 
.A(n_10454),
.B(n_1248),
.Y(n_10741)
);

OR2x2_ASAP7_75t_L g10742 ( 
.A(n_10345),
.B(n_1249),
.Y(n_10742)
);

AOI22xp5_ASAP7_75t_L g10743 ( 
.A1(n_10302),
.A2(n_1251),
.B1(n_1249),
.B2(n_1250),
.Y(n_10743)
);

OR2x2_ASAP7_75t_L g10744 ( 
.A(n_10442),
.B(n_1251),
.Y(n_10744)
);

AOI221xp5_ASAP7_75t_L g10745 ( 
.A1(n_10555),
.A2(n_10565),
.B1(n_10309),
.B2(n_10463),
.C(n_10342),
.Y(n_10745)
);

AND2x2_ASAP7_75t_L g10746 ( 
.A(n_10456),
.B(n_1252),
.Y(n_10746)
);

INVx1_ASAP7_75t_L g10747 ( 
.A(n_10329),
.Y(n_10747)
);

AND2x2_ASAP7_75t_L g10748 ( 
.A(n_10460),
.B(n_1252),
.Y(n_10748)
);

INVx1_ASAP7_75t_L g10749 ( 
.A(n_10330),
.Y(n_10749)
);

HB1xp67_ASAP7_75t_L g10750 ( 
.A(n_10443),
.Y(n_10750)
);

OR2x2_ASAP7_75t_L g10751 ( 
.A(n_10404),
.B(n_1253),
.Y(n_10751)
);

NAND2xp33_ASAP7_75t_L g10752 ( 
.A(n_10428),
.B(n_10335),
.Y(n_10752)
);

HB1xp67_ASAP7_75t_L g10753 ( 
.A(n_10472),
.Y(n_10753)
);

NOR2xp33_ASAP7_75t_L g10754 ( 
.A(n_10392),
.B(n_1254),
.Y(n_10754)
);

A2O1A1Ixp33_ASAP7_75t_L g10755 ( 
.A1(n_10317),
.A2(n_1257),
.B(n_1255),
.C(n_1256),
.Y(n_10755)
);

OR2x6_ASAP7_75t_L g10756 ( 
.A(n_10488),
.B(n_1255),
.Y(n_10756)
);

OAI22xp5_ASAP7_75t_L g10757 ( 
.A1(n_10493),
.A2(n_1258),
.B1(n_1256),
.B2(n_1257),
.Y(n_10757)
);

AOI22xp5_ASAP7_75t_L g10758 ( 
.A1(n_10494),
.A2(n_1260),
.B1(n_1258),
.B2(n_1259),
.Y(n_10758)
);

AND2x4_ASAP7_75t_L g10759 ( 
.A(n_10381),
.B(n_1259),
.Y(n_10759)
);

AND2x2_ASAP7_75t_L g10760 ( 
.A(n_10464),
.B(n_10477),
.Y(n_10760)
);

AND2x2_ASAP7_75t_L g10761 ( 
.A(n_10479),
.B(n_10489),
.Y(n_10761)
);

AOI22xp5_ASAP7_75t_L g10762 ( 
.A1(n_10546),
.A2(n_1262),
.B1(n_1260),
.B2(n_1261),
.Y(n_10762)
);

AND2x2_ASAP7_75t_L g10763 ( 
.A(n_10506),
.B(n_1261),
.Y(n_10763)
);

AND2x6_ASAP7_75t_L g10764 ( 
.A(n_10355),
.B(n_1262),
.Y(n_10764)
);

AND2x2_ASAP7_75t_L g10765 ( 
.A(n_10499),
.B(n_1263),
.Y(n_10765)
);

A2O1A1Ixp33_ASAP7_75t_L g10766 ( 
.A1(n_10566),
.A2(n_10327),
.B(n_10326),
.C(n_10513),
.Y(n_10766)
);

AO32x2_ASAP7_75t_L g10767 ( 
.A1(n_10289),
.A2(n_1266),
.A3(n_1263),
.B1(n_1264),
.B2(n_1267),
.Y(n_10767)
);

AND2x2_ASAP7_75t_L g10768 ( 
.A(n_10426),
.B(n_1266),
.Y(n_10768)
);

AND2x2_ASAP7_75t_L g10769 ( 
.A(n_10484),
.B(n_1267),
.Y(n_10769)
);

NAND2xp33_ASAP7_75t_SL g10770 ( 
.A(n_10519),
.B(n_1268),
.Y(n_10770)
);

OAI21x1_ASAP7_75t_L g10771 ( 
.A1(n_10440),
.A2(n_1268),
.B(n_1269),
.Y(n_10771)
);

OAI21x1_ASAP7_75t_SL g10772 ( 
.A1(n_10511),
.A2(n_1270),
.B(n_1271),
.Y(n_10772)
);

AOI211xp5_ASAP7_75t_L g10773 ( 
.A1(n_10441),
.A2(n_1272),
.B(n_1270),
.C(n_1271),
.Y(n_10773)
);

O2A1O1Ixp5_ASAP7_75t_L g10774 ( 
.A1(n_10363),
.A2(n_1274),
.B(n_1272),
.C(n_1273),
.Y(n_10774)
);

AND2x2_ASAP7_75t_L g10775 ( 
.A(n_10518),
.B(n_1275),
.Y(n_10775)
);

AND2x2_ASAP7_75t_L g10776 ( 
.A(n_10501),
.B(n_1275),
.Y(n_10776)
);

HB1xp67_ASAP7_75t_L g10777 ( 
.A(n_10466),
.Y(n_10777)
);

OAI21xp5_ASAP7_75t_L g10778 ( 
.A1(n_10446),
.A2(n_1276),
.B(n_1277),
.Y(n_10778)
);

AND2x2_ASAP7_75t_L g10779 ( 
.A(n_10508),
.B(n_1276),
.Y(n_10779)
);

A2O1A1Ixp33_ASAP7_75t_L g10780 ( 
.A1(n_10438),
.A2(n_1279),
.B(n_1277),
.C(n_1278),
.Y(n_10780)
);

CKINVDCx6p67_ASAP7_75t_R g10781 ( 
.A(n_10533),
.Y(n_10781)
);

BUFx2_ASAP7_75t_L g10782 ( 
.A(n_10530),
.Y(n_10782)
);

OR2x6_ASAP7_75t_L g10783 ( 
.A(n_10567),
.B(n_1278),
.Y(n_10783)
);

OAI22xp5_ASAP7_75t_L g10784 ( 
.A1(n_10545),
.A2(n_1282),
.B1(n_1279),
.B2(n_1280),
.Y(n_10784)
);

OA21x2_ASAP7_75t_L g10785 ( 
.A1(n_10487),
.A2(n_1280),
.B(n_1282),
.Y(n_10785)
);

NAND2xp5_ASAP7_75t_L g10786 ( 
.A(n_10509),
.B(n_1283),
.Y(n_10786)
);

AND2x2_ASAP7_75t_L g10787 ( 
.A(n_10486),
.B(n_1283),
.Y(n_10787)
);

INVx3_ASAP7_75t_L g10788 ( 
.A(n_10457),
.Y(n_10788)
);

OAI22xp5_ASAP7_75t_L g10789 ( 
.A1(n_10465),
.A2(n_10416),
.B1(n_10490),
.B2(n_10391),
.Y(n_10789)
);

AND2x4_ASAP7_75t_SL g10790 ( 
.A(n_10403),
.B(n_1284),
.Y(n_10790)
);

A2O1A1Ixp33_ASAP7_75t_L g10791 ( 
.A1(n_10448),
.A2(n_1287),
.B(n_1285),
.C(n_1286),
.Y(n_10791)
);

AND2x4_ASAP7_75t_L g10792 ( 
.A(n_10498),
.B(n_1286),
.Y(n_10792)
);

AND2x2_ASAP7_75t_L g10793 ( 
.A(n_10427),
.B(n_1287),
.Y(n_10793)
);

AOI21xp5_ASAP7_75t_L g10794 ( 
.A1(n_10520),
.A2(n_1288),
.B(n_1289),
.Y(n_10794)
);

OR2x2_ASAP7_75t_L g10795 ( 
.A(n_10385),
.B(n_1288),
.Y(n_10795)
);

AND2x2_ASAP7_75t_L g10796 ( 
.A(n_10461),
.B(n_1290),
.Y(n_10796)
);

AND2x2_ASAP7_75t_L g10797 ( 
.A(n_10348),
.B(n_1290),
.Y(n_10797)
);

AO21x2_ASAP7_75t_L g10798 ( 
.A1(n_10571),
.A2(n_1291),
.B(n_1292),
.Y(n_10798)
);

NAND2xp5_ASAP7_75t_L g10799 ( 
.A(n_10470),
.B(n_1291),
.Y(n_10799)
);

OA21x2_ASAP7_75t_L g10800 ( 
.A1(n_10389),
.A2(n_1292),
.B(n_1293),
.Y(n_10800)
);

NAND2x1_ASAP7_75t_L g10801 ( 
.A(n_10298),
.B(n_1294),
.Y(n_10801)
);

OR2x2_ASAP7_75t_L g10802 ( 
.A(n_10431),
.B(n_1295),
.Y(n_10802)
);

NOR2xp33_ASAP7_75t_L g10803 ( 
.A(n_10455),
.B(n_1295),
.Y(n_10803)
);

AO32x2_ASAP7_75t_L g10804 ( 
.A1(n_10394),
.A2(n_1298),
.A3(n_1296),
.B1(n_1297),
.B2(n_1299),
.Y(n_10804)
);

OA21x2_ASAP7_75t_L g10805 ( 
.A1(n_10387),
.A2(n_1298),
.B(n_1299),
.Y(n_10805)
);

OR2x2_ASAP7_75t_L g10806 ( 
.A(n_10365),
.B(n_1300),
.Y(n_10806)
);

INVx2_ASAP7_75t_L g10807 ( 
.A(n_10388),
.Y(n_10807)
);

CKINVDCx16_ASAP7_75t_R g10808 ( 
.A(n_10574),
.Y(n_10808)
);

OAI21xp5_ASAP7_75t_L g10809 ( 
.A1(n_10409),
.A2(n_1300),
.B(n_1301),
.Y(n_10809)
);

NOR2x1_ASAP7_75t_SL g10810 ( 
.A(n_10353),
.B(n_1301),
.Y(n_10810)
);

AND2x2_ASAP7_75t_L g10811 ( 
.A(n_10430),
.B(n_1302),
.Y(n_10811)
);

AOI22xp5_ASAP7_75t_L g10812 ( 
.A1(n_10322),
.A2(n_1305),
.B1(n_1303),
.B2(n_1304),
.Y(n_10812)
);

NOR2x1_ASAP7_75t_SL g10813 ( 
.A(n_10328),
.B(n_1303),
.Y(n_10813)
);

INVx2_ASAP7_75t_L g10814 ( 
.A(n_10306),
.Y(n_10814)
);

INVx1_ASAP7_75t_L g10815 ( 
.A(n_10332),
.Y(n_10815)
);

NOR2xp33_ASAP7_75t_L g10816 ( 
.A(n_10500),
.B(n_1306),
.Y(n_10816)
);

AND2x4_ASAP7_75t_L g10817 ( 
.A(n_10580),
.B(n_1307),
.Y(n_10817)
);

AND2x2_ASAP7_75t_L g10818 ( 
.A(n_10310),
.B(n_1308),
.Y(n_10818)
);

OR2x2_ASAP7_75t_L g10819 ( 
.A(n_10367),
.B(n_1309),
.Y(n_10819)
);

AND2x2_ASAP7_75t_L g10820 ( 
.A(n_10315),
.B(n_1309),
.Y(n_10820)
);

OR2x2_ASAP7_75t_L g10821 ( 
.A(n_10369),
.B(n_10320),
.Y(n_10821)
);

OR2x6_ASAP7_75t_L g10822 ( 
.A(n_10585),
.B(n_1310),
.Y(n_10822)
);

OAI21xp5_ASAP7_75t_L g10823 ( 
.A1(n_10364),
.A2(n_1311),
.B(n_1312),
.Y(n_10823)
);

OA21x2_ASAP7_75t_L g10824 ( 
.A1(n_10366),
.A2(n_1311),
.B(n_1312),
.Y(n_10824)
);

AND2x4_ASAP7_75t_SL g10825 ( 
.A(n_10527),
.B(n_1313),
.Y(n_10825)
);

INVx2_ASAP7_75t_L g10826 ( 
.A(n_10334),
.Y(n_10826)
);

OR2x2_ASAP7_75t_L g10827 ( 
.A(n_10337),
.B(n_1313),
.Y(n_10827)
);

OR2x2_ASAP7_75t_L g10828 ( 
.A(n_10341),
.B(n_1314),
.Y(n_10828)
);

HB1xp67_ASAP7_75t_L g10829 ( 
.A(n_10359),
.Y(n_10829)
);

OR2x2_ASAP7_75t_L g10830 ( 
.A(n_10357),
.B(n_1314),
.Y(n_10830)
);

NOR2x1_ASAP7_75t_R g10831 ( 
.A(n_10396),
.B(n_1315),
.Y(n_10831)
);

INVx1_ASAP7_75t_L g10832 ( 
.A(n_10333),
.Y(n_10832)
);

NAND2xp5_ASAP7_75t_L g10833 ( 
.A(n_10347),
.B(n_1315),
.Y(n_10833)
);

BUFx2_ASAP7_75t_L g10834 ( 
.A(n_10434),
.Y(n_10834)
);

OAI21xp5_ASAP7_75t_L g10835 ( 
.A1(n_10344),
.A2(n_1316),
.B(n_1317),
.Y(n_10835)
);

OA21x2_ASAP7_75t_L g10836 ( 
.A1(n_10361),
.A2(n_1317),
.B(n_1318),
.Y(n_10836)
);

AND2x4_ASAP7_75t_L g10837 ( 
.A(n_10419),
.B(n_1318),
.Y(n_10837)
);

INVx1_ASAP7_75t_L g10838 ( 
.A(n_10338),
.Y(n_10838)
);

NAND2xp5_ASAP7_75t_L g10839 ( 
.A(n_10429),
.B(n_1319),
.Y(n_10839)
);

AND2x2_ASAP7_75t_L g10840 ( 
.A(n_10358),
.B(n_1319),
.Y(n_10840)
);

AOI31xp33_ASAP7_75t_SL g10841 ( 
.A1(n_10379),
.A2(n_1322),
.A3(n_1320),
.B(n_1321),
.Y(n_10841)
);

INVx1_ASAP7_75t_L g10842 ( 
.A(n_10339),
.Y(n_10842)
);

AND2x6_ASAP7_75t_L g10843 ( 
.A(n_10351),
.B(n_1321),
.Y(n_10843)
);

OAI22xp5_ASAP7_75t_L g10844 ( 
.A1(n_10398),
.A2(n_1326),
.B1(n_1323),
.B2(n_1325),
.Y(n_10844)
);

O2A1O1Ixp33_ASAP7_75t_SL g10845 ( 
.A1(n_10400),
.A2(n_10346),
.B(n_10349),
.C(n_10340),
.Y(n_10845)
);

OR2x6_ASAP7_75t_L g10846 ( 
.A(n_10386),
.B(n_1323),
.Y(n_10846)
);

INVx3_ASAP7_75t_L g10847 ( 
.A(n_10377),
.Y(n_10847)
);

AND2x2_ASAP7_75t_L g10848 ( 
.A(n_10383),
.B(n_10362),
.Y(n_10848)
);

O2A1O1Ixp33_ASAP7_75t_L g10849 ( 
.A1(n_10374),
.A2(n_1328),
.B(n_1326),
.C(n_1327),
.Y(n_10849)
);

BUFx5_ASAP7_75t_L g10850 ( 
.A(n_10378),
.Y(n_10850)
);

OAI21xp5_ASAP7_75t_L g10851 ( 
.A1(n_10368),
.A2(n_1327),
.B(n_1328),
.Y(n_10851)
);

AO21x2_ASAP7_75t_L g10852 ( 
.A1(n_10478),
.A2(n_1329),
.B(n_1330),
.Y(n_10852)
);

NOR2xp33_ASAP7_75t_L g10853 ( 
.A(n_10523),
.B(n_1329),
.Y(n_10853)
);

HB1xp67_ASAP7_75t_L g10854 ( 
.A(n_10395),
.Y(n_10854)
);

NAND2xp5_ASAP7_75t_L g10855 ( 
.A(n_10481),
.B(n_1331),
.Y(n_10855)
);

AND2x2_ASAP7_75t_L g10856 ( 
.A(n_10407),
.B(n_1332),
.Y(n_10856)
);

AND2x2_ASAP7_75t_L g10857 ( 
.A(n_10521),
.B(n_1332),
.Y(n_10857)
);

AOI22xp33_ASAP7_75t_L g10858 ( 
.A1(n_10370),
.A2(n_1336),
.B1(n_1334),
.B2(n_1335),
.Y(n_10858)
);

AOI22xp33_ASAP7_75t_SL g10859 ( 
.A1(n_10352),
.A2(n_1337),
.B1(n_1335),
.B2(n_1336),
.Y(n_10859)
);

AOI21xp5_ASAP7_75t_L g10860 ( 
.A1(n_10354),
.A2(n_1337),
.B(n_1338),
.Y(n_10860)
);

OA21x2_ASAP7_75t_L g10861 ( 
.A1(n_10371),
.A2(n_1338),
.B(n_1339),
.Y(n_10861)
);

HB1xp67_ASAP7_75t_L g10862 ( 
.A(n_10568),
.Y(n_10862)
);

AND2x2_ASAP7_75t_L g10863 ( 
.A(n_10569),
.B(n_1339),
.Y(n_10863)
);

AND2x4_ASAP7_75t_L g10864 ( 
.A(n_10572),
.B(n_1340),
.Y(n_10864)
);

OAI21xp5_ASAP7_75t_L g10865 ( 
.A1(n_10376),
.A2(n_1341),
.B(n_1342),
.Y(n_10865)
);

INVx1_ASAP7_75t_L g10866 ( 
.A(n_10573),
.Y(n_10866)
);

AND2x2_ASAP7_75t_L g10867 ( 
.A(n_10575),
.B(n_1342),
.Y(n_10867)
);

AO32x2_ASAP7_75t_L g10868 ( 
.A1(n_10576),
.A2(n_1345),
.A3(n_1343),
.B1(n_1344),
.B2(n_1346),
.Y(n_10868)
);

OR2x2_ASAP7_75t_L g10869 ( 
.A(n_10384),
.B(n_1343),
.Y(n_10869)
);

NAND2xp5_ASAP7_75t_L g10870 ( 
.A(n_10581),
.B(n_1344),
.Y(n_10870)
);

INVx1_ASAP7_75t_L g10871 ( 
.A(n_10582),
.Y(n_10871)
);

AOI22xp5_ASAP7_75t_L g10872 ( 
.A1(n_10583),
.A2(n_1347),
.B1(n_1345),
.B2(n_1346),
.Y(n_10872)
);

AOI21xp5_ASAP7_75t_L g10873 ( 
.A1(n_10549),
.A2(n_1348),
.B(n_1349),
.Y(n_10873)
);

A2O1A1Ixp33_ASAP7_75t_L g10874 ( 
.A1(n_10559),
.A2(n_1352),
.B(n_1350),
.C(n_1351),
.Y(n_10874)
);

A2O1A1Ixp33_ASAP7_75t_L g10875 ( 
.A1(n_10559),
.A2(n_1352),
.B(n_1350),
.C(n_1351),
.Y(n_10875)
);

AND2x4_ASAP7_75t_L g10876 ( 
.A(n_10304),
.B(n_1353),
.Y(n_10876)
);

AND2x2_ASAP7_75t_L g10877 ( 
.A(n_10308),
.B(n_1354),
.Y(n_10877)
);

AND2x2_ASAP7_75t_L g10878 ( 
.A(n_10308),
.B(n_1354),
.Y(n_10878)
);

O2A1O1Ixp33_ASAP7_75t_SL g10879 ( 
.A1(n_10402),
.A2(n_1358),
.B(n_1356),
.C(n_1357),
.Y(n_10879)
);

AND2x2_ASAP7_75t_L g10880 ( 
.A(n_10308),
.B(n_1356),
.Y(n_10880)
);

NOR2xp33_ASAP7_75t_L g10881 ( 
.A(n_10444),
.B(n_1357),
.Y(n_10881)
);

INVx1_ASAP7_75t_L g10882 ( 
.A(n_10399),
.Y(n_10882)
);

A2O1A1Ixp33_ASAP7_75t_L g10883 ( 
.A1(n_10559),
.A2(n_1360),
.B(n_1358),
.C(n_1359),
.Y(n_10883)
);

OAI22xp5_ASAP7_75t_L g10884 ( 
.A1(n_10294),
.A2(n_1362),
.B1(n_1360),
.B2(n_1361),
.Y(n_10884)
);

INVxp67_ASAP7_75t_SL g10885 ( 
.A(n_10308),
.Y(n_10885)
);

AOI21xp5_ASAP7_75t_L g10886 ( 
.A1(n_10549),
.A2(n_1361),
.B(n_1363),
.Y(n_10886)
);

AND2x2_ASAP7_75t_L g10887 ( 
.A(n_10308),
.B(n_1363),
.Y(n_10887)
);

INVx1_ASAP7_75t_L g10888 ( 
.A(n_10399),
.Y(n_10888)
);

NOR2xp33_ASAP7_75t_L g10889 ( 
.A(n_10444),
.B(n_1365),
.Y(n_10889)
);

AND2x4_ASAP7_75t_L g10890 ( 
.A(n_10304),
.B(n_1366),
.Y(n_10890)
);

INVx1_ASAP7_75t_L g10891 ( 
.A(n_10399),
.Y(n_10891)
);

O2A1O1Ixp33_ASAP7_75t_L g10892 ( 
.A1(n_10559),
.A2(n_1368),
.B(n_1366),
.C(n_1367),
.Y(n_10892)
);

AO32x2_ASAP7_75t_L g10893 ( 
.A1(n_10473),
.A2(n_1370),
.A3(n_1368),
.B1(n_1369),
.B2(n_1371),
.Y(n_10893)
);

O2A1O1Ixp33_ASAP7_75t_SL g10894 ( 
.A1(n_10402),
.A2(n_1371),
.B(n_1369),
.C(n_1370),
.Y(n_10894)
);

INVx1_ASAP7_75t_L g10895 ( 
.A(n_10399),
.Y(n_10895)
);

AND2x2_ASAP7_75t_L g10896 ( 
.A(n_10308),
.B(n_1372),
.Y(n_10896)
);

A2O1A1Ixp33_ASAP7_75t_L g10897 ( 
.A1(n_10559),
.A2(n_1374),
.B(n_1372),
.C(n_1373),
.Y(n_10897)
);

AND2x4_ASAP7_75t_L g10898 ( 
.A(n_10304),
.B(n_1373),
.Y(n_10898)
);

AND2x4_ASAP7_75t_L g10899 ( 
.A(n_10304),
.B(n_1374),
.Y(n_10899)
);

OAI22xp5_ASAP7_75t_L g10900 ( 
.A1(n_10294),
.A2(n_1377),
.B1(n_1375),
.B2(n_1376),
.Y(n_10900)
);

NOR2xp33_ASAP7_75t_L g10901 ( 
.A(n_10444),
.B(n_1376),
.Y(n_10901)
);

CKINVDCx5p33_ASAP7_75t_R g10902 ( 
.A(n_10312),
.Y(n_10902)
);

AO22x2_ASAP7_75t_L g10903 ( 
.A1(n_10468),
.A2(n_1379),
.B1(n_1377),
.B2(n_1378),
.Y(n_10903)
);

AOI21xp5_ASAP7_75t_L g10904 ( 
.A1(n_10549),
.A2(n_1378),
.B(n_1379),
.Y(n_10904)
);

AND2x2_ASAP7_75t_L g10905 ( 
.A(n_10308),
.B(n_1380),
.Y(n_10905)
);

INVx3_ASAP7_75t_L g10906 ( 
.A(n_10281),
.Y(n_10906)
);

A2O1A1Ixp33_ASAP7_75t_L g10907 ( 
.A1(n_10559),
.A2(n_1383),
.B(n_1381),
.C(n_1382),
.Y(n_10907)
);

AOI211xp5_ASAP7_75t_L g10908 ( 
.A1(n_10559),
.A2(n_1386),
.B(n_1381),
.C(n_1382),
.Y(n_10908)
);

OAI21xp5_ASAP7_75t_L g10909 ( 
.A1(n_10559),
.A2(n_1387),
.B(n_1388),
.Y(n_10909)
);

INVx3_ASAP7_75t_L g10910 ( 
.A(n_10281),
.Y(n_10910)
);

HB1xp67_ASAP7_75t_L g10911 ( 
.A(n_10399),
.Y(n_10911)
);

NAND2xp5_ASAP7_75t_L g10912 ( 
.A(n_10526),
.B(n_1389),
.Y(n_10912)
);

INVx1_ASAP7_75t_L g10913 ( 
.A(n_10399),
.Y(n_10913)
);

INVx1_ASAP7_75t_L g10914 ( 
.A(n_10399),
.Y(n_10914)
);

AND2x2_ASAP7_75t_L g10915 ( 
.A(n_10308),
.B(n_1390),
.Y(n_10915)
);

NAND2xp5_ASAP7_75t_L g10916 ( 
.A(n_10526),
.B(n_1390),
.Y(n_10916)
);

OAI21x1_ASAP7_75t_L g10917 ( 
.A1(n_10424),
.A2(n_1391),
.B(n_1392),
.Y(n_10917)
);

INVx1_ASAP7_75t_L g10918 ( 
.A(n_10399),
.Y(n_10918)
);

BUFx2_ASAP7_75t_L g10919 ( 
.A(n_10308),
.Y(n_10919)
);

AO21x2_ASAP7_75t_L g10920 ( 
.A1(n_10449),
.A2(n_1391),
.B(n_1392),
.Y(n_10920)
);

AND2x2_ASAP7_75t_L g10921 ( 
.A(n_10308),
.B(n_1393),
.Y(n_10921)
);

AND2x2_ASAP7_75t_L g10922 ( 
.A(n_10308),
.B(n_1393),
.Y(n_10922)
);

INVx1_ASAP7_75t_SL g10923 ( 
.A(n_10324),
.Y(n_10923)
);

INVxp67_ASAP7_75t_L g10924 ( 
.A(n_10469),
.Y(n_10924)
);

OAI21x1_ASAP7_75t_SL g10925 ( 
.A1(n_10511),
.A2(n_1394),
.B(n_1395),
.Y(n_10925)
);

INVx2_ASAP7_75t_L g10926 ( 
.A(n_10782),
.Y(n_10926)
);

NAND2xp5_ASAP7_75t_L g10927 ( 
.A(n_10808),
.B(n_1394),
.Y(n_10927)
);

OAI21xp5_ASAP7_75t_L g10928 ( 
.A1(n_10597),
.A2(n_1396),
.B(n_1397),
.Y(n_10928)
);

AND2x2_ASAP7_75t_L g10929 ( 
.A(n_10630),
.B(n_10600),
.Y(n_10929)
);

INVx2_ASAP7_75t_L g10930 ( 
.A(n_10642),
.Y(n_10930)
);

INVx1_ASAP7_75t_L g10931 ( 
.A(n_10911),
.Y(n_10931)
);

AND2x2_ASAP7_75t_L g10932 ( 
.A(n_10919),
.B(n_10619),
.Y(n_10932)
);

NAND2xp5_ASAP7_75t_L g10933 ( 
.A(n_10885),
.B(n_1398),
.Y(n_10933)
);

INVx1_ASAP7_75t_L g10934 ( 
.A(n_10633),
.Y(n_10934)
);

AOI22xp33_ASAP7_75t_L g10935 ( 
.A1(n_10659),
.A2(n_10909),
.B1(n_10593),
.B2(n_10886),
.Y(n_10935)
);

AND2x2_ASAP7_75t_L g10936 ( 
.A(n_10781),
.B(n_1398),
.Y(n_10936)
);

NAND2xp5_ASAP7_75t_L g10937 ( 
.A(n_10655),
.B(n_1399),
.Y(n_10937)
);

NAND2xp5_ASAP7_75t_L g10938 ( 
.A(n_10743),
.B(n_1400),
.Y(n_10938)
);

INVx2_ASAP7_75t_L g10939 ( 
.A(n_10668),
.Y(n_10939)
);

INVx2_ASAP7_75t_L g10940 ( 
.A(n_10681),
.Y(n_10940)
);

INVx4_ASAP7_75t_L g10941 ( 
.A(n_10609),
.Y(n_10941)
);

HB1xp67_ASAP7_75t_L g10942 ( 
.A(n_10834),
.Y(n_10942)
);

AND2x2_ASAP7_75t_L g10943 ( 
.A(n_10598),
.B(n_1400),
.Y(n_10943)
);

INVx3_ASAP7_75t_L g10944 ( 
.A(n_10683),
.Y(n_10944)
);

INVx1_ASAP7_75t_L g10945 ( 
.A(n_10654),
.Y(n_10945)
);

BUFx2_ASAP7_75t_L g10946 ( 
.A(n_10696),
.Y(n_10946)
);

INVx1_ASAP7_75t_L g10947 ( 
.A(n_10697),
.Y(n_10947)
);

HB1xp67_ASAP7_75t_L g10948 ( 
.A(n_10730),
.Y(n_10948)
);

INVx2_ASAP7_75t_SL g10949 ( 
.A(n_10683),
.Y(n_10949)
);

INVx2_ASAP7_75t_L g10950 ( 
.A(n_10641),
.Y(n_10950)
);

AND2x2_ASAP7_75t_L g10951 ( 
.A(n_10622),
.B(n_1401),
.Y(n_10951)
);

INVx1_ASAP7_75t_L g10952 ( 
.A(n_10708),
.Y(n_10952)
);

INVx1_ASAP7_75t_L g10953 ( 
.A(n_10862),
.Y(n_10953)
);

AND2x2_ASAP7_75t_L g10954 ( 
.A(n_10906),
.B(n_10910),
.Y(n_10954)
);

OAI22xp5_ASAP7_75t_L g10955 ( 
.A1(n_10753),
.A2(n_1405),
.B1(n_1402),
.B2(n_1404),
.Y(n_10955)
);

OR2x2_ASAP7_75t_L g10956 ( 
.A(n_10634),
.B(n_1402),
.Y(n_10956)
);

INVx1_ASAP7_75t_L g10957 ( 
.A(n_10739),
.Y(n_10957)
);

AND2x2_ASAP7_75t_L g10958 ( 
.A(n_10663),
.B(n_1404),
.Y(n_10958)
);

AND2x4_ASAP7_75t_L g10959 ( 
.A(n_10722),
.B(n_1405),
.Y(n_10959)
);

BUFx6f_ASAP7_75t_L g10960 ( 
.A(n_10759),
.Y(n_10960)
);

AND2x2_ASAP7_75t_L g10961 ( 
.A(n_10717),
.B(n_1406),
.Y(n_10961)
);

OR2x2_ASAP7_75t_L g10962 ( 
.A(n_10606),
.B(n_1407),
.Y(n_10962)
);

AND2x2_ASAP7_75t_L g10963 ( 
.A(n_10673),
.B(n_1407),
.Y(n_10963)
);

INVx1_ASAP7_75t_L g10964 ( 
.A(n_10854),
.Y(n_10964)
);

INVx3_ASAP7_75t_L g10965 ( 
.A(n_10788),
.Y(n_10965)
);

AND2x2_ASAP7_75t_L g10966 ( 
.A(n_10662),
.B(n_1408),
.Y(n_10966)
);

AND2x2_ASAP7_75t_L g10967 ( 
.A(n_10678),
.B(n_1408),
.Y(n_10967)
);

AND2x4_ASAP7_75t_L g10968 ( 
.A(n_10693),
.B(n_1409),
.Y(n_10968)
);

INVx1_ASAP7_75t_L g10969 ( 
.A(n_10733),
.Y(n_10969)
);

AND2x2_ASAP7_75t_L g10970 ( 
.A(n_10848),
.B(n_1409),
.Y(n_10970)
);

AND2x2_ASAP7_75t_L g10971 ( 
.A(n_10706),
.B(n_1410),
.Y(n_10971)
);

HB1xp67_ASAP7_75t_L g10972 ( 
.A(n_10631),
.Y(n_10972)
);

NAND2xp5_ASAP7_75t_L g10973 ( 
.A(n_10777),
.B(n_1410),
.Y(n_10973)
);

AND2x2_ASAP7_75t_L g10974 ( 
.A(n_10847),
.B(n_1411),
.Y(n_10974)
);

OR2x2_ASAP7_75t_L g10975 ( 
.A(n_10613),
.B(n_1411),
.Y(n_10975)
);

INVxp67_ASAP7_75t_L g10976 ( 
.A(n_10720),
.Y(n_10976)
);

NAND2xp5_ASAP7_75t_L g10977 ( 
.A(n_10873),
.B(n_1412),
.Y(n_10977)
);

AND2x2_ASAP7_75t_L g10978 ( 
.A(n_10729),
.B(n_1413),
.Y(n_10978)
);

INVx2_ASAP7_75t_L g10979 ( 
.A(n_10923),
.Y(n_10979)
);

AND2x4_ASAP7_75t_SL g10980 ( 
.A(n_10615),
.B(n_1413),
.Y(n_10980)
);

BUFx3_ASAP7_75t_L g10981 ( 
.A(n_10902),
.Y(n_10981)
);

BUFx2_ASAP7_75t_L g10982 ( 
.A(n_10924),
.Y(n_10982)
);

INVx1_ASAP7_75t_L g10983 ( 
.A(n_10624),
.Y(n_10983)
);

AND2x2_ASAP7_75t_L g10984 ( 
.A(n_10761),
.B(n_1414),
.Y(n_10984)
);

OR2x2_ASAP7_75t_L g10985 ( 
.A(n_10882),
.B(n_1415),
.Y(n_10985)
);

INVx1_ASAP7_75t_L g10986 ( 
.A(n_10626),
.Y(n_10986)
);

INVx1_ASAP7_75t_L g10987 ( 
.A(n_10647),
.Y(n_10987)
);

AO21x2_ASAP7_75t_L g10988 ( 
.A1(n_10904),
.A2(n_1415),
.B(n_1416),
.Y(n_10988)
);

INVx1_ASAP7_75t_L g10989 ( 
.A(n_10657),
.Y(n_10989)
);

AND2x2_ASAP7_75t_L g10990 ( 
.A(n_10850),
.B(n_1417),
.Y(n_10990)
);

INVx1_ASAP7_75t_L g10991 ( 
.A(n_10661),
.Y(n_10991)
);

AND2x2_ASAP7_75t_L g10992 ( 
.A(n_10850),
.B(n_10639),
.Y(n_10992)
);

AND2x2_ASAP7_75t_L g10993 ( 
.A(n_10850),
.B(n_1417),
.Y(n_10993)
);

AND2x2_ASAP7_75t_L g10994 ( 
.A(n_10660),
.B(n_1418),
.Y(n_10994)
);

OR2x2_ASAP7_75t_L g10995 ( 
.A(n_10888),
.B(n_1419),
.Y(n_10995)
);

AND2x2_ASAP7_75t_L g10996 ( 
.A(n_10627),
.B(n_1419),
.Y(n_10996)
);

INVxp67_ASAP7_75t_SL g10997 ( 
.A(n_10612),
.Y(n_10997)
);

HB1xp67_ASAP7_75t_L g10998 ( 
.A(n_10750),
.Y(n_10998)
);

BUFx6f_ASAP7_75t_L g10999 ( 
.A(n_10685),
.Y(n_10999)
);

OR2x2_ASAP7_75t_L g11000 ( 
.A(n_10891),
.B(n_1420),
.Y(n_11000)
);

NAND2xp5_ASAP7_75t_L g11001 ( 
.A(n_10766),
.B(n_1420),
.Y(n_11001)
);

INVx1_ASAP7_75t_L g11002 ( 
.A(n_10664),
.Y(n_11002)
);

AND2x2_ASAP7_75t_L g11003 ( 
.A(n_10760),
.B(n_1421),
.Y(n_11003)
);

BUFx3_ASAP7_75t_L g11004 ( 
.A(n_10616),
.Y(n_11004)
);

NAND2xp5_ASAP7_75t_L g11005 ( 
.A(n_10610),
.B(n_1422),
.Y(n_11005)
);

AOI22xp33_ASAP7_75t_L g11006 ( 
.A1(n_10618),
.A2(n_1424),
.B1(n_1422),
.B2(n_1423),
.Y(n_11006)
);

AND2x4_ASAP7_75t_L g11007 ( 
.A(n_10895),
.B(n_10913),
.Y(n_11007)
);

INVxp67_ASAP7_75t_L g11008 ( 
.A(n_10831),
.Y(n_11008)
);

HB1xp67_ASAP7_75t_L g11009 ( 
.A(n_10620),
.Y(n_11009)
);

AND2x4_ASAP7_75t_L g11010 ( 
.A(n_10914),
.B(n_1423),
.Y(n_11010)
);

AND2x2_ASAP7_75t_L g11011 ( 
.A(n_10611),
.B(n_1424),
.Y(n_11011)
);

OAI22xp33_ASAP7_75t_L g11012 ( 
.A1(n_10652),
.A2(n_1428),
.B1(n_1426),
.B2(n_1427),
.Y(n_11012)
);

HB1xp67_ASAP7_75t_L g11013 ( 
.A(n_10620),
.Y(n_11013)
);

INVx1_ASAP7_75t_L g11014 ( 
.A(n_10686),
.Y(n_11014)
);

NOR2xp33_ASAP7_75t_L g11015 ( 
.A(n_10724),
.B(n_1426),
.Y(n_11015)
);

INVx2_ASAP7_75t_L g11016 ( 
.A(n_10629),
.Y(n_11016)
);

HB1xp67_ASAP7_75t_L g11017 ( 
.A(n_10629),
.Y(n_11017)
);

INVx3_ASAP7_75t_L g11018 ( 
.A(n_10876),
.Y(n_11018)
);

AND2x2_ASAP7_75t_SL g11019 ( 
.A(n_10752),
.B(n_10745),
.Y(n_11019)
);

INVx2_ASAP7_75t_SL g11020 ( 
.A(n_10890),
.Y(n_11020)
);

INVx2_ASAP7_75t_SL g11021 ( 
.A(n_10898),
.Y(n_11021)
);

INVx2_ASAP7_75t_L g11022 ( 
.A(n_10795),
.Y(n_11022)
);

INVx2_ASAP7_75t_L g11023 ( 
.A(n_10806),
.Y(n_11023)
);

OAI22xp5_ASAP7_75t_L g11024 ( 
.A1(n_10908),
.A2(n_10874),
.B1(n_10883),
.B2(n_10875),
.Y(n_11024)
);

NAND2xp5_ASAP7_75t_L g11025 ( 
.A(n_10778),
.B(n_1427),
.Y(n_11025)
);

INVx2_ASAP7_75t_L g11026 ( 
.A(n_10819),
.Y(n_11026)
);

AND2x2_ASAP7_75t_L g11027 ( 
.A(n_10918),
.B(n_1428),
.Y(n_11027)
);

BUFx6f_ASAP7_75t_L g11028 ( 
.A(n_10899),
.Y(n_11028)
);

INVx5_ASAP7_75t_SL g11029 ( 
.A(n_10756),
.Y(n_11029)
);

INVx1_ASAP7_75t_L g11030 ( 
.A(n_10704),
.Y(n_11030)
);

INVx2_ASAP7_75t_L g11031 ( 
.A(n_10827),
.Y(n_11031)
);

INVx1_ASAP7_75t_L g11032 ( 
.A(n_10705),
.Y(n_11032)
);

INVx3_ASAP7_75t_L g11033 ( 
.A(n_10649),
.Y(n_11033)
);

INVx4_ASAP7_75t_L g11034 ( 
.A(n_10694),
.Y(n_11034)
);

AND2x4_ASAP7_75t_L g11035 ( 
.A(n_10632),
.B(n_1430),
.Y(n_11035)
);

BUFx6f_ASAP7_75t_L g11036 ( 
.A(n_10817),
.Y(n_11036)
);

AND2x2_ASAP7_75t_L g11037 ( 
.A(n_10725),
.B(n_1431),
.Y(n_11037)
);

HB1xp67_ASAP7_75t_L g11038 ( 
.A(n_10690),
.Y(n_11038)
);

OR2x2_ASAP7_75t_L g11039 ( 
.A(n_10789),
.B(n_10621),
.Y(n_11039)
);

OR2x2_ASAP7_75t_L g11040 ( 
.A(n_10679),
.B(n_1431),
.Y(n_11040)
);

INVx2_ASAP7_75t_L g11041 ( 
.A(n_10828),
.Y(n_11041)
);

OR2x2_ASAP7_75t_L g11042 ( 
.A(n_10821),
.B(n_1432),
.Y(n_11042)
);

INVx1_ASAP7_75t_L g11043 ( 
.A(n_10710),
.Y(n_11043)
);

OR2x2_ASAP7_75t_L g11044 ( 
.A(n_10689),
.B(n_1432),
.Y(n_11044)
);

INVx2_ASAP7_75t_L g11045 ( 
.A(n_10830),
.Y(n_11045)
);

INVx2_ASAP7_75t_L g11046 ( 
.A(n_10734),
.Y(n_11046)
);

AND2x2_ASAP7_75t_L g11047 ( 
.A(n_10594),
.B(n_1434),
.Y(n_11047)
);

INVx1_ASAP7_75t_L g11048 ( 
.A(n_10716),
.Y(n_11048)
);

AND2x4_ASAP7_75t_SL g11049 ( 
.A(n_10731),
.B(n_1434),
.Y(n_11049)
);

INVx1_ASAP7_75t_L g11050 ( 
.A(n_10732),
.Y(n_11050)
);

AND2x2_ASAP7_75t_L g11051 ( 
.A(n_10614),
.B(n_1435),
.Y(n_11051)
);

INVx1_ASAP7_75t_L g11052 ( 
.A(n_10747),
.Y(n_11052)
);

NAND2xp5_ASAP7_75t_L g11053 ( 
.A(n_10721),
.B(n_1435),
.Y(n_11053)
);

INVx2_ASAP7_75t_L g11054 ( 
.A(n_10715),
.Y(n_11054)
);

BUFx6f_ASAP7_75t_L g11055 ( 
.A(n_10756),
.Y(n_11055)
);

HB1xp67_ASAP7_75t_L g11056 ( 
.A(n_10805),
.Y(n_11056)
);

INVx2_ASAP7_75t_L g11057 ( 
.A(n_10605),
.Y(n_11057)
);

OAI21x1_ASAP7_75t_L g11058 ( 
.A1(n_10807),
.A2(n_1437),
.B(n_1438),
.Y(n_11058)
);

INVx1_ASAP7_75t_L g11059 ( 
.A(n_10749),
.Y(n_11059)
);

INVx2_ASAP7_75t_L g11060 ( 
.A(n_10856),
.Y(n_11060)
);

AND2x2_ASAP7_75t_L g11061 ( 
.A(n_10877),
.B(n_1437),
.Y(n_11061)
);

INVx2_ASAP7_75t_L g11062 ( 
.A(n_10751),
.Y(n_11062)
);

AND2x2_ASAP7_75t_L g11063 ( 
.A(n_10878),
.B(n_1438),
.Y(n_11063)
);

INVx1_ASAP7_75t_L g11064 ( 
.A(n_10815),
.Y(n_11064)
);

AOI22xp5_ASAP7_75t_L g11065 ( 
.A1(n_10884),
.A2(n_1441),
.B1(n_1439),
.B2(n_1440),
.Y(n_11065)
);

AND2x2_ASAP7_75t_L g11066 ( 
.A(n_10880),
.B(n_1440),
.Y(n_11066)
);

OR2x2_ASAP7_75t_L g11067 ( 
.A(n_10692),
.B(n_1441),
.Y(n_11067)
);

AND2x2_ASAP7_75t_L g11068 ( 
.A(n_10887),
.B(n_1442),
.Y(n_11068)
);

NOR2x1_ASAP7_75t_L g11069 ( 
.A(n_10920),
.B(n_1442),
.Y(n_11069)
);

NAND2xp5_ASAP7_75t_SL g11070 ( 
.A(n_10737),
.B(n_1443),
.Y(n_11070)
);

OAI221xp5_ASAP7_75t_SL g11071 ( 
.A1(n_10892),
.A2(n_1446),
.B1(n_1444),
.B2(n_1445),
.C(n_1447),
.Y(n_11071)
);

NAND2xp5_ASAP7_75t_L g11072 ( 
.A(n_10798),
.B(n_1444),
.Y(n_11072)
);

INVx2_ASAP7_75t_L g11073 ( 
.A(n_10769),
.Y(n_11073)
);

NAND2xp5_ASAP7_75t_L g11074 ( 
.A(n_10852),
.B(n_1445),
.Y(n_11074)
);

INVx1_ASAP7_75t_L g11075 ( 
.A(n_10832),
.Y(n_11075)
);

INVx1_ASAP7_75t_L g11076 ( 
.A(n_10838),
.Y(n_11076)
);

AND2x2_ASAP7_75t_L g11077 ( 
.A(n_10896),
.B(n_1446),
.Y(n_11077)
);

AND2x2_ASAP7_75t_L g11078 ( 
.A(n_10905),
.B(n_1447),
.Y(n_11078)
);

INVx5_ASAP7_75t_SL g11079 ( 
.A(n_10731),
.Y(n_11079)
);

AND2x2_ASAP7_75t_L g11080 ( 
.A(n_10915),
.B(n_1448),
.Y(n_11080)
);

AND2x2_ASAP7_75t_L g11081 ( 
.A(n_10921),
.B(n_1448),
.Y(n_11081)
);

AND2x2_ASAP7_75t_L g11082 ( 
.A(n_10922),
.B(n_1449),
.Y(n_11082)
);

INVx2_ASAP7_75t_L g11083 ( 
.A(n_10814),
.Y(n_11083)
);

INVxp67_ASAP7_75t_SL g11084 ( 
.A(n_10813),
.Y(n_11084)
);

INVxp67_ASAP7_75t_L g11085 ( 
.A(n_10770),
.Y(n_11085)
);

AND2x2_ASAP7_75t_L g11086 ( 
.A(n_10628),
.B(n_1450),
.Y(n_11086)
);

INVx1_ASAP7_75t_L g11087 ( 
.A(n_10842),
.Y(n_11087)
);

AND2x2_ASAP7_75t_L g11088 ( 
.A(n_10718),
.B(n_1450),
.Y(n_11088)
);

INVx2_ASAP7_75t_L g11089 ( 
.A(n_10826),
.Y(n_11089)
);

HB1xp67_ASAP7_75t_L g11090 ( 
.A(n_10648),
.Y(n_11090)
);

INVx1_ASAP7_75t_L g11091 ( 
.A(n_10866),
.Y(n_11091)
);

INVx1_ASAP7_75t_L g11092 ( 
.A(n_10871),
.Y(n_11092)
);

NAND2xp5_ASAP7_75t_L g11093 ( 
.A(n_10810),
.B(n_1451),
.Y(n_11093)
);

INVx2_ASAP7_75t_SL g11094 ( 
.A(n_10701),
.Y(n_11094)
);

AND2x2_ASAP7_75t_L g11095 ( 
.A(n_10793),
.B(n_1452),
.Y(n_11095)
);

INVx1_ASAP7_75t_L g11096 ( 
.A(n_10829),
.Y(n_11096)
);

INVx1_ASAP7_75t_L g11097 ( 
.A(n_10802),
.Y(n_11097)
);

INVx3_ASAP7_75t_L g11098 ( 
.A(n_10740),
.Y(n_11098)
);

NAND2xp5_ASAP7_75t_L g11099 ( 
.A(n_10794),
.B(n_1452),
.Y(n_11099)
);

BUFx3_ASAP7_75t_L g11100 ( 
.A(n_10764),
.Y(n_11100)
);

AND2x2_ASAP7_75t_L g11101 ( 
.A(n_10765),
.B(n_1453),
.Y(n_11101)
);

AND2x2_ASAP7_75t_L g11102 ( 
.A(n_10763),
.B(n_1454),
.Y(n_11102)
);

AND2x2_ASAP7_75t_L g11103 ( 
.A(n_10601),
.B(n_1457),
.Y(n_11103)
);

HB1xp67_ASAP7_75t_L g11104 ( 
.A(n_10785),
.Y(n_11104)
);

INVx3_ASAP7_75t_L g11105 ( 
.A(n_10792),
.Y(n_11105)
);

AND2x2_ASAP7_75t_L g11106 ( 
.A(n_10651),
.B(n_1457),
.Y(n_11106)
);

INVx1_ASAP7_75t_L g11107 ( 
.A(n_10869),
.Y(n_11107)
);

AND2x2_ASAP7_75t_L g11108 ( 
.A(n_10670),
.B(n_1458),
.Y(n_11108)
);

AND2x2_ASAP7_75t_L g11109 ( 
.A(n_10671),
.B(n_1459),
.Y(n_11109)
);

OR2x2_ASAP7_75t_L g11110 ( 
.A(n_10684),
.B(n_1459),
.Y(n_11110)
);

AND2x2_ASAP7_75t_L g11111 ( 
.A(n_10676),
.B(n_1460),
.Y(n_11111)
);

NAND2xp5_ASAP7_75t_L g11112 ( 
.A(n_10803),
.B(n_1460),
.Y(n_11112)
);

INVx1_ASAP7_75t_L g11113 ( 
.A(n_10744),
.Y(n_11113)
);

INVx1_ASAP7_75t_L g11114 ( 
.A(n_10711),
.Y(n_11114)
);

INVx3_ASAP7_75t_L g11115 ( 
.A(n_10764),
.Y(n_11115)
);

OAI211xp5_ASAP7_75t_L g11116 ( 
.A1(n_10897),
.A2(n_1463),
.B(n_1461),
.C(n_1462),
.Y(n_11116)
);

AND2x2_ASAP7_75t_L g11117 ( 
.A(n_10691),
.B(n_1461),
.Y(n_11117)
);

AND2x4_ASAP7_75t_L g11118 ( 
.A(n_10666),
.B(n_1462),
.Y(n_11118)
);

CKINVDCx5p33_ASAP7_75t_R g11119 ( 
.A(n_10790),
.Y(n_11119)
);

INVx1_ASAP7_75t_L g11120 ( 
.A(n_10712),
.Y(n_11120)
);

AND2x2_ASAP7_75t_L g11121 ( 
.A(n_10695),
.B(n_1463),
.Y(n_11121)
);

INVx2_ASAP7_75t_L g11122 ( 
.A(n_10818),
.Y(n_11122)
);

AOI22xp5_ASAP7_75t_L g11123 ( 
.A1(n_10900),
.A2(n_1466),
.B1(n_1464),
.B2(n_1465),
.Y(n_11123)
);

AND2x4_ASAP7_75t_L g11124 ( 
.A(n_10650),
.B(n_1464),
.Y(n_11124)
);

OAI21xp33_ASAP7_75t_L g11125 ( 
.A1(n_10907),
.A2(n_1465),
.B(n_1466),
.Y(n_11125)
);

AND2x2_ASAP7_75t_L g11126 ( 
.A(n_10665),
.B(n_1467),
.Y(n_11126)
);

INVx2_ASAP7_75t_L g11127 ( 
.A(n_10820),
.Y(n_11127)
);

INVx1_ASAP7_75t_L g11128 ( 
.A(n_10726),
.Y(n_11128)
);

INVx1_ASAP7_75t_L g11129 ( 
.A(n_10840),
.Y(n_11129)
);

INVx1_ASAP7_75t_L g11130 ( 
.A(n_10863),
.Y(n_11130)
);

NAND2xp5_ASAP7_75t_L g11131 ( 
.A(n_10698),
.B(n_10669),
.Y(n_11131)
);

INVx2_ASAP7_75t_L g11132 ( 
.A(n_10735),
.Y(n_11132)
);

INVx11_ASAP7_75t_L g11133 ( 
.A(n_10764),
.Y(n_11133)
);

AND2x2_ASAP7_75t_L g11134 ( 
.A(n_10714),
.B(n_1468),
.Y(n_11134)
);

INVx1_ASAP7_75t_L g11135 ( 
.A(n_10867),
.Y(n_11135)
);

AOI22xp33_ASAP7_75t_L g11136 ( 
.A1(n_10703),
.A2(n_1471),
.B1(n_1469),
.B2(n_1470),
.Y(n_11136)
);

NAND2xp5_ASAP7_75t_L g11137 ( 
.A(n_10903),
.B(n_1469),
.Y(n_11137)
);

INVx2_ASAP7_75t_L g11138 ( 
.A(n_10741),
.Y(n_11138)
);

NAND2xp5_ASAP7_75t_L g11139 ( 
.A(n_10787),
.B(n_10796),
.Y(n_11139)
);

INVx2_ASAP7_75t_L g11140 ( 
.A(n_10746),
.Y(n_11140)
);

OAI21xp5_ASAP7_75t_L g11141 ( 
.A1(n_10603),
.A2(n_1471),
.B(n_1472),
.Y(n_11141)
);

BUFx2_ASAP7_75t_L g11142 ( 
.A(n_10767),
.Y(n_11142)
);

AOI22xp33_ASAP7_75t_L g11143 ( 
.A1(n_10736),
.A2(n_1475),
.B1(n_1472),
.B2(n_1474),
.Y(n_11143)
);

AND2x2_ASAP7_75t_L g11144 ( 
.A(n_10797),
.B(n_10822),
.Y(n_11144)
);

BUFx3_ASAP7_75t_L g11145 ( 
.A(n_10843),
.Y(n_11145)
);

NAND2xp5_ASAP7_75t_L g11146 ( 
.A(n_10816),
.B(n_1474),
.Y(n_11146)
);

HB1xp67_ASAP7_75t_L g11147 ( 
.A(n_10800),
.Y(n_11147)
);

INVx2_ASAP7_75t_L g11148 ( 
.A(n_10748),
.Y(n_11148)
);

INVx2_ASAP7_75t_L g11149 ( 
.A(n_10719),
.Y(n_11149)
);

INVx3_ASAP7_75t_L g11150 ( 
.A(n_10864),
.Y(n_11150)
);

INVx1_ASAP7_75t_L g11151 ( 
.A(n_10824),
.Y(n_11151)
);

AND2x2_ASAP7_75t_L g11152 ( 
.A(n_10822),
.B(n_10811),
.Y(n_11152)
);

INVx3_ASAP7_75t_L g11153 ( 
.A(n_10843),
.Y(n_11153)
);

NAND2xp5_ASAP7_75t_L g11154 ( 
.A(n_10775),
.B(n_10699),
.Y(n_11154)
);

OR2x2_ASAP7_75t_L g11155 ( 
.A(n_10870),
.B(n_1475),
.Y(n_11155)
);

INVx1_ASAP7_75t_L g11156 ( 
.A(n_10836),
.Y(n_11156)
);

INVx1_ASAP7_75t_L g11157 ( 
.A(n_10861),
.Y(n_11157)
);

INVx2_ASAP7_75t_L g11158 ( 
.A(n_10768),
.Y(n_11158)
);

INVx2_ASAP7_75t_L g11159 ( 
.A(n_10707),
.Y(n_11159)
);

AND2x2_ASAP7_75t_L g11160 ( 
.A(n_10645),
.B(n_1476),
.Y(n_11160)
);

NAND2xp5_ASAP7_75t_L g11161 ( 
.A(n_10617),
.B(n_1477),
.Y(n_11161)
);

AOI221xp5_ASAP7_75t_L g11162 ( 
.A1(n_10845),
.A2(n_1480),
.B1(n_1478),
.B2(n_1479),
.C(n_1481),
.Y(n_11162)
);

BUFx6f_ASAP7_75t_L g11163 ( 
.A(n_10658),
.Y(n_11163)
);

INVx1_ASAP7_75t_L g11164 ( 
.A(n_10767),
.Y(n_11164)
);

INVx2_ASAP7_75t_L g11165 ( 
.A(n_10801),
.Y(n_11165)
);

OAI222xp33_ASAP7_75t_L g11166 ( 
.A1(n_10638),
.A2(n_1482),
.B1(n_1484),
.B2(n_1478),
.C1(n_1481),
.C2(n_1483),
.Y(n_11166)
);

AND2x2_ASAP7_75t_L g11167 ( 
.A(n_10667),
.B(n_1482),
.Y(n_11167)
);

INVx1_ASAP7_75t_L g11168 ( 
.A(n_10776),
.Y(n_11168)
);

AND2x2_ASAP7_75t_L g11169 ( 
.A(n_10846),
.B(n_1484),
.Y(n_11169)
);

INVxp67_ASAP7_75t_L g11170 ( 
.A(n_10843),
.Y(n_11170)
);

INVx1_ASAP7_75t_L g11171 ( 
.A(n_10779),
.Y(n_11171)
);

INVx1_ASAP7_75t_L g11172 ( 
.A(n_10786),
.Y(n_11172)
);

INVx1_ASAP7_75t_L g11173 ( 
.A(n_10607),
.Y(n_11173)
);

INVx1_ASAP7_75t_L g11174 ( 
.A(n_10607),
.Y(n_11174)
);

INVx2_ASAP7_75t_L g11175 ( 
.A(n_10713),
.Y(n_11175)
);

NAND2xp5_ASAP7_75t_L g11176 ( 
.A(n_11142),
.B(n_10602),
.Y(n_11176)
);

NAND2xp5_ASAP7_75t_L g11177 ( 
.A(n_10946),
.B(n_10595),
.Y(n_11177)
);

NAND2xp5_ASAP7_75t_L g11178 ( 
.A(n_10982),
.B(n_10640),
.Y(n_11178)
);

AND2x2_ASAP7_75t_L g11179 ( 
.A(n_10929),
.B(n_10846),
.Y(n_11179)
);

INVx1_ASAP7_75t_L g11180 ( 
.A(n_10942),
.Y(n_11180)
);

INVx2_ASAP7_75t_L g11181 ( 
.A(n_10960),
.Y(n_11181)
);

AND2x2_ASAP7_75t_L g11182 ( 
.A(n_10941),
.B(n_10783),
.Y(n_11182)
);

OAI21xp5_ASAP7_75t_SL g11183 ( 
.A1(n_10935),
.A2(n_11024),
.B(n_11085),
.Y(n_11183)
);

NAND3xp33_ASAP7_75t_L g11184 ( 
.A(n_11104),
.B(n_10773),
.C(n_10637),
.Y(n_11184)
);

NAND2xp5_ASAP7_75t_L g11185 ( 
.A(n_11009),
.B(n_11013),
.Y(n_11185)
);

OAI22xp5_ASAP7_75t_L g11186 ( 
.A1(n_11164),
.A2(n_10709),
.B1(n_10727),
.B2(n_10762),
.Y(n_11186)
);

NAND2xp5_ASAP7_75t_L g11187 ( 
.A(n_11017),
.B(n_10656),
.Y(n_11187)
);

AND2x2_ASAP7_75t_L g11188 ( 
.A(n_10932),
.B(n_10783),
.Y(n_11188)
);

INVx1_ASAP7_75t_L g11189 ( 
.A(n_10948),
.Y(n_11189)
);

NAND2xp5_ASAP7_75t_L g11190 ( 
.A(n_11173),
.B(n_10623),
.Y(n_11190)
);

NAND2xp5_ASAP7_75t_L g11191 ( 
.A(n_11174),
.B(n_10881),
.Y(n_11191)
);

AOI21xp5_ASAP7_75t_L g11192 ( 
.A1(n_11001),
.A2(n_10643),
.B(n_10635),
.Y(n_11192)
);

OAI221xp5_ASAP7_75t_SL g11193 ( 
.A1(n_10976),
.A2(n_10653),
.B1(n_10755),
.B2(n_10812),
.C(n_10738),
.Y(n_11193)
);

AOI22xp33_ASAP7_75t_L g11194 ( 
.A1(n_11019),
.A2(n_10636),
.B1(n_10596),
.B2(n_10700),
.Y(n_11194)
);

NAND2xp5_ASAP7_75t_L g11195 ( 
.A(n_11016),
.B(n_10889),
.Y(n_11195)
);

NAND3xp33_ASAP7_75t_L g11196 ( 
.A(n_11147),
.B(n_10680),
.C(n_10774),
.Y(n_11196)
);

NAND2xp5_ASAP7_75t_SL g11197 ( 
.A(n_11055),
.B(n_10772),
.Y(n_11197)
);

AND2x2_ASAP7_75t_L g11198 ( 
.A(n_11029),
.B(n_10638),
.Y(n_11198)
);

NAND2xp5_ASAP7_75t_L g11199 ( 
.A(n_10996),
.B(n_10901),
.Y(n_11199)
);

AND2x2_ASAP7_75t_SL g11200 ( 
.A(n_11055),
.B(n_10825),
.Y(n_11200)
);

NOR2xp33_ASAP7_75t_SL g11201 ( 
.A(n_11119),
.B(n_10925),
.Y(n_11201)
);

NAND3xp33_ASAP7_75t_L g11202 ( 
.A(n_11090),
.B(n_10859),
.C(n_10675),
.Y(n_11202)
);

OAI22xp5_ASAP7_75t_L g11203 ( 
.A1(n_10997),
.A2(n_10644),
.B1(n_10872),
.B2(n_10758),
.Y(n_11203)
);

NAND2xp5_ASAP7_75t_L g11204 ( 
.A(n_11020),
.B(n_10702),
.Y(n_11204)
);

AND2x2_ASAP7_75t_L g11205 ( 
.A(n_11079),
.B(n_10644),
.Y(n_11205)
);

AND2x2_ASAP7_75t_L g11206 ( 
.A(n_10954),
.B(n_10979),
.Y(n_11206)
);

NAND3xp33_ASAP7_75t_L g11207 ( 
.A(n_11162),
.B(n_10865),
.C(n_10851),
.Y(n_11207)
);

NAND2xp5_ASAP7_75t_SL g11208 ( 
.A(n_11028),
.B(n_10849),
.Y(n_11208)
);

OAI22xp5_ASAP7_75t_L g11209 ( 
.A1(n_11071),
.A2(n_10823),
.B1(n_10809),
.B2(n_10791),
.Y(n_11209)
);

OAI21xp5_ASAP7_75t_SL g11210 ( 
.A1(n_11015),
.A2(n_10674),
.B(n_10858),
.Y(n_11210)
);

AND2x2_ASAP7_75t_L g11211 ( 
.A(n_10965),
.B(n_10608),
.Y(n_11211)
);

OAI221xp5_ASAP7_75t_L g11212 ( 
.A1(n_11084),
.A2(n_11131),
.B1(n_10928),
.B2(n_11125),
.C(n_11141),
.Y(n_11212)
);

OAI22xp5_ASAP7_75t_L g11213 ( 
.A1(n_11069),
.A2(n_11038),
.B1(n_10972),
.B2(n_11151),
.Y(n_11213)
);

NAND2xp5_ASAP7_75t_L g11214 ( 
.A(n_11021),
.B(n_10799),
.Y(n_11214)
);

OAI21xp33_ASAP7_75t_SL g11215 ( 
.A1(n_11156),
.A2(n_10771),
.B(n_10912),
.Y(n_11215)
);

AOI22xp33_ASAP7_75t_L g11216 ( 
.A1(n_10926),
.A2(n_10860),
.B1(n_10754),
.B2(n_10835),
.Y(n_11216)
);

NAND2xp5_ASAP7_75t_L g11217 ( 
.A(n_11170),
.B(n_10853),
.Y(n_11217)
);

NAND2xp5_ASAP7_75t_L g11218 ( 
.A(n_11094),
.B(n_10916),
.Y(n_11218)
);

OAI21xp33_ASAP7_75t_L g11219 ( 
.A1(n_10950),
.A2(n_10780),
.B(n_10599),
.Y(n_11219)
);

AOI22xp33_ASAP7_75t_L g11220 ( 
.A1(n_11070),
.A2(n_10784),
.B1(n_10844),
.B2(n_10837),
.Y(n_11220)
);

NAND2xp5_ASAP7_75t_L g11221 ( 
.A(n_11152),
.B(n_10687),
.Y(n_11221)
);

AND2x2_ASAP7_75t_L g11222 ( 
.A(n_11144),
.B(n_10857),
.Y(n_11222)
);

NAND4xp25_ASAP7_75t_L g11223 ( 
.A(n_11039),
.B(n_10677),
.C(n_10604),
.D(n_10839),
.Y(n_11223)
);

AND2x2_ASAP7_75t_L g11224 ( 
.A(n_11145),
.B(n_10672),
.Y(n_11224)
);

AND2x2_ASAP7_75t_L g11225 ( 
.A(n_10960),
.B(n_10682),
.Y(n_11225)
);

NAND3xp33_ASAP7_75t_L g11226 ( 
.A(n_11157),
.B(n_10894),
.C(n_10879),
.Y(n_11226)
);

NAND2xp5_ASAP7_75t_L g11227 ( 
.A(n_11018),
.B(n_10646),
.Y(n_11227)
);

NAND2xp5_ASAP7_75t_L g11228 ( 
.A(n_11153),
.B(n_10742),
.Y(n_11228)
);

NAND2xp5_ASAP7_75t_L g11229 ( 
.A(n_11115),
.B(n_10625),
.Y(n_11229)
);

NAND2xp5_ASAP7_75t_SL g11230 ( 
.A(n_11028),
.B(n_10757),
.Y(n_11230)
);

AND2x2_ASAP7_75t_L g11231 ( 
.A(n_11100),
.B(n_10855),
.Y(n_11231)
);

NAND2xp5_ASAP7_75t_L g11232 ( 
.A(n_11057),
.B(n_11008),
.Y(n_11232)
);

INVx1_ASAP7_75t_L g11233 ( 
.A(n_10998),
.Y(n_11233)
);

NAND2xp5_ASAP7_75t_L g11234 ( 
.A(n_11130),
.B(n_10723),
.Y(n_11234)
);

OAI22xp5_ASAP7_75t_L g11235 ( 
.A1(n_11025),
.A2(n_10841),
.B1(n_10833),
.B2(n_10893),
.Y(n_11235)
);

AND2x2_ASAP7_75t_L g11236 ( 
.A(n_11034),
.B(n_10917),
.Y(n_11236)
);

AND2x2_ASAP7_75t_L g11237 ( 
.A(n_10944),
.B(n_10728),
.Y(n_11237)
);

AND2x2_ASAP7_75t_L g11238 ( 
.A(n_10949),
.B(n_11033),
.Y(n_11238)
);

NAND2xp5_ASAP7_75t_L g11239 ( 
.A(n_11135),
.B(n_1486),
.Y(n_11239)
);

NAND2xp5_ASAP7_75t_L g11240 ( 
.A(n_11129),
.B(n_1486),
.Y(n_11240)
);

NAND2xp5_ASAP7_75t_L g11241 ( 
.A(n_11122),
.B(n_1487),
.Y(n_11241)
);

NAND3xp33_ASAP7_75t_L g11242 ( 
.A(n_11056),
.B(n_10893),
.C(n_10728),
.Y(n_11242)
);

NAND4xp25_ASAP7_75t_L g11243 ( 
.A(n_10931),
.B(n_10688),
.C(n_10804),
.D(n_10868),
.Y(n_11243)
);

NAND2xp5_ASAP7_75t_L g11244 ( 
.A(n_11127),
.B(n_11132),
.Y(n_11244)
);

NAND3xp33_ASAP7_75t_L g11245 ( 
.A(n_11116),
.B(n_10688),
.C(n_10804),
.Y(n_11245)
);

OAI22xp5_ASAP7_75t_L g11246 ( 
.A1(n_11154),
.A2(n_10868),
.B1(n_1490),
.B2(n_1487),
.Y(n_11246)
);

NAND2xp5_ASAP7_75t_L g11247 ( 
.A(n_11138),
.B(n_1489),
.Y(n_11247)
);

NAND3xp33_ASAP7_75t_L g11248 ( 
.A(n_10934),
.B(n_1491),
.C(n_1492),
.Y(n_11248)
);

NAND3xp33_ASAP7_75t_L g11249 ( 
.A(n_10945),
.B(n_10952),
.C(n_10947),
.Y(n_11249)
);

NAND2xp5_ASAP7_75t_L g11250 ( 
.A(n_11140),
.B(n_1491),
.Y(n_11250)
);

NAND2xp5_ASAP7_75t_L g11251 ( 
.A(n_11148),
.B(n_1492),
.Y(n_11251)
);

INVx1_ASAP7_75t_L g11252 ( 
.A(n_10957),
.Y(n_11252)
);

AOI22xp33_ASAP7_75t_SL g11253 ( 
.A1(n_10938),
.A2(n_10988),
.B1(n_11165),
.B2(n_11053),
.Y(n_11253)
);

OAI21xp5_ASAP7_75t_SL g11254 ( 
.A1(n_11006),
.A2(n_1493),
.B(n_1494),
.Y(n_11254)
);

AOI22xp33_ASAP7_75t_L g11255 ( 
.A1(n_11022),
.A2(n_1497),
.B1(n_1493),
.B2(n_1495),
.Y(n_11255)
);

OAI22xp5_ASAP7_75t_L g11256 ( 
.A1(n_11136),
.A2(n_1499),
.B1(n_1495),
.B2(n_1498),
.Y(n_11256)
);

AND2x2_ASAP7_75t_L g11257 ( 
.A(n_10930),
.B(n_1498),
.Y(n_11257)
);

NOR2xp33_ASAP7_75t_L g11258 ( 
.A(n_11133),
.B(n_1499),
.Y(n_11258)
);

NOR3xp33_ASAP7_75t_L g11259 ( 
.A(n_11172),
.B(n_1501),
.C(n_1502),
.Y(n_11259)
);

NAND3xp33_ASAP7_75t_L g11260 ( 
.A(n_11096),
.B(n_1501),
.C(n_1503),
.Y(n_11260)
);

NOR2xp33_ASAP7_75t_SL g11261 ( 
.A(n_11166),
.B(n_1503),
.Y(n_11261)
);

AOI22xp33_ASAP7_75t_L g11262 ( 
.A1(n_11023),
.A2(n_1506),
.B1(n_1504),
.B2(n_1505),
.Y(n_11262)
);

NAND3xp33_ASAP7_75t_L g11263 ( 
.A(n_10964),
.B(n_1504),
.C(n_1505),
.Y(n_11263)
);

OAI21xp5_ASAP7_75t_SL g11264 ( 
.A1(n_11143),
.A2(n_1506),
.B(n_1508),
.Y(n_11264)
);

NAND3xp33_ASAP7_75t_L g11265 ( 
.A(n_11065),
.B(n_1508),
.C(n_1509),
.Y(n_11265)
);

NAND2xp5_ASAP7_75t_L g11266 ( 
.A(n_11158),
.B(n_1509),
.Y(n_11266)
);

NAND2xp5_ASAP7_75t_L g11267 ( 
.A(n_11159),
.B(n_1510),
.Y(n_11267)
);

NAND3xp33_ASAP7_75t_L g11268 ( 
.A(n_11123),
.B(n_1511),
.C(n_1512),
.Y(n_11268)
);

NAND2xp5_ASAP7_75t_L g11269 ( 
.A(n_11175),
.B(n_1511),
.Y(n_11269)
);

NAND2xp5_ASAP7_75t_SL g11270 ( 
.A(n_10999),
.B(n_1513),
.Y(n_11270)
);

AOI22xp5_ASAP7_75t_L g11271 ( 
.A1(n_10939),
.A2(n_1515),
.B1(n_1513),
.B2(n_1514),
.Y(n_11271)
);

AND2x2_ASAP7_75t_L g11272 ( 
.A(n_10940),
.B(n_1514),
.Y(n_11272)
);

AND2x2_ASAP7_75t_L g11273 ( 
.A(n_11098),
.B(n_1515),
.Y(n_11273)
);

OAI22xp5_ASAP7_75t_L g11274 ( 
.A1(n_11105),
.A2(n_1518),
.B1(n_1516),
.B2(n_1517),
.Y(n_11274)
);

OAI221xp5_ASAP7_75t_L g11275 ( 
.A1(n_10977),
.A2(n_1518),
.B1(n_1516),
.B2(n_1517),
.C(n_1519),
.Y(n_11275)
);

AND4x1_ASAP7_75t_L g11276 ( 
.A(n_10927),
.B(n_1521),
.C(n_1519),
.D(n_1520),
.Y(n_11276)
);

AND2x2_ASAP7_75t_L g11277 ( 
.A(n_11150),
.B(n_1520),
.Y(n_11277)
);

NAND3xp33_ASAP7_75t_L g11278 ( 
.A(n_10953),
.B(n_11007),
.C(n_11097),
.Y(n_11278)
);

NAND3xp33_ASAP7_75t_L g11279 ( 
.A(n_11107),
.B(n_1521),
.C(n_1522),
.Y(n_11279)
);

AND2x2_ASAP7_75t_L g11280 ( 
.A(n_10981),
.B(n_1522),
.Y(n_11280)
);

NAND2xp5_ASAP7_75t_L g11281 ( 
.A(n_11168),
.B(n_1523),
.Y(n_11281)
);

AND2x2_ASAP7_75t_L g11282 ( 
.A(n_11004),
.B(n_1524),
.Y(n_11282)
);

NAND2xp5_ASAP7_75t_L g11283 ( 
.A(n_11171),
.B(n_1525),
.Y(n_11283)
);

NAND3xp33_ASAP7_75t_L g11284 ( 
.A(n_11113),
.B(n_1526),
.C(n_1527),
.Y(n_11284)
);

AOI21xp33_ASAP7_75t_L g11285 ( 
.A1(n_11026),
.A2(n_1526),
.B(n_1527),
.Y(n_11285)
);

NOR3xp33_ASAP7_75t_L g11286 ( 
.A(n_11012),
.B(n_1528),
.C(n_1529),
.Y(n_11286)
);

NAND2xp5_ASAP7_75t_L g11287 ( 
.A(n_11060),
.B(n_1531),
.Y(n_11287)
);

AND2x2_ASAP7_75t_L g11288 ( 
.A(n_10999),
.B(n_1531),
.Y(n_11288)
);

AND2x2_ASAP7_75t_L g11289 ( 
.A(n_11036),
.B(n_11163),
.Y(n_11289)
);

OAI21xp33_ASAP7_75t_L g11290 ( 
.A1(n_10992),
.A2(n_1532),
.B(n_1533),
.Y(n_11290)
);

NAND4xp25_ASAP7_75t_L g11291 ( 
.A(n_10969),
.B(n_1535),
.C(n_1532),
.D(n_1534),
.Y(n_11291)
);

OAI22xp5_ASAP7_75t_L g11292 ( 
.A1(n_11139),
.A2(n_1538),
.B1(n_1536),
.B2(n_1537),
.Y(n_11292)
);

NAND3xp33_ASAP7_75t_L g11293 ( 
.A(n_11114),
.B(n_1536),
.C(n_1537),
.Y(n_11293)
);

NAND2xp5_ASAP7_75t_L g11294 ( 
.A(n_11073),
.B(n_1538),
.Y(n_11294)
);

AND2x2_ASAP7_75t_L g11295 ( 
.A(n_11036),
.B(n_1539),
.Y(n_11295)
);

AOI22xp33_ASAP7_75t_L g11296 ( 
.A1(n_11031),
.A2(n_1542),
.B1(n_1540),
.B2(n_1541),
.Y(n_11296)
);

NAND2xp5_ASAP7_75t_L g11297 ( 
.A(n_11149),
.B(n_11062),
.Y(n_11297)
);

INVx1_ASAP7_75t_L g11298 ( 
.A(n_11042),
.Y(n_11298)
);

NAND2xp5_ASAP7_75t_L g11299 ( 
.A(n_11128),
.B(n_1540),
.Y(n_11299)
);

NAND2xp5_ASAP7_75t_L g11300 ( 
.A(n_11041),
.B(n_1541),
.Y(n_11300)
);

AND2x2_ASAP7_75t_SL g11301 ( 
.A(n_11049),
.B(n_1542),
.Y(n_11301)
);

NAND2xp5_ASAP7_75t_L g11302 ( 
.A(n_11045),
.B(n_1543),
.Y(n_11302)
);

AOI221xp5_ASAP7_75t_L g11303 ( 
.A1(n_10955),
.A2(n_1545),
.B1(n_1543),
.B2(n_1544),
.C(n_1546),
.Y(n_11303)
);

NAND2xp5_ASAP7_75t_L g11304 ( 
.A(n_11046),
.B(n_11120),
.Y(n_11304)
);

OAI221xp5_ASAP7_75t_SL g11305 ( 
.A1(n_11072),
.A2(n_1548),
.B1(n_1546),
.B2(n_1547),
.C(n_1549),
.Y(n_11305)
);

AND2x2_ASAP7_75t_L g11306 ( 
.A(n_11163),
.B(n_1548),
.Y(n_11306)
);

NAND3xp33_ASAP7_75t_L g11307 ( 
.A(n_10973),
.B(n_1549),
.C(n_1550),
.Y(n_11307)
);

AND2x2_ASAP7_75t_L g11308 ( 
.A(n_10943),
.B(n_1551),
.Y(n_11308)
);

NAND2xp5_ASAP7_75t_SL g11309 ( 
.A(n_10956),
.B(n_1551),
.Y(n_11309)
);

NAND3xp33_ASAP7_75t_L g11310 ( 
.A(n_11083),
.B(n_1552),
.C(n_1553),
.Y(n_11310)
);

NAND3xp33_ASAP7_75t_L g11311 ( 
.A(n_11089),
.B(n_1553),
.C(n_1554),
.Y(n_11311)
);

AND2x2_ASAP7_75t_L g11312 ( 
.A(n_10936),
.B(n_10966),
.Y(n_11312)
);

AND2x2_ASAP7_75t_L g11313 ( 
.A(n_10970),
.B(n_1555),
.Y(n_11313)
);

AND2x2_ASAP7_75t_L g11314 ( 
.A(n_10984),
.B(n_1555),
.Y(n_11314)
);

AND2x2_ASAP7_75t_L g11315 ( 
.A(n_10971),
.B(n_1556),
.Y(n_11315)
);

NAND3xp33_ASAP7_75t_L g11316 ( 
.A(n_11137),
.B(n_1556),
.C(n_1557),
.Y(n_11316)
);

NAND2xp5_ASAP7_75t_L g11317 ( 
.A(n_10990),
.B(n_1557),
.Y(n_11317)
);

AND2x2_ASAP7_75t_L g11318 ( 
.A(n_11003),
.B(n_1558),
.Y(n_11318)
);

NOR2xp33_ASAP7_75t_L g11319 ( 
.A(n_10933),
.B(n_1558),
.Y(n_11319)
);

NAND3xp33_ASAP7_75t_L g11320 ( 
.A(n_11099),
.B(n_1559),
.C(n_1560),
.Y(n_11320)
);

NAND2xp5_ASAP7_75t_L g11321 ( 
.A(n_10993),
.B(n_1559),
.Y(n_11321)
);

AND2x2_ASAP7_75t_L g11322 ( 
.A(n_11037),
.B(n_1562),
.Y(n_11322)
);

NAND2xp5_ASAP7_75t_L g11323 ( 
.A(n_10994),
.B(n_1562),
.Y(n_11323)
);

OAI221xp5_ASAP7_75t_SL g11324 ( 
.A1(n_11074),
.A2(n_11161),
.B1(n_11093),
.B2(n_10937),
.C(n_11054),
.Y(n_11324)
);

OAI221xp5_ASAP7_75t_L g11325 ( 
.A1(n_11146),
.A2(n_1565),
.B1(n_1563),
.B2(n_1564),
.C(n_1566),
.Y(n_11325)
);

OAI21xp33_ASAP7_75t_L g11326 ( 
.A1(n_10983),
.A2(n_1563),
.B(n_1564),
.Y(n_11326)
);

OAI21xp5_ASAP7_75t_L g11327 ( 
.A1(n_11058),
.A2(n_1565),
.B(n_1566),
.Y(n_11327)
);

AOI22xp33_ASAP7_75t_L g11328 ( 
.A1(n_10986),
.A2(n_1570),
.B1(n_1568),
.B2(n_1569),
.Y(n_11328)
);

OA21x2_ASAP7_75t_L g11329 ( 
.A1(n_10987),
.A2(n_1568),
.B(n_1569),
.Y(n_11329)
);

NAND2xp5_ASAP7_75t_L g11330 ( 
.A(n_11027),
.B(n_1570),
.Y(n_11330)
);

NAND2xp5_ASAP7_75t_L g11331 ( 
.A(n_10951),
.B(n_10967),
.Y(n_11331)
);

AND2x2_ASAP7_75t_SL g11332 ( 
.A(n_10980),
.B(n_1571),
.Y(n_11332)
);

NAND2xp5_ASAP7_75t_SL g11333 ( 
.A(n_10959),
.B(n_1572),
.Y(n_11333)
);

AND2x2_ASAP7_75t_L g11334 ( 
.A(n_11088),
.B(n_1572),
.Y(n_11334)
);

AND2x2_ASAP7_75t_L g11335 ( 
.A(n_11101),
.B(n_1573),
.Y(n_11335)
);

AND2x2_ASAP7_75t_L g11336 ( 
.A(n_11086),
.B(n_1573),
.Y(n_11336)
);

NAND2xp5_ASAP7_75t_L g11337 ( 
.A(n_10974),
.B(n_1574),
.Y(n_11337)
);

NAND2xp5_ASAP7_75t_SL g11338 ( 
.A(n_11010),
.B(n_11118),
.Y(n_11338)
);

AND2x2_ASAP7_75t_L g11339 ( 
.A(n_11011),
.B(n_1574),
.Y(n_11339)
);

OAI22xp5_ASAP7_75t_L g11340 ( 
.A1(n_10962),
.A2(n_1577),
.B1(n_1575),
.B2(n_1576),
.Y(n_11340)
);

AND2x2_ASAP7_75t_L g11341 ( 
.A(n_11051),
.B(n_1575),
.Y(n_11341)
);

NAND3xp33_ASAP7_75t_L g11342 ( 
.A(n_10989),
.B(n_11002),
.C(n_10991),
.Y(n_11342)
);

AND2x2_ASAP7_75t_L g11343 ( 
.A(n_11047),
.B(n_1577),
.Y(n_11343)
);

NAND2xp5_ASAP7_75t_L g11344 ( 
.A(n_10975),
.B(n_1579),
.Y(n_11344)
);

OAI221xp5_ASAP7_75t_L g11345 ( 
.A1(n_11112),
.A2(n_1581),
.B1(n_1579),
.B2(n_1580),
.C(n_1582),
.Y(n_11345)
);

NAND2xp5_ASAP7_75t_L g11346 ( 
.A(n_10985),
.B(n_1580),
.Y(n_11346)
);

AOI22xp33_ASAP7_75t_SL g11347 ( 
.A1(n_11169),
.A2(n_1585),
.B1(n_1581),
.B2(n_1583),
.Y(n_11347)
);

NAND2xp5_ASAP7_75t_L g11348 ( 
.A(n_10995),
.B(n_1585),
.Y(n_11348)
);

AND2x2_ASAP7_75t_L g11349 ( 
.A(n_11061),
.B(n_1586),
.Y(n_11349)
);

NAND2xp5_ASAP7_75t_L g11350 ( 
.A(n_11000),
.B(n_1586),
.Y(n_11350)
);

NAND2xp5_ASAP7_75t_L g11351 ( 
.A(n_11095),
.B(n_1587),
.Y(n_11351)
);

NAND2xp5_ASAP7_75t_SL g11352 ( 
.A(n_11124),
.B(n_1588),
.Y(n_11352)
);

AND2x2_ASAP7_75t_L g11353 ( 
.A(n_11063),
.B(n_1588),
.Y(n_11353)
);

NAND4xp25_ASAP7_75t_L g11354 ( 
.A(n_11014),
.B(n_11030),
.C(n_11043),
.D(n_11032),
.Y(n_11354)
);

NAND2xp5_ASAP7_75t_L g11355 ( 
.A(n_11134),
.B(n_1589),
.Y(n_11355)
);

AND2x2_ASAP7_75t_L g11356 ( 
.A(n_11066),
.B(n_1589),
.Y(n_11356)
);

NAND2xp5_ASAP7_75t_L g11357 ( 
.A(n_10961),
.B(n_1591),
.Y(n_11357)
);

NAND3xp33_ASAP7_75t_L g11358 ( 
.A(n_11048),
.B(n_1591),
.C(n_1592),
.Y(n_11358)
);

INVx1_ASAP7_75t_L g11359 ( 
.A(n_11050),
.Y(n_11359)
);

NAND2xp5_ASAP7_75t_L g11360 ( 
.A(n_10978),
.B(n_1592),
.Y(n_11360)
);

NAND2xp5_ASAP7_75t_SL g11361 ( 
.A(n_11035),
.B(n_1593),
.Y(n_11361)
);

OAI21xp5_ASAP7_75t_SL g11362 ( 
.A1(n_11110),
.A2(n_1593),
.B(n_1594),
.Y(n_11362)
);

NAND3xp33_ASAP7_75t_L g11363 ( 
.A(n_11052),
.B(n_1595),
.C(n_1596),
.Y(n_11363)
);

NAND3xp33_ASAP7_75t_L g11364 ( 
.A(n_11059),
.B(n_1595),
.C(n_1596),
.Y(n_11364)
);

AOI221xp5_ASAP7_75t_L g11365 ( 
.A1(n_11064),
.A2(n_1600),
.B1(n_1598),
.B2(n_1599),
.C(n_1601),
.Y(n_11365)
);

NAND3xp33_ASAP7_75t_L g11366 ( 
.A(n_11075),
.B(n_11087),
.C(n_11076),
.Y(n_11366)
);

OAI21xp33_ASAP7_75t_L g11367 ( 
.A1(n_11091),
.A2(n_1598),
.B(n_1602),
.Y(n_11367)
);

NAND2xp5_ASAP7_75t_L g11368 ( 
.A(n_11068),
.B(n_11077),
.Y(n_11368)
);

NAND2xp33_ASAP7_75t_SL g11369 ( 
.A(n_11040),
.B(n_11078),
.Y(n_11369)
);

NAND2xp5_ASAP7_75t_L g11370 ( 
.A(n_11080),
.B(n_1602),
.Y(n_11370)
);

AND2x2_ASAP7_75t_L g11371 ( 
.A(n_11081),
.B(n_1603),
.Y(n_11371)
);

AND2x2_ASAP7_75t_L g11372 ( 
.A(n_11082),
.B(n_1603),
.Y(n_11372)
);

OR2x2_ASAP7_75t_SL g11373 ( 
.A(n_11044),
.B(n_1604),
.Y(n_11373)
);

NOR2xp33_ASAP7_75t_L g11374 ( 
.A(n_11067),
.B(n_11155),
.Y(n_11374)
);

AND2x2_ASAP7_75t_L g11375 ( 
.A(n_11106),
.B(n_1604),
.Y(n_11375)
);

NAND2xp5_ASAP7_75t_SL g11376 ( 
.A(n_10968),
.B(n_1605),
.Y(n_11376)
);

OAI22xp5_ASAP7_75t_L g11377 ( 
.A1(n_11092),
.A2(n_11005),
.B1(n_10963),
.B2(n_10958),
.Y(n_11377)
);

AND2x2_ASAP7_75t_L g11378 ( 
.A(n_11198),
.B(n_11103),
.Y(n_11378)
);

INVx4_ASAP7_75t_L g11379 ( 
.A(n_11289),
.Y(n_11379)
);

AND2x2_ASAP7_75t_L g11380 ( 
.A(n_11205),
.B(n_11126),
.Y(n_11380)
);

INVx2_ASAP7_75t_L g11381 ( 
.A(n_11200),
.Y(n_11381)
);

INVx2_ASAP7_75t_L g11382 ( 
.A(n_11225),
.Y(n_11382)
);

NOR2xp33_ASAP7_75t_L g11383 ( 
.A(n_11219),
.B(n_11108),
.Y(n_11383)
);

INVxp67_ASAP7_75t_SL g11384 ( 
.A(n_11227),
.Y(n_11384)
);

AND2x2_ASAP7_75t_L g11385 ( 
.A(n_11179),
.B(n_11109),
.Y(n_11385)
);

OR2x2_ASAP7_75t_L g11386 ( 
.A(n_11185),
.B(n_11111),
.Y(n_11386)
);

INVx2_ASAP7_75t_L g11387 ( 
.A(n_11182),
.Y(n_11387)
);

AND2x2_ASAP7_75t_SL g11388 ( 
.A(n_11194),
.B(n_11102),
.Y(n_11388)
);

NAND2xp5_ASAP7_75t_L g11389 ( 
.A(n_11192),
.B(n_11167),
.Y(n_11389)
);

AO21x2_ASAP7_75t_L g11390 ( 
.A1(n_11213),
.A2(n_11121),
.B(n_11117),
.Y(n_11390)
);

NAND3xp33_ASAP7_75t_L g11391 ( 
.A(n_11196),
.B(n_11160),
.C(n_1605),
.Y(n_11391)
);

INVx2_ASAP7_75t_L g11392 ( 
.A(n_11211),
.Y(n_11392)
);

NOR2xp33_ASAP7_75t_SL g11393 ( 
.A(n_11301),
.B(n_1606),
.Y(n_11393)
);

AOI211xp5_ASAP7_75t_L g11394 ( 
.A1(n_11184),
.A2(n_1609),
.B(n_1607),
.C(n_1608),
.Y(n_11394)
);

INVx1_ASAP7_75t_L g11395 ( 
.A(n_11180),
.Y(n_11395)
);

OR2x2_ASAP7_75t_L g11396 ( 
.A(n_11176),
.B(n_1608),
.Y(n_11396)
);

NAND2xp5_ASAP7_75t_L g11397 ( 
.A(n_11237),
.B(n_1609),
.Y(n_11397)
);

INVx2_ASAP7_75t_L g11398 ( 
.A(n_11224),
.Y(n_11398)
);

AND2x2_ASAP7_75t_L g11399 ( 
.A(n_11188),
.B(n_1611),
.Y(n_11399)
);

INVx2_ASAP7_75t_SL g11400 ( 
.A(n_11332),
.Y(n_11400)
);

NOR3xp33_ASAP7_75t_L g11401 ( 
.A(n_11183),
.B(n_1612),
.C(n_1613),
.Y(n_11401)
);

INVx1_ASAP7_75t_SL g11402 ( 
.A(n_11312),
.Y(n_11402)
);

OR2x2_ASAP7_75t_L g11403 ( 
.A(n_11232),
.B(n_1612),
.Y(n_11403)
);

INVx2_ASAP7_75t_L g11404 ( 
.A(n_11206),
.Y(n_11404)
);

AND2x2_ASAP7_75t_L g11405 ( 
.A(n_11238),
.B(n_11222),
.Y(n_11405)
);

NAND2xp5_ASAP7_75t_L g11406 ( 
.A(n_11261),
.B(n_1613),
.Y(n_11406)
);

AND2x2_ASAP7_75t_L g11407 ( 
.A(n_11181),
.B(n_1614),
.Y(n_11407)
);

AND2x2_ASAP7_75t_L g11408 ( 
.A(n_11236),
.B(n_1614),
.Y(n_11408)
);

AOI22xp5_ASAP7_75t_L g11409 ( 
.A1(n_11186),
.A2(n_1617),
.B1(n_1615),
.B2(n_1616),
.Y(n_11409)
);

INVx1_ASAP7_75t_L g11410 ( 
.A(n_11189),
.Y(n_11410)
);

INVx2_ASAP7_75t_L g11411 ( 
.A(n_11288),
.Y(n_11411)
);

INVx2_ASAP7_75t_L g11412 ( 
.A(n_11295),
.Y(n_11412)
);

AOI22xp33_ASAP7_75t_L g11413 ( 
.A1(n_11202),
.A2(n_11242),
.B1(n_11212),
.B2(n_11191),
.Y(n_11413)
);

INVx1_ASAP7_75t_L g11414 ( 
.A(n_11233),
.Y(n_11414)
);

NAND2xp5_ASAP7_75t_L g11415 ( 
.A(n_11253),
.B(n_1615),
.Y(n_11415)
);

HB1xp67_ASAP7_75t_L g11416 ( 
.A(n_11197),
.Y(n_11416)
);

AND2x2_ASAP7_75t_L g11417 ( 
.A(n_11231),
.B(n_1617),
.Y(n_11417)
);

NAND3xp33_ASAP7_75t_L g11418 ( 
.A(n_11226),
.B(n_1618),
.C(n_1619),
.Y(n_11418)
);

INVx2_ASAP7_75t_L g11419 ( 
.A(n_11277),
.Y(n_11419)
);

OAI221xp5_ASAP7_75t_L g11420 ( 
.A1(n_11215),
.A2(n_1620),
.B1(n_1618),
.B2(n_1619),
.C(n_1621),
.Y(n_11420)
);

INVx1_ASAP7_75t_L g11421 ( 
.A(n_11297),
.Y(n_11421)
);

BUFx3_ASAP7_75t_L g11422 ( 
.A(n_11306),
.Y(n_11422)
);

INVxp67_ASAP7_75t_SL g11423 ( 
.A(n_11221),
.Y(n_11423)
);

NOR2xp33_ASAP7_75t_L g11424 ( 
.A(n_11199),
.B(n_1621),
.Y(n_11424)
);

NAND2xp5_ASAP7_75t_L g11425 ( 
.A(n_11235),
.B(n_1622),
.Y(n_11425)
);

AND2x2_ASAP7_75t_L g11426 ( 
.A(n_11201),
.B(n_1622),
.Y(n_11426)
);

OR2x2_ASAP7_75t_L g11427 ( 
.A(n_11178),
.B(n_1623),
.Y(n_11427)
);

OR2x2_ASAP7_75t_L g11428 ( 
.A(n_11177),
.B(n_1624),
.Y(n_11428)
);

OR2x2_ASAP7_75t_L g11429 ( 
.A(n_11187),
.B(n_1624),
.Y(n_11429)
);

INVx1_ASAP7_75t_L g11430 ( 
.A(n_11304),
.Y(n_11430)
);

BUFx3_ASAP7_75t_L g11431 ( 
.A(n_11273),
.Y(n_11431)
);

NOR2xp33_ASAP7_75t_L g11432 ( 
.A(n_11223),
.B(n_1625),
.Y(n_11432)
);

BUFx2_ASAP7_75t_L g11433 ( 
.A(n_11369),
.Y(n_11433)
);

NAND2xp5_ASAP7_75t_L g11434 ( 
.A(n_11220),
.B(n_1625),
.Y(n_11434)
);

NAND3xp33_ASAP7_75t_L g11435 ( 
.A(n_11245),
.B(n_1626),
.C(n_1627),
.Y(n_11435)
);

NAND2xp5_ASAP7_75t_SL g11436 ( 
.A(n_11246),
.B(n_1626),
.Y(n_11436)
);

AND2x2_ASAP7_75t_L g11437 ( 
.A(n_11298),
.B(n_1628),
.Y(n_11437)
);

NAND3xp33_ASAP7_75t_L g11438 ( 
.A(n_11249),
.B(n_1629),
.C(n_1630),
.Y(n_11438)
);

INVx2_ASAP7_75t_L g11439 ( 
.A(n_11257),
.Y(n_11439)
);

INVx1_ASAP7_75t_L g11440 ( 
.A(n_11244),
.Y(n_11440)
);

INVx1_ASAP7_75t_L g11441 ( 
.A(n_11351),
.Y(n_11441)
);

NAND2xp5_ASAP7_75t_SL g11442 ( 
.A(n_11207),
.B(n_1629),
.Y(n_11442)
);

NAND2xp5_ASAP7_75t_L g11443 ( 
.A(n_11374),
.B(n_1630),
.Y(n_11443)
);

INVx1_ASAP7_75t_L g11444 ( 
.A(n_11355),
.Y(n_11444)
);

NOR2xp33_ASAP7_75t_SL g11445 ( 
.A(n_11324),
.B(n_1631),
.Y(n_11445)
);

BUFx6f_ASAP7_75t_L g11446 ( 
.A(n_11280),
.Y(n_11446)
);

INVx1_ASAP7_75t_L g11447 ( 
.A(n_11228),
.Y(n_11447)
);

AOI22xp5_ASAP7_75t_L g11448 ( 
.A1(n_11209),
.A2(n_1633),
.B1(n_1631),
.B2(n_1632),
.Y(n_11448)
);

INVx2_ASAP7_75t_L g11449 ( 
.A(n_11272),
.Y(n_11449)
);

AND2x2_ASAP7_75t_L g11450 ( 
.A(n_11338),
.B(n_1632),
.Y(n_11450)
);

AND2x2_ASAP7_75t_L g11451 ( 
.A(n_11230),
.B(n_1633),
.Y(n_11451)
);

BUFx2_ASAP7_75t_L g11452 ( 
.A(n_11373),
.Y(n_11452)
);

AND2x4_ASAP7_75t_L g11453 ( 
.A(n_11278),
.B(n_1634),
.Y(n_11453)
);

AND2x2_ASAP7_75t_L g11454 ( 
.A(n_11368),
.B(n_1634),
.Y(n_11454)
);

INVx3_ASAP7_75t_L g11455 ( 
.A(n_11282),
.Y(n_11455)
);

INVx1_ASAP7_75t_L g11456 ( 
.A(n_11241),
.Y(n_11456)
);

INVx2_ASAP7_75t_L g11457 ( 
.A(n_11318),
.Y(n_11457)
);

AOI22xp33_ASAP7_75t_L g11458 ( 
.A1(n_11208),
.A2(n_1637),
.B1(n_1635),
.B2(n_1636),
.Y(n_11458)
);

INVx4_ASAP7_75t_L g11459 ( 
.A(n_11336),
.Y(n_11459)
);

INVx5_ASAP7_75t_L g11460 ( 
.A(n_11315),
.Y(n_11460)
);

AND2x2_ASAP7_75t_L g11461 ( 
.A(n_11195),
.B(n_1635),
.Y(n_11461)
);

BUFx3_ASAP7_75t_L g11462 ( 
.A(n_11375),
.Y(n_11462)
);

AND2x2_ASAP7_75t_L g11463 ( 
.A(n_11331),
.B(n_1637),
.Y(n_11463)
);

OR2x2_ASAP7_75t_L g11464 ( 
.A(n_11190),
.B(n_1638),
.Y(n_11464)
);

INVx2_ASAP7_75t_L g11465 ( 
.A(n_11314),
.Y(n_11465)
);

NAND2xp5_ASAP7_75t_L g11466 ( 
.A(n_11362),
.B(n_1639),
.Y(n_11466)
);

OR2x2_ASAP7_75t_L g11467 ( 
.A(n_11234),
.B(n_1639),
.Y(n_11467)
);

INVx1_ASAP7_75t_L g11468 ( 
.A(n_11247),
.Y(n_11468)
);

INVx1_ASAP7_75t_L g11469 ( 
.A(n_11250),
.Y(n_11469)
);

AND2x4_ASAP7_75t_L g11470 ( 
.A(n_11252),
.B(n_1640),
.Y(n_11470)
);

NAND3xp33_ASAP7_75t_L g11471 ( 
.A(n_11193),
.B(n_1640),
.C(n_1641),
.Y(n_11471)
);

AND2x2_ASAP7_75t_SL g11472 ( 
.A(n_11286),
.B(n_1641),
.Y(n_11472)
);

INVx2_ASAP7_75t_L g11473 ( 
.A(n_11322),
.Y(n_11473)
);

INVx2_ASAP7_75t_L g11474 ( 
.A(n_11308),
.Y(n_11474)
);

INVx1_ASAP7_75t_L g11475 ( 
.A(n_11251),
.Y(n_11475)
);

NAND2xp5_ASAP7_75t_L g11476 ( 
.A(n_11210),
.B(n_1642),
.Y(n_11476)
);

INVx1_ASAP7_75t_L g11477 ( 
.A(n_11266),
.Y(n_11477)
);

CKINVDCx16_ASAP7_75t_R g11478 ( 
.A(n_11203),
.Y(n_11478)
);

BUFx3_ASAP7_75t_L g11479 ( 
.A(n_11334),
.Y(n_11479)
);

INVx4_ASAP7_75t_L g11480 ( 
.A(n_11335),
.Y(n_11480)
);

AOI33xp33_ASAP7_75t_L g11481 ( 
.A1(n_11216),
.A2(n_1645),
.A3(n_1648),
.B1(n_1642),
.B2(n_1644),
.B3(n_1647),
.Y(n_11481)
);

AND2x2_ASAP7_75t_L g11482 ( 
.A(n_11217),
.B(n_1644),
.Y(n_11482)
);

BUFx6f_ASAP7_75t_L g11483 ( 
.A(n_11339),
.Y(n_11483)
);

INVx2_ASAP7_75t_L g11484 ( 
.A(n_11313),
.Y(n_11484)
);

BUFx3_ASAP7_75t_L g11485 ( 
.A(n_11341),
.Y(n_11485)
);

AND2x2_ASAP7_75t_L g11486 ( 
.A(n_11214),
.B(n_1648),
.Y(n_11486)
);

NOR3xp33_ASAP7_75t_L g11487 ( 
.A(n_11229),
.B(n_1649),
.C(n_1650),
.Y(n_11487)
);

OAI22xp5_ASAP7_75t_L g11488 ( 
.A1(n_11265),
.A2(n_1651),
.B1(n_1649),
.B2(n_1650),
.Y(n_11488)
);

NAND3xp33_ASAP7_75t_L g11489 ( 
.A(n_11243),
.B(n_1651),
.C(n_1652),
.Y(n_11489)
);

INVx1_ASAP7_75t_L g11490 ( 
.A(n_11267),
.Y(n_11490)
);

NAND3xp33_ASAP7_75t_L g11491 ( 
.A(n_11259),
.B(n_1652),
.C(n_1653),
.Y(n_11491)
);

INVx1_ASAP7_75t_L g11492 ( 
.A(n_11269),
.Y(n_11492)
);

AND2x2_ASAP7_75t_L g11493 ( 
.A(n_11349),
.B(n_1654),
.Y(n_11493)
);

INVx1_ASAP7_75t_L g11494 ( 
.A(n_11287),
.Y(n_11494)
);

AND2x2_ASAP7_75t_SL g11495 ( 
.A(n_11276),
.B(n_1655),
.Y(n_11495)
);

AND2x2_ASAP7_75t_L g11496 ( 
.A(n_11353),
.B(n_1656),
.Y(n_11496)
);

AND2x4_ASAP7_75t_L g11497 ( 
.A(n_11356),
.B(n_1656),
.Y(n_11497)
);

AND2x2_ASAP7_75t_L g11498 ( 
.A(n_11371),
.B(n_1657),
.Y(n_11498)
);

INVx2_ASAP7_75t_L g11499 ( 
.A(n_11372),
.Y(n_11499)
);

INVx3_ASAP7_75t_L g11500 ( 
.A(n_11343),
.Y(n_11500)
);

NOR2x1_ASAP7_75t_SL g11501 ( 
.A(n_11270),
.B(n_1657),
.Y(n_11501)
);

AND2x2_ASAP7_75t_L g11502 ( 
.A(n_11218),
.B(n_1658),
.Y(n_11502)
);

AND2x2_ASAP7_75t_L g11503 ( 
.A(n_11204),
.B(n_1658),
.Y(n_11503)
);

AND2x2_ASAP7_75t_L g11504 ( 
.A(n_11377),
.B(n_1659),
.Y(n_11504)
);

INVx1_ASAP7_75t_L g11505 ( 
.A(n_11294),
.Y(n_11505)
);

BUFx2_ASAP7_75t_L g11506 ( 
.A(n_11329),
.Y(n_11506)
);

INVx2_ASAP7_75t_L g11507 ( 
.A(n_11329),
.Y(n_11507)
);

OAI221xp5_ASAP7_75t_L g11508 ( 
.A1(n_11264),
.A2(n_1662),
.B1(n_1660),
.B2(n_1661),
.C(n_1663),
.Y(n_11508)
);

INVx3_ASAP7_75t_L g11509 ( 
.A(n_11359),
.Y(n_11509)
);

AND2x2_ASAP7_75t_L g11510 ( 
.A(n_11258),
.B(n_1660),
.Y(n_11510)
);

AND2x4_ASAP7_75t_L g11511 ( 
.A(n_11376),
.B(n_1661),
.Y(n_11511)
);

INVx2_ASAP7_75t_SL g11512 ( 
.A(n_11333),
.Y(n_11512)
);

HB1xp67_ASAP7_75t_L g11513 ( 
.A(n_11309),
.Y(n_11513)
);

INVx1_ASAP7_75t_L g11514 ( 
.A(n_11370),
.Y(n_11514)
);

NAND3xp33_ASAP7_75t_L g11515 ( 
.A(n_11365),
.B(n_1664),
.C(n_1665),
.Y(n_11515)
);

NAND2xp5_ASAP7_75t_L g11516 ( 
.A(n_11290),
.B(n_1665),
.Y(n_11516)
);

AND2x4_ASAP7_75t_L g11517 ( 
.A(n_11352),
.B(n_1666),
.Y(n_11517)
);

INVx1_ASAP7_75t_L g11518 ( 
.A(n_11300),
.Y(n_11518)
);

NAND2xp5_ASAP7_75t_L g11519 ( 
.A(n_11319),
.B(n_1666),
.Y(n_11519)
);

AND2x2_ASAP7_75t_L g11520 ( 
.A(n_11302),
.B(n_2799),
.Y(n_11520)
);

AND2x2_ASAP7_75t_L g11521 ( 
.A(n_11240),
.B(n_2799),
.Y(n_11521)
);

AND2x2_ASAP7_75t_L g11522 ( 
.A(n_11281),
.B(n_2800),
.Y(n_11522)
);

INVx11_ASAP7_75t_L g11523 ( 
.A(n_11361),
.Y(n_11523)
);

INVx1_ASAP7_75t_L g11524 ( 
.A(n_11344),
.Y(n_11524)
);

INVx1_ASAP7_75t_L g11525 ( 
.A(n_11346),
.Y(n_11525)
);

AOI221xp5_ASAP7_75t_L g11526 ( 
.A1(n_11354),
.A2(n_1669),
.B1(n_1667),
.B2(n_1668),
.C(n_1670),
.Y(n_11526)
);

AOI33xp33_ASAP7_75t_L g11527 ( 
.A1(n_11347),
.A2(n_1672),
.A3(n_1674),
.B1(n_1668),
.B2(n_1671),
.B3(n_1673),
.Y(n_11527)
);

NOR2x1_ASAP7_75t_L g11528 ( 
.A(n_11316),
.B(n_11320),
.Y(n_11528)
);

NAND2xp5_ASAP7_75t_L g11529 ( 
.A(n_11299),
.B(n_11283),
.Y(n_11529)
);

AND2x2_ASAP7_75t_L g11530 ( 
.A(n_11239),
.B(n_2806),
.Y(n_11530)
);

INVx1_ASAP7_75t_L g11531 ( 
.A(n_11348),
.Y(n_11531)
);

AND2x2_ASAP7_75t_L g11532 ( 
.A(n_11327),
.B(n_2806),
.Y(n_11532)
);

AO21x2_ASAP7_75t_L g11533 ( 
.A1(n_11285),
.A2(n_1671),
.B(n_1672),
.Y(n_11533)
);

INVx2_ASAP7_75t_L g11534 ( 
.A(n_11400),
.Y(n_11534)
);

INVx2_ASAP7_75t_L g11535 ( 
.A(n_11460),
.Y(n_11535)
);

AND2x2_ASAP7_75t_L g11536 ( 
.A(n_11405),
.B(n_11330),
.Y(n_11536)
);

AND2x2_ASAP7_75t_L g11537 ( 
.A(n_11378),
.B(n_11317),
.Y(n_11537)
);

OR2x2_ASAP7_75t_L g11538 ( 
.A(n_11402),
.B(n_11307),
.Y(n_11538)
);

AND2x2_ASAP7_75t_L g11539 ( 
.A(n_11380),
.B(n_11321),
.Y(n_11539)
);

INVx1_ASAP7_75t_L g11540 ( 
.A(n_11506),
.Y(n_11540)
);

INVx1_ASAP7_75t_L g11541 ( 
.A(n_11493),
.Y(n_11541)
);

INVx1_ASAP7_75t_L g11542 ( 
.A(n_11496),
.Y(n_11542)
);

AND2x2_ASAP7_75t_L g11543 ( 
.A(n_11379),
.B(n_11323),
.Y(n_11543)
);

AND2x2_ASAP7_75t_L g11544 ( 
.A(n_11381),
.B(n_11360),
.Y(n_11544)
);

AND2x2_ASAP7_75t_L g11545 ( 
.A(n_11460),
.B(n_11357),
.Y(n_11545)
);

AND2x4_ASAP7_75t_L g11546 ( 
.A(n_11398),
.B(n_11342),
.Y(n_11546)
);

NAND2xp5_ASAP7_75t_L g11547 ( 
.A(n_11452),
.B(n_11350),
.Y(n_11547)
);

AND2x2_ASAP7_75t_L g11548 ( 
.A(n_11385),
.B(n_11337),
.Y(n_11548)
);

NAND2xp5_ASAP7_75t_L g11549 ( 
.A(n_11495),
.B(n_11248),
.Y(n_11549)
);

NAND2xp5_ASAP7_75t_L g11550 ( 
.A(n_11478),
.B(n_11326),
.Y(n_11550)
);

NAND2xp5_ASAP7_75t_L g11551 ( 
.A(n_11433),
.B(n_11367),
.Y(n_11551)
);

NAND2xp5_ASAP7_75t_L g11552 ( 
.A(n_11388),
.B(n_11260),
.Y(n_11552)
);

AND2x2_ASAP7_75t_L g11553 ( 
.A(n_11382),
.B(n_11366),
.Y(n_11553)
);

OR2x2_ASAP7_75t_L g11554 ( 
.A(n_11397),
.B(n_11263),
.Y(n_11554)
);

OR2x2_ASAP7_75t_L g11555 ( 
.A(n_11396),
.B(n_11279),
.Y(n_11555)
);

AND2x2_ASAP7_75t_L g11556 ( 
.A(n_11459),
.B(n_11284),
.Y(n_11556)
);

INVx1_ASAP7_75t_L g11557 ( 
.A(n_11498),
.Y(n_11557)
);

INVx1_ASAP7_75t_L g11558 ( 
.A(n_11437),
.Y(n_11558)
);

INVx2_ASAP7_75t_L g11559 ( 
.A(n_11446),
.Y(n_11559)
);

AND2x2_ASAP7_75t_L g11560 ( 
.A(n_11480),
.B(n_11293),
.Y(n_11560)
);

AND2x2_ASAP7_75t_L g11561 ( 
.A(n_11392),
.B(n_11271),
.Y(n_11561)
);

INVx2_ASAP7_75t_L g11562 ( 
.A(n_11446),
.Y(n_11562)
);

AND2x4_ASAP7_75t_L g11563 ( 
.A(n_11462),
.B(n_11310),
.Y(n_11563)
);

AND2x2_ASAP7_75t_L g11564 ( 
.A(n_11404),
.B(n_11311),
.Y(n_11564)
);

OR2x2_ASAP7_75t_L g11565 ( 
.A(n_11386),
.B(n_11291),
.Y(n_11565)
);

AND2x2_ASAP7_75t_L g11566 ( 
.A(n_11399),
.B(n_11340),
.Y(n_11566)
);

INVx1_ASAP7_75t_L g11567 ( 
.A(n_11450),
.Y(n_11567)
);

AND2x2_ASAP7_75t_L g11568 ( 
.A(n_11451),
.B(n_11358),
.Y(n_11568)
);

NAND2x1_ASAP7_75t_L g11569 ( 
.A(n_11455),
.B(n_11363),
.Y(n_11569)
);

AND2x2_ASAP7_75t_L g11570 ( 
.A(n_11387),
.B(n_11364),
.Y(n_11570)
);

AND2x2_ASAP7_75t_L g11571 ( 
.A(n_11416),
.B(n_11292),
.Y(n_11571)
);

INVx2_ASAP7_75t_L g11572 ( 
.A(n_11483),
.Y(n_11572)
);

INVx1_ASAP7_75t_L g11573 ( 
.A(n_11417),
.Y(n_11573)
);

NAND2xp5_ASAP7_75t_L g11574 ( 
.A(n_11390),
.B(n_11254),
.Y(n_11574)
);

OR2x6_ASAP7_75t_L g11575 ( 
.A(n_11422),
.B(n_11268),
.Y(n_11575)
);

INVx1_ASAP7_75t_L g11576 ( 
.A(n_11457),
.Y(n_11576)
);

INVx2_ASAP7_75t_L g11577 ( 
.A(n_11483),
.Y(n_11577)
);

NAND2xp5_ASAP7_75t_L g11578 ( 
.A(n_11453),
.B(n_11274),
.Y(n_11578)
);

INVx2_ASAP7_75t_L g11579 ( 
.A(n_11479),
.Y(n_11579)
);

AND2x2_ASAP7_75t_L g11580 ( 
.A(n_11485),
.B(n_11255),
.Y(n_11580)
);

NAND2x1_ASAP7_75t_L g11581 ( 
.A(n_11507),
.B(n_11262),
.Y(n_11581)
);

INVx1_ASAP7_75t_L g11582 ( 
.A(n_11465),
.Y(n_11582)
);

AND2x2_ASAP7_75t_L g11583 ( 
.A(n_11500),
.B(n_11296),
.Y(n_11583)
);

AND2x2_ASAP7_75t_L g11584 ( 
.A(n_11431),
.B(n_11328),
.Y(n_11584)
);

AND2x2_ASAP7_75t_L g11585 ( 
.A(n_11411),
.B(n_11412),
.Y(n_11585)
);

NAND2xp5_ASAP7_75t_L g11586 ( 
.A(n_11426),
.B(n_11413),
.Y(n_11586)
);

INVx1_ASAP7_75t_L g11587 ( 
.A(n_11473),
.Y(n_11587)
);

OR2x2_ASAP7_75t_L g11588 ( 
.A(n_11389),
.B(n_11305),
.Y(n_11588)
);

NAND2xp5_ASAP7_75t_L g11589 ( 
.A(n_11383),
.B(n_11275),
.Y(n_11589)
);

INVx2_ASAP7_75t_L g11590 ( 
.A(n_11497),
.Y(n_11590)
);

AND2x2_ASAP7_75t_L g11591 ( 
.A(n_11461),
.B(n_11303),
.Y(n_11591)
);

OR2x2_ASAP7_75t_L g11592 ( 
.A(n_11512),
.B(n_11325),
.Y(n_11592)
);

INVx1_ASAP7_75t_L g11593 ( 
.A(n_11474),
.Y(n_11593)
);

AND2x4_ASAP7_75t_L g11594 ( 
.A(n_11419),
.B(n_11345),
.Y(n_11594)
);

AND2x4_ASAP7_75t_SL g11595 ( 
.A(n_11439),
.B(n_11256),
.Y(n_11595)
);

OAI221xp5_ASAP7_75t_SL g11596 ( 
.A1(n_11489),
.A2(n_1691),
.B1(n_1700),
.B2(n_1683),
.C(n_1673),
.Y(n_11596)
);

AND2x2_ASAP7_75t_L g11597 ( 
.A(n_11484),
.B(n_1675),
.Y(n_11597)
);

NAND2xp5_ASAP7_75t_L g11598 ( 
.A(n_11423),
.B(n_1675),
.Y(n_11598)
);

INVx1_ASAP7_75t_L g11599 ( 
.A(n_11499),
.Y(n_11599)
);

NAND2xp5_ASAP7_75t_L g11600 ( 
.A(n_11408),
.B(n_1676),
.Y(n_11600)
);

AND2x2_ASAP7_75t_L g11601 ( 
.A(n_11513),
.B(n_1676),
.Y(n_11601)
);

NAND2xp5_ASAP7_75t_L g11602 ( 
.A(n_11472),
.B(n_1677),
.Y(n_11602)
);

AND2x2_ASAP7_75t_L g11603 ( 
.A(n_11454),
.B(n_1678),
.Y(n_11603)
);

INVx1_ASAP7_75t_L g11604 ( 
.A(n_11407),
.Y(n_11604)
);

AND2x2_ASAP7_75t_L g11605 ( 
.A(n_11449),
.B(n_1678),
.Y(n_11605)
);

AND2x2_ASAP7_75t_L g11606 ( 
.A(n_11482),
.B(n_1679),
.Y(n_11606)
);

INVx2_ASAP7_75t_L g11607 ( 
.A(n_11501),
.Y(n_11607)
);

AND2x2_ASAP7_75t_L g11608 ( 
.A(n_11463),
.B(n_1679),
.Y(n_11608)
);

INVx1_ASAP7_75t_L g11609 ( 
.A(n_11395),
.Y(n_11609)
);

OR2x2_ASAP7_75t_L g11610 ( 
.A(n_11467),
.B(n_1680),
.Y(n_11610)
);

OR2x2_ASAP7_75t_L g11611 ( 
.A(n_11415),
.B(n_1680),
.Y(n_11611)
);

INVx2_ASAP7_75t_L g11612 ( 
.A(n_11470),
.Y(n_11612)
);

AND2x2_ASAP7_75t_L g11613 ( 
.A(n_11384),
.B(n_1681),
.Y(n_11613)
);

AND2x4_ASAP7_75t_L g11614 ( 
.A(n_11410),
.B(n_1681),
.Y(n_11614)
);

NAND2xp5_ASAP7_75t_L g11615 ( 
.A(n_11393),
.B(n_11445),
.Y(n_11615)
);

OR2x2_ASAP7_75t_L g11616 ( 
.A(n_11476),
.B(n_1683),
.Y(n_11616)
);

NAND2xp5_ASAP7_75t_SL g11617 ( 
.A(n_11391),
.B(n_1684),
.Y(n_11617)
);

NAND2xp5_ASAP7_75t_L g11618 ( 
.A(n_11424),
.B(n_1684),
.Y(n_11618)
);

HB1xp67_ASAP7_75t_L g11619 ( 
.A(n_11523),
.Y(n_11619)
);

INVx1_ASAP7_75t_L g11620 ( 
.A(n_11414),
.Y(n_11620)
);

AND2x2_ASAP7_75t_L g11621 ( 
.A(n_11502),
.B(n_1685),
.Y(n_11621)
);

INVx1_ASAP7_75t_L g11622 ( 
.A(n_11403),
.Y(n_11622)
);

AND2x4_ASAP7_75t_L g11623 ( 
.A(n_11447),
.B(n_1686),
.Y(n_11623)
);

AND3x2_ASAP7_75t_L g11624 ( 
.A(n_11394),
.B(n_2805),
.C(n_1687),
.Y(n_11624)
);

NAND2x1p5_ASAP7_75t_SL g11625 ( 
.A(n_11528),
.B(n_1687),
.Y(n_11625)
);

OR2x2_ASAP7_75t_L g11626 ( 
.A(n_11425),
.B(n_1688),
.Y(n_11626)
);

INVx1_ASAP7_75t_L g11627 ( 
.A(n_11520),
.Y(n_11627)
);

AND2x2_ASAP7_75t_L g11628 ( 
.A(n_11503),
.B(n_1689),
.Y(n_11628)
);

HB1xp67_ASAP7_75t_L g11629 ( 
.A(n_11533),
.Y(n_11629)
);

AND2x2_ASAP7_75t_L g11630 ( 
.A(n_11486),
.B(n_1689),
.Y(n_11630)
);

OR2x2_ASAP7_75t_L g11631 ( 
.A(n_11464),
.B(n_1690),
.Y(n_11631)
);

NAND2x1p5_ASAP7_75t_L g11632 ( 
.A(n_11511),
.B(n_1690),
.Y(n_11632)
);

INVx1_ASAP7_75t_L g11633 ( 
.A(n_11521),
.Y(n_11633)
);

INVx1_ASAP7_75t_L g11634 ( 
.A(n_11522),
.Y(n_11634)
);

INVx1_ASAP7_75t_L g11635 ( 
.A(n_11530),
.Y(n_11635)
);

OR2x2_ASAP7_75t_L g11636 ( 
.A(n_11428),
.B(n_1691),
.Y(n_11636)
);

AND2x4_ASAP7_75t_L g11637 ( 
.A(n_11517),
.B(n_1692),
.Y(n_11637)
);

AND2x4_ASAP7_75t_L g11638 ( 
.A(n_11440),
.B(n_1693),
.Y(n_11638)
);

NAND2xp5_ASAP7_75t_L g11639 ( 
.A(n_11481),
.B(n_1693),
.Y(n_11639)
);

INVx2_ASAP7_75t_L g11640 ( 
.A(n_11510),
.Y(n_11640)
);

INVx2_ASAP7_75t_L g11641 ( 
.A(n_11509),
.Y(n_11641)
);

AND2x2_ASAP7_75t_L g11642 ( 
.A(n_11532),
.B(n_1694),
.Y(n_11642)
);

INVx1_ASAP7_75t_L g11643 ( 
.A(n_11429),
.Y(n_11643)
);

INVx1_ASAP7_75t_L g11644 ( 
.A(n_11427),
.Y(n_11644)
);

AND2x2_ASAP7_75t_L g11645 ( 
.A(n_11504),
.B(n_1696),
.Y(n_11645)
);

INVx1_ASAP7_75t_L g11646 ( 
.A(n_11441),
.Y(n_11646)
);

INVx1_ASAP7_75t_L g11647 ( 
.A(n_11444),
.Y(n_11647)
);

AND2x4_ASAP7_75t_L g11648 ( 
.A(n_11421),
.B(n_1697),
.Y(n_11648)
);

NOR2xp33_ASAP7_75t_L g11649 ( 
.A(n_11435),
.B(n_1697),
.Y(n_11649)
);

INVx1_ASAP7_75t_L g11650 ( 
.A(n_11514),
.Y(n_11650)
);

OR2x2_ASAP7_75t_L g11651 ( 
.A(n_11442),
.B(n_1698),
.Y(n_11651)
);

NAND2x1p5_ASAP7_75t_L g11652 ( 
.A(n_11436),
.B(n_1698),
.Y(n_11652)
);

INVx1_ASAP7_75t_L g11653 ( 
.A(n_11524),
.Y(n_11653)
);

NAND2xp5_ASAP7_75t_L g11654 ( 
.A(n_11401),
.B(n_1699),
.Y(n_11654)
);

INVx2_ASAP7_75t_L g11655 ( 
.A(n_11525),
.Y(n_11655)
);

AND2x2_ASAP7_75t_L g11656 ( 
.A(n_11531),
.B(n_1699),
.Y(n_11656)
);

AND2x4_ASAP7_75t_L g11657 ( 
.A(n_11430),
.B(n_1701),
.Y(n_11657)
);

NOR2xp33_ASAP7_75t_L g11658 ( 
.A(n_11471),
.B(n_1701),
.Y(n_11658)
);

NOR2xp33_ASAP7_75t_L g11659 ( 
.A(n_11420),
.B(n_1702),
.Y(n_11659)
);

AND2x2_ASAP7_75t_L g11660 ( 
.A(n_11518),
.B(n_1702),
.Y(n_11660)
);

NOR2xp33_ASAP7_75t_SL g11661 ( 
.A(n_11418),
.B(n_1703),
.Y(n_11661)
);

NAND2xp5_ASAP7_75t_L g11662 ( 
.A(n_11432),
.B(n_1704),
.Y(n_11662)
);

AND2x2_ASAP7_75t_L g11663 ( 
.A(n_11456),
.B(n_1704),
.Y(n_11663)
);

AND2x2_ASAP7_75t_L g11664 ( 
.A(n_11468),
.B(n_1705),
.Y(n_11664)
);

INVx1_ASAP7_75t_L g11665 ( 
.A(n_11443),
.Y(n_11665)
);

INVx2_ASAP7_75t_L g11666 ( 
.A(n_11535),
.Y(n_11666)
);

BUFx2_ASAP7_75t_L g11667 ( 
.A(n_11607),
.Y(n_11667)
);

INVx1_ASAP7_75t_L g11668 ( 
.A(n_11540),
.Y(n_11668)
);

INVx1_ASAP7_75t_L g11669 ( 
.A(n_11534),
.Y(n_11669)
);

INVx1_ASAP7_75t_L g11670 ( 
.A(n_11606),
.Y(n_11670)
);

OR2x2_ASAP7_75t_L g11671 ( 
.A(n_11625),
.B(n_11529),
.Y(n_11671)
);

OR2x2_ASAP7_75t_L g11672 ( 
.A(n_11549),
.B(n_11438),
.Y(n_11672)
);

INVx2_ASAP7_75t_L g11673 ( 
.A(n_11632),
.Y(n_11673)
);

INVx2_ASAP7_75t_L g11674 ( 
.A(n_11545),
.Y(n_11674)
);

INVx2_ASAP7_75t_L g11675 ( 
.A(n_11572),
.Y(n_11675)
);

NAND2x1p5_ASAP7_75t_L g11676 ( 
.A(n_11637),
.B(n_11543),
.Y(n_11676)
);

INVx1_ASAP7_75t_L g11677 ( 
.A(n_11603),
.Y(n_11677)
);

NAND2xp5_ASAP7_75t_L g11678 ( 
.A(n_11624),
.B(n_11409),
.Y(n_11678)
);

BUFx2_ASAP7_75t_L g11679 ( 
.A(n_11546),
.Y(n_11679)
);

INVx1_ASAP7_75t_L g11680 ( 
.A(n_11608),
.Y(n_11680)
);

AND2x2_ASAP7_75t_L g11681 ( 
.A(n_11619),
.B(n_11469),
.Y(n_11681)
);

AND2x4_ASAP7_75t_L g11682 ( 
.A(n_11579),
.B(n_11475),
.Y(n_11682)
);

AND2x2_ASAP7_75t_L g11683 ( 
.A(n_11566),
.B(n_11477),
.Y(n_11683)
);

AND2x4_ASAP7_75t_SL g11684 ( 
.A(n_11590),
.B(n_11490),
.Y(n_11684)
);

INVx1_ASAP7_75t_L g11685 ( 
.A(n_11621),
.Y(n_11685)
);

O2A1O1Ixp5_ASAP7_75t_L g11686 ( 
.A1(n_11574),
.A2(n_11581),
.B(n_11552),
.C(n_11569),
.Y(n_11686)
);

NAND2xp5_ASAP7_75t_L g11687 ( 
.A(n_11577),
.B(n_11448),
.Y(n_11687)
);

OR2x2_ASAP7_75t_L g11688 ( 
.A(n_11565),
.B(n_11434),
.Y(n_11688)
);

INVx1_ASAP7_75t_L g11689 ( 
.A(n_11628),
.Y(n_11689)
);

AND2x2_ASAP7_75t_L g11690 ( 
.A(n_11556),
.B(n_11492),
.Y(n_11690)
);

INVx1_ASAP7_75t_L g11691 ( 
.A(n_11630),
.Y(n_11691)
);

NAND2xp5_ASAP7_75t_L g11692 ( 
.A(n_11645),
.B(n_11487),
.Y(n_11692)
);

OR2x2_ASAP7_75t_L g11693 ( 
.A(n_11538),
.B(n_11406),
.Y(n_11693)
);

NAND2xp5_ASAP7_75t_L g11694 ( 
.A(n_11563),
.B(n_11526),
.Y(n_11694)
);

INVx2_ASAP7_75t_L g11695 ( 
.A(n_11559),
.Y(n_11695)
);

INVx1_ASAP7_75t_L g11696 ( 
.A(n_11601),
.Y(n_11696)
);

AND2x2_ASAP7_75t_L g11697 ( 
.A(n_11560),
.B(n_11494),
.Y(n_11697)
);

NOR2x1p5_ASAP7_75t_L g11698 ( 
.A(n_11615),
.B(n_11505),
.Y(n_11698)
);

INVx2_ASAP7_75t_L g11699 ( 
.A(n_11562),
.Y(n_11699)
);

NOR2x1_ASAP7_75t_L g11700 ( 
.A(n_11586),
.B(n_11491),
.Y(n_11700)
);

INVxp67_ASAP7_75t_SL g11701 ( 
.A(n_11629),
.Y(n_11701)
);

OAI21xp33_ASAP7_75t_L g11702 ( 
.A1(n_11550),
.A2(n_11515),
.B(n_11458),
.Y(n_11702)
);

AND2x2_ASAP7_75t_L g11703 ( 
.A(n_11537),
.B(n_11539),
.Y(n_11703)
);

NAND2x1_ASAP7_75t_L g11704 ( 
.A(n_11641),
.B(n_11519),
.Y(n_11704)
);

INVx2_ASAP7_75t_L g11705 ( 
.A(n_11612),
.Y(n_11705)
);

NAND2xp5_ASAP7_75t_L g11706 ( 
.A(n_11571),
.B(n_11466),
.Y(n_11706)
);

INVx2_ASAP7_75t_L g11707 ( 
.A(n_11640),
.Y(n_11707)
);

INVx1_ASAP7_75t_SL g11708 ( 
.A(n_11555),
.Y(n_11708)
);

INVx2_ASAP7_75t_L g11709 ( 
.A(n_11610),
.Y(n_11709)
);

AND2x2_ASAP7_75t_L g11710 ( 
.A(n_11553),
.B(n_11516),
.Y(n_11710)
);

INVx1_ASAP7_75t_L g11711 ( 
.A(n_11585),
.Y(n_11711)
);

INVx1_ASAP7_75t_L g11712 ( 
.A(n_11600),
.Y(n_11712)
);

HB1xp67_ASAP7_75t_L g11713 ( 
.A(n_11575),
.Y(n_11713)
);

AND2x2_ASAP7_75t_L g11714 ( 
.A(n_11536),
.B(n_11527),
.Y(n_11714)
);

NOR2xp33_ASAP7_75t_L g11715 ( 
.A(n_11588),
.B(n_11508),
.Y(n_11715)
);

AND2x2_ASAP7_75t_L g11716 ( 
.A(n_11548),
.B(n_11488),
.Y(n_11716)
);

INVx2_ASAP7_75t_L g11717 ( 
.A(n_11636),
.Y(n_11717)
);

OR2x2_ASAP7_75t_L g11718 ( 
.A(n_11547),
.B(n_1705),
.Y(n_11718)
);

AND2x2_ASAP7_75t_L g11719 ( 
.A(n_11570),
.B(n_1706),
.Y(n_11719)
);

INVxp67_ASAP7_75t_SL g11720 ( 
.A(n_11652),
.Y(n_11720)
);

INVx1_ASAP7_75t_L g11721 ( 
.A(n_11631),
.Y(n_11721)
);

AND2x2_ASAP7_75t_L g11722 ( 
.A(n_11568),
.B(n_11575),
.Y(n_11722)
);

AND2x2_ASAP7_75t_L g11723 ( 
.A(n_11544),
.B(n_1706),
.Y(n_11723)
);

INVxp67_ASAP7_75t_L g11724 ( 
.A(n_11661),
.Y(n_11724)
);

INVx1_ASAP7_75t_L g11725 ( 
.A(n_11597),
.Y(n_11725)
);

INVx1_ASAP7_75t_L g11726 ( 
.A(n_11573),
.Y(n_11726)
);

INVx1_ASAP7_75t_L g11727 ( 
.A(n_11541),
.Y(n_11727)
);

AND2x2_ASAP7_75t_L g11728 ( 
.A(n_11561),
.B(n_1707),
.Y(n_11728)
);

INVx1_ASAP7_75t_L g11729 ( 
.A(n_11542),
.Y(n_11729)
);

INVx1_ASAP7_75t_L g11730 ( 
.A(n_11557),
.Y(n_11730)
);

INVx1_ASAP7_75t_L g11731 ( 
.A(n_11605),
.Y(n_11731)
);

OR2x6_ASAP7_75t_L g11732 ( 
.A(n_11567),
.B(n_1707),
.Y(n_11732)
);

INVxp67_ASAP7_75t_SL g11733 ( 
.A(n_11551),
.Y(n_11733)
);

AND2x2_ASAP7_75t_L g11734 ( 
.A(n_11564),
.B(n_1709),
.Y(n_11734)
);

INVx1_ASAP7_75t_L g11735 ( 
.A(n_11558),
.Y(n_11735)
);

NAND2xp5_ASAP7_75t_L g11736 ( 
.A(n_11580),
.B(n_1709),
.Y(n_11736)
);

HB1xp67_ASAP7_75t_L g11737 ( 
.A(n_11613),
.Y(n_11737)
);

AND2x2_ASAP7_75t_L g11738 ( 
.A(n_11583),
.B(n_1710),
.Y(n_11738)
);

AND2x2_ASAP7_75t_L g11739 ( 
.A(n_11584),
.B(n_1711),
.Y(n_11739)
);

NAND2xp5_ASAP7_75t_L g11740 ( 
.A(n_11604),
.B(n_11594),
.Y(n_11740)
);

INVxp67_ASAP7_75t_L g11741 ( 
.A(n_11658),
.Y(n_11741)
);

XNOR2x2_ASAP7_75t_L g11742 ( 
.A(n_11649),
.B(n_1712),
.Y(n_11742)
);

INVx1_ASAP7_75t_L g11743 ( 
.A(n_11642),
.Y(n_11743)
);

AND2x2_ASAP7_75t_L g11744 ( 
.A(n_11595),
.B(n_1712),
.Y(n_11744)
);

INVx1_ASAP7_75t_L g11745 ( 
.A(n_11656),
.Y(n_11745)
);

INVx1_ASAP7_75t_L g11746 ( 
.A(n_11614),
.Y(n_11746)
);

INVx1_ASAP7_75t_L g11747 ( 
.A(n_11660),
.Y(n_11747)
);

INVx1_ASAP7_75t_L g11748 ( 
.A(n_11663),
.Y(n_11748)
);

NAND2xp5_ASAP7_75t_L g11749 ( 
.A(n_11633),
.B(n_11634),
.Y(n_11749)
);

INVx1_ASAP7_75t_L g11750 ( 
.A(n_11664),
.Y(n_11750)
);

INVx1_ASAP7_75t_L g11751 ( 
.A(n_11635),
.Y(n_11751)
);

OR2x2_ASAP7_75t_L g11752 ( 
.A(n_11578),
.B(n_1713),
.Y(n_11752)
);

INVx1_ASAP7_75t_L g11753 ( 
.A(n_11627),
.Y(n_11753)
);

INVx1_ASAP7_75t_L g11754 ( 
.A(n_11576),
.Y(n_11754)
);

NOR2x1_ASAP7_75t_L g11755 ( 
.A(n_11651),
.B(n_1713),
.Y(n_11755)
);

INVx1_ASAP7_75t_L g11756 ( 
.A(n_11582),
.Y(n_11756)
);

NAND2xp5_ASAP7_75t_L g11757 ( 
.A(n_11623),
.B(n_1714),
.Y(n_11757)
);

BUFx3_ASAP7_75t_L g11758 ( 
.A(n_11587),
.Y(n_11758)
);

NAND2xp5_ASAP7_75t_L g11759 ( 
.A(n_11591),
.B(n_11657),
.Y(n_11759)
);

AND2x2_ASAP7_75t_L g11760 ( 
.A(n_11593),
.B(n_1715),
.Y(n_11760)
);

INVx1_ASAP7_75t_L g11761 ( 
.A(n_11599),
.Y(n_11761)
);

NOR2x1_ASAP7_75t_L g11762 ( 
.A(n_11654),
.B(n_11644),
.Y(n_11762)
);

NAND2x1_ASAP7_75t_L g11763 ( 
.A(n_11638),
.B(n_1715),
.Y(n_11763)
);

AND2x4_ASAP7_75t_L g11764 ( 
.A(n_11622),
.B(n_1717),
.Y(n_11764)
);

INVxp67_ASAP7_75t_L g11765 ( 
.A(n_11659),
.Y(n_11765)
);

AND2x2_ASAP7_75t_L g11766 ( 
.A(n_11643),
.B(n_1718),
.Y(n_11766)
);

AND2x2_ASAP7_75t_L g11767 ( 
.A(n_11665),
.B(n_1718),
.Y(n_11767)
);

AND3x2_ASAP7_75t_L g11768 ( 
.A(n_11648),
.B(n_1719),
.C(n_1720),
.Y(n_11768)
);

INVx2_ASAP7_75t_L g11769 ( 
.A(n_11616),
.Y(n_11769)
);

INVx1_ASAP7_75t_L g11770 ( 
.A(n_11602),
.Y(n_11770)
);

OR2x2_ASAP7_75t_L g11771 ( 
.A(n_11592),
.B(n_1719),
.Y(n_11771)
);

AND2x2_ASAP7_75t_L g11772 ( 
.A(n_11554),
.B(n_1720),
.Y(n_11772)
);

AND2x2_ASAP7_75t_L g11773 ( 
.A(n_11655),
.B(n_1721),
.Y(n_11773)
);

NAND2xp5_ASAP7_75t_L g11774 ( 
.A(n_11639),
.B(n_11609),
.Y(n_11774)
);

INVx1_ASAP7_75t_L g11775 ( 
.A(n_11598),
.Y(n_11775)
);

AND2x2_ASAP7_75t_L g11776 ( 
.A(n_11617),
.B(n_1722),
.Y(n_11776)
);

INVx2_ASAP7_75t_L g11777 ( 
.A(n_11626),
.Y(n_11777)
);

OR2x2_ASAP7_75t_L g11778 ( 
.A(n_11611),
.B(n_1722),
.Y(n_11778)
);

AND2x4_ASAP7_75t_L g11779 ( 
.A(n_11646),
.B(n_1723),
.Y(n_11779)
);

INVx1_ASAP7_75t_L g11780 ( 
.A(n_11679),
.Y(n_11780)
);

OR2x2_ASAP7_75t_L g11781 ( 
.A(n_11671),
.B(n_11589),
.Y(n_11781)
);

INVx1_ASAP7_75t_SL g11782 ( 
.A(n_11667),
.Y(n_11782)
);

NAND2xp5_ASAP7_75t_L g11783 ( 
.A(n_11768),
.B(n_11620),
.Y(n_11783)
);

AOI22xp5_ASAP7_75t_L g11784 ( 
.A1(n_11700),
.A2(n_11650),
.B1(n_11647),
.B2(n_11653),
.Y(n_11784)
);

OR2x2_ASAP7_75t_L g11785 ( 
.A(n_11759),
.B(n_11596),
.Y(n_11785)
);

INVx1_ASAP7_75t_L g11786 ( 
.A(n_11737),
.Y(n_11786)
);

INVx2_ASAP7_75t_L g11787 ( 
.A(n_11676),
.Y(n_11787)
);

NAND2xp5_ASAP7_75t_L g11788 ( 
.A(n_11703),
.B(n_11662),
.Y(n_11788)
);

INVx1_ASAP7_75t_SL g11789 ( 
.A(n_11684),
.Y(n_11789)
);

AND2x2_ASAP7_75t_L g11790 ( 
.A(n_11722),
.B(n_11618),
.Y(n_11790)
);

OR2x2_ASAP7_75t_L g11791 ( 
.A(n_11674),
.B(n_1723),
.Y(n_11791)
);

INVx1_ASAP7_75t_L g11792 ( 
.A(n_11713),
.Y(n_11792)
);

INVx2_ASAP7_75t_SL g11793 ( 
.A(n_11763),
.Y(n_11793)
);

AND2x2_ASAP7_75t_L g11794 ( 
.A(n_11683),
.B(n_1724),
.Y(n_11794)
);

AOI32xp33_ASAP7_75t_L g11795 ( 
.A1(n_11715),
.A2(n_1727),
.A3(n_1724),
.B1(n_1725),
.B2(n_1728),
.Y(n_11795)
);

OAI322xp33_ASAP7_75t_L g11796 ( 
.A1(n_11694),
.A2(n_1731),
.A3(n_1730),
.B1(n_1728),
.B2(n_1725),
.C1(n_1727),
.C2(n_1729),
.Y(n_11796)
);

INVx1_ASAP7_75t_L g11797 ( 
.A(n_11744),
.Y(n_11797)
);

HB1xp67_ASAP7_75t_L g11798 ( 
.A(n_11732),
.Y(n_11798)
);

INVxp33_ASAP7_75t_L g11799 ( 
.A(n_11755),
.Y(n_11799)
);

O2A1O1Ixp33_ASAP7_75t_L g11800 ( 
.A1(n_11686),
.A2(n_1732),
.B(n_1730),
.C(n_1731),
.Y(n_11800)
);

OAI322xp33_ASAP7_75t_L g11801 ( 
.A1(n_11701),
.A2(n_1738),
.A3(n_1737),
.B1(n_1735),
.B2(n_1733),
.C1(n_1734),
.C2(n_1736),
.Y(n_11801)
);

OAI33xp33_ASAP7_75t_L g11802 ( 
.A1(n_11668),
.A2(n_2801),
.A3(n_2797),
.B1(n_2802),
.B2(n_2798),
.B3(n_2796),
.Y(n_11802)
);

OR2x2_ASAP7_75t_L g11803 ( 
.A(n_11666),
.B(n_1733),
.Y(n_11803)
);

NAND2x2_ASAP7_75t_L g11804 ( 
.A(n_11698),
.B(n_1735),
.Y(n_11804)
);

BUFx2_ASAP7_75t_L g11805 ( 
.A(n_11732),
.Y(n_11805)
);

INVx2_ASAP7_75t_L g11806 ( 
.A(n_11705),
.Y(n_11806)
);

INVx1_ASAP7_75t_L g11807 ( 
.A(n_11728),
.Y(n_11807)
);

OR2x2_ASAP7_75t_L g11808 ( 
.A(n_11771),
.B(n_1734),
.Y(n_11808)
);

NAND2xp5_ASAP7_75t_L g11809 ( 
.A(n_11711),
.B(n_1736),
.Y(n_11809)
);

INVx2_ASAP7_75t_L g11810 ( 
.A(n_11778),
.Y(n_11810)
);

INVxp67_ASAP7_75t_SL g11811 ( 
.A(n_11692),
.Y(n_11811)
);

AOI22xp33_ASAP7_75t_L g11812 ( 
.A1(n_11702),
.A2(n_1739),
.B1(n_1737),
.B2(n_1738),
.Y(n_11812)
);

INVx1_ASAP7_75t_L g11813 ( 
.A(n_11734),
.Y(n_11813)
);

INVxp67_ASAP7_75t_SL g11814 ( 
.A(n_11742),
.Y(n_11814)
);

OAI22xp5_ASAP7_75t_L g11815 ( 
.A1(n_11708),
.A2(n_1741),
.B1(n_1739),
.B2(n_1740),
.Y(n_11815)
);

INVx1_ASAP7_75t_L g11816 ( 
.A(n_11723),
.Y(n_11816)
);

NOR4xp25_ASAP7_75t_L g11817 ( 
.A(n_11669),
.B(n_1742),
.C(n_1740),
.D(n_1741),
.Y(n_11817)
);

OAI32xp33_ASAP7_75t_L g11818 ( 
.A1(n_11678),
.A2(n_1744),
.A3(n_1747),
.B1(n_1743),
.B2(n_1745),
.Y(n_11818)
);

AOI22xp33_ASAP7_75t_SL g11819 ( 
.A1(n_11720),
.A2(n_1744),
.B1(n_1742),
.B2(n_1743),
.Y(n_11819)
);

AND2x2_ASAP7_75t_L g11820 ( 
.A(n_11738),
.B(n_1745),
.Y(n_11820)
);

NAND2xp5_ASAP7_75t_L g11821 ( 
.A(n_11714),
.B(n_1747),
.Y(n_11821)
);

NAND2x1p5_ASAP7_75t_L g11822 ( 
.A(n_11673),
.B(n_2794),
.Y(n_11822)
);

NAND2xp33_ASAP7_75t_L g11823 ( 
.A(n_11696),
.B(n_1748),
.Y(n_11823)
);

OAI32xp33_ASAP7_75t_L g11824 ( 
.A1(n_11672),
.A2(n_1750),
.A3(n_1752),
.B1(n_1749),
.B2(n_1751),
.Y(n_11824)
);

INVx1_ASAP7_75t_L g11825 ( 
.A(n_11719),
.Y(n_11825)
);

BUFx3_ASAP7_75t_L g11826 ( 
.A(n_11758),
.Y(n_11826)
);

NOR2xp33_ASAP7_75t_L g11827 ( 
.A(n_11746),
.B(n_1748),
.Y(n_11827)
);

AOI22xp5_ASAP7_75t_L g11828 ( 
.A1(n_11724),
.A2(n_1751),
.B1(n_1749),
.B2(n_1750),
.Y(n_11828)
);

OA222x2_ASAP7_75t_L g11829 ( 
.A1(n_11693),
.A2(n_1755),
.B1(n_1757),
.B2(n_1758),
.C1(n_1754),
.C2(n_1756),
.Y(n_11829)
);

AND2x4_ASAP7_75t_L g11830 ( 
.A(n_11681),
.B(n_1753),
.Y(n_11830)
);

AO221x1_ASAP7_75t_L g11831 ( 
.A1(n_11765),
.A2(n_1756),
.B1(n_1754),
.B2(n_1755),
.C(n_1757),
.Y(n_11831)
);

INVx1_ASAP7_75t_L g11832 ( 
.A(n_11740),
.Y(n_11832)
);

OR2x2_ASAP7_75t_L g11833 ( 
.A(n_11706),
.B(n_1758),
.Y(n_11833)
);

OAI32xp33_ASAP7_75t_L g11834 ( 
.A1(n_11688),
.A2(n_1761),
.A3(n_1763),
.B1(n_1760),
.B2(n_1762),
.Y(n_11834)
);

BUFx2_ASAP7_75t_SL g11835 ( 
.A(n_11709),
.Y(n_11835)
);

INVx2_ASAP7_75t_L g11836 ( 
.A(n_11764),
.Y(n_11836)
);

OR2x2_ASAP7_75t_L g11837 ( 
.A(n_11752),
.B(n_1759),
.Y(n_11837)
);

INVx1_ASAP7_75t_L g11838 ( 
.A(n_11739),
.Y(n_11838)
);

OAI32xp33_ASAP7_75t_L g11839 ( 
.A1(n_11687),
.A2(n_1762),
.A3(n_1764),
.B1(n_1761),
.B2(n_1763),
.Y(n_11839)
);

NAND2xp5_ASAP7_75t_SL g11840 ( 
.A(n_11682),
.B(n_1759),
.Y(n_11840)
);

NOR2xp33_ASAP7_75t_L g11841 ( 
.A(n_11743),
.B(n_1764),
.Y(n_11841)
);

AOI211xp5_ASAP7_75t_L g11842 ( 
.A1(n_11726),
.A2(n_2797),
.B(n_2798),
.C(n_2796),
.Y(n_11842)
);

NOR2xp33_ASAP7_75t_L g11843 ( 
.A(n_11670),
.B(n_1765),
.Y(n_11843)
);

AND2x2_ASAP7_75t_L g11844 ( 
.A(n_11710),
.B(n_1765),
.Y(n_11844)
);

NAND2xp5_ASAP7_75t_L g11845 ( 
.A(n_11677),
.B(n_1766),
.Y(n_11845)
);

NAND2xp5_ASAP7_75t_L g11846 ( 
.A(n_11680),
.B(n_1766),
.Y(n_11846)
);

NAND2xp5_ASAP7_75t_L g11847 ( 
.A(n_11685),
.B(n_11689),
.Y(n_11847)
);

INVxp67_ASAP7_75t_L g11848 ( 
.A(n_11716),
.Y(n_11848)
);

NAND2xp5_ASAP7_75t_L g11849 ( 
.A(n_11691),
.B(n_1767),
.Y(n_11849)
);

NAND2xp5_ASAP7_75t_L g11850 ( 
.A(n_11772),
.B(n_1768),
.Y(n_11850)
);

A2O1A1Ixp33_ASAP7_75t_L g11851 ( 
.A1(n_11733),
.A2(n_1777),
.B(n_1786),
.C(n_1769),
.Y(n_11851)
);

INVx1_ASAP7_75t_L g11852 ( 
.A(n_11760),
.Y(n_11852)
);

NAND2xp5_ASAP7_75t_L g11853 ( 
.A(n_11745),
.B(n_1770),
.Y(n_11853)
);

NAND4xp25_ASAP7_75t_L g11854 ( 
.A(n_11774),
.B(n_1772),
.C(n_1770),
.D(n_1771),
.Y(n_11854)
);

AOI22xp5_ASAP7_75t_L g11855 ( 
.A1(n_11675),
.A2(n_1774),
.B1(n_1771),
.B2(n_1773),
.Y(n_11855)
);

INVx1_ASAP7_75t_L g11856 ( 
.A(n_11766),
.Y(n_11856)
);

INVx2_ASAP7_75t_SL g11857 ( 
.A(n_11779),
.Y(n_11857)
);

NAND2xp5_ASAP7_75t_L g11858 ( 
.A(n_11747),
.B(n_11748),
.Y(n_11858)
);

AOI22xp5_ASAP7_75t_L g11859 ( 
.A1(n_11695),
.A2(n_1776),
.B1(n_1774),
.B2(n_1775),
.Y(n_11859)
);

INVx1_ASAP7_75t_L g11860 ( 
.A(n_11718),
.Y(n_11860)
);

INVx1_ASAP7_75t_L g11861 ( 
.A(n_11757),
.Y(n_11861)
);

INVx1_ASAP7_75t_L g11862 ( 
.A(n_11690),
.Y(n_11862)
);

NAND2xp5_ASAP7_75t_L g11863 ( 
.A(n_11750),
.B(n_11725),
.Y(n_11863)
);

OR2x2_ASAP7_75t_L g11864 ( 
.A(n_11707),
.B(n_11736),
.Y(n_11864)
);

AND2x2_ASAP7_75t_L g11865 ( 
.A(n_11697),
.B(n_1776),
.Y(n_11865)
);

NOR2xp33_ASAP7_75t_L g11866 ( 
.A(n_11731),
.B(n_1778),
.Y(n_11866)
);

INVx1_ASAP7_75t_SL g11867 ( 
.A(n_11776),
.Y(n_11867)
);

INVx2_ASAP7_75t_L g11868 ( 
.A(n_11699),
.Y(n_11868)
);

AND2x4_ASAP7_75t_L g11869 ( 
.A(n_11717),
.B(n_1778),
.Y(n_11869)
);

NOR2x1p5_ASAP7_75t_L g11870 ( 
.A(n_11704),
.B(n_2794),
.Y(n_11870)
);

AOI22xp5_ASAP7_75t_L g11871 ( 
.A1(n_11741),
.A2(n_1781),
.B1(n_1779),
.B2(n_1780),
.Y(n_11871)
);

AND2x4_ASAP7_75t_L g11872 ( 
.A(n_11727),
.B(n_1779),
.Y(n_11872)
);

AND2x2_ASAP7_75t_L g11873 ( 
.A(n_11721),
.B(n_1780),
.Y(n_11873)
);

AOI32xp33_ASAP7_75t_L g11874 ( 
.A1(n_11762),
.A2(n_1783),
.A3(n_1781),
.B1(n_1782),
.B2(n_1785),
.Y(n_11874)
);

INVx1_ASAP7_75t_L g11875 ( 
.A(n_11773),
.Y(n_11875)
);

INVx1_ASAP7_75t_L g11876 ( 
.A(n_11729),
.Y(n_11876)
);

INVx1_ASAP7_75t_L g11877 ( 
.A(n_11730),
.Y(n_11877)
);

O2A1O1Ixp5_ASAP7_75t_R g11878 ( 
.A1(n_11749),
.A2(n_11753),
.B(n_11751),
.C(n_11735),
.Y(n_11878)
);

INVx1_ASAP7_75t_L g11879 ( 
.A(n_11767),
.Y(n_11879)
);

INVx2_ASAP7_75t_L g11880 ( 
.A(n_11777),
.Y(n_11880)
);

OA222x2_ASAP7_75t_L g11881 ( 
.A1(n_11754),
.A2(n_1785),
.B1(n_1787),
.B2(n_1788),
.C1(n_1783),
.C2(n_1786),
.Y(n_11881)
);

OR2x2_ASAP7_75t_L g11882 ( 
.A(n_11769),
.B(n_1782),
.Y(n_11882)
);

INVx1_ASAP7_75t_L g11883 ( 
.A(n_11756),
.Y(n_11883)
);

OAI21xp5_ASAP7_75t_SL g11884 ( 
.A1(n_11770),
.A2(n_1787),
.B(n_1788),
.Y(n_11884)
);

NAND2xp5_ASAP7_75t_L g11885 ( 
.A(n_11712),
.B(n_1789),
.Y(n_11885)
);

AND2x2_ASAP7_75t_L g11886 ( 
.A(n_11775),
.B(n_1790),
.Y(n_11886)
);

INVxp67_ASAP7_75t_L g11887 ( 
.A(n_11761),
.Y(n_11887)
);

NAND2xp5_ASAP7_75t_L g11888 ( 
.A(n_11768),
.B(n_1790),
.Y(n_11888)
);

INVx1_ASAP7_75t_L g11889 ( 
.A(n_11679),
.Y(n_11889)
);

INVx1_ASAP7_75t_L g11890 ( 
.A(n_11679),
.Y(n_11890)
);

INVx2_ASAP7_75t_L g11891 ( 
.A(n_11667),
.Y(n_11891)
);

INVx1_ASAP7_75t_L g11892 ( 
.A(n_11679),
.Y(n_11892)
);

OR2x2_ASAP7_75t_L g11893 ( 
.A(n_11671),
.B(n_1791),
.Y(n_11893)
);

OR2x2_ASAP7_75t_L g11894 ( 
.A(n_11671),
.B(n_1791),
.Y(n_11894)
);

NAND2xp5_ASAP7_75t_L g11895 ( 
.A(n_11768),
.B(n_1792),
.Y(n_11895)
);

OAI222xp33_ASAP7_75t_L g11896 ( 
.A1(n_11700),
.A2(n_2792),
.B1(n_2790),
.B2(n_2793),
.C1(n_2791),
.C2(n_2789),
.Y(n_11896)
);

NAND2xp5_ASAP7_75t_L g11897 ( 
.A(n_11768),
.B(n_1792),
.Y(n_11897)
);

AOI211xp5_ASAP7_75t_L g11898 ( 
.A1(n_11702),
.A2(n_2792),
.B(n_2795),
.C(n_2791),
.Y(n_11898)
);

NOR2xp33_ASAP7_75t_L g11899 ( 
.A(n_11667),
.B(n_1793),
.Y(n_11899)
);

O2A1O1Ixp33_ASAP7_75t_L g11900 ( 
.A1(n_11686),
.A2(n_1795),
.B(n_1793),
.C(n_1794),
.Y(n_11900)
);

AND2x2_ASAP7_75t_SL g11901 ( 
.A(n_11679),
.B(n_1794),
.Y(n_11901)
);

AND2x4_ASAP7_75t_L g11902 ( 
.A(n_11679),
.B(n_1796),
.Y(n_11902)
);

INVx1_ASAP7_75t_L g11903 ( 
.A(n_11679),
.Y(n_11903)
);

INVx1_ASAP7_75t_SL g11904 ( 
.A(n_11679),
.Y(n_11904)
);

INVx1_ASAP7_75t_L g11905 ( 
.A(n_11798),
.Y(n_11905)
);

INVx2_ASAP7_75t_L g11906 ( 
.A(n_11793),
.Y(n_11906)
);

INVx2_ASAP7_75t_L g11907 ( 
.A(n_11901),
.Y(n_11907)
);

XNOR2x1_ASAP7_75t_L g11908 ( 
.A(n_11904),
.B(n_2808),
.Y(n_11908)
);

INVxp67_ASAP7_75t_L g11909 ( 
.A(n_11835),
.Y(n_11909)
);

INVx2_ASAP7_75t_L g11910 ( 
.A(n_11870),
.Y(n_11910)
);

INVx1_ASAP7_75t_L g11911 ( 
.A(n_11805),
.Y(n_11911)
);

INVx2_ASAP7_75t_SL g11912 ( 
.A(n_11902),
.Y(n_11912)
);

AND2x2_ASAP7_75t_L g11913 ( 
.A(n_11789),
.B(n_1796),
.Y(n_11913)
);

INVx2_ASAP7_75t_SL g11914 ( 
.A(n_11902),
.Y(n_11914)
);

INVx1_ASAP7_75t_L g11915 ( 
.A(n_11780),
.Y(n_11915)
);

OR2x2_ASAP7_75t_L g11916 ( 
.A(n_11782),
.B(n_1797),
.Y(n_11916)
);

INVx1_ASAP7_75t_L g11917 ( 
.A(n_11889),
.Y(n_11917)
);

XOR2x2_ASAP7_75t_L g11918 ( 
.A(n_11781),
.B(n_1797),
.Y(n_11918)
);

XNOR2x1_ASAP7_75t_L g11919 ( 
.A(n_11785),
.B(n_2811),
.Y(n_11919)
);

CKINVDCx8_ASAP7_75t_R g11920 ( 
.A(n_11830),
.Y(n_11920)
);

XOR2x2_ASAP7_75t_L g11921 ( 
.A(n_11788),
.B(n_1798),
.Y(n_11921)
);

INVx1_ASAP7_75t_L g11922 ( 
.A(n_11890),
.Y(n_11922)
);

OA22x2_ASAP7_75t_L g11923 ( 
.A1(n_11784),
.A2(n_1800),
.B1(n_1801),
.B2(n_1799),
.Y(n_11923)
);

INVxp67_ASAP7_75t_L g11924 ( 
.A(n_11899),
.Y(n_11924)
);

INVx1_ASAP7_75t_L g11925 ( 
.A(n_11892),
.Y(n_11925)
);

AND2x2_ASAP7_75t_SL g11926 ( 
.A(n_11903),
.B(n_1798),
.Y(n_11926)
);

XNOR2xp5_ASAP7_75t_L g11927 ( 
.A(n_11790),
.B(n_1802),
.Y(n_11927)
);

INVx1_ASAP7_75t_SL g11928 ( 
.A(n_11893),
.Y(n_11928)
);

NOR2x1_ASAP7_75t_R g11929 ( 
.A(n_11814),
.B(n_1801),
.Y(n_11929)
);

INVx2_ASAP7_75t_L g11930 ( 
.A(n_11822),
.Y(n_11930)
);

XNOR2xp5_ASAP7_75t_L g11931 ( 
.A(n_11792),
.B(n_1804),
.Y(n_11931)
);

INVx1_ASAP7_75t_L g11932 ( 
.A(n_11794),
.Y(n_11932)
);

INVx1_ASAP7_75t_L g11933 ( 
.A(n_11894),
.Y(n_11933)
);

HB1xp67_ASAP7_75t_L g11934 ( 
.A(n_11830),
.Y(n_11934)
);

AND2x2_ASAP7_75t_L g11935 ( 
.A(n_11891),
.B(n_1802),
.Y(n_11935)
);

INVx1_ASAP7_75t_L g11936 ( 
.A(n_11865),
.Y(n_11936)
);

INVx1_ASAP7_75t_L g11937 ( 
.A(n_11783),
.Y(n_11937)
);

AO22x2_ASAP7_75t_L g11938 ( 
.A1(n_11878),
.A2(n_1808),
.B1(n_1806),
.B2(n_1807),
.Y(n_11938)
);

INVx1_ASAP7_75t_SL g11939 ( 
.A(n_11888),
.Y(n_11939)
);

INVx1_ASAP7_75t_L g11940 ( 
.A(n_11820),
.Y(n_11940)
);

XOR2x2_ASAP7_75t_L g11941 ( 
.A(n_11826),
.B(n_1806),
.Y(n_11941)
);

INVx2_ASAP7_75t_L g11942 ( 
.A(n_11808),
.Y(n_11942)
);

XOR2x2_ASAP7_75t_L g11943 ( 
.A(n_11862),
.B(n_1807),
.Y(n_11943)
);

INVx1_ASAP7_75t_L g11944 ( 
.A(n_11844),
.Y(n_11944)
);

XOR2xp5_ASAP7_75t_L g11945 ( 
.A(n_11838),
.B(n_1808),
.Y(n_11945)
);

XNOR2xp5_ASAP7_75t_L g11946 ( 
.A(n_11797),
.B(n_1811),
.Y(n_11946)
);

NOR3xp33_ASAP7_75t_L g11947 ( 
.A(n_11847),
.B(n_11787),
.C(n_11858),
.Y(n_11947)
);

INVx1_ASAP7_75t_SL g11948 ( 
.A(n_11895),
.Y(n_11948)
);

INVx2_ASAP7_75t_L g11949 ( 
.A(n_11869),
.Y(n_11949)
);

INVx1_ASAP7_75t_L g11950 ( 
.A(n_11897),
.Y(n_11950)
);

INVx1_ASAP7_75t_L g11951 ( 
.A(n_11869),
.Y(n_11951)
);

INVxp33_ASAP7_75t_SL g11952 ( 
.A(n_11867),
.Y(n_11952)
);

INVx1_ASAP7_75t_L g11953 ( 
.A(n_11873),
.Y(n_11953)
);

INVx2_ASAP7_75t_L g11954 ( 
.A(n_11837),
.Y(n_11954)
);

INVxp67_ASAP7_75t_L g11955 ( 
.A(n_11827),
.Y(n_11955)
);

XOR2x2_ASAP7_75t_L g11956 ( 
.A(n_11807),
.B(n_11813),
.Y(n_11956)
);

XNOR2xp5_ASAP7_75t_L g11957 ( 
.A(n_11825),
.B(n_1811),
.Y(n_11957)
);

INVx1_ASAP7_75t_L g11958 ( 
.A(n_11786),
.Y(n_11958)
);

INVx1_ASAP7_75t_L g11959 ( 
.A(n_11804),
.Y(n_11959)
);

INVxp67_ASAP7_75t_L g11960 ( 
.A(n_11841),
.Y(n_11960)
);

INVx1_ASAP7_75t_L g11961 ( 
.A(n_11791),
.Y(n_11961)
);

XNOR2x2_ASAP7_75t_L g11962 ( 
.A(n_11829),
.B(n_1810),
.Y(n_11962)
);

INVx2_ASAP7_75t_L g11963 ( 
.A(n_11857),
.Y(n_11963)
);

XNOR2xp5_ASAP7_75t_L g11964 ( 
.A(n_11898),
.B(n_1812),
.Y(n_11964)
);

NAND2xp5_ASAP7_75t_L g11965 ( 
.A(n_11831),
.B(n_1810),
.Y(n_11965)
);

AND2x2_ASAP7_75t_L g11966 ( 
.A(n_11836),
.B(n_1812),
.Y(n_11966)
);

XNOR2xp5_ASAP7_75t_L g11967 ( 
.A(n_11854),
.B(n_1815),
.Y(n_11967)
);

INVx2_ASAP7_75t_L g11968 ( 
.A(n_11803),
.Y(n_11968)
);

CKINVDCx8_ASAP7_75t_R g11969 ( 
.A(n_11872),
.Y(n_11969)
);

INVx2_ASAP7_75t_L g11970 ( 
.A(n_11882),
.Y(n_11970)
);

OA22x2_ASAP7_75t_L g11971 ( 
.A1(n_11848),
.A2(n_1817),
.B1(n_1818),
.B2(n_1816),
.Y(n_11971)
);

INVxp67_ASAP7_75t_L g11972 ( 
.A(n_11843),
.Y(n_11972)
);

XNOR2xp5_ASAP7_75t_L g11973 ( 
.A(n_11816),
.B(n_1816),
.Y(n_11973)
);

XNOR2xp5_ASAP7_75t_L g11974 ( 
.A(n_11828),
.B(n_1818),
.Y(n_11974)
);

INVx1_ASAP7_75t_SL g11975 ( 
.A(n_11840),
.Y(n_11975)
);

NOR2x1_ASAP7_75t_L g11976 ( 
.A(n_11896),
.B(n_1813),
.Y(n_11976)
);

XNOR2x2_ASAP7_75t_L g11977 ( 
.A(n_11881),
.B(n_1813),
.Y(n_11977)
);

XNOR2xp5_ASAP7_75t_L g11978 ( 
.A(n_11856),
.B(n_1820),
.Y(n_11978)
);

INVx1_ASAP7_75t_L g11979 ( 
.A(n_11850),
.Y(n_11979)
);

NAND2xp5_ASAP7_75t_L g11980 ( 
.A(n_11817),
.B(n_1819),
.Y(n_11980)
);

INVx1_ASAP7_75t_SL g11981 ( 
.A(n_11833),
.Y(n_11981)
);

XOR2x2_ASAP7_75t_L g11982 ( 
.A(n_11821),
.B(n_1819),
.Y(n_11982)
);

HB1xp67_ASAP7_75t_L g11983 ( 
.A(n_11799),
.Y(n_11983)
);

INVx1_ASAP7_75t_L g11984 ( 
.A(n_11823),
.Y(n_11984)
);

INVxp67_ASAP7_75t_L g11985 ( 
.A(n_11866),
.Y(n_11985)
);

INVxp67_ASAP7_75t_L g11986 ( 
.A(n_11845),
.Y(n_11986)
);

INVx1_ASAP7_75t_SL g11987 ( 
.A(n_11886),
.Y(n_11987)
);

INVx1_ASAP7_75t_L g11988 ( 
.A(n_11846),
.Y(n_11988)
);

XNOR2x1_ASAP7_75t_L g11989 ( 
.A(n_11864),
.B(n_2813),
.Y(n_11989)
);

INVx2_ASAP7_75t_L g11990 ( 
.A(n_11806),
.Y(n_11990)
);

XOR2xp5_ASAP7_75t_L g11991 ( 
.A(n_11852),
.B(n_1820),
.Y(n_11991)
);

INVx2_ASAP7_75t_L g11992 ( 
.A(n_11810),
.Y(n_11992)
);

OA22x2_ASAP7_75t_L g11993 ( 
.A1(n_11879),
.A2(n_1823),
.B1(n_1824),
.B2(n_1822),
.Y(n_11993)
);

INVx1_ASAP7_75t_L g11994 ( 
.A(n_11849),
.Y(n_11994)
);

XNOR2xp5_ASAP7_75t_L g11995 ( 
.A(n_11842),
.B(n_1822),
.Y(n_11995)
);

XNOR2xp5_ASAP7_75t_L g11996 ( 
.A(n_11815),
.B(n_1824),
.Y(n_11996)
);

XNOR2xp5_ASAP7_75t_L g11997 ( 
.A(n_11875),
.B(n_1825),
.Y(n_11997)
);

CKINVDCx16_ASAP7_75t_R g11998 ( 
.A(n_11832),
.Y(n_11998)
);

HB1xp67_ASAP7_75t_L g11999 ( 
.A(n_11880),
.Y(n_11999)
);

BUFx3_ASAP7_75t_L g12000 ( 
.A(n_11868),
.Y(n_12000)
);

INVxp67_ASAP7_75t_L g12001 ( 
.A(n_11863),
.Y(n_12001)
);

NOR2xp33_ASAP7_75t_L g12002 ( 
.A(n_11884),
.B(n_1821),
.Y(n_12002)
);

INVx2_ASAP7_75t_L g12003 ( 
.A(n_11860),
.Y(n_12003)
);

XNOR2xp5_ASAP7_75t_L g12004 ( 
.A(n_11819),
.B(n_11855),
.Y(n_12004)
);

INVx1_ASAP7_75t_SL g12005 ( 
.A(n_11809),
.Y(n_12005)
);

XNOR2xp5_ASAP7_75t_L g12006 ( 
.A(n_11859),
.B(n_1825),
.Y(n_12006)
);

NOR2x1_ASAP7_75t_L g12007 ( 
.A(n_11801),
.B(n_1821),
.Y(n_12007)
);

XOR2x2_ASAP7_75t_L g12008 ( 
.A(n_11853),
.B(n_1826),
.Y(n_12008)
);

XOR2x2_ASAP7_75t_L g12009 ( 
.A(n_11812),
.B(n_1826),
.Y(n_12009)
);

INVx1_ASAP7_75t_L g12010 ( 
.A(n_11811),
.Y(n_12010)
);

XOR2x2_ASAP7_75t_L g12011 ( 
.A(n_11871),
.B(n_1828),
.Y(n_12011)
);

INVx1_ASAP7_75t_L g12012 ( 
.A(n_11885),
.Y(n_12012)
);

OAI22xp5_ASAP7_75t_L g12013 ( 
.A1(n_11887),
.A2(n_1831),
.B1(n_1829),
.B2(n_1830),
.Y(n_12013)
);

INVx2_ASAP7_75t_L g12014 ( 
.A(n_11876),
.Y(n_12014)
);

BUFx6f_ASAP7_75t_L g12015 ( 
.A(n_11877),
.Y(n_12015)
);

INVx1_ASAP7_75t_SL g12016 ( 
.A(n_11883),
.Y(n_12016)
);

INVx1_ASAP7_75t_L g12017 ( 
.A(n_11818),
.Y(n_12017)
);

INVx2_ASAP7_75t_SL g12018 ( 
.A(n_11861),
.Y(n_12018)
);

INVx1_ASAP7_75t_L g12019 ( 
.A(n_11800),
.Y(n_12019)
);

INVx2_ASAP7_75t_L g12020 ( 
.A(n_11824),
.Y(n_12020)
);

INVx2_ASAP7_75t_L g12021 ( 
.A(n_11834),
.Y(n_12021)
);

INVx1_ASAP7_75t_SL g12022 ( 
.A(n_11874),
.Y(n_12022)
);

BUFx3_ASAP7_75t_L g12023 ( 
.A(n_11795),
.Y(n_12023)
);

XNOR2xp5_ASAP7_75t_L g12024 ( 
.A(n_11796),
.B(n_1830),
.Y(n_12024)
);

INVx1_ASAP7_75t_SL g12025 ( 
.A(n_11839),
.Y(n_12025)
);

XOR2x2_ASAP7_75t_L g12026 ( 
.A(n_11900),
.B(n_1829),
.Y(n_12026)
);

NOR2xp33_ASAP7_75t_SL g12027 ( 
.A(n_11802),
.B(n_1833),
.Y(n_12027)
);

AOI22xp5_ASAP7_75t_L g12028 ( 
.A1(n_11851),
.A2(n_1835),
.B1(n_1833),
.B2(n_1834),
.Y(n_12028)
);

INVx1_ASAP7_75t_L g12029 ( 
.A(n_11798),
.Y(n_12029)
);

AND2x2_ASAP7_75t_L g12030 ( 
.A(n_11904),
.B(n_1834),
.Y(n_12030)
);

XOR2x2_ASAP7_75t_L g12031 ( 
.A(n_11904),
.B(n_1835),
.Y(n_12031)
);

INVx1_ASAP7_75t_L g12032 ( 
.A(n_11798),
.Y(n_12032)
);

XOR2x2_ASAP7_75t_L g12033 ( 
.A(n_11904),
.B(n_1836),
.Y(n_12033)
);

INVx1_ASAP7_75t_L g12034 ( 
.A(n_11798),
.Y(n_12034)
);

OA22x2_ASAP7_75t_L g12035 ( 
.A1(n_11793),
.A2(n_1838),
.B1(n_1839),
.B2(n_1837),
.Y(n_12035)
);

INVx1_ASAP7_75t_SL g12036 ( 
.A(n_11904),
.Y(n_12036)
);

INVxp67_ASAP7_75t_L g12037 ( 
.A(n_11835),
.Y(n_12037)
);

INVx1_ASAP7_75t_SL g12038 ( 
.A(n_11904),
.Y(n_12038)
);

INVx1_ASAP7_75t_SL g12039 ( 
.A(n_11904),
.Y(n_12039)
);

INVx2_ASAP7_75t_L g12040 ( 
.A(n_11793),
.Y(n_12040)
);

XOR2x2_ASAP7_75t_L g12041 ( 
.A(n_11904),
.B(n_1836),
.Y(n_12041)
);

INVx2_ASAP7_75t_SL g12042 ( 
.A(n_11793),
.Y(n_12042)
);

INVx1_ASAP7_75t_SL g12043 ( 
.A(n_11904),
.Y(n_12043)
);

INVx2_ASAP7_75t_L g12044 ( 
.A(n_11793),
.Y(n_12044)
);

INVx2_ASAP7_75t_L g12045 ( 
.A(n_11793),
.Y(n_12045)
);

INVx1_ASAP7_75t_L g12046 ( 
.A(n_11798),
.Y(n_12046)
);

INVx2_ASAP7_75t_L g12047 ( 
.A(n_11793),
.Y(n_12047)
);

INVx1_ASAP7_75t_L g12048 ( 
.A(n_11798),
.Y(n_12048)
);

XOR2x2_ASAP7_75t_L g12049 ( 
.A(n_11904),
.B(n_1838),
.Y(n_12049)
);

INVx2_ASAP7_75t_SL g12050 ( 
.A(n_11793),
.Y(n_12050)
);

INVx2_ASAP7_75t_SL g12051 ( 
.A(n_11793),
.Y(n_12051)
);

INVxp67_ASAP7_75t_L g12052 ( 
.A(n_11835),
.Y(n_12052)
);

INVx2_ASAP7_75t_SL g12053 ( 
.A(n_11793),
.Y(n_12053)
);

INVx1_ASAP7_75t_L g12054 ( 
.A(n_11934),
.Y(n_12054)
);

INVx1_ASAP7_75t_L g12055 ( 
.A(n_12035),
.Y(n_12055)
);

NAND2xp5_ASAP7_75t_SL g12056 ( 
.A(n_11998),
.B(n_1840),
.Y(n_12056)
);

OAI22xp5_ASAP7_75t_L g12057 ( 
.A1(n_12036),
.A2(n_1843),
.B1(n_1840),
.B2(n_1842),
.Y(n_12057)
);

OAI22xp5_ASAP7_75t_L g12058 ( 
.A1(n_12038),
.A2(n_1846),
.B1(n_1844),
.B2(n_1845),
.Y(n_12058)
);

INVx1_ASAP7_75t_L g12059 ( 
.A(n_11929),
.Y(n_12059)
);

INVx1_ASAP7_75t_L g12060 ( 
.A(n_11993),
.Y(n_12060)
);

NAND2xp5_ASAP7_75t_L g12061 ( 
.A(n_11912),
.B(n_1845),
.Y(n_12061)
);

OAI22xp5_ASAP7_75t_L g12062 ( 
.A1(n_12039),
.A2(n_1849),
.B1(n_1847),
.B2(n_1848),
.Y(n_12062)
);

NAND2xp5_ASAP7_75t_L g12063 ( 
.A(n_11914),
.B(n_1847),
.Y(n_12063)
);

AND2x2_ASAP7_75t_L g12064 ( 
.A(n_11913),
.B(n_1848),
.Y(n_12064)
);

AND2x2_ASAP7_75t_L g12065 ( 
.A(n_11906),
.B(n_1850),
.Y(n_12065)
);

AOI22xp33_ASAP7_75t_L g12066 ( 
.A1(n_11952),
.A2(n_1853),
.B1(n_1850),
.B2(n_1852),
.Y(n_12066)
);

AND2x2_ASAP7_75t_L g12067 ( 
.A(n_12040),
.B(n_1852),
.Y(n_12067)
);

AND2x2_ASAP7_75t_L g12068 ( 
.A(n_12044),
.B(n_1853),
.Y(n_12068)
);

INVx2_ASAP7_75t_L g12069 ( 
.A(n_12042),
.Y(n_12069)
);

INVx1_ASAP7_75t_SL g12070 ( 
.A(n_11962),
.Y(n_12070)
);

AOI22xp33_ASAP7_75t_L g12071 ( 
.A1(n_11911),
.A2(n_12029),
.B1(n_12032),
.B2(n_11905),
.Y(n_12071)
);

INVx1_ASAP7_75t_L g12072 ( 
.A(n_11971),
.Y(n_12072)
);

INVx1_ASAP7_75t_L g12073 ( 
.A(n_11977),
.Y(n_12073)
);

NAND2xp5_ASAP7_75t_L g12074 ( 
.A(n_12050),
.B(n_12051),
.Y(n_12074)
);

OAI22xp5_ASAP7_75t_L g12075 ( 
.A1(n_12043),
.A2(n_1858),
.B1(n_1855),
.B2(n_1856),
.Y(n_12075)
);

INVx1_ASAP7_75t_SL g12076 ( 
.A(n_11908),
.Y(n_12076)
);

INVx2_ASAP7_75t_SL g12077 ( 
.A(n_11949),
.Y(n_12077)
);

OR2x6_ASAP7_75t_L g12078 ( 
.A(n_12053),
.B(n_1855),
.Y(n_12078)
);

INVx4_ASAP7_75t_L g12079 ( 
.A(n_12015),
.Y(n_12079)
);

OR2x2_ASAP7_75t_L g12080 ( 
.A(n_11907),
.B(n_1856),
.Y(n_12080)
);

INVx2_ASAP7_75t_SL g12081 ( 
.A(n_11926),
.Y(n_12081)
);

NOR2xp33_ASAP7_75t_L g12082 ( 
.A(n_11920),
.B(n_1859),
.Y(n_12082)
);

CKINVDCx16_ASAP7_75t_R g12083 ( 
.A(n_12023),
.Y(n_12083)
);

INVx1_ASAP7_75t_L g12084 ( 
.A(n_11927),
.Y(n_12084)
);

AND2x2_ASAP7_75t_L g12085 ( 
.A(n_12045),
.B(n_1859),
.Y(n_12085)
);

NAND2xp5_ASAP7_75t_L g12086 ( 
.A(n_12047),
.B(n_11951),
.Y(n_12086)
);

AND2x2_ASAP7_75t_L g12087 ( 
.A(n_11963),
.B(n_1860),
.Y(n_12087)
);

INVx1_ASAP7_75t_L g12088 ( 
.A(n_11945),
.Y(n_12088)
);

NAND2xp33_ASAP7_75t_R g12089 ( 
.A(n_12030),
.B(n_11980),
.Y(n_12089)
);

NOR2xp33_ASAP7_75t_L g12090 ( 
.A(n_11909),
.B(n_1860),
.Y(n_12090)
);

INVx1_ASAP7_75t_SL g12091 ( 
.A(n_11916),
.Y(n_12091)
);

AND2x4_ASAP7_75t_L g12092 ( 
.A(n_11910),
.B(n_11930),
.Y(n_12092)
);

CKINVDCx16_ASAP7_75t_R g12093 ( 
.A(n_11976),
.Y(n_12093)
);

AND3x2_ASAP7_75t_L g12094 ( 
.A(n_12037),
.B(n_1865),
.C(n_1864),
.Y(n_12094)
);

INVx1_ASAP7_75t_L g12095 ( 
.A(n_11931),
.Y(n_12095)
);

INVx2_ASAP7_75t_L g12096 ( 
.A(n_11956),
.Y(n_12096)
);

INVx2_ASAP7_75t_L g12097 ( 
.A(n_11941),
.Y(n_12097)
);

AND2x2_ASAP7_75t_L g12098 ( 
.A(n_12052),
.B(n_1863),
.Y(n_12098)
);

INVx2_ASAP7_75t_L g12099 ( 
.A(n_12034),
.Y(n_12099)
);

AND2x2_ASAP7_75t_L g12100 ( 
.A(n_12046),
.B(n_1865),
.Y(n_12100)
);

NAND2xp5_ASAP7_75t_L g12101 ( 
.A(n_12048),
.B(n_1866),
.Y(n_12101)
);

INVx1_ASAP7_75t_L g12102 ( 
.A(n_11991),
.Y(n_12102)
);

INVx1_ASAP7_75t_SL g12103 ( 
.A(n_12031),
.Y(n_12103)
);

INVx1_ASAP7_75t_SL g12104 ( 
.A(n_12033),
.Y(n_12104)
);

INVxp67_ASAP7_75t_L g12105 ( 
.A(n_12027),
.Y(n_12105)
);

INVx2_ASAP7_75t_SL g12106 ( 
.A(n_12015),
.Y(n_12106)
);

AOI221xp5_ASAP7_75t_L g12107 ( 
.A1(n_11938),
.A2(n_1868),
.B1(n_1866),
.B2(n_1867),
.C(n_1869),
.Y(n_12107)
);

BUFx2_ASAP7_75t_L g12108 ( 
.A(n_11999),
.Y(n_12108)
);

INVx1_ASAP7_75t_L g12109 ( 
.A(n_11946),
.Y(n_12109)
);

INVx1_ASAP7_75t_L g12110 ( 
.A(n_11957),
.Y(n_12110)
);

INVx1_ASAP7_75t_SL g12111 ( 
.A(n_12041),
.Y(n_12111)
);

INVx3_ASAP7_75t_L g12112 ( 
.A(n_11969),
.Y(n_12112)
);

NAND2xp5_ASAP7_75t_L g12113 ( 
.A(n_11966),
.B(n_11935),
.Y(n_12113)
);

INVxp67_ASAP7_75t_L g12114 ( 
.A(n_11965),
.Y(n_12114)
);

INVx1_ASAP7_75t_L g12115 ( 
.A(n_11973),
.Y(n_12115)
);

NAND2xp5_ASAP7_75t_L g12116 ( 
.A(n_11959),
.B(n_1868),
.Y(n_12116)
);

INVx2_ASAP7_75t_SL g12117 ( 
.A(n_12000),
.Y(n_12117)
);

BUFx3_ASAP7_75t_L g12118 ( 
.A(n_11940),
.Y(n_12118)
);

INVx1_ASAP7_75t_L g12119 ( 
.A(n_11923),
.Y(n_12119)
);

NAND2xp5_ASAP7_75t_L g12120 ( 
.A(n_12025),
.B(n_1869),
.Y(n_12120)
);

HB1xp67_ASAP7_75t_L g12121 ( 
.A(n_12049),
.Y(n_12121)
);

AND2x2_ASAP7_75t_L g12122 ( 
.A(n_12021),
.B(n_1870),
.Y(n_12122)
);

AOI21xp5_ASAP7_75t_L g12123 ( 
.A1(n_11938),
.A2(n_1870),
.B(n_1871),
.Y(n_12123)
);

INVx1_ASAP7_75t_SL g12124 ( 
.A(n_11928),
.Y(n_12124)
);

NAND3xp33_ASAP7_75t_L g12125 ( 
.A(n_11947),
.B(n_1871),
.C(n_1872),
.Y(n_12125)
);

NOR2x1_ASAP7_75t_L g12126 ( 
.A(n_11989),
.B(n_1873),
.Y(n_12126)
);

INVx1_ASAP7_75t_SL g12127 ( 
.A(n_11918),
.Y(n_12127)
);

AND2x4_ASAP7_75t_L g12128 ( 
.A(n_11992),
.B(n_1873),
.Y(n_12128)
);

INVx1_ASAP7_75t_L g12129 ( 
.A(n_11978),
.Y(n_12129)
);

AND2x2_ASAP7_75t_L g12130 ( 
.A(n_12020),
.B(n_1874),
.Y(n_12130)
);

INVx2_ASAP7_75t_L g12131 ( 
.A(n_11943),
.Y(n_12131)
);

INVx2_ASAP7_75t_L g12132 ( 
.A(n_11944),
.Y(n_12132)
);

INVx1_ASAP7_75t_SL g12133 ( 
.A(n_11975),
.Y(n_12133)
);

NAND2x1_ASAP7_75t_SL g12134 ( 
.A(n_11983),
.B(n_1875),
.Y(n_12134)
);

OR2x2_ASAP7_75t_L g12135 ( 
.A(n_12022),
.B(n_1874),
.Y(n_12135)
);

HB1xp67_ASAP7_75t_L g12136 ( 
.A(n_11997),
.Y(n_12136)
);

OR2x2_ASAP7_75t_L g12137 ( 
.A(n_11939),
.B(n_1875),
.Y(n_12137)
);

INVx1_ASAP7_75t_L g12138 ( 
.A(n_11932),
.Y(n_12138)
);

INVx1_ASAP7_75t_L g12139 ( 
.A(n_11936),
.Y(n_12139)
);

NOR3xp33_ASAP7_75t_L g12140 ( 
.A(n_11937),
.B(n_12019),
.C(n_11950),
.Y(n_12140)
);

OA21x2_ASAP7_75t_L g12141 ( 
.A1(n_12017),
.A2(n_1878),
.B(n_1877),
.Y(n_12141)
);

AND2x2_ASAP7_75t_L g12142 ( 
.A(n_11984),
.B(n_1876),
.Y(n_12142)
);

AOI22xp33_ASAP7_75t_L g12143 ( 
.A1(n_11915),
.A2(n_1879),
.B1(n_1876),
.B2(n_1877),
.Y(n_12143)
);

INVx1_ASAP7_75t_L g12144 ( 
.A(n_11982),
.Y(n_12144)
);

OR2x2_ASAP7_75t_L g12145 ( 
.A(n_11948),
.B(n_1879),
.Y(n_12145)
);

INVx3_ASAP7_75t_L g12146 ( 
.A(n_12003),
.Y(n_12146)
);

OR2x6_ASAP7_75t_L g12147 ( 
.A(n_11954),
.B(n_1880),
.Y(n_12147)
);

BUFx2_ASAP7_75t_L g12148 ( 
.A(n_11933),
.Y(n_12148)
);

AND2x2_ASAP7_75t_L g12149 ( 
.A(n_11917),
.B(n_1880),
.Y(n_12149)
);

NAND2xp5_ASAP7_75t_L g12150 ( 
.A(n_11987),
.B(n_11922),
.Y(n_12150)
);

OR2x2_ASAP7_75t_L g12151 ( 
.A(n_11925),
.B(n_11953),
.Y(n_12151)
);

AND2x2_ASAP7_75t_L g12152 ( 
.A(n_11942),
.B(n_1881),
.Y(n_12152)
);

NAND2xp5_ASAP7_75t_L g12153 ( 
.A(n_12007),
.B(n_12024),
.Y(n_12153)
);

NAND2x1p5_ASAP7_75t_L g12154 ( 
.A(n_12016),
.B(n_1883),
.Y(n_12154)
);

AOI222xp33_ASAP7_75t_L g12155 ( 
.A1(n_12004),
.A2(n_1884),
.B1(n_1886),
.B2(n_1882),
.C1(n_1883),
.C2(n_1885),
.Y(n_12155)
);

NAND2xp5_ASAP7_75t_L g12156 ( 
.A(n_11958),
.B(n_1882),
.Y(n_12156)
);

AOI22xp5_ASAP7_75t_L g12157 ( 
.A1(n_12010),
.A2(n_2790),
.B1(n_2803),
.B2(n_2789),
.Y(n_12157)
);

INVx1_ASAP7_75t_L g12158 ( 
.A(n_11996),
.Y(n_12158)
);

NAND2xp5_ASAP7_75t_L g12159 ( 
.A(n_12002),
.B(n_1884),
.Y(n_12159)
);

INVx1_ASAP7_75t_L g12160 ( 
.A(n_12008),
.Y(n_12160)
);

AND2x2_ASAP7_75t_L g12161 ( 
.A(n_11970),
.B(n_1885),
.Y(n_12161)
);

INVx1_ASAP7_75t_SL g12162 ( 
.A(n_11919),
.Y(n_12162)
);

INVx1_ASAP7_75t_L g12163 ( 
.A(n_11967),
.Y(n_12163)
);

CKINVDCx16_ASAP7_75t_R g12164 ( 
.A(n_11981),
.Y(n_12164)
);

NOR2xp33_ASAP7_75t_L g12165 ( 
.A(n_11924),
.B(n_1886),
.Y(n_12165)
);

INVx2_ASAP7_75t_L g12166 ( 
.A(n_11968),
.Y(n_12166)
);

INVx1_ASAP7_75t_SL g12167 ( 
.A(n_11921),
.Y(n_12167)
);

INVxp67_ASAP7_75t_L g12168 ( 
.A(n_11995),
.Y(n_12168)
);

NAND3x1_ASAP7_75t_SL g12169 ( 
.A(n_12026),
.B(n_1896),
.C(n_1887),
.Y(n_12169)
);

OR2x2_ASAP7_75t_L g12170 ( 
.A(n_11990),
.B(n_1887),
.Y(n_12170)
);

NAND2xp5_ASAP7_75t_L g12171 ( 
.A(n_11961),
.B(n_1888),
.Y(n_12171)
);

AND2x2_ASAP7_75t_L g12172 ( 
.A(n_11955),
.B(n_1888),
.Y(n_12172)
);

INVx2_ASAP7_75t_L g12173 ( 
.A(n_12014),
.Y(n_12173)
);

INVx1_ASAP7_75t_L g12174 ( 
.A(n_11964),
.Y(n_12174)
);

AND2x2_ASAP7_75t_L g12175 ( 
.A(n_11960),
.B(n_11972),
.Y(n_12175)
);

INVx1_ASAP7_75t_L g12176 ( 
.A(n_11974),
.Y(n_12176)
);

INVx1_ASAP7_75t_SL g12177 ( 
.A(n_12011),
.Y(n_12177)
);

INVx1_ASAP7_75t_L g12178 ( 
.A(n_12006),
.Y(n_12178)
);

AND2x2_ASAP7_75t_L g12179 ( 
.A(n_11985),
.B(n_1889),
.Y(n_12179)
);

INVx1_ASAP7_75t_L g12180 ( 
.A(n_12013),
.Y(n_12180)
);

INVx2_ASAP7_75t_L g12181 ( 
.A(n_12018),
.Y(n_12181)
);

INVx2_ASAP7_75t_L g12182 ( 
.A(n_11979),
.Y(n_12182)
);

NAND2xp5_ASAP7_75t_L g12183 ( 
.A(n_12028),
.B(n_1889),
.Y(n_12183)
);

OAI22xp5_ASAP7_75t_L g12184 ( 
.A1(n_12001),
.A2(n_1893),
.B1(n_1890),
.B2(n_1892),
.Y(n_12184)
);

NAND2xp5_ASAP7_75t_L g12185 ( 
.A(n_12005),
.B(n_1892),
.Y(n_12185)
);

INVx1_ASAP7_75t_L g12186 ( 
.A(n_12009),
.Y(n_12186)
);

INVx2_ASAP7_75t_L g12187 ( 
.A(n_11988),
.Y(n_12187)
);

AND2x4_ASAP7_75t_L g12188 ( 
.A(n_11994),
.B(n_1893),
.Y(n_12188)
);

AND2x2_ASAP7_75t_L g12189 ( 
.A(n_11986),
.B(n_1894),
.Y(n_12189)
);

AOI222xp33_ASAP7_75t_L g12190 ( 
.A1(n_12012),
.A2(n_1898),
.B1(n_1900),
.B2(n_1895),
.C1(n_1897),
.C2(n_1899),
.Y(n_12190)
);

INVxp67_ASAP7_75t_L g12191 ( 
.A(n_11929),
.Y(n_12191)
);

AND2x4_ASAP7_75t_L g12192 ( 
.A(n_11912),
.B(n_1895),
.Y(n_12192)
);

INVx2_ASAP7_75t_L g12193 ( 
.A(n_11912),
.Y(n_12193)
);

INVx1_ASAP7_75t_L g12194 ( 
.A(n_12134),
.Y(n_12194)
);

OAI22xp5_ASAP7_75t_L g12195 ( 
.A1(n_12071),
.A2(n_12164),
.B1(n_12105),
.B2(n_12070),
.Y(n_12195)
);

OAI221xp5_ASAP7_75t_L g12196 ( 
.A1(n_12073),
.A2(n_2804),
.B1(n_2807),
.B2(n_2788),
.C(n_2787),
.Y(n_12196)
);

OAI21xp33_ASAP7_75t_L g12197 ( 
.A1(n_12074),
.A2(n_1897),
.B(n_1899),
.Y(n_12197)
);

AOI22xp33_ASAP7_75t_L g12198 ( 
.A1(n_12112),
.A2(n_1903),
.B1(n_1901),
.B2(n_1902),
.Y(n_12198)
);

INVx2_ASAP7_75t_L g12199 ( 
.A(n_12154),
.Y(n_12199)
);

INVx1_ASAP7_75t_L g12200 ( 
.A(n_12108),
.Y(n_12200)
);

OAI21xp33_ASAP7_75t_SL g12201 ( 
.A1(n_12081),
.A2(n_1901),
.B(n_1902),
.Y(n_12201)
);

INVx1_ASAP7_75t_L g12202 ( 
.A(n_12078),
.Y(n_12202)
);

INVx1_ASAP7_75t_L g12203 ( 
.A(n_12078),
.Y(n_12203)
);

HB1xp67_ASAP7_75t_L g12204 ( 
.A(n_12147),
.Y(n_12204)
);

INVxp67_ASAP7_75t_L g12205 ( 
.A(n_12082),
.Y(n_12205)
);

NAND2x1_ASAP7_75t_L g12206 ( 
.A(n_12079),
.B(n_1903),
.Y(n_12206)
);

OAI21xp5_ASAP7_75t_L g12207 ( 
.A1(n_12191),
.A2(n_1906),
.B(n_1905),
.Y(n_12207)
);

OR2x2_ASAP7_75t_L g12208 ( 
.A(n_12093),
.B(n_1904),
.Y(n_12208)
);

AOI31xp33_ASAP7_75t_L g12209 ( 
.A1(n_12076),
.A2(n_1913),
.A3(n_1921),
.B(n_1904),
.Y(n_12209)
);

OAI21xp5_ASAP7_75t_SL g12210 ( 
.A1(n_12133),
.A2(n_1905),
.B(n_1906),
.Y(n_12210)
);

AOI211xp5_ASAP7_75t_L g12211 ( 
.A1(n_12054),
.A2(n_1910),
.B(n_1907),
.C(n_1908),
.Y(n_12211)
);

NAND2xp5_ASAP7_75t_L g12212 ( 
.A(n_12094),
.B(n_1907),
.Y(n_12212)
);

INVx1_ASAP7_75t_L g12213 ( 
.A(n_12121),
.Y(n_12213)
);

INVx1_ASAP7_75t_L g12214 ( 
.A(n_12064),
.Y(n_12214)
);

OAI211xp5_ASAP7_75t_SL g12215 ( 
.A1(n_12114),
.A2(n_1911),
.B(n_1908),
.C(n_1910),
.Y(n_12215)
);

AOI221xp5_ASAP7_75t_SL g12216 ( 
.A1(n_12123),
.A2(n_1915),
.B1(n_1912),
.B2(n_1914),
.C(n_1916),
.Y(n_12216)
);

NAND2xp5_ASAP7_75t_L g12217 ( 
.A(n_12192),
.B(n_1914),
.Y(n_12217)
);

AND2x2_ASAP7_75t_L g12218 ( 
.A(n_12193),
.B(n_1915),
.Y(n_12218)
);

AOI21xp33_ASAP7_75t_L g12219 ( 
.A1(n_12124),
.A2(n_12089),
.B(n_12096),
.Y(n_12219)
);

OAI31xp33_ASAP7_75t_L g12220 ( 
.A1(n_12148),
.A2(n_1918),
.A3(n_1916),
.B(n_1917),
.Y(n_12220)
);

AND2x2_ASAP7_75t_L g12221 ( 
.A(n_12122),
.B(n_1917),
.Y(n_12221)
);

INVx1_ASAP7_75t_L g12222 ( 
.A(n_12130),
.Y(n_12222)
);

INVx1_ASAP7_75t_L g12223 ( 
.A(n_12141),
.Y(n_12223)
);

OAI221xp5_ASAP7_75t_L g12224 ( 
.A1(n_12107),
.A2(n_2811),
.B1(n_2812),
.B2(n_2810),
.C(n_2809),
.Y(n_12224)
);

NAND2x1p5_ASAP7_75t_L g12225 ( 
.A(n_12146),
.B(n_1920),
.Y(n_12225)
);

AND2x4_ASAP7_75t_L g12226 ( 
.A(n_12077),
.B(n_1920),
.Y(n_12226)
);

NOR2xp67_ASAP7_75t_L g12227 ( 
.A(n_12117),
.B(n_1921),
.Y(n_12227)
);

INVx1_ASAP7_75t_L g12228 ( 
.A(n_12100),
.Y(n_12228)
);

INVx1_ASAP7_75t_L g12229 ( 
.A(n_12120),
.Y(n_12229)
);

AOI211xp5_ASAP7_75t_L g12230 ( 
.A1(n_12125),
.A2(n_1923),
.B(n_1919),
.C(n_1922),
.Y(n_12230)
);

NAND2xp5_ASAP7_75t_L g12231 ( 
.A(n_12083),
.B(n_1919),
.Y(n_12231)
);

INVx1_ASAP7_75t_L g12232 ( 
.A(n_12086),
.Y(n_12232)
);

INVx1_ASAP7_75t_L g12233 ( 
.A(n_12061),
.Y(n_12233)
);

INVx1_ASAP7_75t_L g12234 ( 
.A(n_12063),
.Y(n_12234)
);

NAND2xp5_ASAP7_75t_L g12235 ( 
.A(n_12103),
.B(n_12104),
.Y(n_12235)
);

AOI22xp5_ASAP7_75t_L g12236 ( 
.A1(n_12069),
.A2(n_1925),
.B1(n_1922),
.B2(n_1924),
.Y(n_12236)
);

AOI222xp33_ASAP7_75t_L g12237 ( 
.A1(n_12111),
.A2(n_12055),
.B1(n_12119),
.B2(n_12059),
.C1(n_12153),
.C2(n_12072),
.Y(n_12237)
);

NAND2xp5_ASAP7_75t_L g12238 ( 
.A(n_12128),
.B(n_1924),
.Y(n_12238)
);

INVx1_ASAP7_75t_L g12239 ( 
.A(n_12065),
.Y(n_12239)
);

NOR2xp33_ASAP7_75t_L g12240 ( 
.A(n_12127),
.B(n_1925),
.Y(n_12240)
);

INVx1_ASAP7_75t_L g12241 ( 
.A(n_12067),
.Y(n_12241)
);

OAI22xp5_ASAP7_75t_L g12242 ( 
.A1(n_12099),
.A2(n_1929),
.B1(n_1927),
.B2(n_1928),
.Y(n_12242)
);

NAND2xp5_ASAP7_75t_SL g12243 ( 
.A(n_12106),
.B(n_1927),
.Y(n_12243)
);

OR3x1_ASAP7_75t_L g12244 ( 
.A(n_12060),
.B(n_12090),
.C(n_12138),
.Y(n_12244)
);

OAI32xp33_ASAP7_75t_L g12245 ( 
.A1(n_12151),
.A2(n_1931),
.A3(n_1929),
.B1(n_1930),
.B2(n_1932),
.Y(n_12245)
);

OAI221xp5_ASAP7_75t_L g12246 ( 
.A1(n_12140),
.A2(n_2788),
.B1(n_2807),
.B2(n_2787),
.C(n_2786),
.Y(n_12246)
);

INVx1_ASAP7_75t_L g12247 ( 
.A(n_12068),
.Y(n_12247)
);

INVx1_ASAP7_75t_L g12248 ( 
.A(n_12085),
.Y(n_12248)
);

NAND2xp5_ASAP7_75t_L g12249 ( 
.A(n_12092),
.B(n_1932),
.Y(n_12249)
);

AND2x2_ASAP7_75t_L g12250 ( 
.A(n_12118),
.B(n_1933),
.Y(n_12250)
);

INVx2_ASAP7_75t_L g12251 ( 
.A(n_12147),
.Y(n_12251)
);

O2A1O1Ixp33_ASAP7_75t_SL g12252 ( 
.A1(n_12056),
.A2(n_1943),
.B(n_1954),
.C(n_1933),
.Y(n_12252)
);

INVx3_ASAP7_75t_L g12253 ( 
.A(n_12188),
.Y(n_12253)
);

INVx2_ASAP7_75t_L g12254 ( 
.A(n_12135),
.Y(n_12254)
);

INVx1_ASAP7_75t_L g12255 ( 
.A(n_12087),
.Y(n_12255)
);

HB1xp67_ASAP7_75t_L g12256 ( 
.A(n_12126),
.Y(n_12256)
);

AOI21xp33_ASAP7_75t_SL g12257 ( 
.A1(n_12080),
.A2(n_12155),
.B(n_12145),
.Y(n_12257)
);

INVx1_ASAP7_75t_L g12258 ( 
.A(n_12142),
.Y(n_12258)
);

AOI21xp33_ASAP7_75t_L g12259 ( 
.A1(n_12150),
.A2(n_1934),
.B(n_1935),
.Y(n_12259)
);

AND2x4_ASAP7_75t_L g12260 ( 
.A(n_12098),
.B(n_1935),
.Y(n_12260)
);

NAND2xp5_ASAP7_75t_SL g12261 ( 
.A(n_12181),
.B(n_1934),
.Y(n_12261)
);

NOR2xp33_ASAP7_75t_SL g12262 ( 
.A(n_12162),
.B(n_1936),
.Y(n_12262)
);

AOI22xp5_ASAP7_75t_L g12263 ( 
.A1(n_12167),
.A2(n_1941),
.B1(n_1938),
.B2(n_1940),
.Y(n_12263)
);

AOI21xp33_ASAP7_75t_L g12264 ( 
.A1(n_12139),
.A2(n_1940),
.B(n_1941),
.Y(n_12264)
);

A2O1A1Ixp33_ASAP7_75t_L g12265 ( 
.A1(n_12165),
.A2(n_1945),
.B(n_1942),
.C(n_1943),
.Y(n_12265)
);

NAND2xp5_ASAP7_75t_L g12266 ( 
.A(n_12149),
.B(n_1942),
.Y(n_12266)
);

NAND2x1p5_ASAP7_75t_L g12267 ( 
.A(n_12091),
.B(n_1946),
.Y(n_12267)
);

AOI22xp5_ASAP7_75t_L g12268 ( 
.A1(n_12177),
.A2(n_1949),
.B1(n_1945),
.B2(n_1948),
.Y(n_12268)
);

AOI22xp5_ASAP7_75t_SL g12269 ( 
.A1(n_12136),
.A2(n_1950),
.B1(n_1948),
.B2(n_1949),
.Y(n_12269)
);

INVx1_ASAP7_75t_L g12270 ( 
.A(n_12152),
.Y(n_12270)
);

AOI222xp33_ASAP7_75t_L g12271 ( 
.A1(n_12168),
.A2(n_1953),
.B1(n_1955),
.B2(n_1950),
.C1(n_1952),
.C2(n_1954),
.Y(n_12271)
);

AOI22xp33_ASAP7_75t_L g12272 ( 
.A1(n_12132),
.A2(n_1956),
.B1(n_1952),
.B2(n_1953),
.Y(n_12272)
);

INVx1_ASAP7_75t_L g12273 ( 
.A(n_12137),
.Y(n_12273)
);

AOI22xp33_ASAP7_75t_L g12274 ( 
.A1(n_12166),
.A2(n_1959),
.B1(n_1957),
.B2(n_1958),
.Y(n_12274)
);

INVx1_ASAP7_75t_L g12275 ( 
.A(n_12161),
.Y(n_12275)
);

INVx1_ASAP7_75t_L g12276 ( 
.A(n_12170),
.Y(n_12276)
);

INVx1_ASAP7_75t_L g12277 ( 
.A(n_12169),
.Y(n_12277)
);

AOI22xp5_ASAP7_75t_L g12278 ( 
.A1(n_12097),
.A2(n_1961),
.B1(n_1958),
.B2(n_1960),
.Y(n_12278)
);

NAND2xp5_ASAP7_75t_L g12279 ( 
.A(n_12066),
.B(n_12172),
.Y(n_12279)
);

O2A1O1Ixp33_ASAP7_75t_SL g12280 ( 
.A1(n_12113),
.A2(n_1969),
.B(n_1977),
.C(n_1960),
.Y(n_12280)
);

AND2x2_ASAP7_75t_L g12281 ( 
.A(n_12131),
.B(n_1961),
.Y(n_12281)
);

AND2x2_ASAP7_75t_L g12282 ( 
.A(n_12144),
.B(n_1962),
.Y(n_12282)
);

INVx1_ASAP7_75t_SL g12283 ( 
.A(n_12179),
.Y(n_12283)
);

NAND2xp5_ASAP7_75t_L g12284 ( 
.A(n_12190),
.B(n_1962),
.Y(n_12284)
);

INVx1_ASAP7_75t_SL g12285 ( 
.A(n_12189),
.Y(n_12285)
);

O2A1O1Ixp5_ASAP7_75t_L g12286 ( 
.A1(n_12173),
.A2(n_1965),
.B(n_1963),
.C(n_1964),
.Y(n_12286)
);

AOI22xp5_ASAP7_75t_L g12287 ( 
.A1(n_12180),
.A2(n_1966),
.B1(n_1963),
.B2(n_1965),
.Y(n_12287)
);

INVx1_ASAP7_75t_L g12288 ( 
.A(n_12101),
.Y(n_12288)
);

NAND2xp5_ASAP7_75t_L g12289 ( 
.A(n_12160),
.B(n_1966),
.Y(n_12289)
);

AOI221xp5_ASAP7_75t_L g12290 ( 
.A1(n_12186),
.A2(n_1971),
.B1(n_1968),
.B2(n_1970),
.C(n_1972),
.Y(n_12290)
);

NOR4xp25_ASAP7_75t_L g12291 ( 
.A(n_12095),
.B(n_1973),
.C(n_1971),
.D(n_1972),
.Y(n_12291)
);

AOI22xp33_ASAP7_75t_L g12292 ( 
.A1(n_12109),
.A2(n_1975),
.B1(n_1973),
.B2(n_1974),
.Y(n_12292)
);

INVx1_ASAP7_75t_L g12293 ( 
.A(n_12116),
.Y(n_12293)
);

OAI22xp5_ASAP7_75t_L g12294 ( 
.A1(n_12110),
.A2(n_1976),
.B1(n_1974),
.B2(n_1975),
.Y(n_12294)
);

HB1xp67_ASAP7_75t_L g12295 ( 
.A(n_12057),
.Y(n_12295)
);

OAI22xp5_ASAP7_75t_L g12296 ( 
.A1(n_12115),
.A2(n_1979),
.B1(n_1976),
.B2(n_1978),
.Y(n_12296)
);

A2O1A1Ixp33_ASAP7_75t_L g12297 ( 
.A1(n_12129),
.A2(n_12084),
.B(n_12102),
.C(n_12088),
.Y(n_12297)
);

INVxp67_ASAP7_75t_L g12298 ( 
.A(n_12156),
.Y(n_12298)
);

NAND2xp5_ASAP7_75t_L g12299 ( 
.A(n_12143),
.B(n_1980),
.Y(n_12299)
);

NOR2xp33_ASAP7_75t_L g12300 ( 
.A(n_12185),
.B(n_12171),
.Y(n_12300)
);

AOI211xp5_ASAP7_75t_SL g12301 ( 
.A1(n_12174),
.A2(n_1982),
.B(n_1980),
.C(n_1981),
.Y(n_12301)
);

NOR2xp33_ASAP7_75t_SL g12302 ( 
.A(n_12058),
.B(n_1983),
.Y(n_12302)
);

NAND2xp5_ASAP7_75t_L g12303 ( 
.A(n_12062),
.B(n_12075),
.Y(n_12303)
);

O2A1O1Ixp33_ASAP7_75t_L g12304 ( 
.A1(n_12184),
.A2(n_1985),
.B(n_1983),
.C(n_1984),
.Y(n_12304)
);

HB1xp67_ASAP7_75t_L g12305 ( 
.A(n_12159),
.Y(n_12305)
);

OAI31xp33_ASAP7_75t_L g12306 ( 
.A1(n_12178),
.A2(n_1987),
.A3(n_1985),
.B(n_1986),
.Y(n_12306)
);

OAI21xp33_ASAP7_75t_L g12307 ( 
.A1(n_12176),
.A2(n_1986),
.B(n_1988),
.Y(n_12307)
);

OAI22xp5_ASAP7_75t_L g12308 ( 
.A1(n_12182),
.A2(n_1990),
.B1(n_1988),
.B2(n_1989),
.Y(n_12308)
);

AOI21xp5_ASAP7_75t_L g12309 ( 
.A1(n_12183),
.A2(n_1989),
.B(n_1990),
.Y(n_12309)
);

NAND2x1_ASAP7_75t_L g12310 ( 
.A(n_12175),
.B(n_12187),
.Y(n_12310)
);

NAND2xp5_ASAP7_75t_L g12311 ( 
.A(n_12157),
.B(n_1991),
.Y(n_12311)
);

AND2x2_ASAP7_75t_L g12312 ( 
.A(n_12163),
.B(n_1991),
.Y(n_12312)
);

AOI22xp5_ASAP7_75t_L g12313 ( 
.A1(n_12158),
.A2(n_1994),
.B1(n_1992),
.B2(n_1993),
.Y(n_12313)
);

HB1xp67_ASAP7_75t_L g12314 ( 
.A(n_12078),
.Y(n_12314)
);

INVx1_ASAP7_75t_L g12315 ( 
.A(n_12134),
.Y(n_12315)
);

OAI22xp5_ASAP7_75t_L g12316 ( 
.A1(n_12071),
.A2(n_1996),
.B1(n_1992),
.B2(n_1994),
.Y(n_12316)
);

OR2x2_ASAP7_75t_L g12317 ( 
.A(n_12164),
.B(n_1996),
.Y(n_12317)
);

NAND2xp5_ASAP7_75t_L g12318 ( 
.A(n_12094),
.B(n_1997),
.Y(n_12318)
);

AOI221xp5_ASAP7_75t_L g12319 ( 
.A1(n_12070),
.A2(n_1999),
.B1(n_1997),
.B2(n_1998),
.C(n_2000),
.Y(n_12319)
);

INVx2_ASAP7_75t_L g12320 ( 
.A(n_12134),
.Y(n_12320)
);

AOI21xp33_ASAP7_75t_SL g12321 ( 
.A1(n_12164),
.A2(n_1998),
.B(n_2001),
.Y(n_12321)
);

AOI21xp5_ASAP7_75t_L g12322 ( 
.A1(n_12081),
.A2(n_2002),
.B(n_2003),
.Y(n_12322)
);

NAND2xp5_ASAP7_75t_L g12323 ( 
.A(n_12094),
.B(n_2002),
.Y(n_12323)
);

INVx1_ASAP7_75t_L g12324 ( 
.A(n_12134),
.Y(n_12324)
);

INVx1_ASAP7_75t_SL g12325 ( 
.A(n_12134),
.Y(n_12325)
);

OAI21xp33_ASAP7_75t_L g12326 ( 
.A1(n_12235),
.A2(n_2810),
.B(n_2786),
.Y(n_12326)
);

INVx2_ASAP7_75t_SL g12327 ( 
.A(n_12206),
.Y(n_12327)
);

INVxp67_ASAP7_75t_SL g12328 ( 
.A(n_12227),
.Y(n_12328)
);

NAND2xp5_ASAP7_75t_L g12329 ( 
.A(n_12226),
.B(n_2003),
.Y(n_12329)
);

AOI22xp5_ASAP7_75t_L g12330 ( 
.A1(n_12195),
.A2(n_2007),
.B1(n_2005),
.B2(n_2006),
.Y(n_12330)
);

AND2x2_ASAP7_75t_L g12331 ( 
.A(n_12281),
.B(n_2005),
.Y(n_12331)
);

INVx1_ASAP7_75t_L g12332 ( 
.A(n_12267),
.Y(n_12332)
);

NOR2xp33_ASAP7_75t_L g12333 ( 
.A(n_12317),
.B(n_2006),
.Y(n_12333)
);

NAND2xp5_ASAP7_75t_SL g12334 ( 
.A(n_12320),
.B(n_2007),
.Y(n_12334)
);

INVx2_ASAP7_75t_L g12335 ( 
.A(n_12226),
.Y(n_12335)
);

AOI21xp5_ASAP7_75t_L g12336 ( 
.A1(n_12310),
.A2(n_2008),
.B(n_2009),
.Y(n_12336)
);

O2A1O1Ixp5_ASAP7_75t_SL g12337 ( 
.A1(n_12219),
.A2(n_2775),
.B(n_2776),
.C(n_2773),
.Y(n_12337)
);

NAND2xp5_ASAP7_75t_L g12338 ( 
.A(n_12314),
.B(n_2009),
.Y(n_12338)
);

AOI322xp5_ASAP7_75t_L g12339 ( 
.A1(n_12213),
.A2(n_2015),
.A3(n_2014),
.B1(n_2012),
.B2(n_2010),
.C1(n_2011),
.C2(n_2013),
.Y(n_12339)
);

NAND2xp5_ASAP7_75t_L g12340 ( 
.A(n_12269),
.B(n_12260),
.Y(n_12340)
);

AOI22xp5_ASAP7_75t_L g12341 ( 
.A1(n_12240),
.A2(n_2012),
.B1(n_2010),
.B2(n_2011),
.Y(n_12341)
);

AND2x4_ASAP7_75t_L g12342 ( 
.A(n_12194),
.B(n_2017),
.Y(n_12342)
);

AOI21xp5_ASAP7_75t_L g12343 ( 
.A1(n_12280),
.A2(n_2018),
.B(n_2019),
.Y(n_12343)
);

AOI22xp5_ASAP7_75t_L g12344 ( 
.A1(n_12200),
.A2(n_2021),
.B1(n_2019),
.B2(n_2020),
.Y(n_12344)
);

NOR2x1_ASAP7_75t_L g12345 ( 
.A(n_12223),
.B(n_2020),
.Y(n_12345)
);

AND2x2_ASAP7_75t_L g12346 ( 
.A(n_12282),
.B(n_2022),
.Y(n_12346)
);

INVx1_ASAP7_75t_L g12347 ( 
.A(n_12204),
.Y(n_12347)
);

OAI22xp5_ASAP7_75t_L g12348 ( 
.A1(n_12268),
.A2(n_2024),
.B1(n_2022),
.B2(n_2023),
.Y(n_12348)
);

NAND2xp5_ASAP7_75t_L g12349 ( 
.A(n_12260),
.B(n_2023),
.Y(n_12349)
);

NAND2xp5_ASAP7_75t_L g12350 ( 
.A(n_12301),
.B(n_2024),
.Y(n_12350)
);

INVx1_ASAP7_75t_SL g12351 ( 
.A(n_12325),
.Y(n_12351)
);

OAI322xp33_ASAP7_75t_L g12352 ( 
.A1(n_12277),
.A2(n_2031),
.A3(n_2029),
.B1(n_2027),
.B2(n_2025),
.C1(n_2026),
.C2(n_2028),
.Y(n_12352)
);

INVx2_ASAP7_75t_L g12353 ( 
.A(n_12225),
.Y(n_12353)
);

INVx1_ASAP7_75t_L g12354 ( 
.A(n_12212),
.Y(n_12354)
);

INVx1_ASAP7_75t_L g12355 ( 
.A(n_12318),
.Y(n_12355)
);

AOI21xp5_ASAP7_75t_L g12356 ( 
.A1(n_12231),
.A2(n_2025),
.B(n_2027),
.Y(n_12356)
);

INVx1_ASAP7_75t_L g12357 ( 
.A(n_12323),
.Y(n_12357)
);

AND2x2_ASAP7_75t_L g12358 ( 
.A(n_12312),
.B(n_2028),
.Y(n_12358)
);

NOR2x1p5_ASAP7_75t_L g12359 ( 
.A(n_12253),
.B(n_2778),
.Y(n_12359)
);

INVx1_ASAP7_75t_L g12360 ( 
.A(n_12208),
.Y(n_12360)
);

OAI21xp5_ASAP7_75t_L g12361 ( 
.A1(n_12201),
.A2(n_2031),
.B(n_2032),
.Y(n_12361)
);

INVx2_ASAP7_75t_L g12362 ( 
.A(n_12250),
.Y(n_12362)
);

O2A1O1Ixp33_ASAP7_75t_SL g12363 ( 
.A1(n_12315),
.A2(n_2036),
.B(n_2032),
.C(n_2035),
.Y(n_12363)
);

AOI21xp33_ASAP7_75t_L g12364 ( 
.A1(n_12237),
.A2(n_2035),
.B(n_2037),
.Y(n_12364)
);

OA21x2_ASAP7_75t_L g12365 ( 
.A1(n_12324),
.A2(n_2038),
.B(n_2039),
.Y(n_12365)
);

INVx1_ASAP7_75t_L g12366 ( 
.A(n_12221),
.Y(n_12366)
);

OR2x2_ASAP7_75t_L g12367 ( 
.A(n_12291),
.B(n_2040),
.Y(n_12367)
);

XNOR2x2_ASAP7_75t_L g12368 ( 
.A(n_12196),
.B(n_2040),
.Y(n_12368)
);

INVx1_ASAP7_75t_L g12369 ( 
.A(n_12249),
.Y(n_12369)
);

INVx1_ASAP7_75t_L g12370 ( 
.A(n_12218),
.Y(n_12370)
);

INVx1_ASAP7_75t_L g12371 ( 
.A(n_12209),
.Y(n_12371)
);

INVx1_ASAP7_75t_L g12372 ( 
.A(n_12217),
.Y(n_12372)
);

OR2x2_ASAP7_75t_L g12373 ( 
.A(n_12202),
.B(n_2041),
.Y(n_12373)
);

OAI21xp33_ASAP7_75t_L g12374 ( 
.A1(n_12302),
.A2(n_2770),
.B(n_2769),
.Y(n_12374)
);

INVx1_ASAP7_75t_L g12375 ( 
.A(n_12256),
.Y(n_12375)
);

AND2x2_ASAP7_75t_L g12376 ( 
.A(n_12199),
.B(n_2041),
.Y(n_12376)
);

INVx1_ASAP7_75t_L g12377 ( 
.A(n_12203),
.Y(n_12377)
);

AO22x1_ASAP7_75t_L g12378 ( 
.A1(n_12253),
.A2(n_12251),
.B1(n_12207),
.B2(n_12214),
.Y(n_12378)
);

AOI22xp33_ASAP7_75t_L g12379 ( 
.A1(n_12232),
.A2(n_2044),
.B1(n_2042),
.B2(n_2043),
.Y(n_12379)
);

AOI21xp5_ASAP7_75t_L g12380 ( 
.A1(n_12252),
.A2(n_2043),
.B(n_2044),
.Y(n_12380)
);

NAND2x1_ASAP7_75t_L g12381 ( 
.A(n_12254),
.B(n_2045),
.Y(n_12381)
);

INVx2_ASAP7_75t_L g12382 ( 
.A(n_12244),
.Y(n_12382)
);

NOR3xp33_ASAP7_75t_SL g12383 ( 
.A(n_12297),
.B(n_12279),
.C(n_12224),
.Y(n_12383)
);

AOI22xp5_ASAP7_75t_L g12384 ( 
.A1(n_12262),
.A2(n_12222),
.B1(n_12283),
.B2(n_12285),
.Y(n_12384)
);

AOI22xp5_ASAP7_75t_L g12385 ( 
.A1(n_12258),
.A2(n_2047),
.B1(n_2045),
.B2(n_2046),
.Y(n_12385)
);

HB1xp67_ASAP7_75t_L g12386 ( 
.A(n_12243),
.Y(n_12386)
);

INVx1_ASAP7_75t_L g12387 ( 
.A(n_12266),
.Y(n_12387)
);

INVx1_ASAP7_75t_L g12388 ( 
.A(n_12238),
.Y(n_12388)
);

INVx1_ASAP7_75t_L g12389 ( 
.A(n_12295),
.Y(n_12389)
);

AOI211xp5_ASAP7_75t_L g12390 ( 
.A1(n_12321),
.A2(n_2048),
.B(n_2046),
.C(n_2047),
.Y(n_12390)
);

OR2x2_ASAP7_75t_L g12391 ( 
.A(n_12284),
.B(n_2049),
.Y(n_12391)
);

AOI22xp5_ASAP7_75t_L g12392 ( 
.A1(n_12228),
.A2(n_2051),
.B1(n_2049),
.B2(n_2050),
.Y(n_12392)
);

INVx1_ASAP7_75t_L g12393 ( 
.A(n_12289),
.Y(n_12393)
);

OAI21xp33_ASAP7_75t_L g12394 ( 
.A1(n_12303),
.A2(n_2784),
.B(n_2783),
.Y(n_12394)
);

INVx1_ASAP7_75t_L g12395 ( 
.A(n_12316),
.Y(n_12395)
);

OAI221xp5_ASAP7_75t_L g12396 ( 
.A1(n_12210),
.A2(n_2053),
.B1(n_2050),
.B2(n_2052),
.C(n_2054),
.Y(n_12396)
);

INVx1_ASAP7_75t_L g12397 ( 
.A(n_12286),
.Y(n_12397)
);

INVx1_ASAP7_75t_L g12398 ( 
.A(n_12299),
.Y(n_12398)
);

OAI321xp33_ASAP7_75t_L g12399 ( 
.A1(n_12205),
.A2(n_2055),
.A3(n_2059),
.B1(n_2053),
.B2(n_2054),
.C(n_2057),
.Y(n_12399)
);

OAI22xp33_ASAP7_75t_L g12400 ( 
.A1(n_12311),
.A2(n_12287),
.B1(n_12263),
.B2(n_12278),
.Y(n_12400)
);

INVx2_ASAP7_75t_L g12401 ( 
.A(n_12239),
.Y(n_12401)
);

AOI22xp33_ASAP7_75t_L g12402 ( 
.A1(n_12273),
.A2(n_2060),
.B1(n_2055),
.B2(n_2057),
.Y(n_12402)
);

INVx2_ASAP7_75t_L g12403 ( 
.A(n_12241),
.Y(n_12403)
);

OAI322xp33_ASAP7_75t_L g12404 ( 
.A1(n_12247),
.A2(n_2065),
.A3(n_2064),
.B1(n_2062),
.B2(n_2060),
.C1(n_2061),
.C2(n_2063),
.Y(n_12404)
);

AOI22xp5_ASAP7_75t_L g12405 ( 
.A1(n_12248),
.A2(n_2063),
.B1(n_2061),
.B2(n_2062),
.Y(n_12405)
);

A2O1A1Ixp33_ASAP7_75t_L g12406 ( 
.A1(n_12304),
.A2(n_12220),
.B(n_12306),
.C(n_12322),
.Y(n_12406)
);

A2O1A1Ixp33_ASAP7_75t_L g12407 ( 
.A1(n_12197),
.A2(n_2066),
.B(n_2064),
.C(n_2065),
.Y(n_12407)
);

INVx1_ASAP7_75t_L g12408 ( 
.A(n_12255),
.Y(n_12408)
);

NAND2xp5_ASAP7_75t_L g12409 ( 
.A(n_12216),
.B(n_2067),
.Y(n_12409)
);

INVx1_ASAP7_75t_L g12410 ( 
.A(n_12261),
.Y(n_12410)
);

AOI22xp5_ASAP7_75t_L g12411 ( 
.A1(n_12270),
.A2(n_2069),
.B1(n_2067),
.B2(n_2068),
.Y(n_12411)
);

INVx1_ASAP7_75t_L g12412 ( 
.A(n_12275),
.Y(n_12412)
);

NAND2xp33_ASAP7_75t_SL g12413 ( 
.A(n_12276),
.B(n_2784),
.Y(n_12413)
);

NOR2xp33_ASAP7_75t_L g12414 ( 
.A(n_12215),
.B(n_2069),
.Y(n_12414)
);

INVx2_ASAP7_75t_L g12415 ( 
.A(n_12229),
.Y(n_12415)
);

INVx2_ASAP7_75t_L g12416 ( 
.A(n_12233),
.Y(n_12416)
);

OAI22xp5_ASAP7_75t_L g12417 ( 
.A1(n_12246),
.A2(n_2072),
.B1(n_2070),
.B2(n_2071),
.Y(n_12417)
);

NAND2xp5_ASAP7_75t_L g12418 ( 
.A(n_12271),
.B(n_2070),
.Y(n_12418)
);

NAND2xp5_ASAP7_75t_L g12419 ( 
.A(n_12319),
.B(n_2071),
.Y(n_12419)
);

INVxp67_ASAP7_75t_SL g12420 ( 
.A(n_12211),
.Y(n_12420)
);

CKINVDCx20_ASAP7_75t_R g12421 ( 
.A(n_12305),
.Y(n_12421)
);

AOI22xp5_ASAP7_75t_L g12422 ( 
.A1(n_12300),
.A2(n_2074),
.B1(n_2072),
.B2(n_2073),
.Y(n_12422)
);

OAI322xp33_ASAP7_75t_L g12423 ( 
.A1(n_12298),
.A2(n_2079),
.A3(n_2078),
.B1(n_2076),
.B2(n_2073),
.C1(n_2075),
.C2(n_2077),
.Y(n_12423)
);

INVx2_ASAP7_75t_L g12424 ( 
.A(n_12234),
.Y(n_12424)
);

INVx1_ASAP7_75t_L g12425 ( 
.A(n_12307),
.Y(n_12425)
);

INVx1_ASAP7_75t_L g12426 ( 
.A(n_12294),
.Y(n_12426)
);

INVxp67_ASAP7_75t_L g12427 ( 
.A(n_12296),
.Y(n_12427)
);

NAND2xp5_ASAP7_75t_L g12428 ( 
.A(n_12292),
.B(n_2075),
.Y(n_12428)
);

INVx1_ASAP7_75t_L g12429 ( 
.A(n_12313),
.Y(n_12429)
);

NAND3xp33_ASAP7_75t_SL g12430 ( 
.A(n_12230),
.B(n_12257),
.C(n_12309),
.Y(n_12430)
);

NAND3xp33_ASAP7_75t_L g12431 ( 
.A(n_12290),
.B(n_12259),
.C(n_12265),
.Y(n_12431)
);

OA21x2_ASAP7_75t_L g12432 ( 
.A1(n_12293),
.A2(n_2077),
.B(n_2080),
.Y(n_12432)
);

INVx1_ASAP7_75t_L g12433 ( 
.A(n_12308),
.Y(n_12433)
);

OR2x2_ASAP7_75t_L g12434 ( 
.A(n_12288),
.B(n_2080),
.Y(n_12434)
);

INVx1_ASAP7_75t_L g12435 ( 
.A(n_12242),
.Y(n_12435)
);

OR3x2_ASAP7_75t_L g12436 ( 
.A(n_12245),
.B(n_12264),
.C(n_12198),
.Y(n_12436)
);

AND3x1_ASAP7_75t_L g12437 ( 
.A(n_12236),
.B(n_2081),
.C(n_2082),
.Y(n_12437)
);

NOR2xp33_ASAP7_75t_L g12438 ( 
.A(n_12274),
.B(n_2081),
.Y(n_12438)
);

INVxp67_ASAP7_75t_L g12439 ( 
.A(n_12272),
.Y(n_12439)
);

OAI22xp5_ASAP7_75t_L g12440 ( 
.A1(n_12200),
.A2(n_2084),
.B1(n_2082),
.B2(n_2083),
.Y(n_12440)
);

INVx1_ASAP7_75t_L g12441 ( 
.A(n_12267),
.Y(n_12441)
);

OAI21xp5_ASAP7_75t_SL g12442 ( 
.A1(n_12237),
.A2(n_2085),
.B(n_2084),
.Y(n_12442)
);

AOI211xp5_ASAP7_75t_L g12443 ( 
.A1(n_12195),
.A2(n_2088),
.B(n_2083),
.C(n_2086),
.Y(n_12443)
);

INVx2_ASAP7_75t_L g12444 ( 
.A(n_12267),
.Y(n_12444)
);

NAND2xp5_ASAP7_75t_L g12445 ( 
.A(n_12227),
.B(n_2089),
.Y(n_12445)
);

OR2x2_ASAP7_75t_L g12446 ( 
.A(n_12327),
.B(n_12367),
.Y(n_12446)
);

NOR2xp33_ASAP7_75t_L g12447 ( 
.A(n_12442),
.B(n_2089),
.Y(n_12447)
);

NAND2xp5_ASAP7_75t_L g12448 ( 
.A(n_12328),
.B(n_2090),
.Y(n_12448)
);

AOI22xp5_ASAP7_75t_L g12449 ( 
.A1(n_12421),
.A2(n_2092),
.B1(n_2090),
.B2(n_2091),
.Y(n_12449)
);

INVx1_ASAP7_75t_L g12450 ( 
.A(n_12365),
.Y(n_12450)
);

INVx2_ASAP7_75t_L g12451 ( 
.A(n_12365),
.Y(n_12451)
);

NAND2xp5_ASAP7_75t_L g12452 ( 
.A(n_12335),
.B(n_2091),
.Y(n_12452)
);

INVx1_ASAP7_75t_L g12453 ( 
.A(n_12345),
.Y(n_12453)
);

NAND2xp5_ASAP7_75t_SL g12454 ( 
.A(n_12444),
.B(n_12343),
.Y(n_12454)
);

NOR2xp33_ASAP7_75t_L g12455 ( 
.A(n_12326),
.B(n_2093),
.Y(n_12455)
);

OAI22xp5_ASAP7_75t_L g12456 ( 
.A1(n_12330),
.A2(n_12351),
.B1(n_12384),
.B2(n_12347),
.Y(n_12456)
);

NAND2xp5_ASAP7_75t_L g12457 ( 
.A(n_12359),
.B(n_2094),
.Y(n_12457)
);

AOI22xp5_ASAP7_75t_L g12458 ( 
.A1(n_12389),
.A2(n_2097),
.B1(n_2094),
.B2(n_2096),
.Y(n_12458)
);

NAND2xp5_ASAP7_75t_L g12459 ( 
.A(n_12346),
.B(n_2097),
.Y(n_12459)
);

NAND2xp5_ASAP7_75t_L g12460 ( 
.A(n_12358),
.B(n_2098),
.Y(n_12460)
);

AND2x2_ASAP7_75t_L g12461 ( 
.A(n_12331),
.B(n_2098),
.Y(n_12461)
);

AND2x2_ASAP7_75t_L g12462 ( 
.A(n_12376),
.B(n_2099),
.Y(n_12462)
);

NOR2xp33_ASAP7_75t_L g12463 ( 
.A(n_12396),
.B(n_2099),
.Y(n_12463)
);

NAND2xp5_ASAP7_75t_L g12464 ( 
.A(n_12378),
.B(n_2100),
.Y(n_12464)
);

HB1xp67_ASAP7_75t_L g12465 ( 
.A(n_12432),
.Y(n_12465)
);

INVx1_ASAP7_75t_SL g12466 ( 
.A(n_12413),
.Y(n_12466)
);

AOI22xp33_ASAP7_75t_L g12467 ( 
.A1(n_12382),
.A2(n_2102),
.B1(n_2100),
.B2(n_2101),
.Y(n_12467)
);

OAI22xp5_ASAP7_75t_L g12468 ( 
.A1(n_12436),
.A2(n_2103),
.B1(n_2101),
.B2(n_2102),
.Y(n_12468)
);

NOR2xp33_ASAP7_75t_L g12469 ( 
.A(n_12364),
.B(n_2103),
.Y(n_12469)
);

AND2x2_ASAP7_75t_L g12470 ( 
.A(n_12371),
.B(n_2104),
.Y(n_12470)
);

NAND2xp5_ASAP7_75t_L g12471 ( 
.A(n_12336),
.B(n_12332),
.Y(n_12471)
);

INVx1_ASAP7_75t_L g12472 ( 
.A(n_12432),
.Y(n_12472)
);

AND2x2_ASAP7_75t_L g12473 ( 
.A(n_12441),
.B(n_2104),
.Y(n_12473)
);

INVx1_ASAP7_75t_L g12474 ( 
.A(n_12373),
.Y(n_12474)
);

NAND2xp5_ASAP7_75t_L g12475 ( 
.A(n_12342),
.B(n_12390),
.Y(n_12475)
);

AND2x2_ASAP7_75t_L g12476 ( 
.A(n_12366),
.B(n_2105),
.Y(n_12476)
);

NAND2xp5_ASAP7_75t_L g12477 ( 
.A(n_12342),
.B(n_12333),
.Y(n_12477)
);

OR2x2_ASAP7_75t_L g12478 ( 
.A(n_12340),
.B(n_2105),
.Y(n_12478)
);

INVx1_ASAP7_75t_SL g12479 ( 
.A(n_12445),
.Y(n_12479)
);

INVx1_ASAP7_75t_L g12480 ( 
.A(n_12329),
.Y(n_12480)
);

AOI22xp33_ASAP7_75t_L g12481 ( 
.A1(n_12375),
.A2(n_2109),
.B1(n_2107),
.B2(n_2108),
.Y(n_12481)
);

INVx1_ASAP7_75t_SL g12482 ( 
.A(n_12350),
.Y(n_12482)
);

NAND2xp5_ASAP7_75t_L g12483 ( 
.A(n_12414),
.B(n_2107),
.Y(n_12483)
);

NOR2xp33_ASAP7_75t_SL g12484 ( 
.A(n_12352),
.B(n_2110),
.Y(n_12484)
);

NOR2xp33_ASAP7_75t_L g12485 ( 
.A(n_12394),
.B(n_2111),
.Y(n_12485)
);

INVx1_ASAP7_75t_L g12486 ( 
.A(n_12381),
.Y(n_12486)
);

NAND2xp5_ASAP7_75t_L g12487 ( 
.A(n_12443),
.B(n_2111),
.Y(n_12487)
);

INVx1_ASAP7_75t_L g12488 ( 
.A(n_12349),
.Y(n_12488)
);

NAND2xp5_ASAP7_75t_L g12489 ( 
.A(n_12380),
.B(n_2112),
.Y(n_12489)
);

AOI21xp33_ASAP7_75t_L g12490 ( 
.A1(n_12377),
.A2(n_12338),
.B(n_12397),
.Y(n_12490)
);

NAND2xp5_ASAP7_75t_L g12491 ( 
.A(n_12353),
.B(n_2113),
.Y(n_12491)
);

INVx1_ASAP7_75t_L g12492 ( 
.A(n_12363),
.Y(n_12492)
);

INVx1_ASAP7_75t_L g12493 ( 
.A(n_12434),
.Y(n_12493)
);

BUFx4f_ASAP7_75t_L g12494 ( 
.A(n_12408),
.Y(n_12494)
);

INVxp67_ASAP7_75t_L g12495 ( 
.A(n_12437),
.Y(n_12495)
);

AO22x1_ASAP7_75t_L g12496 ( 
.A1(n_12361),
.A2(n_2116),
.B1(n_2113),
.B2(n_2115),
.Y(n_12496)
);

INVx1_ASAP7_75t_L g12497 ( 
.A(n_12409),
.Y(n_12497)
);

AND2x2_ASAP7_75t_L g12498 ( 
.A(n_12362),
.B(n_2116),
.Y(n_12498)
);

AOI22xp5_ASAP7_75t_L g12499 ( 
.A1(n_12401),
.A2(n_2119),
.B1(n_2117),
.B2(n_2118),
.Y(n_12499)
);

NAND2xp5_ASAP7_75t_L g12500 ( 
.A(n_12344),
.B(n_2118),
.Y(n_12500)
);

INVx2_ASAP7_75t_L g12501 ( 
.A(n_12391),
.Y(n_12501)
);

INVx2_ASAP7_75t_L g12502 ( 
.A(n_12368),
.Y(n_12502)
);

INVx2_ASAP7_75t_SL g12503 ( 
.A(n_12386),
.Y(n_12503)
);

NAND2xp5_ASAP7_75t_L g12504 ( 
.A(n_12360),
.B(n_2119),
.Y(n_12504)
);

NAND2xp5_ASAP7_75t_L g12505 ( 
.A(n_12341),
.B(n_2120),
.Y(n_12505)
);

INVx1_ASAP7_75t_L g12506 ( 
.A(n_12418),
.Y(n_12506)
);

NAND2xp33_ASAP7_75t_L g12507 ( 
.A(n_12374),
.B(n_2120),
.Y(n_12507)
);

INVx1_ASAP7_75t_L g12508 ( 
.A(n_12419),
.Y(n_12508)
);

INVx2_ASAP7_75t_L g12509 ( 
.A(n_12403),
.Y(n_12509)
);

AND2x2_ASAP7_75t_L g12510 ( 
.A(n_12383),
.B(n_2121),
.Y(n_12510)
);

INVx1_ASAP7_75t_L g12511 ( 
.A(n_12428),
.Y(n_12511)
);

INVx1_ASAP7_75t_L g12512 ( 
.A(n_12334),
.Y(n_12512)
);

NAND2xp5_ASAP7_75t_L g12513 ( 
.A(n_12356),
.B(n_2121),
.Y(n_12513)
);

OR2x2_ASAP7_75t_L g12514 ( 
.A(n_12430),
.B(n_2122),
.Y(n_12514)
);

AND2x4_ASAP7_75t_L g12515 ( 
.A(n_12370),
.B(n_2123),
.Y(n_12515)
);

INVx1_ASAP7_75t_L g12516 ( 
.A(n_12412),
.Y(n_12516)
);

NAND2xp5_ASAP7_75t_L g12517 ( 
.A(n_12402),
.B(n_2123),
.Y(n_12517)
);

OR2x2_ASAP7_75t_L g12518 ( 
.A(n_12348),
.B(n_2124),
.Y(n_12518)
);

INVx2_ASAP7_75t_L g12519 ( 
.A(n_12354),
.Y(n_12519)
);

AOI22xp5_ASAP7_75t_L g12520 ( 
.A1(n_12420),
.A2(n_2128),
.B1(n_2126),
.B2(n_2127),
.Y(n_12520)
);

INVx1_ASAP7_75t_SL g12521 ( 
.A(n_12410),
.Y(n_12521)
);

INVx1_ASAP7_75t_SL g12522 ( 
.A(n_12426),
.Y(n_12522)
);

INVx1_ASAP7_75t_L g12523 ( 
.A(n_12407),
.Y(n_12523)
);

AND2x2_ASAP7_75t_L g12524 ( 
.A(n_12355),
.B(n_2126),
.Y(n_12524)
);

HB1xp67_ASAP7_75t_L g12525 ( 
.A(n_12440),
.Y(n_12525)
);

NAND2x1_ASAP7_75t_L g12526 ( 
.A(n_12425),
.B(n_2127),
.Y(n_12526)
);

INVx1_ASAP7_75t_L g12527 ( 
.A(n_12417),
.Y(n_12527)
);

NAND2xp5_ASAP7_75t_L g12528 ( 
.A(n_12379),
.B(n_2128),
.Y(n_12528)
);

INVx1_ASAP7_75t_L g12529 ( 
.A(n_12357),
.Y(n_12529)
);

NAND2xp5_ASAP7_75t_L g12530 ( 
.A(n_12339),
.B(n_2129),
.Y(n_12530)
);

NAND2xp5_ASAP7_75t_L g12531 ( 
.A(n_12405),
.B(n_2129),
.Y(n_12531)
);

NAND2xp5_ASAP7_75t_L g12532 ( 
.A(n_12411),
.B(n_2130),
.Y(n_12532)
);

AND2x2_ASAP7_75t_L g12533 ( 
.A(n_12427),
.B(n_2130),
.Y(n_12533)
);

NAND2xp5_ASAP7_75t_L g12534 ( 
.A(n_12406),
.B(n_2131),
.Y(n_12534)
);

OR2x2_ASAP7_75t_L g12535 ( 
.A(n_12395),
.B(n_2131),
.Y(n_12535)
);

AND2x2_ASAP7_75t_L g12536 ( 
.A(n_12439),
.B(n_12429),
.Y(n_12536)
);

INVx2_ASAP7_75t_L g12537 ( 
.A(n_12415),
.Y(n_12537)
);

OR2x2_ASAP7_75t_L g12538 ( 
.A(n_12433),
.B(n_2132),
.Y(n_12538)
);

NAND2xp5_ASAP7_75t_L g12539 ( 
.A(n_12438),
.B(n_2132),
.Y(n_12539)
);

AND2x2_ASAP7_75t_L g12540 ( 
.A(n_12435),
.B(n_2133),
.Y(n_12540)
);

INVx2_ASAP7_75t_L g12541 ( 
.A(n_12387),
.Y(n_12541)
);

AOI22xp33_ASAP7_75t_L g12542 ( 
.A1(n_12416),
.A2(n_2135),
.B1(n_2133),
.B2(n_2134),
.Y(n_12542)
);

AND2x2_ASAP7_75t_L g12543 ( 
.A(n_12424),
.B(n_12369),
.Y(n_12543)
);

NAND2xp5_ASAP7_75t_L g12544 ( 
.A(n_12385),
.B(n_12392),
.Y(n_12544)
);

INVxp67_ASAP7_75t_L g12545 ( 
.A(n_12422),
.Y(n_12545)
);

OR2x2_ASAP7_75t_L g12546 ( 
.A(n_12431),
.B(n_2134),
.Y(n_12546)
);

INVx2_ASAP7_75t_L g12547 ( 
.A(n_12372),
.Y(n_12547)
);

NAND2xp5_ASAP7_75t_L g12548 ( 
.A(n_12388),
.B(n_2135),
.Y(n_12548)
);

NOR2xp33_ASAP7_75t_L g12549 ( 
.A(n_12400),
.B(n_2136),
.Y(n_12549)
);

AND2x2_ASAP7_75t_L g12550 ( 
.A(n_12393),
.B(n_2136),
.Y(n_12550)
);

NAND2xp5_ASAP7_75t_L g12551 ( 
.A(n_12398),
.B(n_2137),
.Y(n_12551)
);

NAND2xp5_ASAP7_75t_L g12552 ( 
.A(n_12337),
.B(n_12399),
.Y(n_12552)
);

INVx2_ASAP7_75t_SL g12553 ( 
.A(n_12404),
.Y(n_12553)
);

AOI22x1_ASAP7_75t_L g12554 ( 
.A1(n_12423),
.A2(n_2140),
.B1(n_2138),
.B2(n_2139),
.Y(n_12554)
);

INVx2_ASAP7_75t_L g12555 ( 
.A(n_12365),
.Y(n_12555)
);

INVx3_ASAP7_75t_L g12556 ( 
.A(n_12381),
.Y(n_12556)
);

NAND2xp5_ASAP7_75t_SL g12557 ( 
.A(n_12327),
.B(n_2138),
.Y(n_12557)
);

NAND2xp5_ASAP7_75t_L g12558 ( 
.A(n_12327),
.B(n_2139),
.Y(n_12558)
);

AOI222xp33_ASAP7_75t_L g12559 ( 
.A1(n_12442),
.A2(n_2142),
.B1(n_2144),
.B2(n_2140),
.C1(n_2141),
.C2(n_2143),
.Y(n_12559)
);

AND2x2_ASAP7_75t_L g12560 ( 
.A(n_12346),
.B(n_2141),
.Y(n_12560)
);

INVx1_ASAP7_75t_L g12561 ( 
.A(n_12365),
.Y(n_12561)
);

INVx1_ASAP7_75t_L g12562 ( 
.A(n_12365),
.Y(n_12562)
);

NOR2xp33_ASAP7_75t_L g12563 ( 
.A(n_12327),
.B(n_2142),
.Y(n_12563)
);

INVx1_ASAP7_75t_L g12564 ( 
.A(n_12465),
.Y(n_12564)
);

AO22x1_ASAP7_75t_L g12565 ( 
.A1(n_12450),
.A2(n_2147),
.B1(n_2145),
.B2(n_2146),
.Y(n_12565)
);

INVx1_ASAP7_75t_L g12566 ( 
.A(n_12561),
.Y(n_12566)
);

OA22x2_ASAP7_75t_L g12567 ( 
.A1(n_12492),
.A2(n_2147),
.B1(n_2145),
.B2(n_2146),
.Y(n_12567)
);

NAND4xp75_ASAP7_75t_SL g12568 ( 
.A(n_12510),
.B(n_2150),
.C(n_2148),
.D(n_2149),
.Y(n_12568)
);

AOI22x1_ASAP7_75t_L g12569 ( 
.A1(n_12451),
.A2(n_2151),
.B1(n_2148),
.B2(n_2150),
.Y(n_12569)
);

INVx1_ASAP7_75t_L g12570 ( 
.A(n_12562),
.Y(n_12570)
);

INVx3_ASAP7_75t_L g12571 ( 
.A(n_12556),
.Y(n_12571)
);

NOR2x1_ASAP7_75t_L g12572 ( 
.A(n_12472),
.B(n_12555),
.Y(n_12572)
);

BUFx2_ASAP7_75t_L g12573 ( 
.A(n_12556),
.Y(n_12573)
);

AOI22xp5_ASAP7_75t_L g12574 ( 
.A1(n_12503),
.A2(n_2155),
.B1(n_2152),
.B2(n_2154),
.Y(n_12574)
);

INVx2_ASAP7_75t_SL g12575 ( 
.A(n_12526),
.Y(n_12575)
);

AOI211x1_ASAP7_75t_SL g12576 ( 
.A1(n_12456),
.A2(n_2157),
.B(n_2154),
.C(n_2156),
.Y(n_12576)
);

OA22x2_ASAP7_75t_L g12577 ( 
.A1(n_12466),
.A2(n_2160),
.B1(n_2156),
.B2(n_2159),
.Y(n_12577)
);

OAI322xp33_ASAP7_75t_L g12578 ( 
.A1(n_12484),
.A2(n_2186),
.A3(n_2170),
.B1(n_2195),
.B2(n_2207),
.C1(n_2178),
.C2(n_2160),
.Y(n_12578)
);

INVx2_ASAP7_75t_SL g12579 ( 
.A(n_12494),
.Y(n_12579)
);

INVx1_ASAP7_75t_L g12580 ( 
.A(n_12476),
.Y(n_12580)
);

AOI22xp5_ASAP7_75t_L g12581 ( 
.A1(n_12522),
.A2(n_12549),
.B1(n_12521),
.B2(n_12553),
.Y(n_12581)
);

INVx1_ASAP7_75t_L g12582 ( 
.A(n_12560),
.Y(n_12582)
);

INVx2_ASAP7_75t_L g12583 ( 
.A(n_12515),
.Y(n_12583)
);

INVx1_ASAP7_75t_L g12584 ( 
.A(n_12461),
.Y(n_12584)
);

INVx1_ASAP7_75t_L g12585 ( 
.A(n_12515),
.Y(n_12585)
);

INVx1_ASAP7_75t_L g12586 ( 
.A(n_12498),
.Y(n_12586)
);

NAND4xp25_ASAP7_75t_L g12587 ( 
.A(n_12490),
.B(n_2163),
.C(n_2161),
.D(n_2162),
.Y(n_12587)
);

OA22x2_ASAP7_75t_L g12588 ( 
.A1(n_12486),
.A2(n_2165),
.B1(n_2161),
.B2(n_2163),
.Y(n_12588)
);

AOI22xp5_ASAP7_75t_L g12589 ( 
.A1(n_12509),
.A2(n_2167),
.B1(n_2165),
.B2(n_2166),
.Y(n_12589)
);

INVx1_ASAP7_75t_L g12590 ( 
.A(n_12473),
.Y(n_12590)
);

NOR4xp25_ASAP7_75t_L g12591 ( 
.A(n_12464),
.B(n_2168),
.C(n_2166),
.D(n_2167),
.Y(n_12591)
);

AOI22xp5_ASAP7_75t_L g12592 ( 
.A1(n_12468),
.A2(n_2172),
.B1(n_2170),
.B2(n_2171),
.Y(n_12592)
);

INVx1_ASAP7_75t_L g12593 ( 
.A(n_12462),
.Y(n_12593)
);

OAI322xp33_ASAP7_75t_L g12594 ( 
.A1(n_12495),
.A2(n_2199),
.A3(n_2179),
.B1(n_2210),
.B2(n_2218),
.C1(n_2188),
.C2(n_2171),
.Y(n_12594)
);

INVx1_ASAP7_75t_SL g12595 ( 
.A(n_12478),
.Y(n_12595)
);

AOI22xp5_ASAP7_75t_L g12596 ( 
.A1(n_12536),
.A2(n_2174),
.B1(n_2172),
.B2(n_2173),
.Y(n_12596)
);

AOI22xp5_ASAP7_75t_L g12597 ( 
.A1(n_12502),
.A2(n_12537),
.B1(n_12447),
.B2(n_12533),
.Y(n_12597)
);

AO22x2_ASAP7_75t_L g12598 ( 
.A1(n_12453),
.A2(n_2176),
.B1(n_2174),
.B2(n_2175),
.Y(n_12598)
);

NOR4xp25_ASAP7_75t_L g12599 ( 
.A(n_12454),
.B(n_2178),
.C(n_2176),
.D(n_2177),
.Y(n_12599)
);

INVx1_ASAP7_75t_L g12600 ( 
.A(n_12524),
.Y(n_12600)
);

AOI22xp5_ASAP7_75t_L g12601 ( 
.A1(n_12470),
.A2(n_2181),
.B1(n_2179),
.B2(n_2180),
.Y(n_12601)
);

INVx1_ASAP7_75t_SL g12602 ( 
.A(n_12538),
.Y(n_12602)
);

INVx1_ASAP7_75t_L g12603 ( 
.A(n_12457),
.Y(n_12603)
);

AOI22xp5_ASAP7_75t_SL g12604 ( 
.A1(n_12496),
.A2(n_2182),
.B1(n_2183),
.B2(n_2181),
.Y(n_12604)
);

NAND4xp75_ASAP7_75t_L g12605 ( 
.A(n_12540),
.B(n_2183),
.C(n_2180),
.D(n_2182),
.Y(n_12605)
);

OA22x2_ASAP7_75t_L g12606 ( 
.A1(n_12558),
.A2(n_2187),
.B1(n_2184),
.B2(n_2185),
.Y(n_12606)
);

AOI22xp5_ASAP7_75t_L g12607 ( 
.A1(n_12563),
.A2(n_2189),
.B1(n_2184),
.B2(n_2188),
.Y(n_12607)
);

INVx1_ASAP7_75t_L g12608 ( 
.A(n_12550),
.Y(n_12608)
);

HB1xp67_ASAP7_75t_L g12609 ( 
.A(n_12557),
.Y(n_12609)
);

INVx1_ASAP7_75t_L g12610 ( 
.A(n_12459),
.Y(n_12610)
);

INVxp67_ASAP7_75t_SL g12611 ( 
.A(n_12460),
.Y(n_12611)
);

INVx1_ASAP7_75t_L g12612 ( 
.A(n_12452),
.Y(n_12612)
);

INVx1_ASAP7_75t_L g12613 ( 
.A(n_12535),
.Y(n_12613)
);

INVx1_ASAP7_75t_L g12614 ( 
.A(n_12448),
.Y(n_12614)
);

AOI22xp33_ASAP7_75t_L g12615 ( 
.A1(n_12554),
.A2(n_2191),
.B1(n_2192),
.B2(n_2190),
.Y(n_12615)
);

OAI322xp33_ASAP7_75t_L g12616 ( 
.A1(n_12514),
.A2(n_2219),
.A3(n_2200),
.B1(n_2227),
.B2(n_2235),
.C1(n_2211),
.C2(n_2189),
.Y(n_12616)
);

OAI322xp33_ASAP7_75t_L g12617 ( 
.A1(n_12446),
.A2(n_2221),
.A3(n_2201),
.B1(n_2229),
.B2(n_2238),
.C1(n_2213),
.C2(n_2190),
.Y(n_12617)
);

INVx1_ASAP7_75t_L g12618 ( 
.A(n_12504),
.Y(n_12618)
);

AOI22xp5_ASAP7_75t_L g12619 ( 
.A1(n_12527),
.A2(n_2193),
.B1(n_2191),
.B2(n_2192),
.Y(n_12619)
);

INVx1_ASAP7_75t_L g12620 ( 
.A(n_12534),
.Y(n_12620)
);

BUFx4_ASAP7_75t_R g12621 ( 
.A(n_12501),
.Y(n_12621)
);

AOI22xp5_ASAP7_75t_L g12622 ( 
.A1(n_12455),
.A2(n_12463),
.B1(n_12543),
.B2(n_12507),
.Y(n_12622)
);

AOI22xp5_ASAP7_75t_L g12623 ( 
.A1(n_12523),
.A2(n_2198),
.B1(n_2193),
.B2(n_2195),
.Y(n_12623)
);

INVx1_ASAP7_75t_L g12624 ( 
.A(n_12546),
.Y(n_12624)
);

INVx1_ASAP7_75t_L g12625 ( 
.A(n_12489),
.Y(n_12625)
);

AOI22xp5_ASAP7_75t_L g12626 ( 
.A1(n_12485),
.A2(n_2200),
.B1(n_2198),
.B2(n_2199),
.Y(n_12626)
);

INVx1_ASAP7_75t_L g12627 ( 
.A(n_12530),
.Y(n_12627)
);

INVx1_ASAP7_75t_L g12628 ( 
.A(n_12491),
.Y(n_12628)
);

AOI211xp5_ASAP7_75t_SL g12629 ( 
.A1(n_12469),
.A2(n_2205),
.B(n_2203),
.C(n_2204),
.Y(n_12629)
);

OA22x2_ASAP7_75t_L g12630 ( 
.A1(n_12516),
.A2(n_2209),
.B1(n_2203),
.B2(n_2207),
.Y(n_12630)
);

AOI22xp5_ASAP7_75t_L g12631 ( 
.A1(n_12512),
.A2(n_2212),
.B1(n_2209),
.B2(n_2210),
.Y(n_12631)
);

INVx1_ASAP7_75t_L g12632 ( 
.A(n_12475),
.Y(n_12632)
);

AOI22xp5_ASAP7_75t_L g12633 ( 
.A1(n_12545),
.A2(n_2214),
.B1(n_2212),
.B2(n_2213),
.Y(n_12633)
);

INVx1_ASAP7_75t_L g12634 ( 
.A(n_12525),
.Y(n_12634)
);

INVx1_ASAP7_75t_L g12635 ( 
.A(n_12548),
.Y(n_12635)
);

OAI211xp5_ASAP7_75t_L g12636 ( 
.A1(n_12559),
.A2(n_12552),
.B(n_12517),
.C(n_12528),
.Y(n_12636)
);

NAND5xp2_ASAP7_75t_SL g12637 ( 
.A(n_12467),
.B(n_2216),
.C(n_2214),
.D(n_2215),
.E(n_2217),
.Y(n_12637)
);

OA22x2_ASAP7_75t_L g12638 ( 
.A1(n_12482),
.A2(n_2217),
.B1(n_2215),
.B2(n_2216),
.Y(n_12638)
);

INVx1_ASAP7_75t_L g12639 ( 
.A(n_12471),
.Y(n_12639)
);

INVx1_ASAP7_75t_L g12640 ( 
.A(n_12551),
.Y(n_12640)
);

INVx1_ASAP7_75t_SL g12641 ( 
.A(n_12513),
.Y(n_12641)
);

HB1xp67_ASAP7_75t_L g12642 ( 
.A(n_12474),
.Y(n_12642)
);

OA22x2_ASAP7_75t_L g12643 ( 
.A1(n_12493),
.A2(n_2220),
.B1(n_2218),
.B2(n_2219),
.Y(n_12643)
);

OAI22xp5_ASAP7_75t_L g12644 ( 
.A1(n_12487),
.A2(n_2222),
.B1(n_2220),
.B2(n_2221),
.Y(n_12644)
);

AOI22xp5_ASAP7_75t_L g12645 ( 
.A1(n_12519),
.A2(n_2224),
.B1(n_2222),
.B2(n_2223),
.Y(n_12645)
);

INVx1_ASAP7_75t_L g12646 ( 
.A(n_12483),
.Y(n_12646)
);

INVx1_ASAP7_75t_SL g12647 ( 
.A(n_12518),
.Y(n_12647)
);

INVx2_ASAP7_75t_SL g12648 ( 
.A(n_12477),
.Y(n_12648)
);

INVx2_ASAP7_75t_L g12649 ( 
.A(n_12488),
.Y(n_12649)
);

NOR2xp33_ASAP7_75t_L g12650 ( 
.A(n_12539),
.B(n_2224),
.Y(n_12650)
);

INVx1_ASAP7_75t_L g12651 ( 
.A(n_12500),
.Y(n_12651)
);

OA22x2_ASAP7_75t_L g12652 ( 
.A1(n_12581),
.A2(n_12479),
.B1(n_12532),
.B2(n_12531),
.Y(n_12652)
);

INVx1_ASAP7_75t_L g12653 ( 
.A(n_12567),
.Y(n_12653)
);

NOR2x1_ASAP7_75t_L g12654 ( 
.A(n_12572),
.B(n_12605),
.Y(n_12654)
);

NOR2xp67_ASAP7_75t_L g12655 ( 
.A(n_12575),
.B(n_12458),
.Y(n_12655)
);

NOR2x1_ASAP7_75t_L g12656 ( 
.A(n_12573),
.B(n_12529),
.Y(n_12656)
);

AOI211x1_ASAP7_75t_L g12657 ( 
.A1(n_12636),
.A2(n_12544),
.B(n_12497),
.C(n_12506),
.Y(n_12657)
);

AOI211xp5_ASAP7_75t_L g12658 ( 
.A1(n_12578),
.A2(n_12599),
.B(n_12591),
.C(n_12634),
.Y(n_12658)
);

OAI22xp5_ASAP7_75t_L g12659 ( 
.A1(n_12615),
.A2(n_12547),
.B1(n_12505),
.B2(n_12541),
.Y(n_12659)
);

NAND2xp5_ASAP7_75t_L g12660 ( 
.A(n_12571),
.B(n_12481),
.Y(n_12660)
);

AOI22x1_ASAP7_75t_L g12661 ( 
.A1(n_12604),
.A2(n_12480),
.B1(n_12508),
.B2(n_12511),
.Y(n_12661)
);

NAND2x1_ASAP7_75t_L g12662 ( 
.A(n_12564),
.B(n_12520),
.Y(n_12662)
);

NAND4xp75_ASAP7_75t_L g12663 ( 
.A(n_12579),
.B(n_12449),
.C(n_12499),
.D(n_12542),
.Y(n_12663)
);

OAI22xp5_ASAP7_75t_L g12664 ( 
.A1(n_12592),
.A2(n_2227),
.B1(n_2225),
.B2(n_2226),
.Y(n_12664)
);

NAND4xp75_ASAP7_75t_L g12665 ( 
.A(n_12597),
.B(n_2228),
.C(n_2225),
.D(n_2226),
.Y(n_12665)
);

AOI21xp5_ASAP7_75t_L g12666 ( 
.A1(n_12566),
.A2(n_12570),
.B(n_12642),
.Y(n_12666)
);

INVxp67_ASAP7_75t_L g12667 ( 
.A(n_12585),
.Y(n_12667)
);

NOR3xp33_ASAP7_75t_SL g12668 ( 
.A(n_12582),
.B(n_2228),
.C(n_2230),
.Y(n_12668)
);

INVx1_ASAP7_75t_L g12669 ( 
.A(n_12577),
.Y(n_12669)
);

AO22x1_ASAP7_75t_L g12670 ( 
.A1(n_12583),
.A2(n_2232),
.B1(n_2230),
.B2(n_2231),
.Y(n_12670)
);

AOI22xp5_ASAP7_75t_L g12671 ( 
.A1(n_12648),
.A2(n_2240),
.B1(n_2248),
.B2(n_2231),
.Y(n_12671)
);

AOI21xp5_ASAP7_75t_L g12672 ( 
.A1(n_12609),
.A2(n_2241),
.B(n_2232),
.Y(n_12672)
);

AND2x2_ASAP7_75t_L g12673 ( 
.A(n_12584),
.B(n_2233),
.Y(n_12673)
);

AOI21xp5_ASAP7_75t_L g12674 ( 
.A1(n_12602),
.A2(n_2242),
.B(n_2233),
.Y(n_12674)
);

NOR3xp33_ASAP7_75t_L g12675 ( 
.A(n_12632),
.B(n_2237),
.C(n_2236),
.Y(n_12675)
);

NAND3xp33_ASAP7_75t_L g12676 ( 
.A(n_12629),
.B(n_12569),
.C(n_12650),
.Y(n_12676)
);

INVx1_ASAP7_75t_L g12677 ( 
.A(n_12588),
.Y(n_12677)
);

AOI211xp5_ASAP7_75t_L g12678 ( 
.A1(n_12639),
.A2(n_2238),
.B(n_2234),
.C(n_2237),
.Y(n_12678)
);

NAND2xp5_ASAP7_75t_L g12679 ( 
.A(n_12565),
.B(n_2234),
.Y(n_12679)
);

AOI22xp5_ASAP7_75t_L g12680 ( 
.A1(n_12590),
.A2(n_2248),
.B1(n_2257),
.B2(n_2239),
.Y(n_12680)
);

AOI21xp5_ASAP7_75t_L g12681 ( 
.A1(n_12593),
.A2(n_2250),
.B(n_2239),
.Y(n_12681)
);

INVx3_ASAP7_75t_L g12682 ( 
.A(n_12643),
.Y(n_12682)
);

AO21x1_ASAP7_75t_L g12683 ( 
.A1(n_12580),
.A2(n_2240),
.B(n_2241),
.Y(n_12683)
);

AOI21xp5_ASAP7_75t_SL g12684 ( 
.A1(n_12638),
.A2(n_2243),
.B(n_2244),
.Y(n_12684)
);

OAI21xp33_ASAP7_75t_L g12685 ( 
.A1(n_12622),
.A2(n_2243),
.B(n_2244),
.Y(n_12685)
);

OAI21xp33_ASAP7_75t_L g12686 ( 
.A1(n_12627),
.A2(n_2245),
.B(n_2246),
.Y(n_12686)
);

OAI21xp5_ASAP7_75t_SL g12687 ( 
.A1(n_12576),
.A2(n_2247),
.B(n_2246),
.Y(n_12687)
);

AOI21xp5_ASAP7_75t_L g12688 ( 
.A1(n_12595),
.A2(n_12644),
.B(n_12613),
.Y(n_12688)
);

INVx1_ASAP7_75t_L g12689 ( 
.A(n_12606),
.Y(n_12689)
);

NOR2xp33_ASAP7_75t_SL g12690 ( 
.A(n_12637),
.B(n_2245),
.Y(n_12690)
);

INVx1_ASAP7_75t_L g12691 ( 
.A(n_12630),
.Y(n_12691)
);

INVx1_ASAP7_75t_L g12692 ( 
.A(n_12598),
.Y(n_12692)
);

AOI22xp5_ASAP7_75t_L g12693 ( 
.A1(n_12647),
.A2(n_2257),
.B1(n_2265),
.B2(n_2247),
.Y(n_12693)
);

OA22x2_ASAP7_75t_L g12694 ( 
.A1(n_12626),
.A2(n_2252),
.B1(n_2250),
.B2(n_2251),
.Y(n_12694)
);

OAI21xp5_ASAP7_75t_SL g12695 ( 
.A1(n_12600),
.A2(n_2253),
.B(n_2252),
.Y(n_12695)
);

AOI21xp5_ASAP7_75t_L g12696 ( 
.A1(n_12611),
.A2(n_2262),
.B(n_2251),
.Y(n_12696)
);

NOR3x1_ASAP7_75t_L g12697 ( 
.A(n_12587),
.B(n_2254),
.C(n_2255),
.Y(n_12697)
);

AOI21xp5_ASAP7_75t_L g12698 ( 
.A1(n_12649),
.A2(n_2264),
.B(n_2255),
.Y(n_12698)
);

XNOR2xp5_ASAP7_75t_L g12699 ( 
.A(n_12568),
.B(n_2256),
.Y(n_12699)
);

OAI21xp5_ASAP7_75t_L g12700 ( 
.A1(n_12608),
.A2(n_2267),
.B(n_2258),
.Y(n_12700)
);

NOR3xp33_ASAP7_75t_L g12701 ( 
.A(n_12586),
.B(n_2261),
.C(n_2260),
.Y(n_12701)
);

OAI21xp33_ASAP7_75t_L g12702 ( 
.A1(n_12624),
.A2(n_2259),
.B(n_2262),
.Y(n_12702)
);

AOI22xp5_ASAP7_75t_L g12703 ( 
.A1(n_12620),
.A2(n_2274),
.B1(n_2283),
.B2(n_2263),
.Y(n_12703)
);

AOI21xp5_ASAP7_75t_L g12704 ( 
.A1(n_12616),
.A2(n_2275),
.B(n_2263),
.Y(n_12704)
);

NAND3xp33_ASAP7_75t_L g12705 ( 
.A(n_12619),
.B(n_2265),
.C(n_2266),
.Y(n_12705)
);

AOI211x1_ASAP7_75t_L g12706 ( 
.A1(n_12603),
.A2(n_2269),
.B(n_2266),
.C(n_2267),
.Y(n_12706)
);

NOR3x1_ASAP7_75t_L g12707 ( 
.A(n_12610),
.B(n_2270),
.C(n_2271),
.Y(n_12707)
);

AOI21xp5_ASAP7_75t_L g12708 ( 
.A1(n_12641),
.A2(n_2282),
.B(n_2270),
.Y(n_12708)
);

INVx1_ASAP7_75t_SL g12709 ( 
.A(n_12621),
.Y(n_12709)
);

NOR3x1_ASAP7_75t_L g12710 ( 
.A(n_12625),
.B(n_12614),
.C(n_12651),
.Y(n_12710)
);

INVx1_ASAP7_75t_L g12711 ( 
.A(n_12598),
.Y(n_12711)
);

AOI211xp5_ASAP7_75t_L g12712 ( 
.A1(n_12617),
.A2(n_2276),
.B(n_2272),
.C(n_2275),
.Y(n_12712)
);

NAND2xp5_ASAP7_75t_L g12713 ( 
.A(n_12623),
.B(n_2272),
.Y(n_12713)
);

OAI21xp5_ASAP7_75t_L g12714 ( 
.A1(n_12612),
.A2(n_2285),
.B(n_2276),
.Y(n_12714)
);

NAND2xp5_ASAP7_75t_L g12715 ( 
.A(n_12574),
.B(n_2277),
.Y(n_12715)
);

OA22x2_ASAP7_75t_L g12716 ( 
.A1(n_12596),
.A2(n_2281),
.B1(n_2278),
.B2(n_2279),
.Y(n_12716)
);

NAND3xp33_ASAP7_75t_SL g12717 ( 
.A(n_12658),
.B(n_12628),
.C(n_12618),
.Y(n_12717)
);

NOR3xp33_ASAP7_75t_L g12718 ( 
.A(n_12709),
.B(n_12640),
.C(n_12635),
.Y(n_12718)
);

OR2x2_ASAP7_75t_L g12719 ( 
.A(n_12679),
.B(n_12646),
.Y(n_12719)
);

NAND2xp5_ASAP7_75t_SL g12720 ( 
.A(n_12656),
.B(n_12607),
.Y(n_12720)
);

NOR2xp33_ASAP7_75t_L g12721 ( 
.A(n_12686),
.B(n_12594),
.Y(n_12721)
);

OAI21xp5_ASAP7_75t_L g12722 ( 
.A1(n_12666),
.A2(n_12633),
.B(n_12601),
.Y(n_12722)
);

NAND2xp5_ASAP7_75t_L g12723 ( 
.A(n_12673),
.B(n_12645),
.Y(n_12723)
);

INVx2_ASAP7_75t_SL g12724 ( 
.A(n_12654),
.Y(n_12724)
);

BUFx2_ASAP7_75t_L g12725 ( 
.A(n_12683),
.Y(n_12725)
);

AO22x2_ASAP7_75t_L g12726 ( 
.A1(n_12692),
.A2(n_12589),
.B1(n_12631),
.B2(n_2283),
.Y(n_12726)
);

NOR2x1_ASAP7_75t_L g12727 ( 
.A(n_12711),
.B(n_12665),
.Y(n_12727)
);

NOR2x1_ASAP7_75t_L g12728 ( 
.A(n_12684),
.B(n_2282),
.Y(n_12728)
);

NAND2xp5_ASAP7_75t_L g12729 ( 
.A(n_12699),
.B(n_12682),
.Y(n_12729)
);

XNOR2x2_ASAP7_75t_L g12730 ( 
.A(n_12657),
.B(n_2279),
.Y(n_12730)
);

NAND4xp25_ASAP7_75t_L g12731 ( 
.A(n_12697),
.B(n_2286),
.C(n_2284),
.D(n_2285),
.Y(n_12731)
);

NOR2x1_ASAP7_75t_L g12732 ( 
.A(n_12682),
.B(n_2287),
.Y(n_12732)
);

NOR2xp33_ASAP7_75t_L g12733 ( 
.A(n_12685),
.B(n_2284),
.Y(n_12733)
);

NOR3xp33_ASAP7_75t_L g12734 ( 
.A(n_12667),
.B(n_2287),
.C(n_2288),
.Y(n_12734)
);

NAND2xp5_ASAP7_75t_L g12735 ( 
.A(n_12678),
.B(n_2288),
.Y(n_12735)
);

AOI211xp5_ASAP7_75t_L g12736 ( 
.A1(n_12687),
.A2(n_2292),
.B(n_2289),
.C(n_2290),
.Y(n_12736)
);

NAND4xp75_ASAP7_75t_L g12737 ( 
.A(n_12710),
.B(n_2776),
.C(n_2777),
.D(n_2775),
.Y(n_12737)
);

OAI22xp5_ASAP7_75t_SL g12738 ( 
.A1(n_12706),
.A2(n_2293),
.B1(n_2289),
.B2(n_2292),
.Y(n_12738)
);

NOR3xp33_ASAP7_75t_L g12739 ( 
.A(n_12659),
.B(n_2293),
.C(n_2294),
.Y(n_12739)
);

AND2x2_ASAP7_75t_L g12740 ( 
.A(n_12668),
.B(n_2296),
.Y(n_12740)
);

NOR2xp33_ASAP7_75t_L g12741 ( 
.A(n_12690),
.B(n_2294),
.Y(n_12741)
);

AND2x2_ASAP7_75t_L g12742 ( 
.A(n_12677),
.B(n_2297),
.Y(n_12742)
);

NAND4xp75_ASAP7_75t_L g12743 ( 
.A(n_12655),
.B(n_2812),
.C(n_2785),
.D(n_2298),
.Y(n_12743)
);

INVx1_ASAP7_75t_L g12744 ( 
.A(n_12716),
.Y(n_12744)
);

AOI21xp5_ASAP7_75t_SL g12745 ( 
.A1(n_12700),
.A2(n_2785),
.B(n_2296),
.Y(n_12745)
);

OA21x2_ASAP7_75t_L g12746 ( 
.A1(n_12660),
.A2(n_12669),
.B(n_12653),
.Y(n_12746)
);

NOR3xp33_ASAP7_75t_L g12747 ( 
.A(n_12662),
.B(n_2297),
.C(n_2299),
.Y(n_12747)
);

INVx1_ASAP7_75t_L g12748 ( 
.A(n_12694),
.Y(n_12748)
);

NOR2x1_ASAP7_75t_L g12749 ( 
.A(n_12695),
.B(n_12676),
.Y(n_12749)
);

OA22x2_ASAP7_75t_L g12750 ( 
.A1(n_12691),
.A2(n_2307),
.B1(n_2317),
.B2(n_2299),
.Y(n_12750)
);

NOR2x1_ASAP7_75t_L g12751 ( 
.A(n_12689),
.B(n_2301),
.Y(n_12751)
);

NAND3xp33_ASAP7_75t_L g12752 ( 
.A(n_12712),
.B(n_2300),
.C(n_2302),
.Y(n_12752)
);

NAND2x1p5_ASAP7_75t_L g12753 ( 
.A(n_12707),
.B(n_2767),
.Y(n_12753)
);

AOI21xp5_ASAP7_75t_L g12754 ( 
.A1(n_12688),
.A2(n_2300),
.B(n_2302),
.Y(n_12754)
);

INVx1_ASAP7_75t_L g12755 ( 
.A(n_12702),
.Y(n_12755)
);

NAND5xp2_ASAP7_75t_L g12756 ( 
.A(n_12704),
.B(n_2305),
.C(n_2308),
.D(n_2304),
.E(n_2306),
.Y(n_12756)
);

INVx2_ASAP7_75t_L g12757 ( 
.A(n_12670),
.Y(n_12757)
);

NOR2xp33_ASAP7_75t_L g12758 ( 
.A(n_12705),
.B(n_2303),
.Y(n_12758)
);

NOR2xp33_ASAP7_75t_L g12759 ( 
.A(n_12663),
.B(n_2303),
.Y(n_12759)
);

INVx2_ASAP7_75t_L g12760 ( 
.A(n_12661),
.Y(n_12760)
);

NOR3xp33_ASAP7_75t_L g12761 ( 
.A(n_12664),
.B(n_2305),
.C(n_2306),
.Y(n_12761)
);

NAND4xp75_ASAP7_75t_L g12762 ( 
.A(n_12727),
.B(n_12732),
.C(n_12751),
.D(n_12749),
.Y(n_12762)
);

NAND2xp5_ASAP7_75t_L g12763 ( 
.A(n_12742),
.B(n_12741),
.Y(n_12763)
);

NAND3xp33_ASAP7_75t_SL g12764 ( 
.A(n_12739),
.B(n_12674),
.C(n_12708),
.Y(n_12764)
);

NAND2xp33_ASAP7_75t_L g12765 ( 
.A(n_12747),
.B(n_12701),
.Y(n_12765)
);

OR2x2_ASAP7_75t_L g12766 ( 
.A(n_12731),
.B(n_12715),
.Y(n_12766)
);

NOR2x1_ASAP7_75t_L g12767 ( 
.A(n_12737),
.B(n_12714),
.Y(n_12767)
);

NAND3xp33_ASAP7_75t_SL g12768 ( 
.A(n_12725),
.B(n_12675),
.C(n_12698),
.Y(n_12768)
);

NOR4xp25_ASAP7_75t_L g12769 ( 
.A(n_12717),
.B(n_12713),
.C(n_12652),
.D(n_12696),
.Y(n_12769)
);

OAI22xp5_ASAP7_75t_SL g12770 ( 
.A1(n_12753),
.A2(n_12738),
.B1(n_12728),
.B2(n_12736),
.Y(n_12770)
);

NAND2xp5_ASAP7_75t_L g12771 ( 
.A(n_12759),
.B(n_12681),
.Y(n_12771)
);

NAND4xp75_ASAP7_75t_L g12772 ( 
.A(n_12724),
.B(n_12672),
.C(n_12693),
.D(n_12671),
.Y(n_12772)
);

NOR3x1_ASAP7_75t_L g12773 ( 
.A(n_12743),
.B(n_12680),
.C(n_12703),
.Y(n_12773)
);

INVx2_ASAP7_75t_L g12774 ( 
.A(n_12750),
.Y(n_12774)
);

NAND3xp33_ASAP7_75t_L g12775 ( 
.A(n_12718),
.B(n_2308),
.C(n_2309),
.Y(n_12775)
);

INVx1_ASAP7_75t_SL g12776 ( 
.A(n_12740),
.Y(n_12776)
);

NOR2xp67_ASAP7_75t_L g12777 ( 
.A(n_12756),
.B(n_2312),
.Y(n_12777)
);

NAND3xp33_ASAP7_75t_SL g12778 ( 
.A(n_12754),
.B(n_2310),
.C(n_2312),
.Y(n_12778)
);

INVx1_ASAP7_75t_L g12779 ( 
.A(n_12730),
.Y(n_12779)
);

NAND4xp75_ASAP7_75t_L g12780 ( 
.A(n_12746),
.B(n_12720),
.C(n_12729),
.D(n_12722),
.Y(n_12780)
);

NOR2x1_ASAP7_75t_L g12781 ( 
.A(n_12745),
.B(n_2310),
.Y(n_12781)
);

NAND4xp25_ASAP7_75t_L g12782 ( 
.A(n_12721),
.B(n_12752),
.C(n_12744),
.D(n_12761),
.Y(n_12782)
);

NOR3x1_ASAP7_75t_L g12783 ( 
.A(n_12735),
.B(n_2313),
.C(n_2315),
.Y(n_12783)
);

INVx1_ASAP7_75t_L g12784 ( 
.A(n_12726),
.Y(n_12784)
);

NOR2xp67_ASAP7_75t_L g12785 ( 
.A(n_12757),
.B(n_2316),
.Y(n_12785)
);

NAND4xp75_ASAP7_75t_L g12786 ( 
.A(n_12746),
.B(n_2317),
.C(n_2315),
.D(n_2316),
.Y(n_12786)
);

AOI211xp5_ASAP7_75t_L g12787 ( 
.A1(n_12733),
.A2(n_2320),
.B(n_2318),
.C(n_2319),
.Y(n_12787)
);

NOR3xp33_ASAP7_75t_L g12788 ( 
.A(n_12760),
.B(n_2769),
.C(n_2768),
.Y(n_12788)
);

NAND4xp75_ASAP7_75t_L g12789 ( 
.A(n_12748),
.B(n_2321),
.C(n_2318),
.D(n_2319),
.Y(n_12789)
);

NOR2xp67_ASAP7_75t_L g12790 ( 
.A(n_12758),
.B(n_12723),
.Y(n_12790)
);

NOR3xp33_ASAP7_75t_L g12791 ( 
.A(n_12755),
.B(n_2773),
.C(n_2772),
.Y(n_12791)
);

NOR2x1_ASAP7_75t_L g12792 ( 
.A(n_12719),
.B(n_2322),
.Y(n_12792)
);

NAND2xp5_ASAP7_75t_SL g12793 ( 
.A(n_12734),
.B(n_2322),
.Y(n_12793)
);

AND4x1_ASAP7_75t_L g12794 ( 
.A(n_12726),
.B(n_2331),
.C(n_2340),
.D(n_2323),
.Y(n_12794)
);

OAI22xp5_ASAP7_75t_L g12795 ( 
.A1(n_12724),
.A2(n_2326),
.B1(n_2324),
.B2(n_2325),
.Y(n_12795)
);

NOR3xp33_ASAP7_75t_L g12796 ( 
.A(n_12717),
.B(n_2324),
.C(n_2327),
.Y(n_12796)
);

NAND4xp25_ASAP7_75t_SL g12797 ( 
.A(n_12736),
.B(n_2329),
.C(n_2327),
.D(n_2328),
.Y(n_12797)
);

NOR2x1_ASAP7_75t_L g12798 ( 
.A(n_12732),
.B(n_2329),
.Y(n_12798)
);

NOR3xp33_ASAP7_75t_L g12799 ( 
.A(n_12717),
.B(n_2764),
.C(n_2762),
.Y(n_12799)
);

AOI211xp5_ASAP7_75t_L g12800 ( 
.A1(n_12738),
.A2(n_2332),
.B(n_2330),
.C(n_2331),
.Y(n_12800)
);

NOR3xp33_ASAP7_75t_L g12801 ( 
.A(n_12717),
.B(n_2768),
.C(n_2766),
.Y(n_12801)
);

AOI21xp5_ASAP7_75t_L g12802 ( 
.A1(n_12720),
.A2(n_2333),
.B(n_2335),
.Y(n_12802)
);

AOI22xp5_ASAP7_75t_L g12803 ( 
.A1(n_12759),
.A2(n_2336),
.B1(n_2333),
.B2(n_2335),
.Y(n_12803)
);

HB1xp67_ASAP7_75t_L g12804 ( 
.A(n_12732),
.Y(n_12804)
);

NAND3xp33_ASAP7_75t_SL g12805 ( 
.A(n_12739),
.B(n_2336),
.C(n_2337),
.Y(n_12805)
);

NOR4xp75_ASAP7_75t_L g12806 ( 
.A(n_12720),
.B(n_2339),
.C(n_2337),
.D(n_2338),
.Y(n_12806)
);

AOI22xp33_ASAP7_75t_L g12807 ( 
.A1(n_12796),
.A2(n_12799),
.B1(n_12801),
.B2(n_12779),
.Y(n_12807)
);

BUFx2_ASAP7_75t_L g12808 ( 
.A(n_12798),
.Y(n_12808)
);

OAI211xp5_ASAP7_75t_L g12809 ( 
.A1(n_12800),
.A2(n_2781),
.B(n_2341),
.C(n_2338),
.Y(n_12809)
);

INVx1_ASAP7_75t_SL g12810 ( 
.A(n_12786),
.Y(n_12810)
);

NOR3x1_ASAP7_75t_L g12811 ( 
.A(n_12780),
.B(n_2339),
.C(n_2342),
.Y(n_12811)
);

INVx1_ASAP7_75t_L g12812 ( 
.A(n_12792),
.Y(n_12812)
);

OAI211xp5_ASAP7_75t_L g12813 ( 
.A1(n_12769),
.A2(n_2344),
.B(n_2342),
.C(n_2343),
.Y(n_12813)
);

AOI22xp5_ASAP7_75t_L g12814 ( 
.A1(n_12777),
.A2(n_2346),
.B1(n_2343),
.B2(n_2345),
.Y(n_12814)
);

OAI221xp5_ASAP7_75t_L g12815 ( 
.A1(n_12794),
.A2(n_2348),
.B1(n_2345),
.B2(n_2347),
.C(n_2349),
.Y(n_12815)
);

OAI221xp5_ASAP7_75t_L g12816 ( 
.A1(n_12788),
.A2(n_12785),
.B1(n_12775),
.B2(n_12781),
.C(n_12784),
.Y(n_12816)
);

AOI32xp33_ASAP7_75t_L g12817 ( 
.A1(n_12767),
.A2(n_2349),
.A3(n_2347),
.B1(n_2348),
.B2(n_2350),
.Y(n_12817)
);

O2A1O1Ixp33_ASAP7_75t_L g12818 ( 
.A1(n_12804),
.A2(n_2352),
.B(n_2354),
.C(n_2351),
.Y(n_12818)
);

OAI222xp33_ASAP7_75t_L g12819 ( 
.A1(n_12776),
.A2(n_2352),
.B1(n_2355),
.B2(n_2350),
.C1(n_2351),
.C2(n_2354),
.Y(n_12819)
);

OAI222xp33_ASAP7_75t_L g12820 ( 
.A1(n_12793),
.A2(n_2358),
.B1(n_2360),
.B2(n_2355),
.C1(n_2357),
.C2(n_2359),
.Y(n_12820)
);

AOI22x1_ASAP7_75t_L g12821 ( 
.A1(n_12802),
.A2(n_2362),
.B1(n_2358),
.B2(n_2361),
.Y(n_12821)
);

OAI221xp5_ASAP7_75t_L g12822 ( 
.A1(n_12782),
.A2(n_12803),
.B1(n_12787),
.B2(n_12774),
.C(n_12770),
.Y(n_12822)
);

O2A1O1Ixp5_ASAP7_75t_L g12823 ( 
.A1(n_12771),
.A2(n_12763),
.B(n_12766),
.C(n_12795),
.Y(n_12823)
);

AOI211xp5_ASAP7_75t_L g12824 ( 
.A1(n_12797),
.A2(n_2365),
.B(n_2363),
.C(n_2364),
.Y(n_12824)
);

OAI211xp5_ASAP7_75t_L g12825 ( 
.A1(n_12768),
.A2(n_2782),
.B(n_2760),
.C(n_2367),
.Y(n_12825)
);

AOI222xp33_ASAP7_75t_L g12826 ( 
.A1(n_12765),
.A2(n_2367),
.B1(n_2369),
.B2(n_2363),
.C1(n_2366),
.C2(n_2368),
.Y(n_12826)
);

OAI221xp5_ASAP7_75t_L g12827 ( 
.A1(n_12790),
.A2(n_2370),
.B1(n_2368),
.B2(n_2369),
.C(n_2371),
.Y(n_12827)
);

AOI211xp5_ASAP7_75t_L g12828 ( 
.A1(n_12805),
.A2(n_2375),
.B(n_2373),
.C(n_2374),
.Y(n_12828)
);

XNOR2xp5_ASAP7_75t_L g12829 ( 
.A(n_12806),
.B(n_2374),
.Y(n_12829)
);

AOI22xp33_ASAP7_75t_L g12830 ( 
.A1(n_12778),
.A2(n_2376),
.B1(n_2373),
.B2(n_2375),
.Y(n_12830)
);

AOI22xp5_ASAP7_75t_L g12831 ( 
.A1(n_12772),
.A2(n_2379),
.B1(n_2377),
.B2(n_2378),
.Y(n_12831)
);

OAI221xp5_ASAP7_75t_L g12832 ( 
.A1(n_12791),
.A2(n_2380),
.B1(n_2377),
.B2(n_2378),
.C(n_2381),
.Y(n_12832)
);

NAND2xp5_ASAP7_75t_L g12833 ( 
.A(n_12789),
.B(n_2380),
.Y(n_12833)
);

AOI211xp5_ASAP7_75t_L g12834 ( 
.A1(n_12764),
.A2(n_2386),
.B(n_2383),
.C(n_2385),
.Y(n_12834)
);

OAI22xp5_ASAP7_75t_L g12835 ( 
.A1(n_12762),
.A2(n_2386),
.B1(n_2383),
.B2(n_2385),
.Y(n_12835)
);

NAND3x1_ASAP7_75t_SL g12836 ( 
.A(n_12783),
.B(n_2387),
.C(n_2388),
.Y(n_12836)
);

AOI22xp5_ASAP7_75t_L g12837 ( 
.A1(n_12810),
.A2(n_12773),
.B1(n_2389),
.B2(n_2387),
.Y(n_12837)
);

AOI22xp5_ASAP7_75t_L g12838 ( 
.A1(n_12813),
.A2(n_2390),
.B1(n_2388),
.B2(n_2389),
.Y(n_12838)
);

INVx1_ASAP7_75t_L g12839 ( 
.A(n_12829),
.Y(n_12839)
);

INVx1_ASAP7_75t_L g12840 ( 
.A(n_12833),
.Y(n_12840)
);

NAND2xp5_ASAP7_75t_L g12841 ( 
.A(n_12831),
.B(n_12834),
.Y(n_12841)
);

AOI22xp33_ASAP7_75t_SL g12842 ( 
.A1(n_12821),
.A2(n_2392),
.B1(n_2390),
.B2(n_2391),
.Y(n_12842)
);

NAND2xp5_ASAP7_75t_SL g12843 ( 
.A(n_12814),
.B(n_2392),
.Y(n_12843)
);

INVx1_ASAP7_75t_L g12844 ( 
.A(n_12836),
.Y(n_12844)
);

INVx2_ASAP7_75t_L g12845 ( 
.A(n_12811),
.Y(n_12845)
);

INVx1_ASAP7_75t_L g12846 ( 
.A(n_12815),
.Y(n_12846)
);

NOR2x1_ASAP7_75t_L g12847 ( 
.A(n_12812),
.B(n_2393),
.Y(n_12847)
);

AOI211x1_ASAP7_75t_L g12848 ( 
.A1(n_12816),
.A2(n_12822),
.B(n_12809),
.C(n_12825),
.Y(n_12848)
);

NOR3xp33_ASAP7_75t_L g12849 ( 
.A(n_12823),
.B(n_2393),
.C(n_2395),
.Y(n_12849)
);

INVx1_ASAP7_75t_L g12850 ( 
.A(n_12808),
.Y(n_12850)
);

OAI21xp5_ASAP7_75t_SL g12851 ( 
.A1(n_12830),
.A2(n_2398),
.B(n_2397),
.Y(n_12851)
);

BUFx3_ASAP7_75t_L g12852 ( 
.A(n_12832),
.Y(n_12852)
);

INVx2_ASAP7_75t_L g12853 ( 
.A(n_12827),
.Y(n_12853)
);

INVx1_ASAP7_75t_L g12854 ( 
.A(n_12824),
.Y(n_12854)
);

AOI22xp33_ASAP7_75t_SL g12855 ( 
.A1(n_12835),
.A2(n_2399),
.B1(n_2396),
.B2(n_2397),
.Y(n_12855)
);

NOR3xp33_ASAP7_75t_L g12856 ( 
.A(n_12828),
.B(n_2396),
.C(n_2399),
.Y(n_12856)
);

HB1xp67_ASAP7_75t_L g12857 ( 
.A(n_12820),
.Y(n_12857)
);

OAI22xp5_ASAP7_75t_L g12858 ( 
.A1(n_12807),
.A2(n_2403),
.B1(n_2400),
.B2(n_2402),
.Y(n_12858)
);

INVx1_ASAP7_75t_L g12859 ( 
.A(n_12818),
.Y(n_12859)
);

AND2x2_ASAP7_75t_L g12860 ( 
.A(n_12826),
.B(n_2400),
.Y(n_12860)
);

AOI22xp5_ASAP7_75t_L g12861 ( 
.A1(n_12817),
.A2(n_2405),
.B1(n_2403),
.B2(n_2404),
.Y(n_12861)
);

NOR2x1_ASAP7_75t_L g12862 ( 
.A(n_12819),
.B(n_2404),
.Y(n_12862)
);

NAND2xp5_ASAP7_75t_L g12863 ( 
.A(n_12831),
.B(n_2766),
.Y(n_12863)
);

INVx1_ASAP7_75t_L g12864 ( 
.A(n_12829),
.Y(n_12864)
);

INVxp67_ASAP7_75t_L g12865 ( 
.A(n_12815),
.Y(n_12865)
);

AOI22xp5_ASAP7_75t_L g12866 ( 
.A1(n_12810),
.A2(n_2408),
.B1(n_2406),
.B2(n_2407),
.Y(n_12866)
);

NAND3xp33_ASAP7_75t_L g12867 ( 
.A(n_12849),
.B(n_2407),
.C(n_2408),
.Y(n_12867)
);

NOR3xp33_ASAP7_75t_SL g12868 ( 
.A(n_12850),
.B(n_2409),
.C(n_2410),
.Y(n_12868)
);

AOI22xp33_ASAP7_75t_L g12869 ( 
.A1(n_12856),
.A2(n_2412),
.B1(n_2409),
.B2(n_2411),
.Y(n_12869)
);

BUFx2_ASAP7_75t_L g12870 ( 
.A(n_12847),
.Y(n_12870)
);

AOI31xp33_ASAP7_75t_L g12871 ( 
.A1(n_12844),
.A2(n_2414),
.A3(n_2415),
.B(n_2413),
.Y(n_12871)
);

AOI211xp5_ASAP7_75t_L g12872 ( 
.A1(n_12851),
.A2(n_2414),
.B(n_2411),
.C(n_2413),
.Y(n_12872)
);

NAND2xp5_ASAP7_75t_L g12873 ( 
.A(n_12837),
.B(n_2416),
.Y(n_12873)
);

INVx1_ASAP7_75t_L g12874 ( 
.A(n_12838),
.Y(n_12874)
);

NOR4xp25_ASAP7_75t_L g12875 ( 
.A(n_12859),
.B(n_2782),
.C(n_2758),
.D(n_2419),
.Y(n_12875)
);

XNOR2xp5_ASAP7_75t_L g12876 ( 
.A(n_12848),
.B(n_2415),
.Y(n_12876)
);

INVx2_ASAP7_75t_L g12877 ( 
.A(n_12860),
.Y(n_12877)
);

AND3x4_ASAP7_75t_L g12878 ( 
.A(n_12862),
.B(n_2762),
.C(n_2761),
.Y(n_12878)
);

OAI22xp5_ASAP7_75t_SL g12879 ( 
.A1(n_12842),
.A2(n_2420),
.B1(n_2418),
.B2(n_2419),
.Y(n_12879)
);

NOR4xp25_ASAP7_75t_L g12880 ( 
.A(n_12839),
.B(n_2765),
.C(n_2422),
.D(n_2420),
.Y(n_12880)
);

AOI22xp5_ASAP7_75t_L g12881 ( 
.A1(n_12864),
.A2(n_2424),
.B1(n_2421),
.B2(n_2422),
.Y(n_12881)
);

AOI211x1_ASAP7_75t_L g12882 ( 
.A1(n_12843),
.A2(n_2426),
.B(n_2424),
.C(n_2425),
.Y(n_12882)
);

O2A1O1Ixp33_ASAP7_75t_L g12883 ( 
.A1(n_12857),
.A2(n_2429),
.B(n_2426),
.C(n_2427),
.Y(n_12883)
);

INVx2_ASAP7_75t_L g12884 ( 
.A(n_12845),
.Y(n_12884)
);

NOR2x1_ASAP7_75t_L g12885 ( 
.A(n_12854),
.B(n_2431),
.Y(n_12885)
);

NOR2x1_ASAP7_75t_L g12886 ( 
.A(n_12846),
.B(n_2431),
.Y(n_12886)
);

NAND2xp5_ASAP7_75t_L g12887 ( 
.A(n_12855),
.B(n_2433),
.Y(n_12887)
);

OAI22xp5_ASAP7_75t_L g12888 ( 
.A1(n_12861),
.A2(n_2757),
.B1(n_2758),
.B2(n_2756),
.Y(n_12888)
);

INVx1_ASAP7_75t_L g12889 ( 
.A(n_12863),
.Y(n_12889)
);

NAND2xp5_ASAP7_75t_L g12890 ( 
.A(n_12866),
.B(n_2434),
.Y(n_12890)
);

NOR3xp33_ASAP7_75t_L g12891 ( 
.A(n_12865),
.B(n_2430),
.C(n_2434),
.Y(n_12891)
);

OA22x2_ASAP7_75t_L g12892 ( 
.A1(n_12841),
.A2(n_2437),
.B1(n_2430),
.B2(n_2436),
.Y(n_12892)
);

BUFx2_ASAP7_75t_L g12893 ( 
.A(n_12852),
.Y(n_12893)
);

NOR3xp33_ASAP7_75t_L g12894 ( 
.A(n_12840),
.B(n_2436),
.C(n_2438),
.Y(n_12894)
);

OAI31xp33_ASAP7_75t_L g12895 ( 
.A1(n_12876),
.A2(n_12853),
.A3(n_12858),
.B(n_2440),
.Y(n_12895)
);

AND4x1_ASAP7_75t_L g12896 ( 
.A(n_12868),
.B(n_2440),
.C(n_2438),
.D(n_2439),
.Y(n_12896)
);

NAND3xp33_ASAP7_75t_SL g12897 ( 
.A(n_12878),
.B(n_2439),
.C(n_2441),
.Y(n_12897)
);

NAND2xp5_ASAP7_75t_L g12898 ( 
.A(n_12886),
.B(n_2441),
.Y(n_12898)
);

OAI221xp5_ASAP7_75t_L g12899 ( 
.A1(n_12869),
.A2(n_2444),
.B1(n_2442),
.B2(n_2443),
.C(n_2445),
.Y(n_12899)
);

NOR2x1p5_ASAP7_75t_L g12900 ( 
.A(n_12887),
.B(n_2443),
.Y(n_12900)
);

HB1xp67_ASAP7_75t_L g12901 ( 
.A(n_12892),
.Y(n_12901)
);

AND2x4_ASAP7_75t_L g12902 ( 
.A(n_12874),
.B(n_2444),
.Y(n_12902)
);

AOI21xp5_ASAP7_75t_L g12903 ( 
.A1(n_12870),
.A2(n_2445),
.B(n_2446),
.Y(n_12903)
);

INVx1_ASAP7_75t_L g12904 ( 
.A(n_12885),
.Y(n_12904)
);

NAND4xp75_ASAP7_75t_L g12905 ( 
.A(n_12882),
.B(n_2448),
.C(n_2446),
.D(n_2447),
.Y(n_12905)
);

AOI322xp5_ASAP7_75t_L g12906 ( 
.A1(n_12884),
.A2(n_2454),
.A3(n_2453),
.B1(n_2451),
.B2(n_2447),
.C1(n_2449),
.C2(n_2452),
.Y(n_12906)
);

AND2x4_ASAP7_75t_L g12907 ( 
.A(n_12877),
.B(n_2451),
.Y(n_12907)
);

AOI221xp5_ASAP7_75t_L g12908 ( 
.A1(n_12867),
.A2(n_2455),
.B1(n_2452),
.B2(n_2454),
.C(n_2456),
.Y(n_12908)
);

AOI21xp5_ASAP7_75t_L g12909 ( 
.A1(n_12873),
.A2(n_2455),
.B(n_2457),
.Y(n_12909)
);

AND2x4_ASAP7_75t_L g12910 ( 
.A(n_12893),
.B(n_2457),
.Y(n_12910)
);

AOI221xp5_ASAP7_75t_L g12911 ( 
.A1(n_12879),
.A2(n_2460),
.B1(n_2458),
.B2(n_2459),
.C(n_2463),
.Y(n_12911)
);

NAND3xp33_ASAP7_75t_SL g12912 ( 
.A(n_12872),
.B(n_2463),
.C(n_2464),
.Y(n_12912)
);

AOI221xp5_ASAP7_75t_L g12913 ( 
.A1(n_12888),
.A2(n_12880),
.B1(n_12875),
.B2(n_12890),
.C(n_12883),
.Y(n_12913)
);

OA22x2_ASAP7_75t_L g12914 ( 
.A1(n_12881),
.A2(n_12889),
.B1(n_12891),
.B2(n_12894),
.Y(n_12914)
);

INVx2_ASAP7_75t_L g12915 ( 
.A(n_12871),
.Y(n_12915)
);

NOR2x1_ASAP7_75t_SL g12916 ( 
.A(n_12867),
.B(n_2464),
.Y(n_12916)
);

AND3x2_ASAP7_75t_L g12917 ( 
.A(n_12870),
.B(n_2467),
.C(n_2466),
.Y(n_12917)
);

AOI21xp33_ASAP7_75t_SL g12918 ( 
.A1(n_12876),
.A2(n_2465),
.B(n_2466),
.Y(n_12918)
);

OAI211xp5_ASAP7_75t_L g12919 ( 
.A1(n_12886),
.A2(n_2470),
.B(n_2471),
.C(n_2469),
.Y(n_12919)
);

INVx1_ASAP7_75t_L g12920 ( 
.A(n_12898),
.Y(n_12920)
);

HB1xp67_ASAP7_75t_L g12921 ( 
.A(n_12896),
.Y(n_12921)
);

AO22x1_ASAP7_75t_L g12922 ( 
.A1(n_12904),
.A2(n_2470),
.B1(n_2472),
.B2(n_2469),
.Y(n_12922)
);

NAND4xp75_ASAP7_75t_L g12923 ( 
.A(n_12895),
.B(n_2473),
.C(n_2468),
.D(n_2472),
.Y(n_12923)
);

XNOR2xp5_ASAP7_75t_L g12924 ( 
.A(n_12905),
.B(n_2468),
.Y(n_12924)
);

AND2x2_ASAP7_75t_SL g12925 ( 
.A(n_12915),
.B(n_2473),
.Y(n_12925)
);

INVx1_ASAP7_75t_L g12926 ( 
.A(n_12900),
.Y(n_12926)
);

AND2x2_ASAP7_75t_L g12927 ( 
.A(n_12916),
.B(n_2474),
.Y(n_12927)
);

INVx1_ASAP7_75t_L g12928 ( 
.A(n_12907),
.Y(n_12928)
);

INVxp67_ASAP7_75t_L g12929 ( 
.A(n_12901),
.Y(n_12929)
);

XOR2x1_ASAP7_75t_L g12930 ( 
.A(n_12910),
.B(n_2475),
.Y(n_12930)
);

NAND2x1p5_ASAP7_75t_L g12931 ( 
.A(n_12902),
.B(n_12909),
.Y(n_12931)
);

XNOR2x1_ASAP7_75t_L g12932 ( 
.A(n_12914),
.B(n_2770),
.Y(n_12932)
);

INVx1_ASAP7_75t_L g12933 ( 
.A(n_12919),
.Y(n_12933)
);

INVx2_ASAP7_75t_L g12934 ( 
.A(n_12917),
.Y(n_12934)
);

INVx2_ASAP7_75t_L g12935 ( 
.A(n_12899),
.Y(n_12935)
);

OAI22xp5_ASAP7_75t_SL g12936 ( 
.A1(n_12924),
.A2(n_12897),
.B1(n_12918),
.B2(n_12912),
.Y(n_12936)
);

OAI22x1_ASAP7_75t_L g12937 ( 
.A1(n_12934),
.A2(n_12929),
.B1(n_12933),
.B2(n_12931),
.Y(n_12937)
);

BUFx4f_ASAP7_75t_SL g12938 ( 
.A(n_12920),
.Y(n_12938)
);

OAI22xp5_ASAP7_75t_L g12939 ( 
.A1(n_12932),
.A2(n_12911),
.B1(n_12908),
.B2(n_12913),
.Y(n_12939)
);

INVxp67_ASAP7_75t_SL g12940 ( 
.A(n_12930),
.Y(n_12940)
);

INVx2_ASAP7_75t_L g12941 ( 
.A(n_12925),
.Y(n_12941)
);

AO22x2_ASAP7_75t_L g12942 ( 
.A1(n_12923),
.A2(n_12928),
.B1(n_12926),
.B2(n_12935),
.Y(n_12942)
);

XNOR2xp5_ASAP7_75t_L g12943 ( 
.A(n_12921),
.B(n_12903),
.Y(n_12943)
);

INVx1_ASAP7_75t_L g12944 ( 
.A(n_12927),
.Y(n_12944)
);

OAI22x1_ASAP7_75t_L g12945 ( 
.A1(n_12922),
.A2(n_12906),
.B1(n_2477),
.B2(n_2475),
.Y(n_12945)
);

OAI21xp5_ASAP7_75t_L g12946 ( 
.A1(n_12929),
.A2(n_2476),
.B(n_2478),
.Y(n_12946)
);

AO21x2_ASAP7_75t_L g12947 ( 
.A1(n_12934),
.A2(n_2489),
.B(n_2479),
.Y(n_12947)
);

OAI22xp5_ASAP7_75t_L g12948 ( 
.A1(n_12929),
.A2(n_2481),
.B1(n_2479),
.B2(n_2480),
.Y(n_12948)
);

AND2x4_ASAP7_75t_L g12949 ( 
.A(n_12927),
.B(n_2480),
.Y(n_12949)
);

OAI22xp5_ASAP7_75t_L g12950 ( 
.A1(n_12929),
.A2(n_2483),
.B1(n_2481),
.B2(n_2482),
.Y(n_12950)
);

OAI22x1_ASAP7_75t_L g12951 ( 
.A1(n_12924),
.A2(n_2487),
.B1(n_2482),
.B2(n_2485),
.Y(n_12951)
);

HB1xp67_ASAP7_75t_L g12952 ( 
.A(n_12930),
.Y(n_12952)
);

INVx1_ASAP7_75t_L g12953 ( 
.A(n_12930),
.Y(n_12953)
);

HB1xp67_ASAP7_75t_L g12954 ( 
.A(n_12947),
.Y(n_12954)
);

AOI22xp5_ASAP7_75t_L g12955 ( 
.A1(n_12949),
.A2(n_2496),
.B1(n_2504),
.B2(n_2485),
.Y(n_12955)
);

INVx1_ASAP7_75t_L g12956 ( 
.A(n_12951),
.Y(n_12956)
);

OAI22xp33_ASAP7_75t_L g12957 ( 
.A1(n_12938),
.A2(n_2759),
.B1(n_2764),
.B2(n_2757),
.Y(n_12957)
);

AO22x2_ASAP7_75t_L g12958 ( 
.A1(n_12939),
.A2(n_12953),
.B1(n_12941),
.B2(n_12944),
.Y(n_12958)
);

CKINVDCx20_ASAP7_75t_R g12959 ( 
.A(n_12936),
.Y(n_12959)
);

INVxp67_ASAP7_75t_L g12960 ( 
.A(n_12952),
.Y(n_12960)
);

AO22x2_ASAP7_75t_L g12961 ( 
.A1(n_12940),
.A2(n_2489),
.B1(n_2487),
.B2(n_2488),
.Y(n_12961)
);

OAI22xp5_ASAP7_75t_L g12962 ( 
.A1(n_12943),
.A2(n_2491),
.B1(n_2488),
.B2(n_2490),
.Y(n_12962)
);

INVx1_ASAP7_75t_L g12963 ( 
.A(n_12945),
.Y(n_12963)
);

AOI22xp33_ASAP7_75t_L g12964 ( 
.A1(n_12937),
.A2(n_2494),
.B1(n_2491),
.B2(n_2493),
.Y(n_12964)
);

AOI22xp5_ASAP7_75t_L g12965 ( 
.A1(n_12942),
.A2(n_2503),
.B1(n_2513),
.B2(n_2493),
.Y(n_12965)
);

INVx1_ASAP7_75t_L g12966 ( 
.A(n_12942),
.Y(n_12966)
);

OAI22x1_ASAP7_75t_L g12967 ( 
.A1(n_12946),
.A2(n_2498),
.B1(n_2494),
.B2(n_2497),
.Y(n_12967)
);

INVxp67_ASAP7_75t_SL g12968 ( 
.A(n_12948),
.Y(n_12968)
);

AO22x2_ASAP7_75t_L g12969 ( 
.A1(n_12950),
.A2(n_2500),
.B1(n_2497),
.B2(n_2499),
.Y(n_12969)
);

INVx2_ASAP7_75t_L g12970 ( 
.A(n_12947),
.Y(n_12970)
);

AOI22xp5_ASAP7_75t_L g12971 ( 
.A1(n_12949),
.A2(n_2511),
.B1(n_2519),
.B2(n_2500),
.Y(n_12971)
);

NAND4xp25_ASAP7_75t_L g12972 ( 
.A(n_12966),
.B(n_2505),
.C(n_2501),
.D(n_2502),
.Y(n_12972)
);

OR4x1_ASAP7_75t_L g12973 ( 
.A(n_12963),
.B(n_2506),
.C(n_2501),
.D(n_2505),
.Y(n_12973)
);

OAI222xp33_ASAP7_75t_L g12974 ( 
.A1(n_12960),
.A2(n_2508),
.B1(n_2511),
.B2(n_2506),
.C1(n_2507),
.C2(n_2510),
.Y(n_12974)
);

NOR2x1_ASAP7_75t_L g12975 ( 
.A(n_12970),
.B(n_2507),
.Y(n_12975)
);

OR3x1_ASAP7_75t_L g12976 ( 
.A(n_12956),
.B(n_2513),
.C(n_2512),
.Y(n_12976)
);

XOR2xp5_ASAP7_75t_L g12977 ( 
.A(n_12959),
.B(n_2508),
.Y(n_12977)
);

OR3x1_ASAP7_75t_L g12978 ( 
.A(n_12958),
.B(n_2515),
.C(n_2514),
.Y(n_12978)
);

OAI22xp5_ASAP7_75t_L g12979 ( 
.A1(n_12965),
.A2(n_2516),
.B1(n_2512),
.B2(n_2515),
.Y(n_12979)
);

NAND3xp33_ASAP7_75t_SL g12980 ( 
.A(n_12954),
.B(n_2516),
.C(n_2517),
.Y(n_12980)
);

NOR3xp33_ASAP7_75t_L g12981 ( 
.A(n_12968),
.B(n_2518),
.C(n_2520),
.Y(n_12981)
);

NOR3xp33_ASAP7_75t_L g12982 ( 
.A(n_12957),
.B(n_2520),
.C(n_2521),
.Y(n_12982)
);

OAI221xp5_ASAP7_75t_R g12983 ( 
.A1(n_12964),
.A2(n_2524),
.B1(n_2522),
.B2(n_2523),
.C(n_2525),
.Y(n_12983)
);

NOR3xp33_ASAP7_75t_L g12984 ( 
.A(n_12962),
.B(n_2522),
.C(n_2523),
.Y(n_12984)
);

AND2x2_ASAP7_75t_L g12985 ( 
.A(n_12969),
.B(n_2525),
.Y(n_12985)
);

XOR2x2_ASAP7_75t_L g12986 ( 
.A(n_12975),
.B(n_12955),
.Y(n_12986)
);

AOI21xp33_ASAP7_75t_L g12987 ( 
.A1(n_12985),
.A2(n_12967),
.B(n_12971),
.Y(n_12987)
);

INVx1_ASAP7_75t_L g12988 ( 
.A(n_12978),
.Y(n_12988)
);

INVx1_ASAP7_75t_L g12989 ( 
.A(n_12976),
.Y(n_12989)
);

INVx3_ASAP7_75t_L g12990 ( 
.A(n_12983),
.Y(n_12990)
);

INVx1_ASAP7_75t_L g12991 ( 
.A(n_12982),
.Y(n_12991)
);

INVx1_ASAP7_75t_L g12992 ( 
.A(n_12984),
.Y(n_12992)
);

AOI22x1_ASAP7_75t_L g12993 ( 
.A1(n_12977),
.A2(n_12961),
.B1(n_2529),
.B2(n_2527),
.Y(n_12993)
);

NOR3xp33_ASAP7_75t_L g12994 ( 
.A(n_12980),
.B(n_12961),
.C(n_2527),
.Y(n_12994)
);

AND2x2_ASAP7_75t_L g12995 ( 
.A(n_12979),
.B(n_12981),
.Y(n_12995)
);

XNOR2x1_ASAP7_75t_L g12996 ( 
.A(n_12973),
.B(n_2528),
.Y(n_12996)
);

INVx2_ASAP7_75t_L g12997 ( 
.A(n_12972),
.Y(n_12997)
);

AND2x4_ASAP7_75t_L g12998 ( 
.A(n_12974),
.B(n_2528),
.Y(n_12998)
);

BUFx2_ASAP7_75t_L g12999 ( 
.A(n_12975),
.Y(n_12999)
);

BUFx6f_ASAP7_75t_L g13000 ( 
.A(n_12999),
.Y(n_13000)
);

OAI22xp5_ASAP7_75t_SL g13001 ( 
.A1(n_12989),
.A2(n_2531),
.B1(n_2529),
.B2(n_2530),
.Y(n_13001)
);

OAI22xp5_ASAP7_75t_SL g13002 ( 
.A1(n_12988),
.A2(n_2533),
.B1(n_2531),
.B2(n_2532),
.Y(n_13002)
);

AOI21xp5_ASAP7_75t_L g13003 ( 
.A1(n_12987),
.A2(n_2533),
.B(n_2534),
.Y(n_13003)
);

OAI22xp5_ASAP7_75t_SL g13004 ( 
.A1(n_12997),
.A2(n_2536),
.B1(n_2534),
.B2(n_2535),
.Y(n_13004)
);

OAI22xp5_ASAP7_75t_L g13005 ( 
.A1(n_12993),
.A2(n_2538),
.B1(n_2535),
.B2(n_2537),
.Y(n_13005)
);

OAI22x1_ASAP7_75t_L g13006 ( 
.A1(n_12991),
.A2(n_2539),
.B1(n_2541),
.B2(n_2538),
.Y(n_13006)
);

OAI22xp5_ASAP7_75t_SL g13007 ( 
.A1(n_12992),
.A2(n_2542),
.B1(n_2537),
.B2(n_2541),
.Y(n_13007)
);

CKINVDCx20_ASAP7_75t_R g13008 ( 
.A(n_12986),
.Y(n_13008)
);

XOR2xp5_ASAP7_75t_L g13009 ( 
.A(n_13008),
.B(n_12996),
.Y(n_13009)
);

NAND2xp5_ASAP7_75t_L g13010 ( 
.A(n_13005),
.B(n_12994),
.Y(n_13010)
);

AOI21xp5_ASAP7_75t_SL g13011 ( 
.A1(n_13000),
.A2(n_12998),
.B(n_12995),
.Y(n_13011)
);

OR2x2_ASAP7_75t_L g13012 ( 
.A(n_13000),
.B(n_12990),
.Y(n_13012)
);

INVx1_ASAP7_75t_L g13013 ( 
.A(n_13003),
.Y(n_13013)
);

NOR2xp33_ASAP7_75t_L g13014 ( 
.A(n_13004),
.B(n_2542),
.Y(n_13014)
);

NAND2xp5_ASAP7_75t_L g13015 ( 
.A(n_13014),
.B(n_13006),
.Y(n_13015)
);

XNOR2xp5_ASAP7_75t_L g13016 ( 
.A(n_13009),
.B(n_13001),
.Y(n_13016)
);

OAI22xp5_ASAP7_75t_L g13017 ( 
.A1(n_13012),
.A2(n_13002),
.B1(n_13007),
.B2(n_2545),
.Y(n_13017)
);

XNOR2xp5_ASAP7_75t_L g13018 ( 
.A(n_13010),
.B(n_2543),
.Y(n_13018)
);

AOI22xp5_ASAP7_75t_L g13019 ( 
.A1(n_13013),
.A2(n_2546),
.B1(n_2547),
.B2(n_2544),
.Y(n_13019)
);

XOR2xp5_ASAP7_75t_L g13020 ( 
.A(n_13011),
.B(n_2543),
.Y(n_13020)
);

NAND2xp5_ASAP7_75t_L g13021 ( 
.A(n_13017),
.B(n_2544),
.Y(n_13021)
);

NAND2xp5_ASAP7_75t_SL g13022 ( 
.A(n_13015),
.B(n_13016),
.Y(n_13022)
);

AO21x2_ASAP7_75t_L g13023 ( 
.A1(n_13020),
.A2(n_2546),
.B(n_2547),
.Y(n_13023)
);

AOI21xp5_ASAP7_75t_L g13024 ( 
.A1(n_13018),
.A2(n_2548),
.B(n_2550),
.Y(n_13024)
);

XNOR2xp5_ASAP7_75t_L g13025 ( 
.A(n_13019),
.B(n_2550),
.Y(n_13025)
);

NOR2xp33_ASAP7_75t_L g13026 ( 
.A(n_13022),
.B(n_2548),
.Y(n_13026)
);

OAI21xp5_ASAP7_75t_L g13027 ( 
.A1(n_13025),
.A2(n_2551),
.B(n_2552),
.Y(n_13027)
);

AOI22xp5_ASAP7_75t_SL g13028 ( 
.A1(n_13027),
.A2(n_13021),
.B1(n_13024),
.B2(n_13023),
.Y(n_13028)
);

AOI22xp5_ASAP7_75t_L g13029 ( 
.A1(n_13026),
.A2(n_2553),
.B1(n_2551),
.B2(n_2552),
.Y(n_13029)
);

AO21x2_ASAP7_75t_L g13030 ( 
.A1(n_13028),
.A2(n_2555),
.B(n_2556),
.Y(n_13030)
);

OA21x2_ASAP7_75t_L g13031 ( 
.A1(n_13029),
.A2(n_2555),
.B(n_2557),
.Y(n_13031)
);

AOI22xp5_ASAP7_75t_L g13032 ( 
.A1(n_13031),
.A2(n_2559),
.B1(n_2560),
.B2(n_2558),
.Y(n_13032)
);

AOI21xp33_ASAP7_75t_SL g13033 ( 
.A1(n_13032),
.A2(n_13030),
.B(n_2755),
.Y(n_13033)
);

AOI211xp5_ASAP7_75t_L g13034 ( 
.A1(n_13033),
.A2(n_2559),
.B(n_2557),
.C(n_2558),
.Y(n_13034)
);


endmodule