module fake_jpeg_14702_n_351 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_351);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_351;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx10_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx4f_ASAP7_75t_SL g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_22),
.B(n_7),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_33),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_50),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_53),
.B(n_36),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_25),
.Y(n_54)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_25),
.Y(n_55)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_18),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_57),
.B(n_18),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_30),
.Y(n_58)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_68),
.B(n_19),
.Y(n_100)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_71),
.Y(n_108)
);

INVx2_ASAP7_75t_SL g73 ( 
.A(n_48),
.Y(n_73)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_73),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g76 ( 
.A(n_56),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_76),
.B(n_85),
.Y(n_115)
);

HB1xp67_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_77),
.Y(n_137)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_79),
.Y(n_112)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_80),
.Y(n_111)
);

INVx2_ASAP7_75t_SL g81 ( 
.A(n_66),
.Y(n_81)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_81),
.Y(n_114)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_84),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_64),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_86),
.Y(n_119)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_87),
.Y(n_129)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_88),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_89),
.B(n_100),
.Y(n_110)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_90),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_57),
.A2(n_32),
.B1(n_28),
.B2(n_30),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_93),
.A2(n_33),
.B1(n_21),
.B2(n_24),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_63),
.A2(n_20),
.B(n_29),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_94),
.A2(n_26),
.B(n_18),
.Y(n_120)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_53),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_95),
.B(n_98),
.Y(n_124)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_96),
.Y(n_130)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_60),
.Y(n_97)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_97),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_70),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_65),
.Y(n_99)
);

BUFx4f_ASAP7_75t_SL g123 ( 
.A(n_99),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_62),
.A2(n_32),
.B1(n_41),
.B2(n_39),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_101),
.A2(n_28),
.B1(n_69),
.B2(n_26),
.Y(n_132)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_73),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_102),
.B(n_104),
.Y(n_126)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_60),
.Y(n_103)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_103),
.Y(n_134)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_74),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_61),
.Y(n_105)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_105),
.Y(n_138)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_63),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_106),
.B(n_107),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_69),
.B(n_22),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_94),
.B(n_48),
.C(n_50),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_109),
.B(n_120),
.C(n_118),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_76),
.B(n_48),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_113),
.B(n_122),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_116),
.B(n_136),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_101),
.A2(n_61),
.B1(n_74),
.B2(n_49),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_118),
.A2(n_132),
.B1(n_84),
.B2(n_81),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_120),
.A2(n_26),
.B(n_35),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_91),
.B(n_27),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_75),
.B(n_24),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_127),
.B(n_131),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_106),
.A2(n_28),
.B1(n_32),
.B2(n_33),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_128),
.A2(n_78),
.B1(n_82),
.B2(n_108),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_83),
.B(n_19),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_92),
.B(n_31),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_138),
.Y(n_139)
);

INVxp67_ASAP7_75t_SL g201 ( 
.A(n_139),
.Y(n_201)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_112),
.Y(n_140)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_140),
.Y(n_174)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_112),
.Y(n_141)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_141),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_115),
.B(n_108),
.Y(n_142)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_142),
.Y(n_206)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_129),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_143),
.Y(n_192)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_129),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_144),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_147),
.B(n_152),
.C(n_162),
.Y(n_185)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_123),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_148),
.B(n_155),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_149),
.A2(n_159),
.B1(n_165),
.B2(n_117),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_109),
.B(n_0),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_151),
.A2(n_156),
.B(n_119),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_122),
.B(n_47),
.C(n_51),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_110),
.B(n_31),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_153),
.B(n_157),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_110),
.B(n_80),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_154),
.B(n_158),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_138),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_115),
.B(n_35),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_135),
.B(n_86),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_127),
.B(n_99),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_160),
.B(n_166),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_113),
.A2(n_17),
.B(n_27),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_161),
.A2(n_119),
.B(n_121),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_116),
.B(n_29),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_135),
.B(n_23),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_163),
.B(n_167),
.Y(n_177)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_124),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_164),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_132),
.A2(n_82),
.B1(n_40),
.B2(n_43),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_131),
.B(n_99),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_130),
.B(n_27),
.Y(n_167)
);

MAJx2_ASAP7_75t_L g168 ( 
.A(n_130),
.B(n_29),
.C(n_17),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_168),
.B(n_161),
.C(n_162),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_136),
.B(n_16),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_169),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_126),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_170),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_126),
.B(n_27),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_171),
.B(n_123),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_147),
.B(n_124),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_173),
.B(n_179),
.C(n_200),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_175),
.A2(n_183),
.B1(n_186),
.B2(n_199),
.Y(n_212)
);

AO22x1_ASAP7_75t_L g176 ( 
.A1(n_149),
.A2(n_138),
.B1(n_114),
.B2(n_111),
.Y(n_176)
);

OA21x2_ASAP7_75t_L g229 ( 
.A1(n_176),
.A2(n_182),
.B(n_16),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_178),
.B(n_180),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_150),
.B(n_137),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_150),
.B(n_137),
.Y(n_180)
);

AO22x1_ASAP7_75t_L g182 ( 
.A1(n_168),
.A2(n_114),
.B1(n_111),
.B2(n_40),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_151),
.A2(n_117),
.B1(n_133),
.B2(n_134),
.Y(n_183)
);

AOI32xp33_ASAP7_75t_L g184 ( 
.A1(n_146),
.A2(n_123),
.A3(n_70),
.B1(n_71),
.B2(n_51),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_184),
.B(n_148),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_164),
.A2(n_134),
.B1(n_133),
.B2(n_125),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_187),
.B(n_29),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_190),
.A2(n_193),
.B(n_178),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_191),
.A2(n_193),
.B(n_144),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_158),
.A2(n_123),
.B(n_125),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_154),
.B(n_121),
.Y(n_197)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_197),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_140),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_198),
.B(n_42),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_151),
.A2(n_152),
.B1(n_167),
.B2(n_165),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_163),
.B(n_105),
.C(n_43),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_156),
.B(n_27),
.Y(n_204)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_204),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_171),
.B(n_17),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_205),
.B(n_187),
.C(n_185),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_207),
.A2(n_210),
.B(n_216),
.Y(n_239)
);

NAND3xp33_ASAP7_75t_L g209 ( 
.A(n_203),
.B(n_196),
.C(n_180),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_209),
.B(n_231),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_190),
.A2(n_141),
.B(n_143),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_213),
.B(n_219),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_173),
.B(n_155),
.C(n_139),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_215),
.B(n_217),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_185),
.B(n_145),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_172),
.A2(n_197),
.B(n_204),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_218),
.A2(n_226),
.B1(n_235),
.B2(n_201),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_179),
.B(n_172),
.C(n_205),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_174),
.Y(n_220)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_220),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g244 ( 
.A(n_221),
.B(n_227),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_199),
.B(n_42),
.C(n_17),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_222),
.B(n_230),
.Y(n_245)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_181),
.Y(n_223)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_223),
.Y(n_249)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_224),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_194),
.B(n_16),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_225),
.B(n_228),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_189),
.A2(n_95),
.B1(n_17),
.B2(n_29),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_206),
.B(n_16),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_229),
.B(n_183),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_177),
.B(n_16),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_200),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_189),
.B(n_16),
.Y(n_232)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_232),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_177),
.B(n_14),
.C(n_13),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_233),
.B(n_8),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_202),
.B(n_15),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_234),
.B(n_9),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_176),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_212),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_237),
.B(n_241),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_231),
.A2(n_176),
.B1(n_195),
.B2(n_182),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_238),
.A2(n_246),
.B1(n_251),
.B2(n_254),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g241 ( 
.A(n_226),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_214),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_243),
.B(n_253),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_208),
.A2(n_195),
.B1(n_182),
.B2(n_188),
.Y(n_246)
);

CKINVDCx14_ASAP7_75t_R g272 ( 
.A(n_252),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_214),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_236),
.A2(n_191),
.B1(n_192),
.B2(n_198),
.Y(n_254)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_255),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_212),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_257)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_257),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_233),
.B(n_8),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_258),
.B(n_260),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_218),
.B(n_9),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_261),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_211),
.B(n_219),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_262),
.B(n_213),
.C(n_215),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_240),
.B(n_211),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_263),
.B(n_267),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_264),
.B(n_269),
.C(n_270),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_237),
.A2(n_222),
.B1(n_221),
.B2(n_207),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_265),
.A2(n_241),
.B1(n_238),
.B2(n_255),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_240),
.B(n_217),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_248),
.B(n_262),
.C(n_245),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_248),
.B(n_227),
.C(n_230),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_259),
.B(n_235),
.Y(n_273)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_273),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_245),
.B(n_210),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_275),
.B(n_279),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_249),
.B(n_229),
.Y(n_277)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_277),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_244),
.B(n_239),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_244),
.B(n_229),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_280),
.B(n_257),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_239),
.A2(n_15),
.B(n_14),
.Y(n_282)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_282),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_242),
.B(n_1),
.C(n_3),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_283),
.B(n_260),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_284),
.A2(n_297),
.B1(n_280),
.B2(n_279),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_272),
.B(n_256),
.Y(n_286)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_286),
.Y(n_303)
);

FAx1_ASAP7_75t_SL g289 ( 
.A(n_268),
.B(n_254),
.CI(n_246),
.CON(n_289),
.SN(n_289)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_289),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_290),
.B(n_293),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_291),
.B(n_292),
.Y(n_305)
);

NOR3xp33_ASAP7_75t_SL g292 ( 
.A(n_278),
.B(n_250),
.C(n_283),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_269),
.B(n_247),
.Y(n_293)
);

HB1xp67_ASAP7_75t_L g294 ( 
.A(n_266),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_294),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_271),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_275),
.B(n_10),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_298),
.B(n_290),
.Y(n_313)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_276),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_300),
.B(n_15),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_285),
.B(n_264),
.C(n_263),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_301),
.B(n_310),
.C(n_287),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_299),
.A2(n_284),
.B(n_265),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_302),
.B(n_306),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_296),
.A2(n_274),
.B1(n_281),
.B2(n_270),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_307),
.A2(n_5),
.B1(n_6),
.B2(n_313),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_285),
.B(n_267),
.C(n_4),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_308),
.B(n_311),
.C(n_6),
.Y(n_327)
);

HB1xp67_ASAP7_75t_L g309 ( 
.A(n_295),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_309),
.B(n_289),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_293),
.B(n_13),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_287),
.B(n_288),
.C(n_298),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_313),
.B(n_288),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_314),
.B(n_6),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_317),
.B(n_312),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_318),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_319),
.B(n_320),
.C(n_321),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_315),
.A2(n_292),
.B1(n_4),
.B2(n_5),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_301),
.B(n_3),
.C(n_4),
.Y(n_321)
);

INVx11_ASAP7_75t_L g322 ( 
.A(n_304),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_322),
.B(n_323),
.Y(n_331)
);

INVx13_ASAP7_75t_L g324 ( 
.A(n_304),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_324),
.B(n_325),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_303),
.B(n_3),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_326),
.B(n_327),
.C(n_310),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_321),
.B(n_308),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_328),
.B(n_332),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_325),
.B(n_305),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_333),
.B(n_336),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_334),
.B(n_317),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_327),
.B(n_312),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_335),
.B(n_320),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_338),
.B(n_341),
.C(n_342),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_329),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_340),
.A2(n_331),
.B(n_330),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_329),
.B(n_322),
.Y(n_342)
);

NAND3xp33_ASAP7_75t_L g346 ( 
.A(n_343),
.B(n_344),
.C(n_337),
.Y(n_346)
);

INVxp67_ASAP7_75t_SL g344 ( 
.A(n_340),
.Y(n_344)
);

A2O1A1Ixp33_ASAP7_75t_SL g347 ( 
.A1(n_346),
.A2(n_339),
.B(n_316),
.C(n_324),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_347),
.B(n_345),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_348),
.B(n_319),
.C(n_334),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_349),
.B(n_311),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_350),
.B(n_326),
.Y(n_351)
);


endmodule