module real_jpeg_13862_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_298, n_12, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_298;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_288;
wire n_215;
wire n_166;
wire n_176;
wire n_292;
wire n_221;
wire n_249;
wire n_286;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_105;
wire n_40;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_293;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_294;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_134;
wire n_270;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_195;
wire n_110;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_150;
wire n_70;
wire n_41;
wire n_74;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_225;
wire n_103;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_279;
wire n_216;
wire n_295;
wire n_167;
wire n_128;
wire n_202;
wire n_179;
wire n_133;
wire n_213;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_273;
wire n_96;
wire n_269;
wire n_253;
wire n_89;

BUFx10_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_1),
.A2(n_29),
.B1(n_36),
.B2(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_1),
.A2(n_39),
.B1(n_44),
.B2(n_45),
.Y(n_113)
);

BUFx16f_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_3),
.A2(n_44),
.B1(n_45),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_3),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_3),
.A2(n_29),
.B1(n_36),
.B2(n_54),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_3),
.A2(n_54),
.B1(n_61),
.B2(n_64),
.Y(n_110)
);

BUFx12_ASAP7_75t_L g68 ( 
.A(n_4),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_5),
.A2(n_66),
.B1(n_67),
.B2(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_5),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_5),
.A2(n_61),
.B1(n_64),
.B2(n_72),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_5),
.A2(n_44),
.B1(n_45),
.B2(n_72),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_5),
.A2(n_29),
.B1(n_36),
.B2(n_72),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_7),
.A2(n_66),
.B1(n_67),
.B2(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_7),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_7),
.A2(n_61),
.B1(n_64),
.B2(n_150),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_7),
.A2(n_44),
.B1(n_45),
.B2(n_150),
.Y(n_216)
);

OAI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_7),
.A2(n_29),
.B1(n_36),
.B2(n_150),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_8),
.A2(n_29),
.B1(n_36),
.B2(n_37),
.Y(n_35)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_8),
.A2(n_37),
.B1(n_44),
.B2(n_45),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g289 ( 
.A1(n_8),
.A2(n_37),
.B1(n_61),
.B2(n_64),
.Y(n_289)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_9),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_10),
.A2(n_66),
.B1(n_67),
.B2(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_10),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_10),
.A2(n_61),
.B1(n_64),
.B2(n_104),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_10),
.A2(n_44),
.B1(n_45),
.B2(n_104),
.Y(n_223)
);

OAI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_10),
.A2(n_29),
.B1(n_36),
.B2(n_104),
.Y(n_230)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_11),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_12),
.A2(n_66),
.B1(n_67),
.B2(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_12),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_12),
.A2(n_61),
.B1(n_64),
.B2(n_70),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_12),
.A2(n_44),
.B1(n_45),
.B2(n_70),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_12),
.A2(n_29),
.B1(n_36),
.B2(n_70),
.Y(n_225)
);

BUFx8_ASAP7_75t_L g63 ( 
.A(n_13),
.Y(n_63)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_14),
.Y(n_142)
);

AOI21xp33_ASAP7_75t_L g169 ( 
.A1(n_14),
.A2(n_66),
.B(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_14),
.B(n_153),
.Y(n_184)
);

OAI22xp33_ASAP7_75t_L g215 ( 
.A1(n_14),
.A2(n_44),
.B1(n_45),
.B2(n_142),
.Y(n_215)
);

O2A1O1Ixp33_ASAP7_75t_L g217 ( 
.A1(n_14),
.A2(n_44),
.B(n_50),
.C(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_14),
.B(n_111),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_14),
.B(n_33),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_14),
.B(n_55),
.Y(n_242)
);

A2O1A1Ixp33_ASAP7_75t_L g251 ( 
.A1(n_14),
.A2(n_64),
.B(n_75),
.C(n_252),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_15),
.A2(n_61),
.B1(n_64),
.B2(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_15),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_15),
.A2(n_44),
.B1(n_45),
.B2(n_81),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_15),
.A2(n_66),
.B1(n_67),
.B2(n_81),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_15),
.A2(n_29),
.B1(n_36),
.B2(n_81),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_16),
.A2(n_44),
.B1(n_45),
.B2(n_47),
.Y(n_43)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_16),
.A2(n_47),
.B1(n_61),
.B2(n_64),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_16),
.A2(n_29),
.B1(n_36),
.B2(n_47),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_16),
.A2(n_47),
.B1(n_66),
.B2(n_67),
.Y(n_282)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_273),
.B1(n_295),
.B2(n_296),
.Y(n_19)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_20),
.Y(n_295)
);

OAI21x1_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_126),
.B(n_272),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_105),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_22),
.B(n_105),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_83),
.C(n_89),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_23),
.B(n_83),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_56),
.B2(n_57),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_24),
.B(n_58),
.C(n_73),
.Y(n_125)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_40),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_26),
.A2(n_27),
.B1(n_40),
.B2(n_41),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_33),
.B1(n_34),
.B2(n_38),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_28),
.A2(n_33),
.B(n_38),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_28),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_28),
.A2(n_33),
.B1(n_95),
.B2(n_138),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_28),
.A2(n_33),
.B1(n_138),
.B2(n_186),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_28),
.A2(n_33),
.B1(n_186),
.B2(n_197),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_28),
.A2(n_33),
.B1(n_197),
.B2(n_225),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_28),
.A2(n_33),
.B1(n_142),
.B2(n_237),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_L g241 ( 
.A1(n_28),
.A2(n_33),
.B1(n_230),
.B2(n_237),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_32),
.Y(n_28)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

OA22x2_ASAP7_75t_L g52 ( 
.A1(n_29),
.A2(n_36),
.B1(n_50),
.B2(n_51),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_29),
.B(n_239),
.Y(n_238)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_32),
.A2(n_35),
.B1(n_93),
.B2(n_94),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_32),
.A2(n_93),
.B1(n_229),
.B2(n_231),
.Y(n_228)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

OAI21xp33_ASAP7_75t_L g218 ( 
.A1(n_36),
.A2(n_51),
.B(n_142),
.Y(n_218)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_48),
.B1(n_53),
.B2(n_55),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_43),
.A2(n_52),
.B1(n_97),
.B2(n_99),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_44),
.A2(n_45),
.B1(n_50),
.B2(n_51),
.Y(n_49)
);

OA22x2_ASAP7_75t_L g79 ( 
.A1(n_44),
.A2(n_45),
.B1(n_77),
.B2(n_78),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_44),
.B(n_78),
.Y(n_195)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI32xp33_ASAP7_75t_L g193 ( 
.A1(n_45),
.A2(n_64),
.A3(n_77),
.B1(n_194),
.B2(n_195),
.Y(n_193)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_48),
.A2(n_53),
.B1(n_55),
.B2(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_48),
.A2(n_55),
.B1(n_87),
.B2(n_113),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_48),
.A2(n_55),
.B1(n_98),
.B2(n_165),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_48),
.A2(n_55),
.B1(n_165),
.B2(n_188),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_48),
.A2(n_55),
.B1(n_215),
.B2(n_216),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_48),
.A2(n_55),
.B1(n_216),
.B2(n_223),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_48),
.A2(n_55),
.B(n_113),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_52),
.Y(n_48)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_50),
.Y(n_51)
);

CKINVDCx14_ASAP7_75t_R g55 ( 
.A(n_52),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_52),
.A2(n_99),
.B1(n_189),
.B2(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

XOR2xp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_73),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_69),
.B2(n_71),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_59),
.A2(n_60),
.B1(n_69),
.B2(n_103),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_59),
.A2(n_60),
.B1(n_71),
.B2(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_59),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_59),
.A2(n_60),
.B1(n_149),
.B2(n_169),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_59),
.A2(n_60),
.B1(n_122),
.B2(n_282),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_60),
.B(n_65),
.Y(n_59)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_60),
.Y(n_153)
);

OA22x2_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_62),
.B1(n_63),
.B2(n_64),
.Y(n_60)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_61),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_61),
.A2(n_64),
.B1(n_77),
.B2(n_78),
.Y(n_76)
);

OAI32xp33_ASAP7_75t_L g139 ( 
.A1(n_61),
.A2(n_63),
.A3(n_66),
.B1(n_140),
.B2(n_141),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_61),
.B(n_142),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_62),
.A2(n_63),
.B1(n_66),
.B2(n_67),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_62),
.B(n_64),
.Y(n_140)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_67),
.B(n_142),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_74),
.A2(n_79),
.B1(n_80),
.B2(n_82),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_74),
.A2(n_79),
.B1(n_80),
.B2(n_101),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_74),
.A2(n_79),
.B1(n_145),
.B2(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_75),
.A2(n_109),
.B1(n_110),
.B2(n_111),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_75),
.A2(n_111),
.B1(n_144),
.B2(n_146),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_75),
.A2(n_111),
.B1(n_180),
.B2(n_182),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_75),
.A2(n_110),
.B1(n_111),
.B2(n_288),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_79),
.Y(n_75)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_79),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_79),
.A2(n_181),
.B(n_251),
.Y(n_250)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_82),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_85),
.B1(n_86),
.B2(n_88),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_84),
.B(n_88),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_84),
.A2(n_85),
.B1(n_120),
.B2(n_121),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_85),
.A2(n_121),
.B(n_123),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_86),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_89),
.B(n_155),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_100),
.C(n_102),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_90),
.A2(n_91),
.B1(n_131),
.B2(n_132),
.Y(n_130)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_96),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_92),
.B(n_96),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_100),
.B(n_102),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_101),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_103),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_125),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_115),
.B1(n_116),
.B2(n_124),
.Y(n_106)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_107),
.Y(n_124)
);

OAI21xp33_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_112),
.B(n_114),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_108),
.B(n_112),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_114),
.A2(n_279),
.B1(n_291),
.B2(n_292),
.Y(n_278)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_114),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_115),
.B(n_124),
.C(n_125),
.Y(n_293)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_118),
.B1(n_119),
.B2(n_123),
.Y(n_116)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_117),
.Y(n_123)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

AOI21x1_ASAP7_75t_SL g126 ( 
.A1(n_127),
.A2(n_156),
.B(n_271),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_154),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_128),
.B(n_154),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_133),
.C(n_134),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_129),
.A2(n_130),
.B1(n_133),
.B2(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_133),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_134),
.B(n_172),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_143),
.C(n_147),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_135),
.B(n_160),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_136),
.B(n_139),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_136),
.A2(n_137),
.B1(n_139),
.B2(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_139),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_141),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_143),
.B(n_147),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_151),
.B1(n_152),
.B2(n_153),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

OAI221xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_174),
.B1(n_269),
.B2(n_270),
.C(n_298),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_171),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_158),
.B(n_171),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_161),
.C(n_162),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_159),
.B(n_268),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_161),
.B(n_162),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_166),
.C(n_168),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_163),
.A2(n_164),
.B1(n_166),
.B2(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_166),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_167),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_168),
.B(n_201),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_175),
.B(n_265),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_208),
.B(n_264),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_198),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_177),
.B(n_198),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_187),
.C(n_190),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_178),
.B(n_261),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_SL g178 ( 
.A(n_179),
.B(n_183),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_179),
.B(n_184),
.C(n_185),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_187),
.A2(n_190),
.B1(n_191),
.B2(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_187),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_196),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_192),
.A2(n_193),
.B1(n_196),
.B2(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_194),
.Y(n_252)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_196),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_199),
.A2(n_200),
.B1(n_203),
.B2(n_207),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_199),
.B(n_204),
.C(n_206),
.Y(n_266)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_203),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_204),
.B(n_206),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_258),
.B(n_263),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_210),
.A2(n_246),
.B(n_257),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_226),
.B(n_245),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_219),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_212),
.B(n_219),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_213),
.B(n_217),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_213),
.A2(n_214),
.B1(n_217),
.B2(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_217),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_224),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_221),
.B(n_222),
.C(n_224),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_223),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_225),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_227),
.A2(n_234),
.B(n_244),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_232),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_228),
.B(n_232),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_240),
.B(n_243),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_236),
.B(n_238),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_241),
.B(n_242),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_247),
.B(n_248),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_255),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_253),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_250),
.B(n_253),
.C(n_255),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_259),
.B(n_260),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

OR2x2_ASAP7_75t_L g269 ( 
.A(n_266),
.B(n_267),
.Y(n_269)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_273),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_294),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_276),
.B(n_293),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_276),
.B(n_293),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_279),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_281),
.B1(n_283),
.B2(n_284),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_285),
.A2(n_286),
.B1(n_287),
.B2(n_290),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g290 ( 
.A(n_285),
.Y(n_290)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

CKINVDCx14_ASAP7_75t_R g288 ( 
.A(n_289),
.Y(n_288)
);


endmodule