module fake_jpeg_8793_n_329 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_329);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_329;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

HB1xp67_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx2_ASAP7_75t_SL g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_13),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_34),
.B(n_36),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

OR2x2_ASAP7_75t_L g36 ( 
.A(n_17),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_7),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_38),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_26),
.B(n_7),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_16),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_41),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_39),
.A2(n_29),
.B1(n_26),
.B2(n_30),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_45),
.A2(n_65),
.B1(n_46),
.B2(n_60),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_47),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_34),
.A2(n_29),
.B1(n_26),
.B2(n_18),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_48),
.A2(n_63),
.B1(n_69),
.B2(n_32),
.Y(n_74)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_51),
.B(n_52),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_28),
.Y(n_52)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_36),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_54),
.B(n_55),
.Y(n_79)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_56),
.B(n_59),
.Y(n_82)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_35),
.B(n_30),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_18),
.Y(n_61)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_18),
.Y(n_62)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_43),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_64),
.B(n_27),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_22),
.Y(n_65)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_36),
.B(n_22),
.Y(n_67)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_68),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_39),
.A2(n_29),
.B1(n_20),
.B2(n_17),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g72 ( 
.A(n_67),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_72),
.B(n_95),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_74),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_61),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_76),
.B(n_86),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_51),
.A2(n_20),
.B1(n_32),
.B2(n_27),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_78),
.A2(n_85),
.B1(n_94),
.B2(n_68),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_53),
.B(n_56),
.C(n_64),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_81),
.B(n_57),
.C(n_59),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_83),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_54),
.A2(n_12),
.B1(n_13),
.B2(n_10),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_62),
.Y(n_86)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_70),
.A2(n_55),
.B1(n_60),
.B2(n_66),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_89),
.B(n_19),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_70),
.A2(n_24),
.B(n_23),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_90),
.A2(n_49),
.B(n_63),
.Y(n_99)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_92),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_46),
.A2(n_19),
.B1(n_27),
.B2(n_25),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_99),
.A2(n_102),
.B(n_76),
.Y(n_125)
);

A2O1A1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_90),
.A2(n_72),
.B(n_75),
.C(n_82),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_100),
.B(n_121),
.Y(n_131)
);

OAI21xp33_ASAP7_75t_L g101 ( 
.A1(n_82),
.A2(n_49),
.B(n_59),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_101),
.A2(n_114),
.B1(n_77),
.B2(n_86),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_1),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_87),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_104),
.B(n_105),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_75),
.B(n_52),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_74),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_106),
.B(n_107),
.Y(n_145)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_79),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_79),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_108),
.B(n_109),
.Y(n_140)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_110),
.B(n_99),
.C(n_80),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_93),
.B(n_52),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g143 ( 
.A(n_112),
.B(n_12),
.Y(n_143)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_95),
.Y(n_113)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_113),
.Y(n_127)
);

AOI22x1_ASAP7_75t_SL g114 ( 
.A1(n_77),
.A2(n_23),
.B1(n_27),
.B2(n_25),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_116),
.A2(n_84),
.B1(n_88),
.B2(n_73),
.Y(n_130)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_91),
.Y(n_117)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_117),
.Y(n_148)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_83),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_119),
.A2(n_96),
.B1(n_50),
.B2(n_83),
.Y(n_137)
);

INVxp33_ASAP7_75t_L g120 ( 
.A(n_92),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_120),
.Y(n_135)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_91),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_122),
.B(n_80),
.Y(n_128)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_73),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_123),
.Y(n_141)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_85),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_124),
.B(n_19),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_125),
.A2(n_138),
.B(n_142),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_126),
.A2(n_100),
.B1(n_118),
.B2(n_107),
.Y(n_158)
);

AOI21xp33_ASAP7_75t_L g172 ( 
.A1(n_128),
.A2(n_21),
.B(n_33),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_129),
.B(n_132),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_130),
.A2(n_25),
.B1(n_71),
.B2(n_33),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_110),
.B(n_84),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_122),
.B(n_93),
.C(n_88),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_133),
.B(n_152),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_123),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_134),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_113),
.A2(n_50),
.B1(n_73),
.B2(n_57),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_136),
.A2(n_121),
.B1(n_119),
.B2(n_115),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_137),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_97),
.A2(n_106),
.B1(n_124),
.B2(n_109),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_143),
.B(n_144),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_111),
.Y(n_144)
);

OA22x2_ASAP7_75t_L g146 ( 
.A1(n_114),
.A2(n_71),
.B1(n_33),
.B2(n_21),
.Y(n_146)
);

AO21x2_ASAP7_75t_SL g162 ( 
.A1(n_146),
.A2(n_71),
.B(n_31),
.Y(n_162)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_103),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_147),
.B(n_103),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_97),
.A2(n_96),
.B1(n_25),
.B2(n_33),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_149),
.Y(n_175)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_105),
.B(n_10),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_150),
.B(n_151),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_117),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_118),
.B(n_71),
.Y(n_152)
);

OR2x2_ASAP7_75t_L g153 ( 
.A(n_140),
.B(n_108),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_153),
.B(n_154),
.Y(n_184)
);

OR2x2_ASAP7_75t_L g154 ( 
.A(n_131),
.B(n_104),
.Y(n_154)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_136),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_157),
.B(n_164),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_158),
.A2(n_166),
.B(n_172),
.Y(n_195)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_160),
.Y(n_182)
);

OA21x2_ASAP7_75t_L g185 ( 
.A1(n_162),
.A2(n_146),
.B(n_149),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_127),
.A2(n_98),
.B1(n_102),
.B2(n_112),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_163),
.A2(n_176),
.B(n_178),
.Y(n_190)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_131),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_145),
.A2(n_98),
.B(n_102),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_148),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_167),
.B(n_169),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_168),
.A2(n_177),
.B1(n_58),
.B2(n_2),
.Y(n_204)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_148),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_141),
.B(n_115),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_170),
.B(n_173),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_171),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_141),
.B(n_47),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_127),
.A2(n_47),
.B(n_31),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_138),
.A2(n_58),
.B1(n_47),
.B2(n_31),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_142),
.A2(n_47),
.B(n_31),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_139),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_180),
.B(n_150),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_128),
.B(n_152),
.Y(n_181)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_181),
.Y(n_187)
);

AOI322xp5_ASAP7_75t_L g183 ( 
.A1(n_165),
.A2(n_128),
.A3(n_129),
.B1(n_126),
.B2(n_125),
.C1(n_133),
.C2(n_132),
.Y(n_183)
);

AO21x1_ASAP7_75t_L g219 ( 
.A1(n_183),
.A2(n_195),
.B(n_187),
.Y(n_219)
);

AOI22x1_ASAP7_75t_L g226 ( 
.A1(n_185),
.A2(n_175),
.B1(n_159),
.B2(n_155),
.Y(n_226)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_186),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_161),
.B(n_147),
.C(n_134),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_188),
.B(n_198),
.C(n_199),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_153),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_189),
.B(n_194),
.Y(n_229)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_168),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_191),
.B(n_202),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_153),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_161),
.B(n_135),
.C(n_146),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_196),
.B(n_177),
.C(n_162),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_154),
.B(n_143),
.Y(n_197)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_197),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_174),
.B(n_135),
.C(n_146),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_174),
.B(n_58),
.C(n_21),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_154),
.B(n_21),
.Y(n_201)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_201),
.Y(n_215)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_176),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_164),
.B(n_1),
.Y(n_203)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_203),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_204),
.A2(n_208),
.B(n_6),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_162),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_205),
.A2(n_162),
.B1(n_157),
.B2(n_179),
.Y(n_210)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_167),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_207),
.B(n_169),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_165),
.A2(n_181),
.B(n_175),
.Y(n_208)
);

CKINVDCx14_ASAP7_75t_R g245 ( 
.A(n_210),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_184),
.A2(n_178),
.B(n_180),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_212),
.A2(n_226),
.B(n_227),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_208),
.B(n_166),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_213),
.B(n_225),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_188),
.B(n_163),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_214),
.B(n_218),
.C(n_231),
.Y(n_235)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_193),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_217),
.B(n_221),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_219),
.B(n_195),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_193),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_220),
.B(n_233),
.Y(n_242)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_184),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_200),
.Y(n_222)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_222),
.Y(n_243)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_224),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_199),
.B(n_156),
.Y(n_225)
);

OA21x2_ASAP7_75t_L g227 ( 
.A1(n_202),
.A2(n_159),
.B(n_155),
.Y(n_227)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_228),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_189),
.B(n_1),
.Y(n_230)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_230),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_187),
.B(n_198),
.C(n_196),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_201),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_232),
.B(n_192),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_200),
.Y(n_233)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_236),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_239),
.B(n_247),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_224),
.Y(n_240)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_240),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_234),
.B(n_190),
.C(n_183),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_241),
.B(n_234),
.C(n_231),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_209),
.A2(n_191),
.B1(n_194),
.B2(n_192),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_244),
.A2(n_246),
.B1(n_253),
.B2(n_211),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_209),
.A2(n_229),
.B1(n_223),
.B2(n_218),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_214),
.B(n_190),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_230),
.B(n_203),
.Y(n_250)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_250),
.Y(n_272)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_226),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_251),
.B(n_228),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_226),
.A2(n_206),
.B1(n_204),
.B2(n_205),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_252),
.A2(n_232),
.B1(n_212),
.B2(n_215),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_223),
.A2(n_207),
.B1(n_197),
.B2(n_185),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_225),
.B(n_186),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_254),
.B(n_249),
.Y(n_267)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_257),
.Y(n_276)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_258),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_236),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_260),
.B(n_267),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_261),
.A2(n_264),
.B1(n_268),
.B2(n_273),
.Y(n_279)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_245),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_263),
.B(n_274),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_246),
.A2(n_210),
.B1(n_227),
.B2(n_216),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_265),
.B(n_235),
.C(n_255),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_251),
.A2(n_182),
.B1(n_227),
.B2(n_185),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_255),
.B(n_213),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_269),
.B(n_259),
.Y(n_275)
);

OR2x2_ASAP7_75t_L g270 ( 
.A(n_242),
.B(n_253),
.Y(n_270)
);

OAI322xp33_ASAP7_75t_L g286 ( 
.A1(n_270),
.A2(n_256),
.A3(n_250),
.B1(n_185),
.B2(n_5),
.C1(n_6),
.C2(n_8),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_235),
.B(n_219),
.C(n_182),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_271),
.B(n_239),
.C(n_241),
.Y(n_283)
);

XOR2x2_ASAP7_75t_L g273 ( 
.A(n_238),
.B(n_244),
.Y(n_273)
);

OA21x2_ASAP7_75t_L g278 ( 
.A1(n_273),
.A2(n_238),
.B(n_237),
.Y(n_278)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_243),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_275),
.B(n_281),
.C(n_284),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_278),
.B(n_287),
.Y(n_290)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_279),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_270),
.B(n_248),
.Y(n_280)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_280),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_283),
.B(n_285),
.C(n_289),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_265),
.B(n_271),
.C(n_237),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_269),
.B(n_247),
.Y(n_285)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_286),
.Y(n_295)
);

CKINVDCx14_ASAP7_75t_R g287 ( 
.A(n_258),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_262),
.B(n_259),
.C(n_266),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_278),
.B(n_274),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_292),
.B(n_293),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_277),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_278),
.B(n_272),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_294),
.B(n_296),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_276),
.B(n_264),
.Y(n_296)
);

INVx6_ASAP7_75t_L g297 ( 
.A(n_282),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_297),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_288),
.B(n_6),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_298),
.B(n_300),
.Y(n_308)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_289),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_301),
.B(n_283),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_303),
.B(n_306),
.C(n_309),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_SL g306 ( 
.A(n_290),
.B(n_285),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_301),
.B(n_284),
.Y(n_309)
);

INVx1_ASAP7_75t_SL g310 ( 
.A(n_290),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_310),
.B(n_307),
.Y(n_319)
);

OAI21x1_ASAP7_75t_SL g311 ( 
.A1(n_295),
.A2(n_275),
.B(n_8),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_311),
.A2(n_9),
.B(n_12),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_293),
.B(n_8),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_312),
.B(n_304),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_310),
.A2(n_302),
.B1(n_291),
.B2(n_297),
.Y(n_313)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_313),
.Y(n_323)
);

BUFx4f_ASAP7_75t_SL g314 ( 
.A(n_305),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_314),
.A2(n_316),
.B(n_317),
.Y(n_324)
);

BUFx24_ASAP7_75t_SL g321 ( 
.A(n_315),
.Y(n_321)
);

NOR2x1_ASAP7_75t_L g317 ( 
.A(n_306),
.B(n_299),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_319),
.A2(n_320),
.B(n_5),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_308),
.B(n_299),
.Y(n_320)
);

OAI21x1_ASAP7_75t_L g325 ( 
.A1(n_322),
.A2(n_319),
.B(n_314),
.Y(n_325)
);

AOI311xp33_ASAP7_75t_L g327 ( 
.A1(n_325),
.A2(n_326),
.A3(n_321),
.B(n_323),
.C(n_9),
.Y(n_327)
);

NAND2x1_ASAP7_75t_SL g326 ( 
.A(n_324),
.B(n_318),
.Y(n_326)
);

A2O1A1O1Ixp25_ASAP7_75t_L g328 ( 
.A1(n_327),
.A2(n_10),
.B(n_3),
.C(n_4),
.D(n_2),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_328),
.B(n_4),
.Y(n_329)
);


endmodule