module fake_jpeg_12236_n_99 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_29, n_12, n_8, n_15, n_7, n_99);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_99;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_30),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_27),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_18),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

BUFx16f_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx2_ASAP7_75t_R g42 ( 
.A(n_38),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_46),
.Y(n_50)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_32),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_39),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_49),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_2),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_40),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_53),
.B(n_58),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_36),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_54),
.B(n_55),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_39),
.Y(n_55)
);

NAND2x1p5_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_41),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_60),
.C(n_41),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_3),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_4),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_51),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_62),
.B(n_64),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_73),
.Y(n_75)
);

INVx6_ASAP7_75t_SL g64 ( 
.A(n_56),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_50),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_67),
.B(n_71),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_52),
.A2(n_35),
.B1(n_4),
.B2(n_7),
.Y(n_68)
);

AND2x2_ASAP7_75t_SL g76 ( 
.A(n_68),
.B(n_72),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_52),
.A2(n_35),
.B1(n_8),
.B2(n_9),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_69),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g70 ( 
.A(n_50),
.B(n_35),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_19),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_59),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_52),
.A2(n_6),
.B1(n_11),
.B2(n_12),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_54),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_74),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_78),
.Y(n_87)
);

A2O1A1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_67),
.A2(n_13),
.B(n_14),
.C(n_17),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_SL g88 ( 
.A(n_80),
.B(n_24),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_20),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_83),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_84),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_88),
.B(n_89),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_86),
.A2(n_76),
.B1(n_82),
.B2(n_85),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_92),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_91),
.A2(n_75),
.B(n_82),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_93),
.A2(n_87),
.B(n_79),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_95),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_96),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_94),
.C(n_90),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_98),
.B(n_76),
.Y(n_99)
);


endmodule