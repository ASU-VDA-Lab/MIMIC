module fake_jpeg_1962_n_674 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_674);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_674;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_6),
.B(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_10),
.B(n_19),
.Y(n_25)
);

BUFx4f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_10),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_14),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

BUFx10_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_6),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

CKINVDCx5p33_ASAP7_75t_R g54 ( 
.A(n_15),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_2),
.Y(n_55)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_12),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_16),
.Y(n_58)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_10),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_25),
.B(n_0),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_60),
.B(n_62),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g154 ( 
.A(n_61),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_25),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g156 ( 
.A(n_63),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_30),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_64),
.B(n_70),
.Y(n_168)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_65),
.Y(n_163)
);

BUFx24_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

BUFx24_ASAP7_75t_L g165 ( 
.A(n_66),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_67),
.Y(n_132)
);

BUFx10_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g176 ( 
.A(n_68),
.Y(n_176)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

INVx11_ASAP7_75t_L g207 ( 
.A(n_69),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_30),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_30),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_71),
.B(n_80),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_72),
.Y(n_151)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

INVx8_ASAP7_75t_L g171 ( 
.A(n_73),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_20),
.B(n_0),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_74),
.B(n_103),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_23),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_75),
.Y(n_153)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_76),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_33),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_77),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_33),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_78),
.Y(n_161)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_33),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_79),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_47),
.Y(n_80)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_34),
.Y(n_81)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_81),
.Y(n_152)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_82),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_47),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_83),
.B(n_88),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_47),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_84)
);

OA22x2_ASAP7_75t_L g147 ( 
.A1(n_84),
.A2(n_27),
.B1(n_39),
.B2(n_40),
.Y(n_147)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_24),
.Y(n_85)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_85),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_86),
.Y(n_184)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_87),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_51),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_20),
.B(n_24),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_89),
.B(n_104),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_90),
.Y(n_185)
);

INVx2_ASAP7_75t_SL g91 ( 
.A(n_58),
.Y(n_91)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_91),
.Y(n_170)
);

BUFx12_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g140 ( 
.A(n_92),
.Y(n_140)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_93),
.Y(n_139)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_31),
.Y(n_94)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_94),
.Y(n_137)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_29),
.Y(n_95)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_95),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_28),
.Y(n_96)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_96),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_57),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_97),
.Y(n_192)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_26),
.Y(n_98)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_98),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_57),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_99),
.Y(n_197)
);

INVx2_ASAP7_75t_SL g100 ( 
.A(n_34),
.Y(n_100)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_100),
.Y(n_189)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_53),
.Y(n_101)
);

INVx8_ASAP7_75t_L g220 ( 
.A(n_101),
.Y(n_220)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_26),
.Y(n_102)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_102),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_54),
.B(n_17),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_31),
.B(n_36),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_21),
.B(n_17),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_105),
.B(n_121),
.Y(n_162)
);

INVx11_ASAP7_75t_L g106 ( 
.A(n_34),
.Y(n_106)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_106),
.Y(n_193)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_29),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g145 ( 
.A(n_107),
.Y(n_145)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_38),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_108),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_57),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_109),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_53),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_110),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_37),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_111),
.B(n_112),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_36),
.B(n_3),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g113 ( 
.A(n_56),
.Y(n_113)
);

INVx8_ASAP7_75t_L g148 ( 
.A(n_113),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_41),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_114),
.B(n_115),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_41),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_26),
.Y(n_116)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_116),
.Y(n_150)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_56),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_117),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_21),
.B(n_3),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_118),
.B(n_130),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_41),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_119),
.Y(n_221)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_38),
.Y(n_120)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_120),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_22),
.B(n_4),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_59),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_122),
.Y(n_225)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_52),
.Y(n_123)
);

BUFx12f_ASAP7_75t_L g159 ( 
.A(n_123),
.Y(n_159)
);

BUFx4f_ASAP7_75t_L g124 ( 
.A(n_51),
.Y(n_124)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_124),
.Y(n_160)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_52),
.Y(n_125)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_125),
.Y(n_169)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_26),
.Y(n_126)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_126),
.Y(n_174)
);

BUFx5_ASAP7_75t_L g127 ( 
.A(n_51),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_127),
.Y(n_211)
);

BUFx12f_ASAP7_75t_L g128 ( 
.A(n_56),
.Y(n_128)
);

INVx8_ASAP7_75t_L g217 ( 
.A(n_128),
.Y(n_217)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_27),
.Y(n_129)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_129),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_59),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_59),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_131),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_89),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_135),
.B(n_187),
.Y(n_233)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_67),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_138),
.Y(n_236)
);

OA22x2_ASAP7_75t_L g230 ( 
.A1(n_147),
.A2(n_84),
.B1(n_95),
.B2(n_107),
.Y(n_230)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_87),
.Y(n_149)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_149),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_72),
.A2(n_46),
.B1(n_44),
.B2(n_43),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_157),
.A2(n_128),
.B1(n_73),
.B2(n_113),
.Y(n_257)
);

FAx1_ASAP7_75t_L g164 ( 
.A(n_92),
.B(n_51),
.CI(n_52),
.CON(n_164),
.SN(n_164)
);

OR2x2_ASAP7_75t_L g304 ( 
.A(n_164),
.B(n_172),
.Y(n_304)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_91),
.Y(n_166)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_166),
.Y(n_239)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_75),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_167),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_100),
.B(n_52),
.Y(n_172)
);

AND2x2_ASAP7_75t_SL g178 ( 
.A(n_76),
.B(n_52),
.Y(n_178)
);

NAND2x1_ASAP7_75t_SL g249 ( 
.A(n_178),
.B(n_183),
.Y(n_249)
);

INVx6_ASAP7_75t_SL g179 ( 
.A(n_92),
.Y(n_179)
);

INVx6_ASAP7_75t_SL g308 ( 
.A(n_179),
.Y(n_308)
);

INVx13_ASAP7_75t_L g180 ( 
.A(n_66),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g305 ( 
.A(n_180),
.Y(n_305)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_102),
.Y(n_182)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_182),
.Y(n_228)
);

INVx6_ASAP7_75t_SL g183 ( 
.A(n_66),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_119),
.Y(n_187)
);

INVx6_ASAP7_75t_L g190 ( 
.A(n_77),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_190),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_122),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_191),
.B(n_200),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_123),
.B(n_44),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_194),
.B(n_203),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_79),
.A2(n_46),
.B1(n_49),
.B2(n_48),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_L g240 ( 
.A1(n_195),
.A2(n_32),
.B1(n_55),
.B2(n_49),
.Y(n_240)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_65),
.Y(n_198)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_198),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_125),
.B(n_46),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_124),
.B(n_40),
.Y(n_203)
);

INVx13_ASAP7_75t_L g204 ( 
.A(n_68),
.Y(n_204)
);

BUFx16f_ASAP7_75t_L g238 ( 
.A(n_204),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_117),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_205),
.B(n_215),
.Y(n_292)
);

INVx6_ASAP7_75t_L g208 ( 
.A(n_78),
.Y(n_208)
);

INVx5_ASAP7_75t_L g272 ( 
.A(n_208),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_124),
.B(n_42),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_209),
.B(n_210),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_82),
.B(n_42),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_86),
.B(n_39),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_212),
.B(n_16),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_90),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_131),
.Y(n_216)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_216),
.Y(n_244)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_97),
.Y(n_219)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_219),
.Y(n_247)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_99),
.Y(n_222)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_222),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_109),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_128),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_61),
.B(n_55),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_224),
.B(n_120),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_227),
.B(n_241),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_172),
.B(n_178),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g313 ( 
.A(n_229),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_SL g316 ( 
.A1(n_230),
.A2(n_231),
.B1(n_258),
.B2(n_265),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_164),
.A2(n_110),
.B1(n_43),
.B2(n_108),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_162),
.B(n_35),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_235),
.B(n_252),
.Y(n_324)
);

CKINVDCx14_ASAP7_75t_R g331 ( 
.A(n_237),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_240),
.A2(n_255),
.B1(n_132),
.B2(n_161),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_177),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_196),
.B(n_96),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_242),
.B(n_246),
.Y(n_317)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_189),
.Y(n_245)
);

INVx4_ASAP7_75t_L g362 ( 
.A(n_245),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_196),
.B(n_188),
.Y(n_246)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_136),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_248),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_188),
.B(n_63),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_250),
.B(n_266),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_206),
.B(n_22),
.Y(n_252)
);

NAND2x1_ASAP7_75t_SL g254 ( 
.A(n_180),
.B(n_68),
.Y(n_254)
);

AO21x1_ASAP7_75t_L g336 ( 
.A1(n_254),
.A2(n_259),
.B(n_260),
.Y(n_336)
);

AOI22xp33_ASAP7_75t_L g255 ( 
.A1(n_202),
.A2(n_32),
.B1(n_35),
.B2(n_48),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_257),
.A2(n_220),
.B1(n_151),
.B2(n_153),
.Y(n_343)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_186),
.A2(n_113),
.B1(n_101),
.B2(n_73),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_186),
.B(n_101),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_170),
.B(n_4),
.Y(n_260)
);

OAI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_202),
.A2(n_106),
.B1(n_81),
.B2(n_69),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_261),
.A2(n_278),
.B1(n_176),
.B2(n_156),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_206),
.B(n_134),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_262),
.B(n_264),
.Y(n_349)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_148),
.Y(n_263)
);

INVx3_ASAP7_75t_L g320 ( 
.A(n_263),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_224),
.B(n_4),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_145),
.A2(n_127),
.B1(n_7),
.B2(n_8),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_144),
.B(n_6),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_200),
.B(n_6),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_267),
.B(n_301),
.C(n_185),
.Y(n_363)
);

INVx4_ASAP7_75t_L g268 ( 
.A(n_148),
.Y(n_268)
);

INVx3_ASAP7_75t_L g326 ( 
.A(n_268),
.Y(n_326)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_137),
.Y(n_271)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_271),
.Y(n_311)
);

AND2x4_ASAP7_75t_SL g273 ( 
.A(n_133),
.B(n_7),
.Y(n_273)
);

MAJx3_ASAP7_75t_L g325 ( 
.A(n_273),
.B(n_165),
.C(n_154),
.Y(n_325)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_146),
.Y(n_274)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_274),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_144),
.B(n_9),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_275),
.B(n_283),
.Y(n_321)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_145),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_276),
.B(n_281),
.Y(n_366)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_160),
.Y(n_277)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_277),
.Y(n_319)
);

OAI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_168),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_218),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g328 ( 
.A1(n_279),
.A2(n_291),
.B1(n_176),
.B2(n_156),
.Y(n_328)
);

INVx5_ASAP7_75t_L g280 ( 
.A(n_217),
.Y(n_280)
);

INVx3_ASAP7_75t_L g365 ( 
.A(n_280),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_177),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_141),
.Y(n_282)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_282),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_142),
.B(n_11),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_139),
.B(n_11),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_284),
.B(n_298),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_168),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_285),
.B(n_286),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_140),
.B(n_12),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_150),
.Y(n_287)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_287),
.Y(n_347)
);

INVx4_ASAP7_75t_L g288 ( 
.A(n_217),
.Y(n_288)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_288),
.Y(n_369)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_174),
.Y(n_289)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_289),
.Y(n_312)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_169),
.Y(n_290)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_290),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_SL g291 ( 
.A1(n_218),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_291)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_199),
.Y(n_293)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_293),
.Y(n_329)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_163),
.Y(n_294)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_294),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_173),
.A2(n_13),
.B(n_15),
.Y(n_295)
);

OR2x2_ASAP7_75t_L g345 ( 
.A(n_295),
.B(n_296),
.Y(n_345)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_143),
.Y(n_297)
);

INVx5_ASAP7_75t_L g334 ( 
.A(n_297),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_147),
.B(n_158),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_147),
.B(n_16),
.Y(n_299)
);

OAI32xp33_ASAP7_75t_L g314 ( 
.A1(n_299),
.A2(n_306),
.A3(n_165),
.B1(n_204),
.B2(n_211),
.Y(n_314)
);

INVx3_ASAP7_75t_L g300 ( 
.A(n_171),
.Y(n_300)
);

INVx5_ASAP7_75t_L g337 ( 
.A(n_300),
.Y(n_337)
);

AND2x2_ASAP7_75t_SL g301 ( 
.A(n_140),
.B(n_16),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_154),
.B(n_17),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_302),
.B(n_305),
.Y(n_353)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_175),
.Y(n_303)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_303),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_214),
.B(n_181),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_159),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_307),
.Y(n_322)
);

INVx8_ASAP7_75t_L g310 ( 
.A(n_238),
.Y(n_310)
);

INVx4_ASAP7_75t_L g390 ( 
.A(n_310),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_314),
.B(n_249),
.Y(n_373)
);

CKINVDCx14_ASAP7_75t_R g412 ( 
.A(n_325),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_328),
.Y(n_376)
);

AND2x2_ASAP7_75t_L g377 ( 
.A(n_330),
.B(n_332),
.Y(n_377)
);

AO22x1_ASAP7_75t_L g332 ( 
.A1(n_229),
.A2(n_207),
.B1(n_214),
.B2(n_213),
.Y(n_332)
);

OAI32xp33_ASAP7_75t_L g333 ( 
.A1(n_299),
.A2(n_181),
.A3(n_175),
.B1(n_213),
.B2(n_193),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_333),
.B(n_352),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_298),
.A2(n_226),
.B1(n_152),
.B2(n_225),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g394 ( 
.A1(n_339),
.A2(n_325),
.B(n_343),
.Y(n_394)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_247),
.Y(n_341)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_341),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_343),
.A2(n_351),
.B1(n_355),
.B2(n_368),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_304),
.A2(n_225),
.B1(n_221),
.B2(n_153),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g397 ( 
.A1(n_344),
.A2(n_346),
.B1(n_357),
.B2(n_272),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_304),
.A2(n_221),
.B1(n_151),
.B2(n_155),
.Y(n_346)
);

O2A1O1Ixp33_ASAP7_75t_L g350 ( 
.A1(n_230),
.A2(n_159),
.B(n_226),
.C(n_155),
.Y(n_350)
);

AOI21xp5_ASAP7_75t_L g378 ( 
.A1(n_350),
.A2(n_308),
.B(n_254),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_251),
.A2(n_243),
.B1(n_230),
.B2(n_229),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_353),
.B(n_356),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_233),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_354),
.B(n_359),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_230),
.A2(n_132),
.B1(n_161),
.B2(n_184),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_292),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_257),
.A2(n_306),
.B1(n_273),
.B2(n_284),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_247),
.Y(n_358)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_358),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_252),
.B(n_184),
.Y(n_359)
);

AOI22xp33_ASAP7_75t_SL g360 ( 
.A1(n_259),
.A2(n_305),
.B1(n_227),
.B2(n_297),
.Y(n_360)
);

AOI22xp33_ASAP7_75t_SL g380 ( 
.A1(n_360),
.A2(n_308),
.B1(n_238),
.B2(n_263),
.Y(n_380)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_256),
.Y(n_361)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_361),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_363),
.B(n_273),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_262),
.B(n_235),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_364),
.B(n_367),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_264),
.B(n_239),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_270),
.A2(n_185),
.B1(n_192),
.B2(n_197),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_338),
.B(n_259),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_SL g428 ( 
.A(n_370),
.B(n_400),
.Y(n_428)
);

INVx13_ASAP7_75t_L g371 ( 
.A(n_310),
.Y(n_371)
);

INVx4_ASAP7_75t_L g440 ( 
.A(n_371),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_373),
.A2(n_311),
.B1(n_320),
.B2(n_369),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_313),
.B(n_232),
.C(n_249),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_374),
.B(n_363),
.C(n_348),
.Y(n_421)
);

INVx13_ASAP7_75t_L g375 ( 
.A(n_325),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_375),
.Y(n_423)
);

OAI22xp33_ASAP7_75t_SL g420 ( 
.A1(n_378),
.A2(n_330),
.B1(n_336),
.B2(n_314),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_SL g426 ( 
.A1(n_380),
.A2(n_394),
.B(n_365),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_315),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_383),
.B(n_395),
.Y(n_425)
);

INVx8_ASAP7_75t_L g384 ( 
.A(n_350),
.Y(n_384)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_384),
.Y(n_448)
);

AND2x6_ASAP7_75t_L g386 ( 
.A(n_351),
.B(n_238),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_386),
.B(n_407),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_387),
.B(n_267),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_357),
.A2(n_295),
.B1(n_301),
.B2(n_201),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_388),
.A2(n_397),
.B1(n_405),
.B2(n_332),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_338),
.B(n_301),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_389),
.B(n_398),
.Y(n_439)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_335),
.Y(n_392)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_392),
.Y(n_435)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_335),
.Y(n_393)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_393),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_334),
.Y(n_395)
);

INVx3_ASAP7_75t_L g396 ( 
.A(n_334),
.Y(n_396)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_396),
.Y(n_446)
);

OAI32xp33_ASAP7_75t_L g398 ( 
.A1(n_349),
.A2(n_324),
.A3(n_313),
.B1(n_317),
.B2(n_318),
.Y(n_398)
);

INVx13_ASAP7_75t_L g399 ( 
.A(n_337),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_399),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_356),
.B(n_267),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_349),
.B(n_260),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_401),
.B(n_404),
.Y(n_442)
);

AOI22xp33_ASAP7_75t_SL g403 ( 
.A1(n_355),
.A2(n_300),
.B1(n_268),
.B2(n_288),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_403),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_345),
.B(n_260),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_316),
.A2(n_345),
.B1(n_339),
.B2(n_344),
.Y(n_405)
);

INVx3_ASAP7_75t_L g406 ( 
.A(n_337),
.Y(n_406)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_406),
.Y(n_452)
);

AND2x6_ASAP7_75t_L g407 ( 
.A(n_331),
.B(n_280),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_340),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_408),
.B(n_411),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_327),
.B(n_245),
.Y(n_409)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_409),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_366),
.B(n_294),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g453 ( 
.A(n_410),
.Y(n_453)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_340),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_322),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_413),
.B(n_347),
.Y(n_454)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_323),
.Y(n_414)
);

INVxp67_ASAP7_75t_L g456 ( 
.A(n_414),
.Y(n_456)
);

INVx8_ASAP7_75t_L g415 ( 
.A(n_322),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_415),
.Y(n_430)
);

CKINVDCx16_ASAP7_75t_R g416 ( 
.A(n_336),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_416),
.B(n_341),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_418),
.A2(n_431),
.B1(n_438),
.B2(n_445),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_417),
.A2(n_346),
.B1(n_332),
.B2(n_333),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_419),
.A2(n_424),
.B1(n_384),
.B2(n_415),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_420),
.B(n_405),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_421),
.B(n_432),
.C(n_441),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_422),
.B(n_400),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_417),
.A2(n_324),
.B1(n_321),
.B2(n_311),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_SL g458 ( 
.A1(n_426),
.A2(n_427),
.B(n_450),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_372),
.A2(n_303),
.B1(n_272),
.B2(n_269),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_370),
.B(n_329),
.C(n_323),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g438 ( 
.A1(n_372),
.A2(n_236),
.B1(n_269),
.B2(n_253),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_389),
.B(n_329),
.C(n_312),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_382),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_443),
.B(n_383),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_SL g444 ( 
.A(n_398),
.B(n_312),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_444),
.B(n_447),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_417),
.A2(n_253),
.B1(n_236),
.B2(n_201),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_SL g447 ( 
.A(n_401),
.B(n_274),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_382),
.B(n_391),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_SL g487 ( 
.A(n_451),
.B(n_379),
.Y(n_487)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_454),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_413),
.B(n_320),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_455),
.B(n_395),
.Y(n_467)
);

OR2x2_ASAP7_75t_L g457 ( 
.A(n_373),
.B(n_365),
.Y(n_457)
);

CKINVDCx16_ASAP7_75t_R g475 ( 
.A(n_457),
.Y(n_475)
);

OAI21xp5_ASAP7_75t_SL g459 ( 
.A1(n_423),
.A2(n_378),
.B(n_375),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_L g499 ( 
.A1(n_459),
.A2(n_480),
.B(n_482),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_SL g514 ( 
.A(n_460),
.B(n_466),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_421),
.B(n_412),
.C(n_387),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_464),
.B(n_465),
.C(n_481),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_422),
.B(n_374),
.C(n_416),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_453),
.B(n_402),
.Y(n_466)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_467),
.Y(n_504)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_435),
.Y(n_468)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_468),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_443),
.B(n_404),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_SL g517 ( 
.A(n_469),
.B(n_477),
.Y(n_517)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_470),
.B(n_471),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_442),
.B(n_388),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_455),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_472),
.B(n_479),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_430),
.B(n_392),
.Y(n_473)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_473),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_L g513 ( 
.A1(n_474),
.A2(n_487),
.B1(n_384),
.B2(n_448),
.Y(n_513)
);

OR2x2_ASAP7_75t_L g476 ( 
.A(n_427),
.B(n_375),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_476),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_437),
.B(n_415),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_451),
.B(n_390),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_478),
.B(n_486),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_454),
.Y(n_479)
);

OAI21xp5_ASAP7_75t_L g480 ( 
.A1(n_423),
.A2(n_394),
.B(n_376),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_439),
.B(n_393),
.C(n_386),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_L g482 ( 
.A1(n_457),
.A2(n_376),
.B(n_377),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_430),
.B(n_425),
.Y(n_483)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_483),
.Y(n_519)
);

AND2x6_ASAP7_75t_L g485 ( 
.A(n_434),
.B(n_407),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_485),
.B(n_491),
.Y(n_498)
);

NOR3xp33_ASAP7_75t_SL g486 ( 
.A(n_439),
.B(n_377),
.C(n_414),
.Y(n_486)
);

OAI21xp5_ASAP7_75t_SL g488 ( 
.A1(n_457),
.A2(n_377),
.B(n_397),
.Y(n_488)
);

INVxp67_ASAP7_75t_L g500 ( 
.A(n_488),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_428),
.B(n_390),
.Y(n_489)
);

CKINVDCx16_ASAP7_75t_R g495 ( 
.A(n_489),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_SL g490 ( 
.A(n_428),
.B(n_385),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g518 ( 
.A(n_490),
.Y(n_518)
);

INVxp67_ASAP7_75t_L g491 ( 
.A(n_425),
.Y(n_491)
);

OAI21xp5_ASAP7_75t_SL g492 ( 
.A1(n_426),
.A2(n_450),
.B(n_434),
.Y(n_492)
);

INVxp67_ASAP7_75t_L g505 ( 
.A(n_492),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g524 ( 
.A1(n_493),
.A2(n_445),
.B1(n_431),
.B2(n_436),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_442),
.B(n_379),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g511 ( 
.A(n_494),
.B(n_470),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g501 ( 
.A(n_482),
.B(n_448),
.Y(n_501)
);

OAI21xp33_ASAP7_75t_SL g557 ( 
.A1(n_501),
.A2(n_513),
.B(n_406),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_462),
.B(n_444),
.C(n_441),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_502),
.B(n_522),
.C(n_484),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_477),
.B(n_449),
.Y(n_503)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_503),
.Y(n_542)
);

MAJx2_ASAP7_75t_L g507 ( 
.A(n_464),
.B(n_432),
.C(n_447),
.Y(n_507)
);

MAJx2_ASAP7_75t_L g532 ( 
.A(n_507),
.B(n_511),
.C(n_512),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_SL g509 ( 
.A1(n_474),
.A2(n_418),
.B1(n_424),
.B2(n_419),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g549 ( 
.A1(n_509),
.A2(n_528),
.B1(n_475),
.B2(n_476),
.Y(n_549)
);

XOR2xp5_ASAP7_75t_L g512 ( 
.A(n_462),
.B(n_447),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_483),
.B(n_449),
.Y(n_520)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_520),
.Y(n_545)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_473),
.Y(n_521)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_521),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_465),
.B(n_456),
.C(n_435),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_L g523 ( 
.A1(n_461),
.A2(n_438),
.B1(n_433),
.B2(n_436),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_L g548 ( 
.A1(n_523),
.A2(n_524),
.B1(n_527),
.B2(n_475),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_494),
.B(n_429),
.Y(n_525)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_525),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_460),
.B(n_467),
.Y(n_526)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_526),
.Y(n_551)
);

OAI22xp33_ASAP7_75t_SL g527 ( 
.A1(n_461),
.A2(n_429),
.B1(n_446),
.B2(n_452),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_SL g528 ( 
.A1(n_474),
.A2(n_452),
.B1(n_446),
.B2(n_440),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_491),
.B(n_381),
.Y(n_529)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_529),
.Y(n_555)
);

CKINVDCx20_ASAP7_75t_R g530 ( 
.A(n_487),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_530),
.B(n_490),
.Y(n_531)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_531),
.Y(n_563)
);

AO221x1_ASAP7_75t_L g533 ( 
.A1(n_495),
.A2(n_485),
.B1(n_486),
.B2(n_371),
.C(n_472),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_533),
.B(n_559),
.Y(n_564)
);

XNOR2xp5_ASAP7_75t_L g569 ( 
.A(n_534),
.B(n_508),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_512),
.B(n_484),
.C(n_481),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g574 ( 
.A(n_536),
.B(n_539),
.C(n_543),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_518),
.B(n_479),
.Y(n_537)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_537),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_518),
.B(n_463),
.Y(n_538)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_538),
.Y(n_587)
);

MAJIxp5_ASAP7_75t_SL g539 ( 
.A(n_498),
.B(n_492),
.C(n_493),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_530),
.B(n_469),
.Y(n_540)
);

INVxp67_ASAP7_75t_SL g573 ( 
.A(n_540),
.Y(n_573)
);

XOR2xp5_ASAP7_75t_L g541 ( 
.A(n_502),
.B(n_471),
.Y(n_541)
);

XOR2xp5_ASAP7_75t_L g571 ( 
.A(n_541),
.B(n_560),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_522),
.B(n_476),
.C(n_463),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_514),
.B(n_510),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_544),
.B(n_546),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_514),
.B(n_396),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_526),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_547),
.B(n_553),
.Y(n_565)
);

OAI22xp5_ASAP7_75t_L g578 ( 
.A1(n_548),
.A2(n_549),
.B1(n_515),
.B2(n_521),
.Y(n_578)
);

OAI22xp5_ASAP7_75t_SL g552 ( 
.A1(n_504),
.A2(n_480),
.B1(n_488),
.B2(n_458),
.Y(n_552)
);

AOI22xp5_ASAP7_75t_SL g576 ( 
.A1(n_552),
.A2(n_500),
.B1(n_516),
.B2(n_509),
.Y(n_576)
);

AOI21xp5_ASAP7_75t_L g553 ( 
.A1(n_499),
.A2(n_459),
.B(n_458),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_496),
.B(n_468),
.C(n_326),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_554),
.B(n_556),
.C(n_562),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_496),
.B(n_326),
.C(n_369),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_557),
.B(n_501),
.Y(n_579)
);

OAI21xp5_ASAP7_75t_SL g558 ( 
.A1(n_505),
.A2(n_371),
.B(n_411),
.Y(n_558)
);

CKINVDCx14_ASAP7_75t_R g582 ( 
.A(n_558),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_517),
.B(n_505),
.Y(n_559)
);

XOR2xp5_ASAP7_75t_L g560 ( 
.A(n_508),
.B(n_381),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_520),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_561),
.B(n_517),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g562 ( 
.A(n_507),
.B(n_385),
.C(n_408),
.Y(n_562)
);

OAI22xp5_ASAP7_75t_SL g567 ( 
.A1(n_549),
.A2(n_498),
.B1(n_504),
.B2(n_519),
.Y(n_567)
);

AOI22xp5_ASAP7_75t_L g601 ( 
.A1(n_567),
.A2(n_568),
.B1(n_578),
.B2(n_535),
.Y(n_601)
);

OAI22xp5_ASAP7_75t_SL g568 ( 
.A1(n_537),
.A2(n_555),
.B1(n_545),
.B2(n_538),
.Y(n_568)
);

XNOR2xp5_ASAP7_75t_L g606 ( 
.A(n_569),
.B(n_572),
.Y(n_606)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_570),
.Y(n_591)
);

XNOR2xp5_ASAP7_75t_L g572 ( 
.A(n_541),
.B(n_511),
.Y(n_572)
);

OAI22xp5_ASAP7_75t_SL g594 ( 
.A1(n_576),
.A2(n_553),
.B1(n_516),
.B2(n_501),
.Y(n_594)
);

XOR2xp5_ASAP7_75t_L g577 ( 
.A(n_536),
.B(n_543),
.Y(n_577)
);

MAJIxp5_ASAP7_75t_L g596 ( 
.A(n_577),
.B(n_581),
.C(n_586),
.Y(n_596)
);

AOI21xp5_ASAP7_75t_L g593 ( 
.A1(n_579),
.A2(n_558),
.B(n_500),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_531),
.B(n_529),
.Y(n_580)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_580),
.Y(n_589)
);

XOR2xp5_ASAP7_75t_L g581 ( 
.A(n_532),
.B(n_499),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_554),
.B(n_503),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_583),
.B(n_584),
.Y(n_597)
);

MAJIxp5_ASAP7_75t_L g584 ( 
.A(n_556),
.B(n_515),
.C(n_525),
.Y(n_584)
);

XOR2xp5_ASAP7_75t_L g586 ( 
.A(n_532),
.B(n_519),
.Y(n_586)
);

XOR2xp5_ASAP7_75t_L g588 ( 
.A(n_562),
.B(n_497),
.Y(n_588)
);

MAJIxp5_ASAP7_75t_L g609 ( 
.A(n_588),
.B(n_440),
.C(n_362),
.Y(n_609)
);

OAI22xp5_ASAP7_75t_L g590 ( 
.A1(n_573),
.A2(n_563),
.B1(n_564),
.B2(n_566),
.Y(n_590)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_590),
.Y(n_626)
);

NOR3xp33_ASAP7_75t_SL g592 ( 
.A(n_585),
.B(n_545),
.C(n_551),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_592),
.B(n_600),
.Y(n_615)
);

AOI21x1_ASAP7_75t_L g624 ( 
.A1(n_593),
.A2(n_589),
.B(n_600),
.Y(n_624)
);

XNOR2xp5_ASAP7_75t_L g611 ( 
.A(n_594),
.B(n_609),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_580),
.B(n_568),
.Y(n_595)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_595),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_587),
.B(n_555),
.Y(n_598)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_598),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_567),
.B(n_497),
.Y(n_599)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_599),
.Y(n_627)
);

BUFx12_ASAP7_75t_L g600 ( 
.A(n_582),
.Y(n_600)
);

OAI22xp5_ASAP7_75t_SL g620 ( 
.A1(n_601),
.A2(n_589),
.B1(n_598),
.B2(n_608),
.Y(n_620)
);

OAI22xp5_ASAP7_75t_SL g602 ( 
.A1(n_576),
.A2(n_551),
.B1(n_542),
.B2(n_524),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_602),
.B(n_603),
.Y(n_618)
);

OAI22xp5_ASAP7_75t_SL g603 ( 
.A1(n_565),
.A2(n_542),
.B1(n_539),
.B2(n_550),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_588),
.B(n_534),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_SL g616 ( 
.A(n_604),
.B(n_605),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_584),
.B(n_550),
.Y(n_605)
);

AOI322xp5_ASAP7_75t_L g607 ( 
.A1(n_579),
.A2(n_506),
.A3(n_528),
.B1(n_552),
.B2(n_560),
.C1(n_399),
.C2(n_440),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_607),
.B(n_571),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_575),
.B(n_506),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_608),
.B(n_610),
.Y(n_622)
);

OAI22xp5_ASAP7_75t_SL g610 ( 
.A1(n_574),
.A2(n_586),
.B1(n_581),
.B2(n_577),
.Y(n_610)
);

AOI21xp5_ASAP7_75t_L g613 ( 
.A1(n_603),
.A2(n_593),
.B(n_594),
.Y(n_613)
);

AOI21xp5_ASAP7_75t_L g638 ( 
.A1(n_613),
.A2(n_617),
.B(n_619),
.Y(n_638)
);

OAI21xp5_ASAP7_75t_SL g617 ( 
.A1(n_599),
.A2(n_574),
.B(n_575),
.Y(n_617)
);

AOI21xp5_ASAP7_75t_L g619 ( 
.A1(n_595),
.A2(n_571),
.B(n_572),
.Y(n_619)
);

AOI22xp5_ASAP7_75t_L g634 ( 
.A1(n_620),
.A2(n_621),
.B1(n_614),
.B2(n_627),
.Y(n_634)
);

OAI21xp5_ASAP7_75t_SL g623 ( 
.A1(n_601),
.A2(n_569),
.B(n_399),
.Y(n_623)
);

OAI21xp5_ASAP7_75t_SL g631 ( 
.A1(n_623),
.A2(n_597),
.B(n_600),
.Y(n_631)
);

OAI21xp5_ASAP7_75t_L g640 ( 
.A1(n_624),
.A2(n_319),
.B(n_244),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_592),
.B(n_591),
.Y(n_625)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_625),
.Y(n_629)
);

MAJIxp5_ASAP7_75t_L g628 ( 
.A(n_606),
.B(n_361),
.C(n_358),
.Y(n_628)
);

MAJIxp5_ASAP7_75t_L g630 ( 
.A(n_628),
.B(n_606),
.C(n_596),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_630),
.B(n_632),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_631),
.B(n_634),
.Y(n_646)
);

MAJIxp5_ASAP7_75t_L g632 ( 
.A(n_617),
.B(n_596),
.C(n_610),
.Y(n_632)
);

OAI22xp5_ASAP7_75t_L g633 ( 
.A1(n_625),
.A2(n_602),
.B1(n_609),
.B2(n_362),
.Y(n_633)
);

MAJIxp5_ASAP7_75t_L g644 ( 
.A(n_633),
.B(n_635),
.C(n_641),
.Y(n_644)
);

MAJIxp5_ASAP7_75t_L g635 ( 
.A(n_622),
.B(n_309),
.C(n_342),
.Y(n_635)
);

OAI22xp5_ASAP7_75t_SL g636 ( 
.A1(n_613),
.A2(n_192),
.B1(n_197),
.B2(n_309),
.Y(n_636)
);

AOI22xp5_ASAP7_75t_SL g649 ( 
.A1(n_636),
.A2(n_620),
.B1(n_612),
.B2(n_627),
.Y(n_649)
);

XNOR2xp5_ASAP7_75t_SL g637 ( 
.A(n_619),
.B(n_347),
.Y(n_637)
);

MAJIxp5_ASAP7_75t_L g654 ( 
.A(n_637),
.B(n_612),
.C(n_228),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_616),
.B(n_342),
.Y(n_639)
);

AOI21xp5_ASAP7_75t_SL g652 ( 
.A1(n_639),
.A2(n_628),
.B(n_623),
.Y(n_652)
);

CKINVDCx20_ASAP7_75t_R g653 ( 
.A(n_640),
.Y(n_653)
);

XNOR2xp5_ASAP7_75t_L g641 ( 
.A(n_611),
.B(n_319),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_615),
.Y(n_642)
);

NOR4xp25_ASAP7_75t_L g647 ( 
.A(n_642),
.B(n_614),
.C(n_626),
.D(n_618),
.Y(n_647)
);

MAJIxp5_ASAP7_75t_L g643 ( 
.A(n_622),
.B(n_244),
.C(n_256),
.Y(n_643)
);

MAJIxp5_ASAP7_75t_L g648 ( 
.A(n_643),
.B(n_630),
.C(n_641),
.Y(n_648)
);

OAI21xp5_ASAP7_75t_SL g645 ( 
.A1(n_638),
.A2(n_615),
.B(n_624),
.Y(n_645)
);

AOI21xp5_ASAP7_75t_L g660 ( 
.A1(n_645),
.A2(n_647),
.B(n_638),
.Y(n_660)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_648),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_649),
.B(n_651),
.Y(n_656)
);

MAJIxp5_ASAP7_75t_L g651 ( 
.A(n_632),
.B(n_611),
.C(n_618),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_652),
.B(n_654),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_650),
.B(n_629),
.Y(n_655)
);

OR2x2_ASAP7_75t_L g666 ( 
.A(n_655),
.B(n_658),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_646),
.B(n_634),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_660),
.B(n_661),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_644),
.B(n_635),
.Y(n_661)
);

AOI22xp5_ASAP7_75t_SL g662 ( 
.A1(n_653),
.A2(n_636),
.B1(n_637),
.B2(n_640),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_662),
.B(n_228),
.Y(n_667)
);

MAJIxp5_ASAP7_75t_L g663 ( 
.A(n_657),
.B(n_656),
.C(n_659),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_663),
.B(n_664),
.Y(n_669)
);

MAJIxp5_ASAP7_75t_L g664 ( 
.A(n_661),
.B(n_643),
.C(n_653),
.Y(n_664)
);

AOI22xp5_ASAP7_75t_L g668 ( 
.A1(n_667),
.A2(n_282),
.B1(n_287),
.B2(n_289),
.Y(n_668)
);

OAI21xp5_ASAP7_75t_L g670 ( 
.A1(n_668),
.A2(n_665),
.B(n_666),
.Y(n_670)
);

AOI21xp5_ASAP7_75t_L g671 ( 
.A1(n_670),
.A2(n_669),
.B(n_234),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_671),
.B(n_277),
.Y(n_672)
);

BUFx24_ASAP7_75t_SL g673 ( 
.A(n_672),
.Y(n_673)
);

XNOR2xp5_ASAP7_75t_L g674 ( 
.A(n_673),
.B(n_234),
.Y(n_674)
);


endmodule