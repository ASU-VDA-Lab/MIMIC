module fake_jpeg_218_n_244 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_244);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_244;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_118;
wire n_128;
wire n_82;
wire n_96;

BUFx5_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_15),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_15),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

INVx11_ASAP7_75t_SL g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_3),
.B(n_4),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_14),
.B(n_3),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_7),
.B(n_9),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_11),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_9),
.Y(n_38)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_42),
.Y(n_111)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_43),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_0),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_44),
.B(n_58),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_10),
.Y(n_45)
);

A2O1A1Ixp33_ASAP7_75t_L g114 ( 
.A1(n_45),
.A2(n_49),
.B(n_55),
.C(n_65),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_27),
.B(n_0),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_46),
.B(n_60),
.Y(n_80)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_47),
.Y(n_98)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_48),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_31),
.B(n_10),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_53),
.Y(n_118)
);

INVx6_ASAP7_75t_SL g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx8_ASAP7_75t_L g106 ( 
.A(n_54),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_30),
.B(n_0),
.Y(n_55)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_57),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_19),
.B(n_26),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_59),
.Y(n_109)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_61),
.B(n_67),
.Y(n_84)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_62),
.B(n_63),
.Y(n_86)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_64),
.B(n_21),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_38),
.B(n_1),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_17),
.Y(n_66)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_17),
.Y(n_68)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_68),
.Y(n_110)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_69),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_70),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g117 ( 
.A(n_71),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_18),
.B(n_5),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_72),
.B(n_65),
.Y(n_85)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_28),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_73),
.B(n_77),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_32),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_74),
.Y(n_105)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_75),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_39),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_76),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_32),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_78),
.B(n_19),
.Y(n_101)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_32),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_79),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_85),
.B(n_89),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_88),
.B(n_91),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_45),
.B(n_21),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_49),
.B(n_46),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_72),
.B(n_35),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_93),
.B(n_96),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_55),
.B(n_29),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_66),
.B(n_35),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_97),
.B(n_100),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_71),
.A2(n_29),
.B(n_24),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_99),
.B(n_114),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_50),
.B(n_24),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_101),
.B(n_5),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_76),
.B(n_18),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_103),
.B(n_104),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_77),
.B(n_20),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_44),
.A2(n_20),
.B1(n_26),
.B2(n_22),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_115),
.A2(n_22),
.B1(n_32),
.B2(n_7),
.Y(n_123)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_111),
.Y(n_120)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_120),
.Y(n_169)
);

NOR2x1_ASAP7_75t_L g156 ( 
.A(n_123),
.B(n_131),
.Y(n_156)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_86),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_124),
.B(n_135),
.Y(n_172)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_84),
.Y(n_125)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_125),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_106),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_126),
.B(n_132),
.Y(n_159)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_107),
.Y(n_127)
);

INVx5_ASAP7_75t_L g175 ( 
.A(n_127),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_128),
.B(n_145),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_84),
.A2(n_32),
.B1(n_6),
.B2(n_8),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_129),
.A2(n_152),
.B1(n_149),
.B2(n_151),
.Y(n_177)
);

AND2x4_ASAP7_75t_SL g131 ( 
.A(n_108),
.B(n_8),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_106),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_81),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_133),
.B(n_139),
.Y(n_166)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_113),
.Y(n_134)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_107),
.Y(n_135)
);

NOR2x1_ASAP7_75t_L g163 ( 
.A(n_136),
.B(n_142),
.Y(n_163)
);

BUFx24_ASAP7_75t_L g137 ( 
.A(n_107),
.Y(n_137)
);

INVx13_ASAP7_75t_L g138 ( 
.A(n_102),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_138),
.Y(n_167)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_119),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_92),
.A2(n_80),
.B1(n_98),
.B2(n_95),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_140),
.A2(n_146),
.B1(n_123),
.B2(n_153),
.Y(n_162)
);

MAJx2_ASAP7_75t_L g141 ( 
.A(n_81),
.B(n_112),
.C(n_87),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_141),
.B(n_154),
.Y(n_168)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_119),
.Y(n_143)
);

OR2x2_ASAP7_75t_L g174 ( 
.A(n_143),
.B(n_150),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_118),
.A2(n_112),
.B(n_90),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_144),
.A2(n_148),
.B(n_149),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_110),
.B(n_116),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_82),
.A2(n_110),
.B1(n_83),
.B2(n_117),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_117),
.A2(n_83),
.B(n_109),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_109),
.B(n_116),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_94),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_94),
.B(n_117),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_151),
.A2(n_153),
.B(n_144),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_102),
.A2(n_23),
.B1(n_84),
.B2(n_67),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_82),
.A2(n_84),
.B(n_99),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_105),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_105),
.B(n_91),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_155),
.B(n_121),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_128),
.B(n_105),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_158),
.B(n_160),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_128),
.B(n_142),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_162),
.A2(n_164),
.B1(n_161),
.B2(n_158),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_163),
.A2(n_177),
.B(n_178),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_140),
.A2(n_125),
.B1(n_136),
.B2(n_141),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_130),
.B(n_120),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_165),
.B(n_176),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_171),
.B(n_131),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_122),
.B(n_147),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_173),
.B(n_179),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_134),
.B(n_148),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_150),
.B(n_149),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_180),
.B(n_183),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g181 ( 
.A(n_164),
.B(n_131),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_181),
.B(n_182),
.Y(n_206)
);

FAx1_ASAP7_75t_SL g182 ( 
.A(n_163),
.B(n_151),
.CI(n_138),
.CON(n_182),
.SN(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_166),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_176),
.A2(n_143),
.B1(n_127),
.B2(n_135),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_185),
.A2(n_186),
.B(n_174),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_168),
.A2(n_137),
.B1(n_162),
.B2(n_170),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_169),
.Y(n_187)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_187),
.Y(n_202)
);

INVx13_ASAP7_75t_L g188 ( 
.A(n_167),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_188),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_163),
.B(n_137),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_192),
.B(n_156),
.Y(n_199)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_169),
.Y(n_193)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_193),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_160),
.B(n_170),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_194),
.B(n_195),
.C(n_197),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_178),
.B(n_165),
.C(n_157),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_196),
.A2(n_161),
.B1(n_156),
.B2(n_171),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_157),
.B(n_172),
.C(n_177),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_159),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_198),
.B(n_173),
.Y(n_200)
);

OR2x2_ASAP7_75t_L g213 ( 
.A(n_199),
.B(n_208),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_200),
.B(n_190),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_201),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_203),
.A2(n_192),
.B1(n_191),
.B2(n_184),
.Y(n_212)
);

AOI22x1_ASAP7_75t_SL g205 ( 
.A1(n_191),
.A2(n_156),
.B1(n_174),
.B2(n_172),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_205),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_189),
.A2(n_167),
.B(n_174),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_195),
.B(n_175),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_210),
.B(n_197),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_212),
.A2(n_220),
.B1(n_201),
.B2(n_205),
.Y(n_222)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_202),
.Y(n_214)
);

NAND3xp33_ASAP7_75t_L g228 ( 
.A(n_214),
.B(n_216),
.C(n_219),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_215),
.B(n_204),
.C(n_210),
.Y(n_223)
);

OR2x2_ASAP7_75t_L g216 ( 
.A(n_208),
.B(n_186),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_199),
.A2(n_196),
.B1(n_185),
.B2(n_184),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_207),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_221),
.B(n_211),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_222),
.B(n_223),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_224),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_215),
.B(n_204),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_225),
.B(n_226),
.Y(n_233)
);

MAJx2_ASAP7_75t_L g226 ( 
.A(n_212),
.B(n_206),
.C(n_189),
.Y(n_226)
);

XNOR2x1_ASAP7_75t_L g227 ( 
.A(n_213),
.B(n_206),
.Y(n_227)
);

AOI321xp33_ASAP7_75t_L g232 ( 
.A1(n_227),
.A2(n_181),
.A3(n_217),
.B1(n_182),
.B2(n_220),
.C(n_213),
.Y(n_232)
);

BUFx24_ASAP7_75t_SL g231 ( 
.A(n_228),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_231),
.B(n_223),
.Y(n_236)
);

OAI221xp5_ASAP7_75t_L g235 ( 
.A1(n_232),
.A2(n_226),
.B1(n_218),
.B2(n_227),
.C(n_182),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_230),
.A2(n_216),
.B(n_209),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_234),
.B(n_235),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_236),
.B(n_237),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_229),
.B(n_194),
.Y(n_237)
);

AOI211xp5_ASAP7_75t_L g240 ( 
.A1(n_234),
.A2(n_218),
.B(n_233),
.C(n_188),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_240),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_238),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_241),
.B(n_242),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_243),
.A2(n_239),
.B(n_240),
.Y(n_244)
);


endmodule