module real_aes_17361_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_800;
wire n_778;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_852;
wire n_766;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_886;
wire n_856;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_889;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_860;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_880;
wire n_146;
wire n_432;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_891;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_193;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_481;
wire n_148;
wire n_498;
wire n_765;
wire n_691;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_888;
wire n_198;
wire n_152;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
wire n_869;
AND2x4_ASAP7_75t_L g877 ( .A(n_0), .B(n_878), .Y(n_877) );
AOI22xp5_ASAP7_75t_L g613 ( .A1(n_1), .A2(n_4), .B1(n_137), .B2(n_614), .Y(n_613) );
AOI22xp33_ASAP7_75t_L g197 ( .A1(n_2), .A2(n_42), .B1(n_144), .B2(n_198), .Y(n_197) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_3), .A2(n_23), .B1(n_198), .B2(n_233), .Y(n_602) );
AOI22xp5_ASAP7_75t_L g253 ( .A1(n_5), .A2(n_16), .B1(n_134), .B2(n_254), .Y(n_253) );
AOI22xp5_ASAP7_75t_L g508 ( .A1(n_6), .A2(n_30), .B1(n_509), .B2(n_510), .Y(n_508) );
INVx1_ASAP7_75t_L g510 ( .A(n_6), .Y(n_510) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_7), .A2(n_60), .B1(n_178), .B2(n_235), .Y(n_559) );
AOI22xp5_ASAP7_75t_L g523 ( .A1(n_8), .A2(n_17), .B1(n_144), .B2(n_182), .Y(n_523) );
INVx1_ASAP7_75t_L g878 ( .A(n_9), .Y(n_878) );
CKINVDCx5p33_ASAP7_75t_R g597 ( .A(n_10), .Y(n_597) );
CKINVDCx5p33_ASAP7_75t_R g219 ( .A(n_11), .Y(n_219) );
AOI22xp5_ASAP7_75t_L g176 ( .A1(n_12), .A2(n_18), .B1(n_177), .B2(n_180), .Y(n_176) );
OR2x2_ASAP7_75t_L g489 ( .A(n_13), .B(n_39), .Y(n_489) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_14), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g257 ( .A(n_15), .Y(n_257) );
AOI22xp5_ASAP7_75t_L g133 ( .A1(n_19), .A2(n_100), .B1(n_134), .B2(n_137), .Y(n_133) );
AOI22xp33_ASAP7_75t_L g250 ( .A1(n_20), .A2(n_38), .B1(n_223), .B2(n_251), .Y(n_250) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_21), .B(n_135), .Y(n_220) );
OAI21x1_ASAP7_75t_L g152 ( .A1(n_22), .A2(n_58), .B(n_153), .Y(n_152) );
CKINVDCx5p33_ASAP7_75t_R g155 ( .A(n_24), .Y(n_155) );
CKINVDCx5p33_ASAP7_75t_R g605 ( .A(n_25), .Y(n_605) );
INVx4_ASAP7_75t_R g550 ( .A(n_26), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_27), .B(n_141), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g199 ( .A1(n_28), .A2(n_48), .B1(n_161), .B2(n_164), .Y(n_199) );
AOI22xp33_ASAP7_75t_L g163 ( .A1(n_29), .A2(n_54), .B1(n_134), .B2(n_164), .Y(n_163) );
INVx1_ASAP7_75t_L g509 ( .A(n_30), .Y(n_509) );
CKINVDCx5p33_ASAP7_75t_R g238 ( .A(n_31), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_32), .B(n_223), .Y(n_222) );
CKINVDCx5p33_ASAP7_75t_R g212 ( .A(n_33), .Y(n_212) );
NAND2xp5_ASAP7_75t_SL g582 ( .A(n_34), .B(n_198), .Y(n_582) );
INVx1_ASAP7_75t_L g616 ( .A(n_35), .Y(n_616) );
A2O1A1Ixp33_ASAP7_75t_SL g595 ( .A1(n_36), .A2(n_140), .B(n_144), .C(n_596), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_37), .A2(n_55), .B1(n_144), .B2(n_164), .Y(n_603) );
AOI22xp5_ASAP7_75t_L g231 ( .A1(n_40), .A2(n_87), .B1(n_144), .B2(n_232), .Y(n_231) );
AOI22xp33_ASAP7_75t_L g181 ( .A1(n_41), .A2(n_47), .B1(n_144), .B2(n_182), .Y(n_181) );
OAI22xp5_ASAP7_75t_L g506 ( .A1(n_43), .A2(n_507), .B1(n_508), .B2(n_511), .Y(n_506) );
CKINVDCx5p33_ASAP7_75t_R g511 ( .A(n_43), .Y(n_511) );
CKINVDCx5p33_ASAP7_75t_R g593 ( .A(n_44), .Y(n_593) );
OAI22xp5_ASAP7_75t_L g115 ( .A1(n_45), .A2(n_68), .B1(n_116), .B2(n_117), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_45), .Y(n_117) );
AOI22xp33_ASAP7_75t_L g142 ( .A1(n_46), .A2(n_59), .B1(n_134), .B2(n_143), .Y(n_142) );
INVx1_ASAP7_75t_L g579 ( .A(n_49), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_50), .B(n_144), .Y(n_581) );
CKINVDCx5p33_ASAP7_75t_R g532 ( .A(n_51), .Y(n_532) );
INVx2_ASAP7_75t_L g109 ( .A(n_52), .Y(n_109) );
INVx1_ASAP7_75t_L g487 ( .A(n_53), .Y(n_487) );
BUFx3_ASAP7_75t_L g503 ( .A(n_53), .Y(n_503) );
CKINVDCx5p33_ASAP7_75t_R g551 ( .A(n_56), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g524 ( .A1(n_57), .A2(n_88), .B1(n_144), .B2(n_164), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g160 ( .A1(n_61), .A2(n_75), .B1(n_143), .B2(n_161), .Y(n_160) );
CKINVDCx5p33_ASAP7_75t_R g526 ( .A(n_62), .Y(n_526) );
AOI22xp33_ASAP7_75t_L g210 ( .A1(n_63), .A2(n_77), .B1(n_144), .B2(n_182), .Y(n_210) );
AOI22xp5_ASAP7_75t_L g209 ( .A1(n_64), .A2(n_97), .B1(n_134), .B2(n_180), .Y(n_209) );
AND2x4_ASAP7_75t_L g130 ( .A(n_65), .B(n_131), .Y(n_130) );
INVx1_ASAP7_75t_L g153 ( .A(n_66), .Y(n_153) );
CKINVDCx5p33_ASAP7_75t_R g865 ( .A(n_67), .Y(n_865) );
INVx1_ASAP7_75t_L g116 ( .A(n_68), .Y(n_116) );
AOI22xp33_ASAP7_75t_L g612 ( .A1(n_69), .A2(n_90), .B1(n_161), .B2(n_164), .Y(n_612) );
AO22x1_ASAP7_75t_L g562 ( .A1(n_70), .A2(n_76), .B1(n_251), .B2(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g131 ( .A(n_71), .Y(n_131) );
AND2x2_ASAP7_75t_L g598 ( .A(n_72), .B(n_201), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_73), .B(n_235), .Y(n_538) );
CKINVDCx5p33_ASAP7_75t_R g591 ( .A(n_74), .Y(n_591) );
CKINVDCx14_ASAP7_75t_R g111 ( .A(n_78), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_78), .B(n_492), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_79), .B(n_198), .Y(n_533) );
INVx2_ASAP7_75t_L g141 ( .A(n_80), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g547 ( .A(n_81), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_82), .B(n_201), .Y(n_572) );
AOI22xp33_ASAP7_75t_L g234 ( .A1(n_83), .A2(n_98), .B1(n_164), .B2(n_235), .Y(n_234) );
CKINVDCx5p33_ASAP7_75t_R g168 ( .A(n_84), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_85), .B(n_151), .Y(n_560) );
CKINVDCx5p33_ASAP7_75t_R g204 ( .A(n_86), .Y(n_204) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_89), .B(n_201), .Y(n_226) );
CKINVDCx5p33_ASAP7_75t_R g188 ( .A(n_91), .Y(n_188) );
NAND2xp5_ASAP7_75t_SL g529 ( .A(n_92), .B(n_201), .Y(n_529) );
NOR2xp33_ASAP7_75t_L g485 ( .A(n_93), .B(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g859 ( .A(n_93), .Y(n_859) );
NAND2xp33_ASAP7_75t_L g224 ( .A(n_94), .B(n_135), .Y(n_224) );
A2O1A1Ixp33_ASAP7_75t_L g545 ( .A1(n_95), .A2(n_184), .B(n_235), .C(n_546), .Y(n_545) );
CKINVDCx5p33_ASAP7_75t_R g496 ( .A(n_96), .Y(n_496) );
AND2x2_ASAP7_75t_L g552 ( .A(n_99), .B(n_553), .Y(n_552) );
NAND2xp33_ASAP7_75t_L g537 ( .A(n_101), .B(n_162), .Y(n_537) );
AOI21xp33_ASAP7_75t_L g102 ( .A1(n_103), .A2(n_872), .B(n_880), .Y(n_102) );
OAI21x1_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_110), .B(n_497), .Y(n_103) );
INVx4_ASAP7_75t_SL g104 ( .A(n_105), .Y(n_104) );
BUFx6f_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
CKINVDCx11_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
BUFx6f_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g887 ( .A(n_108), .B(n_888), .Y(n_887) );
INVx3_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g500 ( .A(n_109), .Y(n_500) );
NOR2xp33_ASAP7_75t_L g868 ( .A(n_109), .B(n_869), .Y(n_868) );
NOR2xp33_ASAP7_75t_L g894 ( .A(n_109), .B(n_890), .Y(n_894) );
OAI22xp5_ASAP7_75t_L g880 ( .A1(n_110), .A2(n_111), .B1(n_881), .B2(n_891), .Y(n_880) );
AOI21x1_ASAP7_75t_L g110 ( .A1(n_111), .A2(n_112), .B(n_490), .Y(n_110) );
INVx1_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_114), .B(n_481), .Y(n_113) );
OAI21xp33_ASAP7_75t_SL g490 ( .A1(n_114), .A2(n_491), .B(n_494), .Y(n_490) );
XNOR2x1_ASAP7_75t_L g114 ( .A(n_115), .B(n_118), .Y(n_114) );
OAI22x1_ASAP7_75t_L g512 ( .A1(n_118), .A2(n_513), .B1(n_856), .B2(n_860), .Y(n_512) );
AND3x4_ASAP7_75t_L g118 ( .A(n_119), .B(n_343), .C(n_397), .Y(n_118) );
NOR2x1_ASAP7_75t_L g119 ( .A(n_120), .B(n_303), .Y(n_119) );
NAND3xp33_ASAP7_75t_L g120 ( .A(n_121), .B(n_239), .C(n_285), .Y(n_120) );
OAI21xp33_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_169), .B(n_190), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
HB1xp67_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
OR2x2_ASAP7_75t_L g335 ( .A(n_124), .B(n_243), .Y(n_335) );
INVx2_ASAP7_75t_L g361 ( .A(n_124), .Y(n_361) );
OR2x2_ASAP7_75t_L g124 ( .A(n_125), .B(n_157), .Y(n_124) );
INVx1_ASAP7_75t_L g260 ( .A(n_125), .Y(n_260) );
INVx2_ASAP7_75t_L g375 ( .A(n_125), .Y(n_375) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx2_ASAP7_75t_L g172 ( .A(n_126), .Y(n_172) );
AND2x4_ASAP7_75t_L g318 ( .A(n_126), .B(n_280), .Y(n_318) );
AO31x2_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_132), .A3(n_148), .B(n_154), .Y(n_126) );
AO31x2_ASAP7_75t_L g207 ( .A1(n_127), .A2(n_185), .A3(n_208), .B(n_211), .Y(n_207) );
INVx1_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
AOI21xp5_ASAP7_75t_L g544 ( .A1(n_128), .A2(n_545), .B(n_548), .Y(n_544) );
INVx2_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
AO31x2_ASAP7_75t_L g174 ( .A1(n_129), .A2(n_175), .A3(n_185), .B(n_187), .Y(n_174) );
AO31x2_ASAP7_75t_L g195 ( .A1(n_129), .A2(n_196), .A3(n_200), .B(n_203), .Y(n_195) );
AO31x2_ASAP7_75t_L g248 ( .A1(n_129), .A2(n_229), .A3(n_249), .B(n_256), .Y(n_248) );
AO31x2_ASAP7_75t_L g521 ( .A1(n_129), .A2(n_156), .A3(n_522), .B(n_525), .Y(n_521) );
BUFx10_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx1_ASAP7_75t_L g166 ( .A(n_130), .Y(n_166) );
BUFx10_ASAP7_75t_L g541 ( .A(n_130), .Y(n_541) );
INVx1_ASAP7_75t_L g566 ( .A(n_130), .Y(n_566) );
OAI22xp5_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_139), .B1(n_142), .B2(n_145), .Y(n_132) );
INVx3_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVxp67_ASAP7_75t_SL g563 ( .A(n_135), .Y(n_563) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx1_ASAP7_75t_L g138 ( .A(n_136), .Y(n_138) );
INVx3_ASAP7_75t_L g144 ( .A(n_136), .Y(n_144) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_136), .Y(n_162) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_136), .Y(n_164) );
INVx1_ASAP7_75t_L g179 ( .A(n_136), .Y(n_179) );
BUFx6f_ASAP7_75t_L g198 ( .A(n_136), .Y(n_198) );
INVx2_ASAP7_75t_L g233 ( .A(n_136), .Y(n_233) );
INVx1_ASAP7_75t_L g235 ( .A(n_136), .Y(n_235) );
INVx1_ASAP7_75t_L g252 ( .A(n_136), .Y(n_252) );
INVx1_ASAP7_75t_L g255 ( .A(n_136), .Y(n_255) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
NOR2xp33_ASAP7_75t_L g592 ( .A(n_138), .B(n_593), .Y(n_592) );
OAI22xp5_ASAP7_75t_L g159 ( .A1(n_139), .A2(n_145), .B1(n_160), .B2(n_163), .Y(n_159) );
OAI22xp5_ASAP7_75t_L g175 ( .A1(n_139), .A2(n_176), .B1(n_181), .B2(n_183), .Y(n_175) );
OAI22xp5_ASAP7_75t_L g196 ( .A1(n_139), .A2(n_145), .B1(n_197), .B2(n_199), .Y(n_196) );
OAI22xp5_ASAP7_75t_L g208 ( .A1(n_139), .A2(n_183), .B1(n_209), .B2(n_210), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_139), .A2(n_222), .B(n_224), .Y(n_221) );
OAI22xp5_ASAP7_75t_L g230 ( .A1(n_139), .A2(n_231), .B1(n_234), .B2(n_236), .Y(n_230) );
OAI22xp5_ASAP7_75t_L g249 ( .A1(n_139), .A2(n_145), .B1(n_250), .B2(n_253), .Y(n_249) );
OAI22x1_ASAP7_75t_L g522 ( .A1(n_139), .A2(n_236), .B1(n_523), .B2(n_524), .Y(n_522) );
OAI22xp5_ASAP7_75t_L g601 ( .A1(n_139), .A2(n_558), .B1(n_602), .B2(n_603), .Y(n_601) );
OAI22xp5_ASAP7_75t_L g611 ( .A1(n_139), .A2(n_236), .B1(n_612), .B2(n_613), .Y(n_611) );
INVx6_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
O2A1O1Ixp5_ASAP7_75t_L g218 ( .A1(n_140), .A2(n_182), .B(n_219), .C(n_220), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_140), .A2(n_537), .B(n_538), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_140), .B(n_562), .Y(n_561) );
A2O1A1Ixp33_ASAP7_75t_L g646 ( .A1(n_140), .A2(n_557), .B(n_562), .C(n_565), .Y(n_646) );
BUFx8_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx2_ASAP7_75t_L g147 ( .A(n_141), .Y(n_147) );
INVx1_ASAP7_75t_L g184 ( .A(n_141), .Y(n_184) );
INVx1_ASAP7_75t_L g578 ( .A(n_141), .Y(n_578) );
INVx1_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx1_ASAP7_75t_L g180 ( .A(n_144), .Y(n_180) );
INVx4_ASAP7_75t_L g182 ( .A(n_144), .Y(n_182) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g558 ( .A(n_146), .Y(n_558) );
BUFx3_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx2_ASAP7_75t_L g535 ( .A(n_147), .Y(n_535) );
AO31x2_ASAP7_75t_L g158 ( .A1(n_148), .A2(n_159), .A3(n_165), .B(n_167), .Y(n_158) );
AO21x2_ASAP7_75t_L g543 ( .A1(n_148), .A2(n_544), .B(n_552), .Y(n_543) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
NOR2xp33_ASAP7_75t_SL g187 ( .A(n_150), .B(n_188), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g237 ( .A(n_150), .B(n_238), .Y(n_237) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g156 ( .A(n_151), .Y(n_156) );
INVx2_ASAP7_75t_L g186 ( .A(n_151), .Y(n_186) );
OAI21xp33_ASAP7_75t_L g565 ( .A1(n_151), .A2(n_560), .B(n_566), .Y(n_565) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
BUFx6f_ASAP7_75t_L g202 ( .A(n_152), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g154 ( .A(n_155), .B(n_156), .Y(n_154) );
NOR2xp33_ASAP7_75t_L g167 ( .A(n_156), .B(n_168), .Y(n_167) );
INVx1_ASAP7_75t_L g371 ( .A(n_157), .Y(n_371) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx1_ASAP7_75t_L g189 ( .A(n_158), .Y(n_189) );
AND2x4_ASAP7_75t_L g246 ( .A(n_158), .B(n_247), .Y(n_246) );
HB1xp67_ASAP7_75t_L g277 ( .A(n_158), .Y(n_277) );
INVx2_ASAP7_75t_L g280 ( .A(n_158), .Y(n_280) );
OR2x2_ASAP7_75t_L g294 ( .A(n_158), .B(n_248), .Y(n_294) );
AND2x2_ASAP7_75t_L g396 ( .A(n_158), .B(n_174), .Y(n_396) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx1_ASAP7_75t_L g223 ( .A(n_162), .Y(n_223) );
OAI22xp33_ASAP7_75t_L g549 ( .A1(n_162), .A2(n_255), .B1(n_550), .B2(n_551), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_164), .B(n_577), .Y(n_576) );
INVx2_ASAP7_75t_L g614 ( .A(n_164), .Y(n_614) );
AO31x2_ASAP7_75t_L g228 ( .A1(n_165), .A2(n_229), .A3(n_230), .B(n_237), .Y(n_228) );
AO31x2_ASAP7_75t_L g610 ( .A1(n_165), .A2(n_185), .A3(n_611), .B(n_615), .Y(n_610) );
INVx2_ASAP7_75t_SL g165 ( .A(n_166), .Y(n_165) );
INVx2_ASAP7_75t_SL g225 ( .A(n_166), .Y(n_225) );
INVx1_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
NAND2xp5_ASAP7_75t_SL g451 ( .A(n_170), .B(n_452), .Y(n_451) );
OR2x2_ASAP7_75t_L g170 ( .A(n_171), .B(n_173), .Y(n_170) );
OR2x2_ASAP7_75t_L g278 ( .A(n_171), .B(n_279), .Y(n_278) );
NAND2xp5_ASAP7_75t_SL g342 ( .A(n_171), .B(n_297), .Y(n_342) );
AND2x2_ASAP7_75t_L g407 ( .A(n_171), .B(n_383), .Y(n_407) );
INVx4_ASAP7_75t_L g441 ( .A(n_171), .Y(n_441) );
INVx3_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
AND2x2_ASAP7_75t_L g276 ( .A(n_172), .B(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g314 ( .A(n_172), .B(n_245), .Y(n_314) );
AND2x2_ASAP7_75t_L g424 ( .A(n_172), .B(n_248), .Y(n_424) );
AND2x2_ASAP7_75t_L g458 ( .A(n_172), .B(n_280), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_174), .B(n_189), .Y(n_173) );
INVx4_ASAP7_75t_SL g245 ( .A(n_174), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_174), .B(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g359 ( .A(n_174), .B(n_248), .Y(n_359) );
BUFx2_ASAP7_75t_L g377 ( .A(n_174), .Y(n_377) );
INVx1_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g546 ( .A(n_179), .B(n_547), .Y(n_546) );
O2A1O1Ixp33_ASAP7_75t_L g531 ( .A1(n_182), .A2(n_532), .B(n_533), .C(n_534), .Y(n_531) );
INVx1_ASAP7_75t_SL g183 ( .A(n_184), .Y(n_183) );
INVx1_ASAP7_75t_L g236 ( .A(n_184), .Y(n_236) );
AOI21x1_ASAP7_75t_L g587 ( .A1(n_185), .A2(n_588), .B(n_598), .Y(n_587) );
BUFx2_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_186), .B(n_526), .Y(n_525) );
INVx2_ASAP7_75t_L g553 ( .A(n_186), .Y(n_553) );
NOR2xp33_ASAP7_75t_L g604 ( .A(n_186), .B(n_605), .Y(n_604) );
NOR2xp33_ASAP7_75t_L g615 ( .A(n_186), .B(n_616), .Y(n_615) );
AOI222xp33_ASAP7_75t_L g285 ( .A1(n_189), .A2(n_286), .B1(n_291), .B2(n_292), .C1(n_295), .C2(n_299), .Y(n_285) );
INVx1_ASAP7_75t_L g416 ( .A(n_189), .Y(n_416) );
AND2x2_ASAP7_75t_L g190 ( .A(n_191), .B(n_205), .Y(n_190) );
AND2x2_ASAP7_75t_L g453 ( .A(n_191), .B(n_265), .Y(n_453) );
INVx1_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
AND2x2_ASAP7_75t_L g474 ( .A(n_192), .B(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
AND2x4_ASAP7_75t_L g283 ( .A(n_193), .B(n_284), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_193), .B(n_266), .Y(n_422) );
INVx2_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_194), .B(n_270), .Y(n_312) );
AND2x2_ASAP7_75t_L g340 ( .A(n_194), .B(n_214), .Y(n_340) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
AND2x2_ASAP7_75t_L g269 ( .A(n_195), .B(n_270), .Y(n_269) );
OR2x2_ASAP7_75t_L g302 ( .A(n_195), .B(n_228), .Y(n_302) );
INVx1_ASAP7_75t_L g330 ( .A(n_195), .Y(n_330) );
HB1xp67_ASAP7_75t_L g436 ( .A(n_195), .Y(n_436) );
NOR2xp33_ASAP7_75t_L g590 ( .A(n_198), .B(n_591), .Y(n_590) );
AO31x2_ASAP7_75t_L g600 ( .A1(n_200), .A2(n_541), .A3(n_601), .B(n_604), .Y(n_600) );
INVx2_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
NOR2x1_ASAP7_75t_L g539 ( .A(n_201), .B(n_540), .Y(n_539) );
INVx4_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_202), .B(n_204), .Y(n_203) );
NOR2xp33_ASAP7_75t_L g211 ( .A(n_202), .B(n_212), .Y(n_211) );
INVx2_ASAP7_75t_SL g216 ( .A(n_202), .Y(n_216) );
BUFx3_ASAP7_75t_L g229 ( .A(n_202), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g256 ( .A(n_202), .B(n_257), .Y(n_256) );
AND2x2_ASAP7_75t_L g583 ( .A(n_202), .B(n_541), .Y(n_583) );
AOI222xp33_ASAP7_75t_L g385 ( .A1(n_205), .A2(n_328), .B1(n_386), .B2(n_387), .C1(n_389), .C2(n_391), .Y(n_385) );
AND2x4_ASAP7_75t_L g205 ( .A(n_206), .B(n_213), .Y(n_205) );
INVx1_ASAP7_75t_L g320 ( .A(n_206), .Y(n_320) );
BUFx2_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
INVx3_ASAP7_75t_L g266 ( .A(n_207), .Y(n_266) );
AND2x2_ASAP7_75t_L g271 ( .A(n_207), .B(n_228), .Y(n_271) );
AND2x2_ASAP7_75t_L g331 ( .A(n_207), .B(n_227), .Y(n_331) );
AND2x2_ASAP7_75t_L g319 ( .A(n_213), .B(n_320), .Y(n_319) );
AND2x4_ASAP7_75t_L g414 ( .A(n_213), .B(n_330), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_213), .B(n_421), .Y(n_420) );
AND3x1_ASAP7_75t_L g479 ( .A(n_213), .B(n_246), .C(n_480), .Y(n_479) );
AND2x4_ASAP7_75t_L g213 ( .A(n_214), .B(n_227), .Y(n_213) );
AND2x2_ASAP7_75t_L g300 ( .A(n_214), .B(n_266), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_214), .B(n_402), .Y(n_449) );
INVx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
BUFx2_ASAP7_75t_L g263 ( .A(n_215), .Y(n_263) );
OAI21x1_ASAP7_75t_L g215 ( .A1(n_216), .A2(n_217), .B(n_226), .Y(n_215) );
OAI21x1_ASAP7_75t_L g270 ( .A1(n_216), .A2(n_217), .B(n_226), .Y(n_270) );
OAI21x1_ASAP7_75t_L g217 ( .A1(n_218), .A2(n_221), .B(n_225), .Y(n_217) );
INVx2_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
AND2x4_ASAP7_75t_L g265 ( .A(n_228), .B(n_266), .Y(n_265) );
OR2x2_ASAP7_75t_L g298 ( .A(n_228), .B(n_284), .Y(n_298) );
INVx1_ASAP7_75t_L g308 ( .A(n_228), .Y(n_308) );
BUFx2_ASAP7_75t_L g402 ( .A(n_228), .Y(n_402) );
INVx2_ASAP7_75t_SL g232 ( .A(n_233), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g596 ( .A(n_233), .B(n_597), .Y(n_596) );
NAND2xp5_ASAP7_75t_SL g548 ( .A(n_236), .B(n_549), .Y(n_548) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_240), .A2(n_261), .B(n_267), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
NAND2x1_ASAP7_75t_L g241 ( .A(n_242), .B(n_258), .Y(n_241) );
AOI221xp5_ASAP7_75t_SL g325 ( .A1(n_242), .A2(n_326), .B1(n_332), .B2(n_336), .C(n_341), .Y(n_325) );
AND2x4_ASAP7_75t_L g242 ( .A(n_243), .B(n_246), .Y(n_242) );
INVx2_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_244), .B(n_260), .Y(n_446) );
INVx2_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_245), .B(n_280), .Y(n_279) );
AND2x4_ASAP7_75t_L g288 ( .A(n_245), .B(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g324 ( .A(n_245), .Y(n_324) );
INVx1_ASAP7_75t_L g334 ( .A(n_245), .Y(n_334) );
AND2x2_ASAP7_75t_L g353 ( .A(n_245), .B(n_354), .Y(n_353) );
OR2x2_ASAP7_75t_L g365 ( .A(n_245), .B(n_366), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_245), .B(n_371), .Y(n_478) );
INVx2_ASAP7_75t_L g313 ( .A(n_246), .Y(n_313) );
AND2x2_ASAP7_75t_L g323 ( .A(n_246), .B(n_324), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_246), .B(n_334), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_246), .B(n_467), .Y(n_466) );
INVx2_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
INVx1_ASAP7_75t_L g274 ( .A(n_248), .Y(n_274) );
HB1xp67_ASAP7_75t_L g317 ( .A(n_248), .Y(n_317) );
INVx1_ASAP7_75t_L g354 ( .A(n_248), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_248), .B(n_371), .Y(n_370) );
OAI21xp33_ASAP7_75t_SL g574 ( .A1(n_251), .A2(n_575), .B(n_576), .Y(n_574) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
OR2x2_ASAP7_75t_L g293 ( .A(n_259), .B(n_294), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_259), .B(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
HB1xp67_ASAP7_75t_L g352 ( .A(n_260), .Y(n_352) );
NOR2xp33_ASAP7_75t_R g261 ( .A(n_262), .B(n_264), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
NOR3xp33_ASAP7_75t_L g341 ( .A(n_263), .B(n_333), .C(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_L g364 ( .A(n_263), .B(n_271), .Y(n_364) );
AND2x2_ASAP7_75t_L g393 ( .A(n_263), .B(n_363), .Y(n_393) );
OR2x2_ASAP7_75t_L g460 ( .A(n_263), .B(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
AND2x4_ASAP7_75t_L g386 ( .A(n_265), .B(n_269), .Y(n_386) );
INVx2_ASAP7_75t_SL g470 ( .A(n_265), .Y(n_470) );
INVx2_ASAP7_75t_L g297 ( .A(n_266), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_266), .B(n_311), .Y(n_310) );
INVx3_ASAP7_75t_L g339 ( .A(n_266), .Y(n_339) );
HB1xp67_ASAP7_75t_L g412 ( .A(n_266), .Y(n_412) );
OAI32xp33_ASAP7_75t_L g267 ( .A1(n_268), .A2(n_272), .A3(n_275), .B1(n_278), .B2(n_281), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_269), .B(n_271), .Y(n_268) );
AND2x2_ASAP7_75t_L g291 ( .A(n_269), .B(n_271), .Y(n_291) );
AND2x2_ASAP7_75t_L g349 ( .A(n_269), .B(n_331), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_269), .B(n_331), .Y(n_357) );
INVx1_ASAP7_75t_L g284 ( .A(n_270), .Y(n_284) );
AND2x4_ASAP7_75t_SL g282 ( .A(n_271), .B(n_283), .Y(n_282) );
INVx1_ASAP7_75t_SL g426 ( .A(n_271), .Y(n_426) );
INVx2_ASAP7_75t_L g461 ( .A(n_271), .Y(n_461) );
AND2x2_ASAP7_75t_L g473 ( .A(n_271), .B(n_340), .Y(n_473) );
NOR3xp33_ASAP7_75t_L g403 ( .A(n_272), .B(n_394), .C(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
INVx1_ASAP7_75t_L g289 ( .A(n_274), .Y(n_289) );
AOI321xp33_ASAP7_75t_L g472 ( .A1(n_275), .A2(n_334), .A3(n_473), .B1(n_474), .B2(n_476), .C(n_479), .Y(n_472) );
INVx2_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
INVx1_ASAP7_75t_L g290 ( .A(n_277), .Y(n_290) );
OAI22xp5_ASAP7_75t_L g476 ( .A1(n_279), .A2(n_298), .B1(n_477), .B2(n_478), .Y(n_476) );
INVx3_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g379 ( .A(n_283), .B(n_338), .Y(n_379) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
NAND2xp5_ASAP7_75t_SL g287 ( .A(n_288), .B(n_290), .Y(n_287) );
INVx1_ASAP7_75t_L g413 ( .A(n_288), .Y(n_413) );
NAND2x1_ASAP7_75t_L g440 ( .A(n_288), .B(n_441), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_288), .B(n_458), .Y(n_457) );
AND2x2_ASAP7_75t_L g438 ( .A(n_290), .B(n_424), .Y(n_438) );
INVx2_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
INVx2_ASAP7_75t_L g378 ( .A(n_294), .Y(n_378) );
OR2x2_ASAP7_75t_L g445 ( .A(n_294), .B(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
OR2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
NOR2xp33_ASAP7_75t_L g322 ( .A(n_297), .B(n_298), .Y(n_322) );
NOR2x1p5_ASAP7_75t_L g363 ( .A(n_297), .B(n_302), .Y(n_363) );
INVx1_ASAP7_75t_L g433 ( .A(n_297), .Y(n_433) );
NOR2x1_ASAP7_75t_L g434 ( .A(n_298), .B(n_435), .Y(n_434) );
AND2x2_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
INVxp67_ASAP7_75t_SL g477 ( .A(n_300), .Y(n_477) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
NAND3xp33_ASAP7_75t_L g303 ( .A(n_304), .B(n_315), .C(n_325), .Y(n_303) );
NAND3xp33_ASAP7_75t_L g304 ( .A(n_305), .B(n_313), .C(n_314), .Y(n_304) );
AND2x4_ASAP7_75t_L g305 ( .A(n_306), .B(n_309), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
BUFx2_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g455 ( .A(n_309), .Y(n_455) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVxp67_ASAP7_75t_SL g311 ( .A(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g347 ( .A(n_312), .Y(n_347) );
INVx1_ASAP7_75t_L g383 ( .A(n_312), .Y(n_383) );
NAND2xp33_ASAP7_75t_L g387 ( .A(n_313), .B(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g391 ( .A(n_313), .Y(n_391) );
INVx1_ASAP7_75t_L g417 ( .A(n_314), .Y(n_417) );
AOI21xp5_ASAP7_75t_L g315 ( .A1(n_316), .A2(n_319), .B(n_321), .Y(n_315) );
AND2x4_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
INVx3_ASAP7_75t_L g366 ( .A(n_318), .Y(n_366) );
AND2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
INVxp67_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g328 ( .A(n_329), .B(n_331), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g443 ( .A(n_330), .B(n_433), .Y(n_443) );
AND2x2_ASAP7_75t_L g346 ( .A(n_331), .B(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g411 ( .A(n_331), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_333), .B(n_335), .Y(n_332) );
OR2x2_ASAP7_75t_L g369 ( .A(n_334), .B(n_370), .Y(n_369) );
INVx2_ASAP7_75t_L g348 ( .A(n_335), .Y(n_348) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_338), .B(n_340), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
AND2x4_ASAP7_75t_L g382 ( .A(n_339), .B(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g471 ( .A(n_340), .Y(n_471) );
NOR2xp67_ASAP7_75t_L g343 ( .A(n_344), .B(n_380), .Y(n_343) );
NAND3xp33_ASAP7_75t_SL g344 ( .A(n_345), .B(n_355), .C(n_367), .Y(n_344) );
AOI22xp33_ASAP7_75t_L g345 ( .A1(n_346), .A2(n_348), .B1(n_349), .B2(n_350), .Y(n_345) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_352), .B(n_353), .Y(n_351) );
INVx1_ASAP7_75t_L g388 ( .A(n_353), .Y(n_388) );
AND2x2_ASAP7_75t_L g463 ( .A(n_353), .B(n_374), .Y(n_463) );
INVx1_ASAP7_75t_L g410 ( .A(n_354), .Y(n_410) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
OAI32xp33_ASAP7_75t_L g356 ( .A1(n_357), .A2(n_358), .A3(n_360), .B1(n_362), .B2(n_365), .Y(n_356) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx2_ASAP7_75t_L g390 ( .A(n_359), .Y(n_390) );
NAND2x1_ASAP7_75t_L g428 ( .A(n_359), .B(n_429), .Y(n_428) );
HB1xp67_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g389 ( .A(n_361), .B(n_390), .Y(n_389) );
NOR2x1_ASAP7_75t_L g362 ( .A(n_363), .B(n_364), .Y(n_362) );
OAI211xp5_ASAP7_75t_SL g415 ( .A1(n_366), .A2(n_409), .B(n_416), .C(n_417), .Y(n_415) );
INVx2_ASAP7_75t_L g429 ( .A(n_366), .Y(n_429) );
OAI21xp5_ASAP7_75t_L g367 ( .A1(n_368), .A2(n_372), .B(n_379), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_373), .Y(n_384) );
NAND2x1_ASAP7_75t_L g373 ( .A(n_374), .B(n_376), .Y(n_373) );
INVx2_ASAP7_75t_L g467 ( .A(n_374), .Y(n_467) );
INVx3_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g475 ( .A(n_375), .B(n_410), .Y(n_475) );
AND2x2_ASAP7_75t_L g480 ( .A(n_375), .B(n_436), .Y(n_480) );
AND2x4_ASAP7_75t_L g376 ( .A(n_377), .B(n_378), .Y(n_376) );
INVx1_ASAP7_75t_L g405 ( .A(n_378), .Y(n_405) );
OAI211xp5_ASAP7_75t_L g380 ( .A1(n_381), .A2(n_384), .B(n_385), .C(n_392), .Y(n_380) );
INVxp67_ASAP7_75t_SL g381 ( .A(n_382), .Y(n_381) );
NAND2x1p5_ASAP7_75t_L g399 ( .A(n_382), .B(n_400), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_393), .B(n_394), .Y(n_392) );
INVx2_ASAP7_75t_SL g394 ( .A(n_395), .Y(n_394) );
NOR3xp33_ASAP7_75t_L g397 ( .A(n_398), .B(n_430), .C(n_459), .Y(n_397) );
OAI211xp5_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_403), .B(n_406), .C(n_418), .Y(n_398) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
AOI22xp5_ASAP7_75t_L g442 ( .A1(n_404), .A2(n_443), .B1(n_444), .B2(n_447), .Y(n_442) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
AOI22xp5_ASAP7_75t_L g406 ( .A1(n_407), .A2(n_408), .B1(n_414), .B2(n_415), .Y(n_406) );
OAI22xp33_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_411), .B1(n_412), .B2(n_413), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_409), .B(n_441), .Y(n_452) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
AND2x2_ASAP7_75t_L g423 ( .A(n_416), .B(n_424), .Y(n_423) );
AOI22xp5_ASAP7_75t_L g418 ( .A1(n_419), .A2(n_423), .B1(n_425), .B2(n_427), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
OR2x2_ASAP7_75t_L g448 ( .A(n_422), .B(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
OAI211xp5_ASAP7_75t_SL g430 ( .A1(n_431), .A2(n_437), .B(n_442), .C(n_450), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_433), .B(n_434), .Y(n_432) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
NOR2xp33_ASAP7_75t_L g437 ( .A(n_438), .B(n_439), .Y(n_437) );
INVx2_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx2_ASAP7_75t_SL g447 ( .A(n_448), .Y(n_447) );
AOI22xp5_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_453), .B1(n_454), .B2(n_456), .Y(n_450) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
OAI211xp5_ASAP7_75t_SL g459 ( .A1(n_460), .A2(n_462), .B(n_464), .C(n_472), .Y(n_459) );
INVxp67_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_465), .B(n_468), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
OR2x2_ASAP7_75t_L g469 ( .A(n_470), .B(n_471), .Y(n_469) );
INVx3_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx3_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
CKINVDCx8_ASAP7_75t_R g483 ( .A(n_484), .Y(n_483) );
INVx4_ASAP7_75t_L g493 ( .A(n_484), .Y(n_493) );
INVx5_ASAP7_75t_L g879 ( .A(n_484), .Y(n_879) );
INVx3_ASAP7_75t_L g890 ( .A(n_484), .Y(n_890) );
AND2x6_ASAP7_75t_SL g484 ( .A(n_485), .B(n_488), .Y(n_484) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_488), .B(n_502), .Y(n_501) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
NOR2x1_ASAP7_75t_L g871 ( .A(n_489), .B(n_503), .Y(n_871) );
BUFx12f_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
NOR2x1_ASAP7_75t_R g495 ( .A(n_493), .B(n_496), .Y(n_495) );
INVxp67_ASAP7_75t_SL g494 ( .A(n_495), .Y(n_494) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_498), .A2(n_504), .B(n_864), .Y(n_497) );
BUFx6f_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
AND2x6_ASAP7_75t_SL g499 ( .A(n_500), .B(n_501), .Y(n_499) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
OAI22xp33_ASAP7_75t_SL g504 ( .A1(n_505), .A2(n_506), .B1(n_512), .B2(n_863), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx2_ASAP7_75t_L g863 ( .A(n_512), .Y(n_863) );
AND2x2_ASAP7_75t_L g513 ( .A(n_514), .B(n_765), .Y(n_513) );
NOR3xp33_ASAP7_75t_L g514 ( .A(n_515), .B(n_681), .C(n_712), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_516), .B(n_647), .Y(n_515) );
AOI211x1_ASAP7_75t_SL g516 ( .A1(n_517), .A2(n_567), .B(n_606), .C(n_633), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_519), .B(n_542), .Y(n_518) );
AND2x2_ASAP7_75t_L g788 ( .A(n_519), .B(n_663), .Y(n_788) );
AND2x2_ASAP7_75t_L g519 ( .A(n_520), .B(n_527), .Y(n_519) );
INVx1_ASAP7_75t_L g673 ( .A(n_520), .Y(n_673) );
OR2x2_ASAP7_75t_L g794 ( .A(n_520), .B(n_645), .Y(n_794) );
INVx2_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
AND2x2_ASAP7_75t_L g630 ( .A(n_521), .B(n_528), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_521), .B(n_645), .Y(n_644) );
INVx2_ASAP7_75t_L g662 ( .A(n_521), .Y(n_662) );
OR2x2_ASAP7_75t_L g693 ( .A(n_521), .B(n_543), .Y(n_693) );
AND2x2_ASAP7_75t_L g707 ( .A(n_521), .B(n_543), .Y(n_707) );
AND2x2_ASAP7_75t_L g744 ( .A(n_521), .B(n_700), .Y(n_744) );
BUFx2_ASAP7_75t_L g624 ( .A(n_527), .Y(n_624) );
AND2x2_ASAP7_75t_L g675 ( .A(n_527), .B(n_554), .Y(n_675) );
AND2x2_ASAP7_75t_L g818 ( .A(n_527), .B(n_543), .Y(n_818) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
BUFx3_ASAP7_75t_L g642 ( .A(n_528), .Y(n_642) );
AND2x2_ASAP7_75t_L g661 ( .A(n_528), .B(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g698 ( .A(n_528), .Y(n_698) );
AND2x2_ASAP7_75t_L g722 ( .A(n_528), .B(n_543), .Y(n_722) );
NAND2x1p5_ASAP7_75t_L g528 ( .A(n_529), .B(n_530), .Y(n_528) );
OAI21x1_ASAP7_75t_L g530 ( .A1(n_531), .A2(n_536), .B(n_539), .Y(n_530) );
INVx2_ASAP7_75t_SL g534 ( .A(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
HB1xp67_ASAP7_75t_L g622 ( .A(n_542), .Y(n_622) );
AND2x2_ASAP7_75t_L g683 ( .A(n_542), .B(n_672), .Y(n_683) );
INVx2_ASAP7_75t_L g815 ( .A(n_542), .Y(n_815) );
AND2x2_ASAP7_75t_L g542 ( .A(n_543), .B(n_554), .Y(n_542) );
INVx1_ASAP7_75t_L g620 ( .A(n_543), .Y(n_620) );
AND2x4_ASAP7_75t_L g632 ( .A(n_543), .B(n_555), .Y(n_632) );
INVx2_ASAP7_75t_L g700 ( .A(n_543), .Y(n_700) );
AND2x2_ASAP7_75t_L g699 ( .A(n_554), .B(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g706 ( .A(n_554), .Y(n_706) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g784 ( .A(n_555), .B(n_700), .Y(n_784) );
AOI21x1_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_561), .B(n_564), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
OAI21x1_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_559), .B(n_560), .Y(n_557) );
AOI21xp5_ASAP7_75t_L g580 ( .A1(n_558), .A2(n_581), .B(n_582), .Y(n_580) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
AOI21xp5_ASAP7_75t_L g588 ( .A1(n_566), .A2(n_589), .B(n_595), .Y(n_588) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_569), .B(n_584), .Y(n_568) );
OR2x2_ASAP7_75t_L g689 ( .A(n_569), .B(n_585), .Y(n_689) );
AND2x2_ASAP7_75t_L g827 ( .A(n_569), .B(n_771), .Y(n_827) );
INVx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
AND2x4_ASAP7_75t_L g608 ( .A(n_570), .B(n_609), .Y(n_608) );
OR2x2_ASAP7_75t_L g709 ( .A(n_570), .B(n_710), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_570), .B(n_651), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g764 ( .A(n_570), .B(n_627), .Y(n_764) );
INVx3_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g621 ( .A(n_571), .Y(n_621) );
AND2x2_ASAP7_75t_L g637 ( .A(n_571), .B(n_638), .Y(n_637) );
NAND2x1p5_ASAP7_75t_SL g650 ( .A(n_571), .B(n_651), .Y(n_650) );
OR2x2_ASAP7_75t_L g658 ( .A(n_571), .B(n_659), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_571), .B(n_627), .Y(n_729) );
AND2x2_ASAP7_75t_L g777 ( .A(n_571), .B(n_610), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g820 ( .A(n_571), .B(n_609), .Y(n_820) );
BUFx2_ASAP7_75t_L g839 ( .A(n_571), .Y(n_839) );
AND2x4_ASAP7_75t_L g571 ( .A(n_572), .B(n_573), .Y(n_571) );
OAI21xp5_ASAP7_75t_L g573 ( .A1(n_574), .A2(n_580), .B(n_583), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g577 ( .A(n_578), .B(n_579), .Y(n_577) );
BUFx4f_ASAP7_75t_L g594 ( .A(n_578), .Y(n_594) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
OR2x2_ASAP7_75t_L g623 ( .A(n_585), .B(n_624), .Y(n_623) );
INVx2_ASAP7_75t_L g736 ( .A(n_585), .Y(n_736) );
OR2x2_ASAP7_75t_L g585 ( .A(n_586), .B(n_599), .Y(n_585) );
NOR2xp33_ASAP7_75t_L g639 ( .A(n_586), .B(n_610), .Y(n_639) );
INVx2_ASAP7_75t_L g651 ( .A(n_586), .Y(n_651) );
AND2x2_ASAP7_75t_L g687 ( .A(n_586), .B(n_600), .Y(n_687) );
INVx2_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g627 ( .A(n_587), .Y(n_627) );
OAI21xp5_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_592), .B(n_594), .Y(n_589) );
INVx1_ASAP7_75t_L g711 ( .A(n_599), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_599), .B(n_610), .Y(n_728) );
INVx2_ASAP7_75t_SL g599 ( .A(n_600), .Y(n_599) );
BUFx2_ASAP7_75t_L g638 ( .A(n_600), .Y(n_638) );
OR2x2_ASAP7_75t_L g670 ( .A(n_600), .B(n_610), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_600), .B(n_610), .Y(n_748) );
OAI22xp5_ASAP7_75t_L g606 ( .A1(n_607), .A2(n_623), .B1(n_625), .B2(n_629), .Y(n_606) );
AOI22xp5_ASAP7_75t_L g607 ( .A1(n_608), .A2(n_617), .B1(n_621), .B2(n_622), .Y(n_607) );
INVx2_ASAP7_75t_L g628 ( .A(n_608), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_608), .B(n_687), .Y(n_701) );
AND2x2_ASAP7_75t_L g735 ( .A(n_608), .B(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx1_ASAP7_75t_L g653 ( .A(n_610), .Y(n_653) );
INVx1_ASAP7_75t_L g659 ( .A(n_610), .Y(n_659) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
OR2x2_ASAP7_75t_L g793 ( .A(n_619), .B(n_794), .Y(n_793) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g674 ( .A(n_620), .Y(n_674) );
AND3x1_ASAP7_75t_L g778 ( .A(n_620), .B(n_641), .C(n_779), .Y(n_778) );
INVx1_ASAP7_75t_L g734 ( .A(n_621), .Y(n_734) );
AND2x4_ASAP7_75t_L g770 ( .A(n_621), .B(n_771), .Y(n_770) );
INVx1_ASAP7_75t_L g808 ( .A(n_624), .Y(n_808) );
INVx1_ASAP7_75t_L g812 ( .A(n_625), .Y(n_812) );
OR2x2_ASAP7_75t_L g625 ( .A(n_626), .B(n_628), .Y(n_625) );
OR2x2_ASAP7_75t_L g785 ( .A(n_626), .B(n_786), .Y(n_785) );
INVxp67_ASAP7_75t_SL g833 ( .A(n_626), .Y(n_833) );
INVxp67_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
OR2x2_ASAP7_75t_L g733 ( .A(n_627), .B(n_711), .Y(n_733) );
AND2x2_ASAP7_75t_L g775 ( .A(n_627), .B(n_642), .Y(n_775) );
HB1xp67_ASAP7_75t_L g779 ( .A(n_627), .Y(n_779) );
NAND2xp5_ASAP7_75t_SL g629 ( .A(n_630), .B(n_631), .Y(n_629) );
O2A1O1Ixp33_ASAP7_75t_L g694 ( .A1(n_630), .A2(n_631), .B(n_695), .C(n_701), .Y(n_694) );
NAND2x1_ASAP7_75t_L g738 ( .A(n_630), .B(n_739), .Y(n_738) );
NOR2xp33_ASAP7_75t_L g834 ( .A(n_630), .B(n_788), .Y(n_834) );
INVx3_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_632), .B(n_661), .Y(n_680) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
NAND2xp5_ASAP7_75t_SL g634 ( .A(n_635), .B(n_640), .Y(n_634) );
INVx2_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_637), .B(n_639), .Y(n_636) );
INVx2_ASAP7_75t_L g656 ( .A(n_638), .Y(n_656) );
HB1xp67_ASAP7_75t_L g717 ( .A(n_639), .Y(n_717) );
NOR2xp33_ASAP7_75t_L g781 ( .A(n_640), .B(n_782), .Y(n_781) );
AND2x2_ASAP7_75t_L g640 ( .A(n_641), .B(n_643), .Y(n_640) );
AND2x2_ASAP7_75t_L g690 ( .A(n_641), .B(n_691), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_641), .B(n_707), .Y(n_754) );
NAND2x1p5_ASAP7_75t_L g760 ( .A(n_641), .B(n_761), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g855 ( .A(n_641), .B(n_699), .Y(n_855) );
INVx3_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
BUFx2_ASAP7_75t_L g838 ( .A(n_642), .Y(n_838) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx2_ASAP7_75t_L g664 ( .A(n_645), .Y(n_664) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
AOI21xp5_ASAP7_75t_L g647 ( .A1(n_648), .A2(n_660), .B(n_665), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_649), .B(n_654), .Y(n_648) );
OR2x2_ASAP7_75t_L g649 ( .A(n_650), .B(n_652), .Y(n_649) );
OAI33xp33_ASAP7_75t_L g714 ( .A1(n_650), .A2(n_655), .A3(n_715), .B1(n_716), .B2(n_718), .B3(n_719), .Y(n_714) );
OR2x2_ASAP7_75t_L g846 ( .A(n_650), .B(n_670), .Y(n_846) );
INVx2_ASAP7_75t_L g848 ( .A(n_650), .Y(n_848) );
INVx1_ASAP7_75t_L g669 ( .A(n_651), .Y(n_669) );
OR2x2_ASAP7_75t_L g710 ( .A(n_651), .B(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_655), .B(n_657), .Y(n_654) );
INVx1_ASAP7_75t_L g718 ( .A(n_655), .Y(n_718) );
NOR3xp33_ASAP7_75t_L g836 ( .A(n_655), .B(n_837), .C(n_839), .Y(n_836) );
INVx2_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
NOR2xp33_ASAP7_75t_L g795 ( .A(n_656), .B(n_796), .Y(n_795) );
NOR2xp33_ASAP7_75t_L g824 ( .A(n_656), .B(n_820), .Y(n_824) );
AND2x4_ASAP7_75t_L g853 ( .A(n_656), .B(n_854), .Y(n_853) );
INVxp67_ASAP7_75t_SL g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g679 ( .A(n_658), .Y(n_679) );
OR2x2_ASAP7_75t_L g685 ( .A(n_658), .B(n_686), .Y(n_685) );
OR2x2_ASAP7_75t_L g798 ( .A(n_658), .B(n_733), .Y(n_798) );
INVx1_ASAP7_75t_L g854 ( .A(n_658), .Y(n_854) );
AND2x4_ASAP7_75t_SL g660 ( .A(n_661), .B(n_663), .Y(n_660) );
INVx1_ASAP7_75t_L g677 ( .A(n_661), .Y(n_677) );
INVx1_ASAP7_75t_L g720 ( .A(n_662), .Y(n_720) );
AND2x2_ASAP7_75t_L g761 ( .A(n_662), .B(n_664), .Y(n_761) );
INVx1_ASAP7_75t_L g801 ( .A(n_663), .Y(n_801) );
INVx2_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
OR2x2_ASAP7_75t_L g692 ( .A(n_664), .B(n_693), .Y(n_692) );
OAI22xp33_ASAP7_75t_L g665 ( .A1(n_666), .A2(n_671), .B1(n_678), .B2(n_680), .Y(n_665) );
INVx2_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx2_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
OR2x2_ASAP7_75t_L g668 ( .A(n_669), .B(n_670), .Y(n_668) );
INVx2_ASAP7_75t_L g757 ( .A(n_670), .Y(n_757) );
INVx2_ASAP7_75t_L g771 ( .A(n_670), .Y(n_771) );
AOI211xp5_ASAP7_75t_L g671 ( .A1(n_672), .A2(n_674), .B(n_675), .C(n_676), .Y(n_671) );
INVx1_ASAP7_75t_L g715 ( .A(n_672), .Y(n_715) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_673), .B(n_698), .Y(n_800) );
OR2x2_ASAP7_75t_L g816 ( .A(n_673), .B(n_817), .Y(n_816) );
INVx1_ASAP7_75t_L g829 ( .A(n_673), .Y(n_829) );
NAND2xp5_ASAP7_75t_L g804 ( .A(n_675), .B(n_743), .Y(n_804) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
NAND2xp5_ASAP7_75t_SL g681 ( .A(n_682), .B(n_702), .Y(n_681) );
AOI221xp5_ASAP7_75t_L g682 ( .A1(n_683), .A2(n_684), .B1(n_688), .B2(n_690), .C(n_694), .Y(n_682) );
INVx2_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
OAI32xp33_ASAP7_75t_L g851 ( .A1(n_685), .A2(n_782), .A3(n_800), .B1(n_852), .B2(n_855), .Y(n_851) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g821 ( .A(n_687), .Y(n_821) );
INVx2_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
OAI21xp5_ASAP7_75t_L g702 ( .A1(n_690), .A2(n_703), .B(n_708), .Y(n_702) );
NAND2x1_ASAP7_75t_L g850 ( .A(n_691), .B(n_838), .Y(n_850) );
INVx2_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx2_ASAP7_75t_L g725 ( .A(n_693), .Y(n_725) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
AND2x2_ASAP7_75t_L g696 ( .A(n_697), .B(n_699), .Y(n_696) );
AND2x2_ASAP7_75t_L g844 ( .A(n_697), .B(n_725), .Y(n_844) );
INVx2_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g792 ( .A(n_698), .Y(n_792) );
INVx2_ASAP7_75t_L g745 ( .A(n_699), .Y(n_745) );
INVx2_ASAP7_75t_SL g703 ( .A(n_704), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_705), .B(n_707), .Y(n_704) );
AND2x2_ASAP7_75t_L g721 ( .A(n_705), .B(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx2_ASAP7_75t_L g740 ( .A(n_706), .Y(n_740) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
NAND4xp25_ASAP7_75t_L g712 ( .A(n_713), .B(n_730), .C(n_741), .D(n_752), .Y(n_712) );
AOI22xp5_ASAP7_75t_L g713 ( .A1(n_714), .A2(n_721), .B1(n_723), .B2(n_726), .Y(n_713) );
OAI22xp5_ASAP7_75t_L g842 ( .A1(n_715), .A2(n_843), .B1(n_845), .B2(n_846), .Y(n_842) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
AND2x2_ASAP7_75t_L g825 ( .A(n_720), .B(n_784), .Y(n_825) );
AND2x2_ASAP7_75t_L g828 ( .A(n_722), .B(n_829), .Y(n_828) );
AOI22xp5_ASAP7_75t_L g741 ( .A1(n_723), .A2(n_742), .B1(n_746), .B2(n_749), .Y(n_741) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx2_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
OR2x2_ASAP7_75t_L g727 ( .A(n_728), .B(n_729), .Y(n_727) );
OR2x2_ASAP7_75t_L g763 ( .A(n_728), .B(n_764), .Y(n_763) );
OR2x2_ASAP7_75t_L g747 ( .A(n_729), .B(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g758 ( .A(n_729), .Y(n_758) );
OAI21xp5_ASAP7_75t_L g730 ( .A1(n_731), .A2(n_735), .B(n_737), .Y(n_730) );
O2A1O1Ixp33_ASAP7_75t_L g835 ( .A1(n_731), .A2(n_836), .B(n_840), .C(n_842), .Y(n_835) );
AND2x2_ASAP7_75t_L g731 ( .A(n_732), .B(n_734), .Y(n_731) );
INVxp67_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g810 ( .A(n_733), .Y(n_810) );
AND2x4_ASAP7_75t_L g803 ( .A(n_736), .B(n_777), .Y(n_803) );
INVx2_ASAP7_75t_SL g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_743), .B(n_745), .Y(n_742) );
OAI21xp33_ASAP7_75t_L g768 ( .A1(n_743), .A2(n_769), .B(n_772), .Y(n_768) );
INVx2_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
AND2x2_ASAP7_75t_L g774 ( .A(n_744), .B(n_775), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g807 ( .A(n_744), .B(n_808), .Y(n_807) );
INVx2_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
OR2x2_ASAP7_75t_L g750 ( .A(n_748), .B(n_751), .Y(n_750) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
OAI22xp5_ASAP7_75t_L g780 ( .A1(n_750), .A2(n_781), .B1(n_785), .B2(n_787), .Y(n_780) );
AOI22xp33_ASAP7_75t_L g752 ( .A1(n_753), .A2(n_755), .B1(n_759), .B2(n_762), .Y(n_752) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_757), .B(n_758), .Y(n_756) );
HB1xp67_ASAP7_75t_L g773 ( .A(n_757), .Y(n_773) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
NOR2xp33_ASAP7_75t_L g765 ( .A(n_766), .B(n_830), .Y(n_765) );
NAND4xp25_ASAP7_75t_L g766 ( .A(n_767), .B(n_789), .C(n_805), .D(n_822), .Y(n_766) );
NOR2xp33_ASAP7_75t_L g767 ( .A(n_768), .B(n_780), .Y(n_767) );
INVx2_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
AND2x2_ASAP7_75t_L g832 ( .A(n_770), .B(n_833), .Y(n_832) );
AOI22xp5_ASAP7_75t_L g772 ( .A1(n_773), .A2(n_774), .B1(n_776), .B2(n_778), .Y(n_772) );
INVxp67_ASAP7_75t_L g796 ( .A(n_776), .Y(n_796) );
BUFx2_ASAP7_75t_SL g776 ( .A(n_777), .Y(n_776) );
INVx1_ASAP7_75t_L g786 ( .A(n_777), .Y(n_786) );
AND2x2_ASAP7_75t_L g809 ( .A(n_777), .B(n_810), .Y(n_809) );
INVx3_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
INVx2_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
INVx1_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
AOI21xp5_ASAP7_75t_L g789 ( .A1(n_790), .A2(n_795), .B(n_797), .Y(n_789) );
NOR2x1_ASAP7_75t_L g790 ( .A(n_791), .B(n_793), .Y(n_790) );
INVx1_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
OR2x6_ASAP7_75t_L g814 ( .A(n_792), .B(n_815), .Y(n_814) );
INVx3_ASAP7_75t_L g811 ( .A(n_793), .Y(n_811) );
OAI32xp33_ASAP7_75t_L g797 ( .A1(n_798), .A2(n_799), .A3(n_801), .B1(n_802), .B2(n_804), .Y(n_797) );
INVx2_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
INVx1_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
AOI221xp5_ASAP7_75t_L g805 ( .A1(n_806), .A2(n_809), .B1(n_811), .B2(n_812), .C(n_813), .Y(n_805) );
INVx1_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
AOI21xp5_ASAP7_75t_L g813 ( .A1(n_814), .A2(n_816), .B(n_819), .Y(n_813) );
INVx2_ASAP7_75t_SL g817 ( .A(n_818), .Y(n_817) );
OR2x2_ASAP7_75t_L g819 ( .A(n_820), .B(n_821), .Y(n_819) );
NOR2x1_ASAP7_75t_L g822 ( .A(n_823), .B(n_826), .Y(n_822) );
AND2x2_ASAP7_75t_L g823 ( .A(n_824), .B(n_825), .Y(n_823) );
INVx1_ASAP7_75t_L g845 ( .A(n_824), .Y(n_845) );
INVx1_ASAP7_75t_L g841 ( .A(n_825), .Y(n_841) );
AND2x2_ASAP7_75t_L g826 ( .A(n_827), .B(n_828), .Y(n_826) );
OAI211xp5_ASAP7_75t_SL g830 ( .A1(n_831), .A2(n_834), .B(n_835), .C(n_847), .Y(n_830) );
INVx1_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
INVx1_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
INVxp67_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
INVx1_ASAP7_75t_SL g843 ( .A(n_844), .Y(n_843) );
AOI21xp33_ASAP7_75t_L g847 ( .A1(n_848), .A2(n_849), .B(n_851), .Y(n_847) );
INVx2_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
INVx2_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
CKINVDCx5p33_ASAP7_75t_R g856 ( .A(n_857), .Y(n_856) );
BUFx8_ASAP7_75t_SL g857 ( .A(n_858), .Y(n_857) );
AND2x2_ASAP7_75t_L g870 ( .A(n_858), .B(n_871), .Y(n_870) );
INVx2_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
BUFx2_ASAP7_75t_L g862 ( .A(n_859), .Y(n_862) );
INVx4_ASAP7_75t_L g860 ( .A(n_861), .Y(n_860) );
BUFx6f_ASAP7_75t_L g861 ( .A(n_862), .Y(n_861) );
NOR2xp33_ASAP7_75t_L g864 ( .A(n_865), .B(n_866), .Y(n_864) );
INVx2_ASAP7_75t_L g866 ( .A(n_867), .Y(n_866) );
BUFx10_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
INVx1_ASAP7_75t_L g869 ( .A(n_870), .Y(n_869) );
CKINVDCx20_ASAP7_75t_R g872 ( .A(n_873), .Y(n_872) );
CKINVDCx20_ASAP7_75t_R g873 ( .A(n_874), .Y(n_873) );
CKINVDCx5p33_ASAP7_75t_R g874 ( .A(n_875), .Y(n_874) );
CKINVDCx16_ASAP7_75t_R g875 ( .A(n_876), .Y(n_875) );
AND2x2_ASAP7_75t_L g876 ( .A(n_877), .B(n_879), .Y(n_876) );
INVx2_ASAP7_75t_SL g889 ( .A(n_877), .Y(n_889) );
CKINVDCx20_ASAP7_75t_R g881 ( .A(n_882), .Y(n_881) );
CKINVDCx20_ASAP7_75t_R g882 ( .A(n_883), .Y(n_882) );
CKINVDCx20_ASAP7_75t_R g883 ( .A(n_884), .Y(n_883) );
CKINVDCx20_ASAP7_75t_R g884 ( .A(n_885), .Y(n_884) );
OR2x6_ASAP7_75t_L g885 ( .A(n_886), .B(n_890), .Y(n_885) );
INVx1_ASAP7_75t_L g886 ( .A(n_887), .Y(n_886) );
OR2x4_ASAP7_75t_L g893 ( .A(n_888), .B(n_894), .Y(n_893) );
BUFx2_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
CKINVDCx6p67_ASAP7_75t_R g891 ( .A(n_892), .Y(n_891) );
BUFx3_ASAP7_75t_L g892 ( .A(n_893), .Y(n_892) );
endmodule