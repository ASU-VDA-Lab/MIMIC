module fake_jpeg_12001_n_55 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_55);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_55;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

INVx1_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

BUFx12f_ASAP7_75t_L g9 ( 
.A(n_6),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_5),
.B(n_1),
.Y(n_10)
);

INVx6_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

INVx8_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_2),
.B(n_4),
.Y(n_13)
);

BUFx10_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

BUFx4f_ASAP7_75t_SL g18 ( 
.A(n_14),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_18),
.B(n_19),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_20),
.B(n_21),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_10),
.B(n_0),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_23),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_9),
.B(n_0),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_15),
.A2(n_11),
.B1(n_16),
.B2(n_14),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_24),
.B(n_23),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_23),
.B(n_13),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_30),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_26),
.A2(n_17),
.B1(n_11),
.B2(n_12),
.Y(n_34)
);

XNOR2xp5_ASAP7_75t_L g27 ( 
.A(n_24),
.B(n_14),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_18),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_20),
.B(n_8),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_L g33 ( 
.A1(n_32),
.A2(n_19),
.B(n_8),
.Y(n_33)
);

XNOR2xp5_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_34),
.Y(n_41)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_36),
.B(n_38),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_28),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_34),
.A2(n_26),
.B1(n_29),
.B2(n_27),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_9),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_37),
.A2(n_9),
.B1(n_12),
.B2(n_18),
.Y(n_40)
);

XOR2xp5_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_1),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_42),
.B(n_33),
.C(n_9),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_45),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_SL g45 ( 
.A(n_41),
.B(n_3),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_46),
.A2(n_47),
.B(n_48),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_40),
.C(n_43),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_46),
.A2(n_1),
.B(n_3),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_L g53 ( 
.A1(n_50),
.A2(n_7),
.B(n_51),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_49),
.B(n_7),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g54 ( 
.A(n_52),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g55 ( 
.A(n_54),
.B(n_53),
.Y(n_55)
);


endmodule