module real_aes_9075_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_504;
wire n_310;
wire n_455;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_404;
wire n_147;
wire n_288;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_193;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g429 ( .A(n_0), .Y(n_429) );
INVx1_ASAP7_75t_L g464 ( .A(n_1), .Y(n_464) );
INVx1_ASAP7_75t_L g238 ( .A(n_2), .Y(n_238) );
AOI22xp33_ASAP7_75t_L g539 ( .A1(n_3), .A2(n_37), .B1(n_188), .B2(n_503), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_4), .B(n_432), .Y(n_431) );
AOI21xp33_ASAP7_75t_L g199 ( .A1(n_5), .A2(n_121), .B(n_200), .Y(n_199) );
AOI222xp33_ASAP7_75t_L g103 ( .A1(n_6), .A2(n_104), .B1(n_434), .B2(n_443), .C1(n_741), .C2(n_746), .Y(n_103) );
XNOR2xp5_ASAP7_75t_L g105 ( .A(n_6), .B(n_106), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_6), .B(n_143), .Y(n_489) );
AND2x6_ASAP7_75t_L g126 ( .A(n_7), .B(n_127), .Y(n_126) );
AOI21xp5_ASAP7_75t_L g119 ( .A1(n_8), .A2(n_120), .B(n_128), .Y(n_119) );
NOR2xp33_ASAP7_75t_L g430 ( .A(n_9), .B(n_38), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_10), .B(n_186), .Y(n_185) );
INVx1_ASAP7_75t_L g205 ( .A(n_11), .Y(n_205) );
INVx1_ASAP7_75t_L g118 ( .A(n_12), .Y(n_118) );
INVx1_ASAP7_75t_L g458 ( .A(n_13), .Y(n_458) );
INVx1_ASAP7_75t_L g138 ( .A(n_14), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_15), .B(n_212), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_16), .B(n_144), .Y(n_491) );
AO32x2_ASAP7_75t_L g537 ( .A1(n_17), .A2(n_143), .A3(n_159), .B1(n_477), .B2(n_538), .Y(n_537) );
NAND2xp5_ASAP7_75t_SL g523 ( .A(n_18), .B(n_188), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_19), .B(n_155), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_20), .B(n_144), .Y(n_467) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_21), .A2(n_49), .B1(n_188), .B2(n_503), .Y(n_540) );
NAND2xp5_ASAP7_75t_SL g148 ( .A(n_22), .B(n_121), .Y(n_148) );
AOI22xp33_ASAP7_75t_SL g504 ( .A1(n_23), .A2(n_77), .B1(n_188), .B2(n_212), .Y(n_504) );
NAND2xp5_ASAP7_75t_SL g513 ( .A(n_24), .B(n_188), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_25), .B(n_198), .Y(n_228) );
A2O1A1Ixp33_ASAP7_75t_L g134 ( .A1(n_26), .A2(n_135), .B(n_137), .C(n_139), .Y(n_134) );
BUFx6f_ASAP7_75t_L g125 ( .A(n_27), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_28), .B(n_114), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_29), .B(n_170), .Y(n_239) );
OAI22xp5_ASAP7_75t_L g730 ( .A1(n_30), .A2(n_101), .B1(n_731), .B2(n_732), .Y(n_730) );
INVx1_ASAP7_75t_L g732 ( .A(n_30), .Y(n_732) );
INVx1_ASAP7_75t_L g217 ( .A(n_31), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_32), .B(n_114), .Y(n_515) );
INVx2_ASAP7_75t_L g124 ( .A(n_33), .Y(n_124) );
NAND2xp5_ASAP7_75t_SL g472 ( .A(n_34), .B(n_188), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_35), .B(n_114), .Y(n_525) );
A2O1A1Ixp33_ASAP7_75t_L g149 ( .A1(n_36), .A2(n_126), .B(n_131), .C(n_150), .Y(n_149) );
INVx1_ASAP7_75t_L g215 ( .A(n_39), .Y(n_215) );
NAND2xp5_ASAP7_75t_SL g169 ( .A(n_40), .B(n_170), .Y(n_169) );
AOI22xp5_ASAP7_75t_L g726 ( .A1(n_41), .A2(n_727), .B1(n_728), .B2(n_729), .Y(n_726) );
CKINVDCx20_ASAP7_75t_R g727 ( .A(n_41), .Y(n_727) );
NAND2xp5_ASAP7_75t_SL g484 ( .A(n_42), .B(n_188), .Y(n_484) );
AOI22xp33_ASAP7_75t_L g502 ( .A1(n_43), .A2(n_87), .B1(n_140), .B2(n_503), .Y(n_502) );
NAND2xp5_ASAP7_75t_SL g487 ( .A(n_44), .B(n_188), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_45), .B(n_188), .Y(n_459) );
CKINVDCx16_ASAP7_75t_R g218 ( .A(n_46), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_47), .B(n_463), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_48), .B(n_121), .Y(n_189) );
AOI22xp33_ASAP7_75t_SL g495 ( .A1(n_50), .A2(n_60), .B1(n_188), .B2(n_212), .Y(n_495) );
OAI22xp5_ASAP7_75t_SL g416 ( .A1(n_51), .A2(n_417), .B1(n_420), .B2(n_421), .Y(n_416) );
CKINVDCx20_ASAP7_75t_R g420 ( .A(n_51), .Y(n_420) );
AOI22xp5_ASAP7_75t_L g211 ( .A1(n_52), .A2(n_131), .B1(n_212), .B2(n_214), .Y(n_211) );
CKINVDCx20_ASAP7_75t_R g161 ( .A(n_53), .Y(n_161) );
NAND2xp5_ASAP7_75t_SL g476 ( .A(n_54), .B(n_188), .Y(n_476) );
CKINVDCx16_ASAP7_75t_R g235 ( .A(n_55), .Y(n_235) );
NAND2xp5_ASAP7_75t_SL g519 ( .A(n_56), .B(n_188), .Y(n_519) );
A2O1A1Ixp33_ASAP7_75t_L g202 ( .A1(n_57), .A2(n_203), .B(n_204), .C(n_206), .Y(n_202) );
CKINVDCx20_ASAP7_75t_R g174 ( .A(n_58), .Y(n_174) );
INVx1_ASAP7_75t_L g201 ( .A(n_59), .Y(n_201) );
INVx1_ASAP7_75t_L g127 ( .A(n_61), .Y(n_127) );
OAI22xp5_ASAP7_75t_SL g729 ( .A1(n_62), .A2(n_730), .B1(n_733), .B2(n_734), .Y(n_729) );
CKINVDCx20_ASAP7_75t_R g734 ( .A(n_62), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_63), .B(n_188), .Y(n_465) );
INVx1_ASAP7_75t_L g117 ( .A(n_64), .Y(n_117) );
OAI22xp5_ASAP7_75t_SL g417 ( .A1(n_65), .A2(n_76), .B1(n_418), .B2(n_419), .Y(n_417) );
CKINVDCx20_ASAP7_75t_R g418 ( .A(n_65), .Y(n_418) );
CKINVDCx20_ASAP7_75t_R g439 ( .A(n_66), .Y(n_439) );
AO32x2_ASAP7_75t_L g500 ( .A1(n_67), .A2(n_143), .A3(n_180), .B1(n_477), .B2(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g475 ( .A(n_68), .Y(n_475) );
INVx1_ASAP7_75t_L g510 ( .A(n_69), .Y(n_510) );
A2O1A1Ixp33_ASAP7_75t_SL g225 ( .A1(n_70), .A2(n_155), .B(n_206), .C(n_226), .Y(n_225) );
INVxp67_ASAP7_75t_L g227 ( .A(n_71), .Y(n_227) );
NAND2xp5_ASAP7_75t_SL g511 ( .A(n_72), .B(n_212), .Y(n_511) );
INVx1_ASAP7_75t_L g442 ( .A(n_73), .Y(n_442) );
CKINVDCx20_ASAP7_75t_R g220 ( .A(n_74), .Y(n_220) );
INVx1_ASAP7_75t_L g165 ( .A(n_75), .Y(n_165) );
CKINVDCx20_ASAP7_75t_R g419 ( .A(n_76), .Y(n_419) );
A2O1A1Ixp33_ASAP7_75t_L g167 ( .A1(n_78), .A2(n_126), .B(n_131), .C(n_168), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_79), .B(n_503), .Y(n_524) );
NAND2xp5_ASAP7_75t_SL g514 ( .A(n_80), .B(n_212), .Y(n_514) );
NAND2xp5_ASAP7_75t_SL g151 ( .A(n_81), .B(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g115 ( .A(n_82), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_83), .B(n_155), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_84), .B(n_212), .Y(n_485) );
A2O1A1Ixp33_ASAP7_75t_L g236 ( .A1(n_85), .A2(n_126), .B(n_131), .C(n_237), .Y(n_236) );
OR2x2_ASAP7_75t_L g426 ( .A(n_86), .B(n_427), .Y(n_426) );
OR2x2_ASAP7_75t_L g446 ( .A(n_86), .B(n_428), .Y(n_446) );
INVx2_ASAP7_75t_L g724 ( .A(n_86), .Y(n_724) );
AOI22xp33_ASAP7_75t_L g494 ( .A1(n_88), .A2(n_102), .B1(n_212), .B2(n_213), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_89), .B(n_114), .Y(n_207) );
CKINVDCx20_ASAP7_75t_R g242 ( .A(n_90), .Y(n_242) );
A2O1A1Ixp33_ASAP7_75t_L g182 ( .A1(n_91), .A2(n_126), .B(n_131), .C(n_183), .Y(n_182) );
CKINVDCx20_ASAP7_75t_R g191 ( .A(n_92), .Y(n_191) );
INVx1_ASAP7_75t_L g224 ( .A(n_93), .Y(n_224) );
CKINVDCx16_ASAP7_75t_R g129 ( .A(n_94), .Y(n_129) );
NAND2xp5_ASAP7_75t_SL g184 ( .A(n_95), .B(n_152), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_96), .B(n_212), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_97), .B(n_143), .Y(n_142) );
AOI222xp33_ASAP7_75t_L g444 ( .A1(n_98), .A2(n_445), .B1(n_725), .B2(n_726), .C1(n_735), .C2(n_738), .Y(n_444) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_99), .A2(n_121), .B(n_223), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_100), .B(n_442), .Y(n_441) );
CKINVDCx20_ASAP7_75t_R g731 ( .A(n_101), .Y(n_731) );
OAI21xp5_ASAP7_75t_SL g104 ( .A1(n_105), .A2(n_423), .B(n_431), .Y(n_104) );
OAI22xp5_ASAP7_75t_SL g106 ( .A1(n_107), .A2(n_415), .B1(n_416), .B2(n_422), .Y(n_106) );
INVx2_ASAP7_75t_SL g422 ( .A(n_107), .Y(n_422) );
OAI22xp5_ASAP7_75t_L g735 ( .A1(n_107), .A2(n_446), .B1(n_448), .B2(n_736), .Y(n_735) );
OR4x2_ASAP7_75t_L g107 ( .A(n_108), .B(n_311), .C(n_370), .D(n_397), .Y(n_107) );
NAND3xp33_ASAP7_75t_SL g108 ( .A(n_109), .B(n_253), .C(n_278), .Y(n_108) );
O2A1O1Ixp33_ASAP7_75t_L g109 ( .A1(n_110), .A2(n_176), .B(n_196), .C(n_229), .Y(n_109) );
AOI211xp5_ASAP7_75t_SL g401 ( .A1(n_110), .A2(n_402), .B(n_404), .C(n_407), .Y(n_401) );
AND2x2_ASAP7_75t_L g110 ( .A(n_111), .B(n_145), .Y(n_110) );
INVx1_ASAP7_75t_L g276 ( .A(n_111), .Y(n_276) );
INVx1_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
OR2x2_ASAP7_75t_L g251 ( .A(n_112), .B(n_252), .Y(n_251) );
INVx2_ASAP7_75t_L g283 ( .A(n_112), .Y(n_283) );
AND2x2_ASAP7_75t_L g338 ( .A(n_112), .B(n_307), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_112), .B(n_194), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_112), .B(n_195), .Y(n_396) );
INVx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
INVx1_ASAP7_75t_L g257 ( .A(n_113), .Y(n_257) );
AND2x2_ASAP7_75t_L g300 ( .A(n_113), .B(n_163), .Y(n_300) );
AND2x2_ASAP7_75t_L g318 ( .A(n_113), .B(n_195), .Y(n_318) );
OA21x2_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_119), .B(n_142), .Y(n_113) );
INVx1_ASAP7_75t_L g175 ( .A(n_114), .Y(n_175) );
INVx2_ASAP7_75t_L g180 ( .A(n_114), .Y(n_180) );
OA21x2_ASAP7_75t_L g507 ( .A1(n_114), .A2(n_508), .B(n_515), .Y(n_507) );
OA21x2_ASAP7_75t_L g516 ( .A1(n_114), .A2(n_517), .B(n_525), .Y(n_516) );
AND2x2_ASAP7_75t_SL g114 ( .A(n_115), .B(n_116), .Y(n_114) );
AND2x2_ASAP7_75t_L g144 ( .A(n_115), .B(n_116), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_117), .B(n_118), .Y(n_116) );
BUFx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
AND2x4_ASAP7_75t_L g121 ( .A(n_122), .B(n_126), .Y(n_121) );
NAND2x1p5_ASAP7_75t_L g166 ( .A(n_122), .B(n_126), .Y(n_166) );
AND2x2_ASAP7_75t_L g122 ( .A(n_123), .B(n_125), .Y(n_122) );
INVx1_ASAP7_75t_L g463 ( .A(n_123), .Y(n_463) );
INVx1_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
INVx2_ASAP7_75t_L g132 ( .A(n_124), .Y(n_132) );
INVx1_ASAP7_75t_L g213 ( .A(n_124), .Y(n_213) );
INVx1_ASAP7_75t_L g133 ( .A(n_125), .Y(n_133) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_125), .Y(n_136) );
INVx3_ASAP7_75t_L g153 ( .A(n_125), .Y(n_153) );
INVx1_ASAP7_75t_L g155 ( .A(n_125), .Y(n_155) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_125), .Y(n_170) );
INVx4_ASAP7_75t_SL g141 ( .A(n_126), .Y(n_141) );
OAI21xp5_ASAP7_75t_L g456 ( .A1(n_126), .A2(n_457), .B(n_461), .Y(n_456) );
BUFx3_ASAP7_75t_L g477 ( .A(n_126), .Y(n_477) );
OAI21xp5_ASAP7_75t_L g482 ( .A1(n_126), .A2(n_483), .B(n_486), .Y(n_482) );
OAI21xp5_ASAP7_75t_L g508 ( .A1(n_126), .A2(n_509), .B(n_512), .Y(n_508) );
OAI21xp5_ASAP7_75t_L g517 ( .A1(n_126), .A2(n_518), .B(n_522), .Y(n_517) );
O2A1O1Ixp33_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_130), .B(n_134), .C(n_141), .Y(n_128) );
O2A1O1Ixp33_ASAP7_75t_L g200 ( .A1(n_130), .A2(n_141), .B(n_201), .C(n_202), .Y(n_200) );
O2A1O1Ixp33_ASAP7_75t_L g223 ( .A1(n_130), .A2(n_141), .B(n_224), .C(n_225), .Y(n_223) );
INVx5_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
AND2x6_ASAP7_75t_L g131 ( .A(n_132), .B(n_133), .Y(n_131) );
BUFx3_ASAP7_75t_L g140 ( .A(n_132), .Y(n_140) );
BUFx6f_ASAP7_75t_L g188 ( .A(n_132), .Y(n_188) );
INVx1_ASAP7_75t_L g503 ( .A(n_132), .Y(n_503) );
NOR2xp33_ASAP7_75t_L g137 ( .A(n_135), .B(n_138), .Y(n_137) );
INVx1_ASAP7_75t_L g460 ( .A(n_135), .Y(n_460) );
AOI21xp5_ASAP7_75t_L g512 ( .A1(n_135), .A2(n_513), .B(n_514), .Y(n_512) );
INVx4_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
OAI22xp5_ASAP7_75t_SL g214 ( .A1(n_136), .A2(n_215), .B1(n_216), .B2(n_217), .Y(n_214) );
INVx2_ASAP7_75t_L g216 ( .A(n_136), .Y(n_216) );
INVx1_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx2_ASAP7_75t_L g157 ( .A(n_140), .Y(n_157) );
OAI22xp33_ASAP7_75t_L g210 ( .A1(n_141), .A2(n_166), .B1(n_211), .B2(n_218), .Y(n_210) );
INVx4_ASAP7_75t_L g162 ( .A(n_143), .Y(n_162) );
OA21x2_ASAP7_75t_L g221 ( .A1(n_143), .A2(n_222), .B(n_228), .Y(n_221) );
OA21x2_ASAP7_75t_L g481 ( .A1(n_143), .A2(n_482), .B(n_489), .Y(n_481) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx1_ASAP7_75t_L g159 ( .A(n_144), .Y(n_159) );
INVx4_ASAP7_75t_L g250 ( .A(n_145), .Y(n_250) );
OAI21xp5_ASAP7_75t_L g305 ( .A1(n_145), .A2(n_306), .B(n_308), .Y(n_305) );
AND2x2_ASAP7_75t_L g386 ( .A(n_145), .B(n_387), .Y(n_386) );
AND2x2_ASAP7_75t_L g145 ( .A(n_146), .B(n_163), .Y(n_145) );
INVx1_ASAP7_75t_L g193 ( .A(n_146), .Y(n_193) );
AND2x2_ASAP7_75t_L g255 ( .A(n_146), .B(n_195), .Y(n_255) );
OR2x2_ASAP7_75t_L g284 ( .A(n_146), .B(n_285), .Y(n_284) );
INVx2_ASAP7_75t_L g298 ( .A(n_146), .Y(n_298) );
INVx3_ASAP7_75t_L g307 ( .A(n_146), .Y(n_307) );
AND2x2_ASAP7_75t_L g317 ( .A(n_146), .B(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g350 ( .A(n_146), .B(n_256), .Y(n_350) );
AND2x2_ASAP7_75t_L g374 ( .A(n_146), .B(n_330), .Y(n_374) );
OR2x6_ASAP7_75t_L g146 ( .A(n_147), .B(n_160), .Y(n_146) );
AOI21xp5_ASAP7_75t_SL g147 ( .A1(n_148), .A2(n_149), .B(n_158), .Y(n_147) );
AOI21xp5_ASAP7_75t_L g150 ( .A1(n_151), .A2(n_154), .B(n_156), .Y(n_150) );
O2A1O1Ixp33_ASAP7_75t_L g237 ( .A1(n_152), .A2(n_238), .B(n_239), .C(n_240), .Y(n_237) );
INVx2_ASAP7_75t_L g466 ( .A(n_152), .Y(n_466) );
AOI21xp5_ASAP7_75t_L g471 ( .A1(n_152), .A2(n_472), .B(n_473), .Y(n_471) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_152), .A2(n_484), .B(n_485), .Y(n_483) );
O2A1O1Ixp5_ASAP7_75t_SL g509 ( .A1(n_152), .A2(n_206), .B(n_510), .C(n_511), .Y(n_509) );
INVx5_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
NOR2xp33_ASAP7_75t_L g204 ( .A(n_153), .B(n_205), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_153), .B(n_227), .Y(n_226) );
OAI22xp5_ASAP7_75t_SL g501 ( .A1(n_153), .A2(n_170), .B1(n_502), .B2(n_504), .Y(n_501) );
INVx1_ASAP7_75t_L g521 ( .A(n_155), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g168 ( .A1(n_156), .A2(n_169), .B(n_171), .Y(n_168) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx1_ASAP7_75t_L g172 ( .A(n_158), .Y(n_172) );
OA21x2_ASAP7_75t_L g455 ( .A1(n_158), .A2(n_456), .B(n_467), .Y(n_455) );
OA21x2_ASAP7_75t_L g469 ( .A1(n_158), .A2(n_470), .B(n_478), .Y(n_469) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
AO21x2_ASAP7_75t_L g209 ( .A1(n_159), .A2(n_210), .B(n_219), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_159), .B(n_220), .Y(n_219) );
AO21x2_ASAP7_75t_L g233 ( .A1(n_159), .A2(n_234), .B(n_241), .Y(n_233) );
NOR2xp33_ASAP7_75t_SL g160 ( .A(n_161), .B(n_162), .Y(n_160) );
INVx3_ASAP7_75t_L g198 ( .A(n_162), .Y(n_198) );
NAND3xp33_ASAP7_75t_L g492 ( .A(n_162), .B(n_477), .C(n_493), .Y(n_492) );
AO21x1_ASAP7_75t_L g571 ( .A1(n_162), .A2(n_493), .B(n_572), .Y(n_571) );
INVx2_ASAP7_75t_L g195 ( .A(n_163), .Y(n_195) );
AND2x2_ASAP7_75t_L g410 ( .A(n_163), .B(n_252), .Y(n_410) );
AO21x2_ASAP7_75t_L g163 ( .A1(n_164), .A2(n_172), .B(n_173), .Y(n_163) );
OAI21xp5_ASAP7_75t_L g164 ( .A1(n_165), .A2(n_166), .B(n_167), .Y(n_164) );
OAI21xp5_ASAP7_75t_L g234 ( .A1(n_166), .A2(n_235), .B(n_236), .Y(n_234) );
INVx4_ASAP7_75t_L g186 ( .A(n_170), .Y(n_186) );
INVx2_ASAP7_75t_L g203 ( .A(n_170), .Y(n_203) );
OAI22xp5_ASAP7_75t_L g493 ( .A1(n_170), .A2(n_466), .B1(n_494), .B2(n_495), .Y(n_493) );
OAI22xp5_ASAP7_75t_L g538 ( .A1(n_170), .A2(n_466), .B1(n_539), .B2(n_540), .Y(n_538) );
NOR2xp33_ASAP7_75t_L g173 ( .A(n_174), .B(n_175), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g190 ( .A(n_175), .B(n_191), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_175), .B(n_242), .Y(n_241) );
AND2x2_ASAP7_75t_L g176 ( .A(n_177), .B(n_192), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g306 ( .A(n_178), .B(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g330 ( .A(n_178), .B(n_318), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_178), .B(n_307), .Y(n_392) );
INVx1_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
INVx2_ASAP7_75t_L g252 ( .A(n_179), .Y(n_252) );
AND2x2_ASAP7_75t_L g256 ( .A(n_179), .B(n_257), .Y(n_256) );
AND2x2_ASAP7_75t_L g297 ( .A(n_179), .B(n_298), .Y(n_297) );
AO21x2_ASAP7_75t_L g179 ( .A1(n_180), .A2(n_181), .B(n_190), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_182), .B(n_189), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g183 ( .A1(n_184), .A2(n_185), .B(n_187), .Y(n_183) );
HB1xp67_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx3_ASAP7_75t_L g206 ( .A(n_188), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_192), .B(n_293), .Y(n_315) );
INVx1_ASAP7_75t_L g354 ( .A(n_192), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_192), .B(n_281), .Y(n_398) );
AND2x2_ASAP7_75t_L g192 ( .A(n_193), .B(n_194), .Y(n_192) );
AND2x2_ASAP7_75t_L g261 ( .A(n_193), .B(n_256), .Y(n_261) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_195), .B(n_252), .Y(n_285) );
INVx1_ASAP7_75t_L g364 ( .A(n_195), .Y(n_364) );
AOI322xp5_ASAP7_75t_L g388 ( .A1(n_196), .A2(n_303), .A3(n_363), .B1(n_389), .B2(n_391), .C1(n_393), .C2(n_395), .Y(n_388) );
AND2x2_ASAP7_75t_SL g196 ( .A(n_197), .B(n_208), .Y(n_196) );
AND2x2_ASAP7_75t_L g243 ( .A(n_197), .B(n_221), .Y(n_243) );
INVx1_ASAP7_75t_SL g246 ( .A(n_197), .Y(n_246) );
AND2x2_ASAP7_75t_L g248 ( .A(n_197), .B(n_209), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_197), .B(n_265), .Y(n_271) );
INVx2_ASAP7_75t_L g290 ( .A(n_197), .Y(n_290) );
AND2x2_ASAP7_75t_L g303 ( .A(n_197), .B(n_304), .Y(n_303) );
OR2x2_ASAP7_75t_L g341 ( .A(n_197), .B(n_265), .Y(n_341) );
BUFx2_ASAP7_75t_L g358 ( .A(n_197), .Y(n_358) );
AND2x2_ASAP7_75t_L g372 ( .A(n_197), .B(n_232), .Y(n_372) );
OA21x2_ASAP7_75t_L g197 ( .A1(n_198), .A2(n_199), .B(n_207), .Y(n_197) );
O2A1O1Ixp5_ASAP7_75t_L g474 ( .A1(n_203), .A2(n_462), .B(n_475), .C(n_476), .Y(n_474) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_203), .A2(n_523), .B(n_524), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_208), .B(n_260), .Y(n_287) );
AND2x2_ASAP7_75t_L g414 ( .A(n_208), .B(n_290), .Y(n_414) );
AND2x2_ASAP7_75t_L g208 ( .A(n_209), .B(n_221), .Y(n_208) );
OR2x2_ASAP7_75t_L g259 ( .A(n_209), .B(n_260), .Y(n_259) );
INVx3_ASAP7_75t_L g265 ( .A(n_209), .Y(n_265) );
AND2x2_ASAP7_75t_L g310 ( .A(n_209), .B(n_233), .Y(n_310) );
NOR2xp33_ASAP7_75t_L g357 ( .A(n_209), .B(n_358), .Y(n_357) );
HB1xp67_ASAP7_75t_L g394 ( .A(n_209), .Y(n_394) );
INVx2_ASAP7_75t_L g240 ( .A(n_212), .Y(n_240) );
INVx3_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
AND2x2_ASAP7_75t_L g245 ( .A(n_221), .B(n_246), .Y(n_245) );
INVx1_ASAP7_75t_L g267 ( .A(n_221), .Y(n_267) );
BUFx2_ASAP7_75t_L g273 ( .A(n_221), .Y(n_273) );
AND2x2_ASAP7_75t_L g292 ( .A(n_221), .B(n_265), .Y(n_292) );
INVx3_ASAP7_75t_L g304 ( .A(n_221), .Y(n_304) );
OR2x2_ASAP7_75t_L g314 ( .A(n_221), .B(n_265), .Y(n_314) );
AOI31xp33_ASAP7_75t_SL g229 ( .A1(n_230), .A2(n_244), .A3(n_247), .B(n_249), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_231), .B(n_243), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_231), .B(n_266), .Y(n_277) );
OR2x2_ASAP7_75t_L g301 ( .A(n_231), .B(n_271), .Y(n_301) );
INVx1_ASAP7_75t_SL g231 ( .A(n_232), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_232), .B(n_245), .Y(n_244) );
OR2x2_ASAP7_75t_L g322 ( .A(n_232), .B(n_314), .Y(n_322) );
NOR2xp33_ASAP7_75t_L g332 ( .A(n_232), .B(n_304), .Y(n_332) );
AND2x2_ASAP7_75t_L g339 ( .A(n_232), .B(n_340), .Y(n_339) );
NAND2x1_ASAP7_75t_L g367 ( .A(n_232), .B(n_303), .Y(n_367) );
NOR2xp33_ASAP7_75t_L g368 ( .A(n_232), .B(n_358), .Y(n_368) );
AND2x2_ASAP7_75t_L g380 ( .A(n_232), .B(n_265), .Y(n_380) );
INVx3_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
INVx3_ASAP7_75t_L g260 ( .A(n_233), .Y(n_260) );
O2A1O1Ixp33_ASAP7_75t_L g457 ( .A1(n_240), .A2(n_458), .B(n_459), .C(n_460), .Y(n_457) );
INVx1_ASAP7_75t_L g326 ( .A(n_243), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_243), .B(n_380), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_245), .B(n_321), .Y(n_355) );
AND2x4_ASAP7_75t_L g266 ( .A(n_246), .B(n_267), .Y(n_266) );
CKINVDCx16_ASAP7_75t_R g247 ( .A(n_248), .Y(n_247) );
OR2x2_ASAP7_75t_L g249 ( .A(n_250), .B(n_251), .Y(n_249) );
INVx2_ASAP7_75t_L g345 ( .A(n_251), .Y(n_345) );
NOR2xp33_ASAP7_75t_L g362 ( .A(n_251), .B(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_L g293 ( .A(n_252), .B(n_283), .Y(n_293) );
AND2x2_ASAP7_75t_L g387 ( .A(n_252), .B(n_257), .Y(n_387) );
INVx1_ASAP7_75t_L g412 ( .A(n_252), .Y(n_412) );
AOI221xp5_ASAP7_75t_L g253 ( .A1(n_254), .A2(n_258), .B1(n_261), .B2(n_262), .C(n_268), .Y(n_253) );
CKINVDCx14_ASAP7_75t_R g274 ( .A(n_254), .Y(n_274) );
AND2x2_ASAP7_75t_L g254 ( .A(n_255), .B(n_256), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_255), .B(n_276), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_258), .B(n_309), .Y(n_328) );
INVx3_ASAP7_75t_SL g258 ( .A(n_259), .Y(n_258) );
OR2x2_ASAP7_75t_L g377 ( .A(n_259), .B(n_273), .Y(n_377) );
AND2x2_ASAP7_75t_L g291 ( .A(n_260), .B(n_292), .Y(n_291) );
INVx1_ASAP7_75t_L g321 ( .A(n_260), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_260), .B(n_304), .Y(n_349) );
NOR3xp33_ASAP7_75t_L g391 ( .A(n_260), .B(n_361), .C(n_392), .Y(n_391) );
AOI211xp5_ASAP7_75t_SL g324 ( .A1(n_261), .A2(n_325), .B(n_327), .C(n_335), .Y(n_324) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
OAI22xp33_ASAP7_75t_L g313 ( .A1(n_263), .A2(n_314), .B1(n_315), .B2(n_316), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_264), .B(n_266), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_264), .B(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_264), .B(n_348), .Y(n_347) );
BUFx2_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
AND2x2_ASAP7_75t_L g406 ( .A(n_266), .B(n_380), .Y(n_406) );
OAI22xp5_ASAP7_75t_L g268 ( .A1(n_269), .A2(n_274), .B1(n_275), .B2(n_277), .Y(n_268) );
NOR2xp33_ASAP7_75t_SL g269 ( .A(n_270), .B(n_272), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_272), .B(n_321), .Y(n_352) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
OAI22xp5_ASAP7_75t_L g404 ( .A1(n_275), .A2(n_367), .B1(n_398), .B2(n_405), .Y(n_404) );
AOI221xp5_ASAP7_75t_L g278 ( .A1(n_279), .A2(n_286), .B1(n_288), .B2(n_293), .C(n_294), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
OR2x2_ASAP7_75t_L g280 ( .A(n_281), .B(n_284), .Y(n_280) );
HB1xp67_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVxp67_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
OAI221xp5_ASAP7_75t_L g294 ( .A1(n_284), .A2(n_295), .B1(n_301), .B2(n_302), .C(n_305), .Y(n_294) );
INVx1_ASAP7_75t_L g337 ( .A(n_285), .Y(n_337) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
INVx1_ASAP7_75t_SL g309 ( .A(n_290), .Y(n_309) );
OR2x2_ASAP7_75t_L g382 ( .A(n_290), .B(n_314), .Y(n_382) );
AND2x2_ASAP7_75t_L g384 ( .A(n_290), .B(n_292), .Y(n_384) );
INVx1_ASAP7_75t_L g323 ( .A(n_293), .Y(n_323) );
OR2x2_ASAP7_75t_L g295 ( .A(n_296), .B(n_299), .Y(n_295) );
AOI21xp33_ASAP7_75t_SL g353 ( .A1(n_296), .A2(n_354), .B(n_355), .Y(n_353) );
OR2x2_ASAP7_75t_L g360 ( .A(n_296), .B(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g334 ( .A(n_297), .B(n_318), .Y(n_334) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
NAND2xp33_ASAP7_75t_SL g351 ( .A(n_302), .B(n_352), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_303), .B(n_321), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_304), .B(n_340), .Y(n_403) );
O2A1O1Ixp33_ASAP7_75t_L g319 ( .A1(n_307), .A2(n_320), .B(n_322), .C(n_323), .Y(n_319) );
NAND2x1_ASAP7_75t_SL g344 ( .A(n_307), .B(n_345), .Y(n_344) );
AOI22xp5_ASAP7_75t_L g356 ( .A1(n_308), .A2(n_357), .B1(n_359), .B2(n_362), .Y(n_356) );
AND2x2_ASAP7_75t_L g308 ( .A(n_309), .B(n_310), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_310), .B(n_400), .Y(n_399) );
NAND5xp2_ASAP7_75t_L g311 ( .A(n_312), .B(n_324), .C(n_342), .D(n_356), .E(n_365), .Y(n_311) );
NOR2xp33_ASAP7_75t_L g312 ( .A(n_313), .B(n_319), .Y(n_312) );
INVx1_ASAP7_75t_L g369 ( .A(n_315), .Y(n_369) );
INVx1_ASAP7_75t_SL g316 ( .A(n_317), .Y(n_316) );
AOI221xp5_ASAP7_75t_L g375 ( .A1(n_317), .A2(n_336), .B1(n_376), .B2(n_378), .C(n_381), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_318), .B(n_412), .Y(n_411) );
NOR2xp33_ASAP7_75t_L g325 ( .A(n_321), .B(n_326), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_321), .B(n_387), .Y(n_390) );
OAI22xp5_ASAP7_75t_L g327 ( .A1(n_328), .A2(n_329), .B1(n_331), .B2(n_333), .Y(n_327) );
INVx1_ASAP7_75t_SL g329 ( .A(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
AND2x2_ASAP7_75t_L g335 ( .A(n_336), .B(n_339), .Y(n_335) );
AND2x2_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
AND2x2_ASAP7_75t_L g409 ( .A(n_338), .B(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
AOI221xp5_ASAP7_75t_L g342 ( .A1(n_343), .A2(n_346), .B1(n_350), .B2(n_351), .C(n_353), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g393 ( .A(n_348), .B(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_SL g400 ( .A(n_358), .Y(n_400) );
INVx1_ASAP7_75t_SL g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
OAI21xp5_ASAP7_75t_SL g365 ( .A1(n_366), .A2(n_368), .B(n_369), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
OAI211xp5_ASAP7_75t_SL g370 ( .A1(n_371), .A2(n_373), .B(n_375), .C(n_388), .Y(n_370) );
INVx1_ASAP7_75t_SL g371 ( .A(n_372), .Y(n_371) );
A2O1A1Ixp33_ASAP7_75t_L g397 ( .A1(n_373), .A2(n_398), .B(n_399), .C(n_401), .Y(n_397) );
INVx1_ASAP7_75t_SL g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
NAND2xp5_ASAP7_75t_SL g378 ( .A(n_377), .B(n_379), .Y(n_378) );
AOI21xp33_ASAP7_75t_L g381 ( .A1(n_382), .A2(n_383), .B(n_385), .Y(n_381) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx2_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
AOI21xp33_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_411), .B(n_413), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx2_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
CKINVDCx20_ASAP7_75t_R g415 ( .A(n_416), .Y(n_415) );
CKINVDCx14_ASAP7_75t_R g421 ( .A(n_417), .Y(n_421) );
OAI22xp5_ASAP7_75t_SL g445 ( .A1(n_422), .A2(n_446), .B1(n_447), .B2(n_723), .Y(n_445) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_SL g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_SL g425 ( .A(n_426), .Y(n_425) );
HB1xp67_ASAP7_75t_L g433 ( .A(n_426), .Y(n_433) );
INVx1_ASAP7_75t_SL g745 ( .A(n_426), .Y(n_745) );
BUFx2_ASAP7_75t_L g748 ( .A(n_426), .Y(n_748) );
NOR2x2_ASAP7_75t_L g740 ( .A(n_427), .B(n_724), .Y(n_740) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
OR2x2_ASAP7_75t_L g723 ( .A(n_428), .B(n_724), .Y(n_723) );
AND2x2_ASAP7_75t_L g428 ( .A(n_429), .B(n_430), .Y(n_428) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
CKINVDCx20_ASAP7_75t_R g434 ( .A(n_435), .Y(n_434) );
CKINVDCx6p67_ASAP7_75t_R g435 ( .A(n_436), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_437), .B(n_440), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
NOR2xp33_ASAP7_75t_SL g743 ( .A(n_439), .B(n_441), .Y(n_743) );
OA21x2_ASAP7_75t_L g747 ( .A1(n_439), .A2(n_440), .B(n_748), .Y(n_747) );
INVx1_ASAP7_75t_SL g440 ( .A(n_441), .Y(n_440) );
INVxp67_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
OR5x1_ASAP7_75t_L g450 ( .A(n_451), .B(n_614), .C(n_672), .D(n_708), .E(n_715), .Y(n_450) );
NAND3xp33_ASAP7_75t_SL g451 ( .A(n_452), .B(n_560), .C(n_584), .Y(n_451) );
AOI221xp5_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_496), .B1(n_526), .B2(n_531), .C(n_541), .Y(n_452) );
OAI21xp5_ASAP7_75t_SL g694 ( .A1(n_453), .A2(n_695), .B(n_697), .Y(n_694) );
AND2x2_ASAP7_75t_L g453 ( .A(n_454), .B(n_479), .Y(n_453) );
NAND2x1p5_ASAP7_75t_L g684 ( .A(n_454), .B(n_685), .Y(n_684) );
AND2x2_ASAP7_75t_L g454 ( .A(n_455), .B(n_468), .Y(n_454) );
INVx2_ASAP7_75t_L g530 ( .A(n_455), .Y(n_530) );
AND2x2_ASAP7_75t_L g543 ( .A(n_455), .B(n_481), .Y(n_543) );
AND2x2_ASAP7_75t_L g597 ( .A(n_455), .B(n_480), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_455), .B(n_469), .Y(n_612) );
O2A1O1Ixp33_ASAP7_75t_L g461 ( .A1(n_462), .A2(n_464), .B(n_465), .C(n_466), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
AOI21xp5_ASAP7_75t_L g486 ( .A1(n_466), .A2(n_487), .B(n_488), .Y(n_486) );
AND2x2_ASAP7_75t_L g630 ( .A(n_468), .B(n_571), .Y(n_630) );
AND2x2_ASAP7_75t_L g663 ( .A(n_468), .B(n_481), .Y(n_663) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
OR2x2_ASAP7_75t_L g570 ( .A(n_469), .B(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g583 ( .A(n_469), .B(n_481), .Y(n_583) );
AND2x2_ASAP7_75t_L g590 ( .A(n_469), .B(n_571), .Y(n_590) );
HB1xp67_ASAP7_75t_L g599 ( .A(n_469), .Y(n_599) );
AND2x2_ASAP7_75t_L g606 ( .A(n_469), .B(n_480), .Y(n_606) );
INVx1_ASAP7_75t_L g637 ( .A(n_469), .Y(n_637) );
OAI21xp5_ASAP7_75t_L g470 ( .A1(n_471), .A2(n_474), .B(n_477), .Y(n_470) );
INVx1_ASAP7_75t_L g613 ( .A(n_479), .Y(n_613) );
AND2x2_ASAP7_75t_L g479 ( .A(n_480), .B(n_490), .Y(n_479) );
INVx2_ASAP7_75t_L g569 ( .A(n_480), .Y(n_569) );
AND2x2_ASAP7_75t_L g591 ( .A(n_480), .B(n_530), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_480), .B(n_637), .Y(n_642) );
INVx3_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_481), .B(n_530), .Y(n_529) );
AND2x2_ASAP7_75t_L g714 ( .A(n_481), .B(n_678), .Y(n_714) );
INVx2_ASAP7_75t_L g528 ( .A(n_490), .Y(n_528) );
INVx3_ASAP7_75t_L g629 ( .A(n_490), .Y(n_629) );
OR2x2_ASAP7_75t_L g659 ( .A(n_490), .B(n_660), .Y(n_659) );
NOR2x1_ASAP7_75t_L g685 ( .A(n_490), .B(n_569), .Y(n_685) );
AND2x4_ASAP7_75t_L g490 ( .A(n_491), .B(n_492), .Y(n_490) );
INVx1_ASAP7_75t_L g572 ( .A(n_491), .Y(n_572) );
AOI33xp33_ASAP7_75t_L g705 ( .A1(n_496), .A2(n_543), .A3(n_557), .B1(n_629), .B2(n_706), .B3(n_707), .Y(n_705) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
OR2x2_ASAP7_75t_L g497 ( .A(n_498), .B(n_505), .Y(n_497) );
OR2x2_ASAP7_75t_L g558 ( .A(n_498), .B(n_559), .Y(n_558) );
NOR2xp33_ASAP7_75t_L g617 ( .A(n_498), .B(n_555), .Y(n_617) );
OR2x2_ASAP7_75t_L g670 ( .A(n_498), .B(n_671), .Y(n_670) );
INVx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
AND2x2_ASAP7_75t_L g596 ( .A(n_499), .B(n_597), .Y(n_596) );
OR2x2_ASAP7_75t_L g621 ( .A(n_499), .B(n_505), .Y(n_621) );
AND2x2_ASAP7_75t_L g688 ( .A(n_499), .B(n_533), .Y(n_688) );
AOI21xp5_ASAP7_75t_L g713 ( .A1(n_499), .A2(n_588), .B(n_714), .Y(n_713) );
BUFx6f_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g535 ( .A(n_500), .Y(n_535) );
INVx1_ASAP7_75t_L g548 ( .A(n_500), .Y(n_548) );
AND2x2_ASAP7_75t_L g567 ( .A(n_500), .B(n_537), .Y(n_567) );
AND2x2_ASAP7_75t_L g616 ( .A(n_500), .B(n_536), .Y(n_616) );
INVx2_ASAP7_75t_SL g658 ( .A(n_505), .Y(n_658) );
OR2x2_ASAP7_75t_L g505 ( .A(n_506), .B(n_516), .Y(n_505) );
INVx2_ASAP7_75t_L g578 ( .A(n_506), .Y(n_578) );
INVx1_ASAP7_75t_L g709 ( .A(n_506), .Y(n_709) );
AND2x2_ASAP7_75t_L g722 ( .A(n_506), .B(n_603), .Y(n_722) );
INVx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx2_ASAP7_75t_L g549 ( .A(n_507), .Y(n_549) );
OR2x2_ASAP7_75t_L g555 ( .A(n_507), .B(n_556), .Y(n_555) );
HB1xp67_ASAP7_75t_L g566 ( .A(n_507), .Y(n_566) );
HB1xp67_ASAP7_75t_L g533 ( .A(n_516), .Y(n_533) );
AND2x2_ASAP7_75t_L g550 ( .A(n_516), .B(n_536), .Y(n_550) );
INVx1_ASAP7_75t_L g556 ( .A(n_516), .Y(n_556) );
INVx1_ASAP7_75t_L g563 ( .A(n_516), .Y(n_563) );
AND2x2_ASAP7_75t_L g588 ( .A(n_516), .B(n_537), .Y(n_588) );
INVx2_ASAP7_75t_L g604 ( .A(n_516), .Y(n_604) );
AND2x2_ASAP7_75t_L g697 ( .A(n_516), .B(n_698), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_516), .B(n_578), .Y(n_718) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_519), .A2(n_520), .B(n_521), .Y(n_518) );
INVx1_ASAP7_75t_SL g526 ( .A(n_527), .Y(n_526) );
OR2x2_ASAP7_75t_L g527 ( .A(n_528), .B(n_529), .Y(n_527) );
INVx2_ASAP7_75t_L g552 ( .A(n_528), .Y(n_552) );
INVx1_ASAP7_75t_L g581 ( .A(n_528), .Y(n_581) );
NOR2xp33_ASAP7_75t_L g678 ( .A(n_528), .B(n_612), .Y(n_678) );
INVx1_ASAP7_75t_SL g638 ( .A(n_529), .Y(n_638) );
INVx2_ASAP7_75t_L g559 ( .A(n_530), .Y(n_559) );
AND2x2_ASAP7_75t_L g628 ( .A(n_530), .B(n_629), .Y(n_628) );
AND2x2_ASAP7_75t_L g644 ( .A(n_530), .B(n_645), .Y(n_644) );
AND2x2_ASAP7_75t_L g531 ( .A(n_532), .B(n_534), .Y(n_531) );
INVx1_ASAP7_75t_L g706 ( .A(n_532), .Y(n_706) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
AND2x2_ASAP7_75t_L g561 ( .A(n_534), .B(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_L g664 ( .A(n_534), .B(n_654), .Y(n_664) );
AOI21xp5_ASAP7_75t_L g716 ( .A1(n_534), .A2(n_675), .B(n_717), .Y(n_716) );
AND2x2_ASAP7_75t_L g534 ( .A(n_535), .B(n_536), .Y(n_534) );
AND2x2_ASAP7_75t_L g577 ( .A(n_535), .B(n_578), .Y(n_577) );
BUFx2_ASAP7_75t_L g602 ( .A(n_535), .Y(n_602) );
INVx1_ASAP7_75t_L g626 ( .A(n_535), .Y(n_626) );
OR2x2_ASAP7_75t_L g690 ( .A(n_536), .B(n_549), .Y(n_690) );
NOR2xp67_ASAP7_75t_L g698 ( .A(n_536), .B(n_699), .Y(n_698) );
INVx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
AND2x2_ASAP7_75t_L g603 ( .A(n_537), .B(n_604), .Y(n_603) );
BUFx2_ASAP7_75t_L g610 ( .A(n_537), .Y(n_610) );
OAI22xp5_ASAP7_75t_L g541 ( .A1(n_542), .A2(n_544), .B1(n_551), .B2(n_553), .Y(n_541) );
OR2x2_ASAP7_75t_L g620 ( .A(n_542), .B(n_570), .Y(n_620) );
INVx1_ASAP7_75t_SL g542 ( .A(n_543), .Y(n_542) );
AOI222xp33_ASAP7_75t_L g661 ( .A1(n_543), .A2(n_662), .B1(n_664), .B2(n_665), .C1(n_666), .C2(n_669), .Y(n_661) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_546), .B(n_550), .Y(n_545) );
INVx1_ASAP7_75t_SL g546 ( .A(n_547), .Y(n_546) );
OR2x2_ASAP7_75t_L g608 ( .A(n_547), .B(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_548), .B(n_549), .Y(n_547) );
AND2x2_ASAP7_75t_SL g562 ( .A(n_549), .B(n_563), .Y(n_562) );
HB1xp67_ASAP7_75t_L g633 ( .A(n_549), .Y(n_633) );
AND2x2_ASAP7_75t_L g681 ( .A(n_549), .B(n_550), .Y(n_681) );
INVx1_ASAP7_75t_L g699 ( .A(n_549), .Y(n_699) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g665 ( .A(n_552), .B(n_591), .Y(n_665) );
AND2x2_ASAP7_75t_L g707 ( .A(n_552), .B(n_583), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_554), .B(n_557), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_554), .B(n_602), .Y(n_689) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
NAND2xp5_ASAP7_75t_SL g586 ( .A(n_555), .B(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
AND2x2_ASAP7_75t_L g582 ( .A(n_559), .B(n_583), .Y(n_582) );
INVx3_ASAP7_75t_L g650 ( .A(n_559), .Y(n_650) );
O2A1O1Ixp33_ASAP7_75t_L g560 ( .A1(n_561), .A2(n_564), .B(n_568), .C(n_573), .Y(n_560) );
INVxp67_ASAP7_75t_L g574 ( .A(n_561), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_562), .B(n_626), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_562), .B(n_609), .Y(n_704) );
BUFx3_ASAP7_75t_L g668 ( .A(n_563), .Y(n_668) );
INVx1_ASAP7_75t_L g575 ( .A(n_564), .Y(n_575) );
AND2x2_ASAP7_75t_L g564 ( .A(n_565), .B(n_567), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g594 ( .A(n_566), .B(n_588), .Y(n_594) );
INVx1_ASAP7_75t_SL g634 ( .A(n_567), .Y(n_634) );
NOR2xp33_ASAP7_75t_L g568 ( .A(n_569), .B(n_570), .Y(n_568) );
INVx1_ASAP7_75t_L g624 ( .A(n_569), .Y(n_624) );
AND2x2_ASAP7_75t_L g647 ( .A(n_569), .B(n_630), .Y(n_647) );
INVx1_ASAP7_75t_SL g618 ( .A(n_570), .Y(n_618) );
INVx1_ASAP7_75t_L g645 ( .A(n_571), .Y(n_645) );
AOI31xp33_ASAP7_75t_L g573 ( .A1(n_574), .A2(n_575), .A3(n_576), .B(n_579), .Y(n_573) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g666 ( .A(n_577), .B(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g640 ( .A(n_578), .Y(n_640) );
BUFx2_ASAP7_75t_L g654 ( .A(n_578), .Y(n_654) );
AND2x2_ASAP7_75t_L g682 ( .A(n_578), .B(n_603), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_580), .B(n_582), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx1_ASAP7_75t_SL g655 ( .A(n_582), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_583), .B(n_650), .Y(n_696) );
AND2x2_ASAP7_75t_L g703 ( .A(n_583), .B(n_629), .Y(n_703) );
AOI211xp5_ASAP7_75t_L g584 ( .A1(n_585), .A2(n_589), .B(n_592), .C(n_607), .Y(n_584) );
INVxp67_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVx2_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
AOI221xp5_ASAP7_75t_L g615 ( .A1(n_589), .A2(n_616), .B1(n_617), .B2(n_618), .C(n_619), .Y(n_615) );
AND2x2_ASAP7_75t_L g589 ( .A(n_590), .B(n_591), .Y(n_589) );
AND2x2_ASAP7_75t_L g623 ( .A(n_590), .B(n_624), .Y(n_623) );
INVx2_ASAP7_75t_L g660 ( .A(n_591), .Y(n_660) );
OAI32xp33_ASAP7_75t_L g592 ( .A1(n_593), .A2(n_595), .A3(n_598), .B1(n_600), .B2(n_605), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
O2A1O1Ixp33_ASAP7_75t_L g646 ( .A1(n_594), .A2(n_647), .B(n_648), .C(n_651), .Y(n_646) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_602), .B(n_603), .Y(n_601) );
OAI21xp5_ASAP7_75t_SL g710 ( .A1(n_602), .A2(n_711), .B(n_712), .Y(n_710) );
INVx1_ASAP7_75t_L g671 ( .A(n_603), .Y(n_671) );
INVxp67_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
NOR2xp33_ASAP7_75t_L g607 ( .A(n_608), .B(n_611), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_609), .B(n_640), .Y(n_639) );
AND2x2_ASAP7_75t_L g657 ( .A(n_609), .B(n_658), .Y(n_657) );
INVx2_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx1_ASAP7_75t_L g674 ( .A(n_611), .Y(n_674) );
OR2x2_ASAP7_75t_L g611 ( .A(n_612), .B(n_613), .Y(n_611) );
NAND4xp25_ASAP7_75t_SL g614 ( .A(n_615), .B(n_627), .C(n_646), .D(n_661), .Y(n_614) );
AND2x2_ASAP7_75t_L g653 ( .A(n_616), .B(n_654), .Y(n_653) );
AND2x4_ASAP7_75t_L g675 ( .A(n_616), .B(n_668), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_618), .B(n_650), .Y(n_649) );
OAI22xp5_ASAP7_75t_L g619 ( .A1(n_620), .A2(n_621), .B1(n_622), .B2(n_625), .Y(n_619) );
OAI22xp5_ASAP7_75t_L g701 ( .A1(n_620), .A2(n_671), .B1(n_702), .B2(n_704), .Y(n_701) );
O2A1O1Ixp33_ASAP7_75t_L g708 ( .A1(n_620), .A2(n_709), .B(n_710), .C(n_713), .Y(n_708) );
INVx2_ASAP7_75t_L g679 ( .A(n_621), .Y(n_679) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
AOI222xp33_ASAP7_75t_L g673 ( .A1(n_623), .A2(n_657), .B1(n_674), .B2(n_675), .C1(n_676), .C2(n_679), .Y(n_673) );
O2A1O1Ixp33_ASAP7_75t_L g627 ( .A1(n_628), .A2(n_630), .B(n_631), .C(n_635), .Y(n_627) );
INVx1_ASAP7_75t_L g693 ( .A(n_628), .Y(n_693) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
OAI22xp33_ASAP7_75t_L g635 ( .A1(n_632), .A2(n_636), .B1(n_639), .B2(n_641), .Y(n_635) );
OR2x2_ASAP7_75t_L g632 ( .A(n_633), .B(n_634), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_637), .B(n_638), .Y(n_636) );
OR2x2_ASAP7_75t_L g641 ( .A(n_642), .B(n_643), .Y(n_641) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g662 ( .A(n_644), .B(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g720 ( .A(n_647), .Y(n_720) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
OAI22xp33_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_655), .B1(n_656), .B2(n_659), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_654), .B(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g711 ( .A(n_659), .Y(n_711) );
INVx1_ASAP7_75t_L g692 ( .A(n_663), .Y(n_692) );
CKINVDCx16_ASAP7_75t_R g719 ( .A(n_665), .Y(n_719) );
INVxp67_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
NAND5xp2_ASAP7_75t_L g672 ( .A(n_673), .B(n_680), .C(n_694), .D(n_700), .E(n_705), .Y(n_672) );
INVx1_ASAP7_75t_SL g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
O2A1O1Ixp33_ASAP7_75t_L g680 ( .A1(n_681), .A2(n_682), .B(n_683), .C(n_686), .Y(n_680) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
AOI31xp33_ASAP7_75t_L g686 ( .A1(n_687), .A2(n_689), .A3(n_690), .B(n_691), .Y(n_686) );
INVx1_ASAP7_75t_L g712 ( .A(n_688), .Y(n_712) );
OR2x2_ASAP7_75t_L g691 ( .A(n_692), .B(n_693), .Y(n_691) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
OAI222xp33_ASAP7_75t_L g715 ( .A1(n_702), .A2(n_704), .B1(n_716), .B2(n_719), .C1(n_720), .C2(n_721), .Y(n_715) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx2_ASAP7_75t_SL g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g737 ( .A(n_723), .Y(n_737) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g733 ( .A(n_730), .Y(n_733) );
INVx2_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_SL g738 ( .A(n_739), .Y(n_738) );
INVx3_ASAP7_75t_SL g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_SL g741 ( .A(n_742), .Y(n_741) );
NAND2xp33_ASAP7_75t_L g742 ( .A(n_743), .B(n_744), .Y(n_742) );
INVx1_ASAP7_75t_SL g744 ( .A(n_745), .Y(n_744) );
INVx1_ASAP7_75t_SL g746 ( .A(n_747), .Y(n_746) );
endmodule