module fake_aes_8008_n_1237 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_267, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_262, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_272, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_16, n_13, n_198, n_169, n_193, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_265, n_191, n_264, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_266, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_263, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_268, n_231, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_261, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_271, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_270, n_246, n_153, n_61, n_259, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_269, n_225, n_39, n_1237);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_267;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_262;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_272;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_265;
input n_191;
input n_264;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_266;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_263;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_268;
input n_231;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_261;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_271;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_270;
input n_246;
input n_153;
input n_61;
input n_259;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_269;
input n_225;
input n_39;
output n_1237;
wire n_963;
wire n_1034;
wire n_949;
wire n_858;
wire n_646;
wire n_829;
wire n_1198;
wire n_667;
wire n_988;
wire n_311;
wire n_655;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_545;
wire n_896;
wire n_334;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_387;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_860;
wire n_1208;
wire n_305;
wire n_1201;
wire n_340;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_830;
wire n_1112;
wire n_517;
wire n_502;
wire n_543;
wire n_312;
wire n_1159;
wire n_1002;
wire n_915;
wire n_367;
wire n_314;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1018;
wire n_979;
wire n_319;
wire n_499;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_613;
wire n_648;
wire n_304;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_331;
wire n_746;
wire n_619;
wire n_501;
wire n_299;
wire n_699;
wire n_338;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1209;
wire n_926;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1099;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_954;
wire n_574;
wire n_822;
wire n_706;
wire n_823;
wire n_1181;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1199;
wire n_883;
wire n_573;
wire n_673;
wire n_1071;
wire n_1079;
wire n_315;
wire n_409;
wire n_295;
wire n_677;
wire n_283;
wire n_756;
wire n_1139;
wire n_577;
wire n_870;
wire n_790;
wire n_761;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_327;
wire n_1102;
wire n_723;
wire n_972;
wire n_997;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_359;
wire n_1189;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_930;
wire n_994;
wire n_410;
wire n_774;
wire n_1207;
wire n_377;
wire n_510;
wire n_1075;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1164;
wire n_281;
wire n_487;
wire n_451;
wire n_748;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_483;
wire n_280;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_925;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_958;
wire n_468;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_275;
wire n_1048;
wire n_973;
wire n_587;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_796;
wire n_1216;
wire n_927;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_586;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_293;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_294;
wire n_459;
wire n_907;
wire n_310;
wire n_1062;
wire n_708;
wire n_307;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_519;
wire n_329;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_308;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_557;
wire n_842;
wire n_439;
wire n_614;
wire n_1107;
wire n_446;
wire n_423;
wire n_342;
wire n_799;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_273;
wire n_970;
wire n_984;
wire n_720;
wire n_806;
wire n_1157;
wire n_539;
wire n_1153;
wire n_317;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_721;
wire n_1060;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_306;
wire n_1007;
wire n_1117;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_867;
wire n_1070;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_323;
wire n_347;
wire n_515;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_713;
wire n_457;
wire n_736;
wire n_287;
wire n_606;
wire n_332;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_885;
wire n_284;
wire n_278;
wire n_500;
wire n_607;
wire n_496;
wire n_801;
wire n_1059;
wire n_309;
wire n_701;
wire n_612;
wire n_1032;
wire n_336;
wire n_464;
wire n_1196;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_532;
wire n_400;
wire n_386;
wire n_432;
wire n_659;
wire n_316;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_330;
wire n_1087;
wire n_662;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_301;
wire n_609;
wire n_909;
wire n_366;
wire n_596;
wire n_1215;
wire n_286;
wire n_951;
wire n_321;
wire n_1024;
wire n_1016;
wire n_652;
wire n_333;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_764;
wire n_426;
wire n_282;
wire n_969;
wire n_417;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_381;
wire n_313;
wire n_322;
wire n_427;
wire n_703;
wire n_415;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_729;
wire n_805;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_788;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_285;
wire n_420;
wire n_1089;
wire n_1058;
wire n_388;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_416;
wire n_536;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_615;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_835;
wire n_778;
wire n_1156;
wire n_300;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1043;
wire n_346;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_341;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_473;
wire n_991;
wire n_843;
wire n_538;
wire n_492;
wire n_1150;
wire n_368;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_290;
wire n_385;
wire n_1127;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_998;
wire n_604;
wire n_755;
wire n_848;
wire n_1031;
wire n_292;
wire n_1158;
wire n_328;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1224;
wire n_288;
wire n_383;
wire n_762;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_296;
wire n_765;
wire n_1177;
wire n_462;
wire n_783;
wire n_1074;
wire n_463;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_628;
wire n_812;
wire n_777;
wire n_351;
wire n_401;
wire n_360;
wire n_345;
wire n_481;
wire n_443;
wire n_694;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_279;
wire n_303;
wire n_326;
wire n_289;
wire n_1081;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_455;
wire n_529;
wire n_1025;
wire n_1132;
wire n_630;
wire n_1180;
wire n_647;
wire n_844;
wire n_1160;
wire n_274;
wire n_1195;
wire n_895;
wire n_798;
wire n_318;
wire n_887;
wire n_471;
wire n_1014;
wire n_665;
wire n_1154;
wire n_863;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_910;
wire n_935;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1113;
wire n_760;
wire n_941;
wire n_302;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_601;
wire n_1176;
wire n_649;
wire n_526;
wire n_276;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_374;
wire n_718;
wire n_1114;
wire n_948;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_639;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_398;
wire n_445;
wire n_656;
wire n_1230;
wire n_553;
wire n_325;
wire n_349;
wire n_1021;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_924;
wire n_378;
wire n_441;
wire n_335;
wire n_700;
wire n_534;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_297;
wire n_1053;
wire n_1223;
wire n_967;
wire n_291;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_929;
wire n_1111;
wire n_976;
wire n_695;
wire n_1104;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_405;
wire n_491;
INVx1_ASAP7_75t_L g273 ( .A(n_200), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_88), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_161), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_69), .Y(n_276) );
CKINVDCx16_ASAP7_75t_R g277 ( .A(n_191), .Y(n_277) );
CKINVDCx5p33_ASAP7_75t_R g278 ( .A(n_74), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_218), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_177), .Y(n_280) );
CKINVDCx16_ASAP7_75t_R g281 ( .A(n_166), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_121), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_107), .Y(n_283) );
INVxp33_ASAP7_75t_L g284 ( .A(n_108), .Y(n_284) );
BUFx6f_ASAP7_75t_L g285 ( .A(n_246), .Y(n_285) );
BUFx3_ASAP7_75t_L g286 ( .A(n_257), .Y(n_286) );
CKINVDCx14_ASAP7_75t_R g287 ( .A(n_226), .Y(n_287) );
CKINVDCx20_ASAP7_75t_R g288 ( .A(n_221), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_21), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_174), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_37), .Y(n_291) );
CKINVDCx14_ASAP7_75t_R g292 ( .A(n_37), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_262), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_64), .Y(n_294) );
CKINVDCx20_ASAP7_75t_R g295 ( .A(n_230), .Y(n_295) );
CKINVDCx5p33_ASAP7_75t_R g296 ( .A(n_133), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_10), .Y(n_297) );
INVxp67_ASAP7_75t_SL g298 ( .A(n_222), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_170), .Y(n_299) );
CKINVDCx5p33_ASAP7_75t_R g300 ( .A(n_81), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_217), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_271), .Y(n_302) );
BUFx5_ASAP7_75t_L g303 ( .A(n_231), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_189), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_160), .Y(n_305) );
CKINVDCx5p33_ASAP7_75t_R g306 ( .A(n_233), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_5), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_56), .Y(n_308) );
NOR2xp67_ASAP7_75t_L g309 ( .A(n_77), .B(n_53), .Y(n_309) );
INVxp33_ASAP7_75t_SL g310 ( .A(n_114), .Y(n_310) );
CKINVDCx16_ASAP7_75t_R g311 ( .A(n_250), .Y(n_311) );
HB1xp67_ASAP7_75t_L g312 ( .A(n_5), .Y(n_312) );
CKINVDCx20_ASAP7_75t_R g313 ( .A(n_153), .Y(n_313) );
CKINVDCx5p33_ASAP7_75t_R g314 ( .A(n_40), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_136), .Y(n_315) );
CKINVDCx5p33_ASAP7_75t_R g316 ( .A(n_103), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_234), .B(n_42), .Y(n_317) );
CKINVDCx5p33_ASAP7_75t_R g318 ( .A(n_268), .Y(n_318) );
INVxp33_ASAP7_75t_L g319 ( .A(n_20), .Y(n_319) );
BUFx6f_ASAP7_75t_L g320 ( .A(n_206), .Y(n_320) );
CKINVDCx16_ASAP7_75t_R g321 ( .A(n_165), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_141), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_40), .Y(n_323) );
BUFx3_ASAP7_75t_L g324 ( .A(n_15), .Y(n_324) );
HB1xp67_ASAP7_75t_L g325 ( .A(n_96), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_16), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_70), .Y(n_327) );
CKINVDCx16_ASAP7_75t_R g328 ( .A(n_245), .Y(n_328) );
INVxp67_ASAP7_75t_SL g329 ( .A(n_50), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_169), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_131), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_86), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_97), .Y(n_333) );
CKINVDCx5p33_ASAP7_75t_R g334 ( .A(n_29), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_4), .Y(n_335) );
CKINVDCx5p33_ASAP7_75t_R g336 ( .A(n_185), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_269), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_54), .Y(n_338) );
CKINVDCx20_ASAP7_75t_R g339 ( .A(n_220), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_242), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_83), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_25), .Y(n_342) );
CKINVDCx5p33_ASAP7_75t_R g343 ( .A(n_101), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_80), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_123), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_60), .Y(n_346) );
HB1xp67_ASAP7_75t_L g347 ( .A(n_194), .Y(n_347) );
BUFx6f_ASAP7_75t_L g348 ( .A(n_142), .Y(n_348) );
INVxp67_ASAP7_75t_L g349 ( .A(n_182), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_248), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_175), .Y(n_351) );
CKINVDCx16_ASAP7_75t_R g352 ( .A(n_127), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_227), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_84), .Y(n_354) );
CKINVDCx5p33_ASAP7_75t_R g355 ( .A(n_90), .Y(n_355) );
CKINVDCx20_ASAP7_75t_R g356 ( .A(n_149), .Y(n_356) );
INVxp33_ASAP7_75t_SL g357 ( .A(n_85), .Y(n_357) );
INVxp67_ASAP7_75t_SL g358 ( .A(n_239), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_3), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_48), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_7), .Y(n_361) );
CKINVDCx20_ASAP7_75t_R g362 ( .A(n_18), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_159), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_148), .Y(n_364) );
CKINVDCx5p33_ASAP7_75t_R g365 ( .A(n_168), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_58), .Y(n_366) );
CKINVDCx5p33_ASAP7_75t_R g367 ( .A(n_176), .Y(n_367) );
CKINVDCx20_ASAP7_75t_R g368 ( .A(n_25), .Y(n_368) );
CKINVDCx5p33_ASAP7_75t_R g369 ( .A(n_162), .Y(n_369) );
CKINVDCx14_ASAP7_75t_R g370 ( .A(n_249), .Y(n_370) );
CKINVDCx5p33_ASAP7_75t_R g371 ( .A(n_260), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_240), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_155), .Y(n_373) );
NOR2xp33_ASAP7_75t_L g374 ( .A(n_78), .B(n_135), .Y(n_374) );
CKINVDCx5p33_ASAP7_75t_R g375 ( .A(n_71), .Y(n_375) );
CKINVDCx20_ASAP7_75t_R g376 ( .A(n_109), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_43), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_60), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_50), .Y(n_379) );
NOR2xp67_ASAP7_75t_L g380 ( .A(n_54), .B(n_6), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_164), .Y(n_381) );
CKINVDCx20_ASAP7_75t_R g382 ( .A(n_229), .Y(n_382) );
INVx1_ASAP7_75t_SL g383 ( .A(n_263), .Y(n_383) );
INVx2_ASAP7_75t_SL g384 ( .A(n_144), .Y(n_384) );
CKINVDCx5p33_ASAP7_75t_R g385 ( .A(n_36), .Y(n_385) );
CKINVDCx14_ASAP7_75t_R g386 ( .A(n_104), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_87), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_205), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_172), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_244), .Y(n_390) );
CKINVDCx5p33_ASAP7_75t_R g391 ( .A(n_251), .Y(n_391) );
CKINVDCx5p33_ASAP7_75t_R g392 ( .A(n_184), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_261), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_255), .Y(n_394) );
CKINVDCx20_ASAP7_75t_R g395 ( .A(n_66), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_186), .Y(n_396) );
INVxp33_ASAP7_75t_SL g397 ( .A(n_15), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_111), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_12), .Y(n_399) );
CKINVDCx5p33_ASAP7_75t_R g400 ( .A(n_181), .Y(n_400) );
INVx3_ASAP7_75t_L g401 ( .A(n_93), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_115), .Y(n_402) );
INVxp67_ASAP7_75t_SL g403 ( .A(n_118), .Y(n_403) );
INVxp33_ASAP7_75t_SL g404 ( .A(n_211), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_30), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_132), .Y(n_406) );
CKINVDCx5p33_ASAP7_75t_R g407 ( .A(n_82), .Y(n_407) );
CKINVDCx20_ASAP7_75t_R g408 ( .A(n_152), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_151), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_34), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_134), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_171), .Y(n_412) );
CKINVDCx5p33_ASAP7_75t_R g413 ( .A(n_46), .Y(n_413) );
INVxp67_ASAP7_75t_L g414 ( .A(n_0), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_187), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_335), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_335), .Y(n_417) );
AND2x4_ASAP7_75t_L g418 ( .A(n_401), .B(n_0), .Y(n_418) );
AND2x4_ASAP7_75t_L g419 ( .A(n_401), .B(n_1), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_319), .B(n_1), .Y(n_420) );
AND3x2_ASAP7_75t_L g421 ( .A(n_325), .B(n_2), .C(n_3), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_360), .Y(n_422) );
INVx3_ASAP7_75t_L g423 ( .A(n_324), .Y(n_423) );
CKINVDCx5p33_ASAP7_75t_R g424 ( .A(n_277), .Y(n_424) );
INVx6_ASAP7_75t_L g425 ( .A(n_303), .Y(n_425) );
INVx3_ASAP7_75t_L g426 ( .A(n_324), .Y(n_426) );
HB1xp67_ASAP7_75t_L g427 ( .A(n_292), .Y(n_427) );
INVxp67_ASAP7_75t_L g428 ( .A(n_347), .Y(n_428) );
AND2x4_ASAP7_75t_L g429 ( .A(n_360), .B(n_2), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_366), .Y(n_430) );
BUFx3_ASAP7_75t_L g431 ( .A(n_286), .Y(n_431) );
BUFx6f_ASAP7_75t_L g432 ( .A(n_285), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_366), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_273), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_274), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_275), .Y(n_436) );
CKINVDCx5p33_ASAP7_75t_R g437 ( .A(n_281), .Y(n_437) );
INVx3_ASAP7_75t_L g438 ( .A(n_282), .Y(n_438) );
CKINVDCx5p33_ASAP7_75t_R g439 ( .A(n_311), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_319), .B(n_4), .Y(n_440) );
CKINVDCx20_ASAP7_75t_R g441 ( .A(n_292), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_276), .Y(n_442) );
OR2x6_ASAP7_75t_L g443 ( .A(n_309), .B(n_72), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_279), .Y(n_444) );
BUFx6f_ASAP7_75t_L g445 ( .A(n_285), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_284), .B(n_6), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_280), .Y(n_447) );
INVx3_ASAP7_75t_L g448 ( .A(n_282), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_384), .B(n_7), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_429), .Y(n_450) );
INVx3_ASAP7_75t_L g451 ( .A(n_419), .Y(n_451) );
INVx4_ASAP7_75t_SL g452 ( .A(n_425), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_428), .B(n_284), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_428), .B(n_321), .Y(n_454) );
INVx3_ASAP7_75t_L g455 ( .A(n_419), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_429), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_418), .Y(n_457) );
NAND2xp5_ASAP7_75t_SL g458 ( .A(n_427), .B(n_328), .Y(n_458) );
AO22x2_ASAP7_75t_L g459 ( .A1(n_418), .A2(n_329), .B1(n_289), .B2(n_294), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_418), .Y(n_460) );
INVx2_ASAP7_75t_SL g461 ( .A(n_425), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_427), .B(n_352), .Y(n_462) );
NAND2xp5_ASAP7_75t_SL g463 ( .A(n_419), .B(n_349), .Y(n_463) );
BUFx6f_ASAP7_75t_L g464 ( .A(n_432), .Y(n_464) );
BUFx10_ASAP7_75t_L g465 ( .A(n_418), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_446), .B(n_287), .Y(n_466) );
NAND2xp5_ASAP7_75t_SL g467 ( .A(n_419), .B(n_310), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_425), .Y(n_468) );
NOR2xp33_ASAP7_75t_L g469 ( .A(n_434), .B(n_310), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_429), .Y(n_470) );
BUFx10_ASAP7_75t_L g471 ( .A(n_418), .Y(n_471) );
NAND2x1p5_ASAP7_75t_L g472 ( .A(n_429), .B(n_283), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_425), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_429), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_446), .B(n_287), .Y(n_475) );
INVx1_ASAP7_75t_SL g476 ( .A(n_441), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_446), .B(n_420), .Y(n_477) );
NOR2xp33_ASAP7_75t_R g478 ( .A(n_424), .B(n_370), .Y(n_478) );
BUFx6f_ASAP7_75t_L g479 ( .A(n_432), .Y(n_479) );
BUFx10_ASAP7_75t_L g480 ( .A(n_437), .Y(n_480) );
BUFx4f_ASAP7_75t_L g481 ( .A(n_443), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_434), .B(n_370), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_435), .B(n_386), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_435), .B(n_386), .Y(n_484) );
BUFx10_ASAP7_75t_L g485 ( .A(n_439), .Y(n_485) );
CKINVDCx5p33_ASAP7_75t_R g486 ( .A(n_420), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_420), .B(n_312), .Y(n_487) );
BUFx4_ASAP7_75t_L g488 ( .A(n_440), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_436), .B(n_314), .Y(n_489) );
NOR2xp33_ASAP7_75t_L g490 ( .A(n_436), .B(n_357), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_440), .Y(n_491) );
BUFx3_ASAP7_75t_L g492 ( .A(n_431), .Y(n_492) );
INVx1_ASAP7_75t_SL g493 ( .A(n_449), .Y(n_493) );
INVx4_ASAP7_75t_SL g494 ( .A(n_425), .Y(n_494) );
INVxp67_ASAP7_75t_L g495 ( .A(n_449), .Y(n_495) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_442), .B(n_357), .Y(n_496) );
INVx1_ASAP7_75t_SL g497 ( .A(n_493), .Y(n_497) );
CKINVDCx20_ASAP7_75t_R g498 ( .A(n_478), .Y(n_498) );
CKINVDCx5p33_ASAP7_75t_R g499 ( .A(n_480), .Y(n_499) );
BUFx6f_ASAP7_75t_L g500 ( .A(n_465), .Y(n_500) );
OR2x6_ASAP7_75t_L g501 ( .A(n_459), .B(n_443), .Y(n_501) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_481), .B(n_442), .Y(n_502) );
AOI22xp5_ASAP7_75t_SL g503 ( .A1(n_486), .A2(n_368), .B1(n_395), .B2(n_362), .Y(n_503) );
INVx3_ASAP7_75t_L g504 ( .A(n_465), .Y(n_504) );
INVx8_ASAP7_75t_L g505 ( .A(n_475), .Y(n_505) );
INVx5_ASAP7_75t_L g506 ( .A(n_465), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_477), .Y(n_507) );
BUFx2_ASAP7_75t_L g508 ( .A(n_486), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_495), .B(n_444), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_477), .Y(n_510) );
BUFx6f_ASAP7_75t_L g511 ( .A(n_471), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_491), .B(n_444), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_475), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_453), .B(n_447), .Y(n_514) );
AOI22xp5_ASAP7_75t_L g515 ( .A1(n_459), .A2(n_397), .B1(n_443), .B2(n_288), .Y(n_515) );
NAND2xp5_ASAP7_75t_SL g516 ( .A(n_481), .B(n_471), .Y(n_516) );
AOI22xp5_ASAP7_75t_L g517 ( .A1(n_459), .A2(n_397), .B1(n_443), .B2(n_288), .Y(n_517) );
INVx2_ASAP7_75t_SL g518 ( .A(n_488), .Y(n_518) );
INVx2_ASAP7_75t_SL g519 ( .A(n_488), .Y(n_519) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_457), .A2(n_443), .B(n_447), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_492), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_496), .B(n_431), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_469), .B(n_423), .Y(n_523) );
NOR3xp33_ASAP7_75t_SL g524 ( .A(n_458), .B(n_385), .C(n_334), .Y(n_524) );
AND2x4_ASAP7_75t_L g525 ( .A(n_487), .B(n_443), .Y(n_525) );
NAND2xp5_ASAP7_75t_SL g526 ( .A(n_481), .B(n_293), .Y(n_526) );
O2A1O1Ixp33_ASAP7_75t_L g527 ( .A1(n_450), .A2(n_417), .B(n_422), .C(n_416), .Y(n_527) );
BUFx2_ASAP7_75t_L g528 ( .A(n_459), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_492), .Y(n_529) );
HB1xp67_ASAP7_75t_L g530 ( .A(n_472), .Y(n_530) );
CKINVDCx20_ASAP7_75t_R g531 ( .A(n_480), .Y(n_531) );
INVx3_ASAP7_75t_L g532 ( .A(n_471), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_472), .Y(n_533) );
INVx2_ASAP7_75t_SL g534 ( .A(n_487), .Y(n_534) );
NOR3xp33_ASAP7_75t_SL g535 ( .A(n_467), .B(n_413), .C(n_296), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_472), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_490), .B(n_423), .Y(n_537) );
NOR2xp33_ASAP7_75t_SL g538 ( .A(n_480), .B(n_295), .Y(n_538) );
INVx2_ASAP7_75t_L g539 ( .A(n_451), .Y(n_539) );
NAND2xp5_ASAP7_75t_SL g540 ( .A(n_457), .B(n_299), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_466), .B(n_423), .Y(n_541) );
INVx5_ASAP7_75t_L g542 ( .A(n_451), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_482), .B(n_423), .Y(n_543) );
HB1xp67_ASAP7_75t_L g544 ( .A(n_460), .Y(n_544) );
NOR2xp33_ASAP7_75t_L g545 ( .A(n_463), .B(n_404), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_454), .B(n_414), .Y(n_546) );
AND2x4_ASAP7_75t_L g547 ( .A(n_489), .B(n_421), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_483), .B(n_426), .Y(n_548) );
AND2x4_ASAP7_75t_L g549 ( .A(n_456), .B(n_421), .Y(n_549) );
HB1xp67_ASAP7_75t_L g550 ( .A(n_460), .Y(n_550) );
OR2x6_ASAP7_75t_L g551 ( .A(n_462), .B(n_380), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_485), .B(n_426), .Y(n_552) );
INVx2_ASAP7_75t_L g553 ( .A(n_451), .Y(n_553) );
INVx2_ASAP7_75t_L g554 ( .A(n_455), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_470), .Y(n_555) );
AOI22xp5_ASAP7_75t_L g556 ( .A1(n_474), .A2(n_313), .B1(n_339), .B2(n_295), .Y(n_556) );
INVx2_ASAP7_75t_L g557 ( .A(n_455), .Y(n_557) );
AOI21xp5_ASAP7_75t_L g558 ( .A1(n_455), .A2(n_426), .B(n_301), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_484), .Y(n_559) );
INVxp67_ASAP7_75t_L g560 ( .A(n_485), .Y(n_560) );
AOI22xp5_ASAP7_75t_L g561 ( .A1(n_485), .A2(n_339), .B1(n_356), .B2(n_313), .Y(n_561) );
CKINVDCx5p33_ASAP7_75t_R g562 ( .A(n_476), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_452), .B(n_426), .Y(n_563) );
NOR2xp33_ASAP7_75t_L g564 ( .A(n_473), .B(n_404), .Y(n_564) );
CKINVDCx5p33_ASAP7_75t_R g565 ( .A(n_452), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_473), .Y(n_566) );
INVx2_ASAP7_75t_L g567 ( .A(n_468), .Y(n_567) );
CKINVDCx11_ASAP7_75t_R g568 ( .A(n_452), .Y(n_568) );
HB1xp67_ASAP7_75t_L g569 ( .A(n_494), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_468), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_494), .B(n_438), .Y(n_571) );
NAND2xp5_ASAP7_75t_SL g572 ( .A(n_494), .B(n_302), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_494), .B(n_438), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_461), .B(n_438), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_461), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_464), .B(n_448), .Y(n_576) );
BUFx3_ASAP7_75t_L g577 ( .A(n_464), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_464), .B(n_448), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_464), .Y(n_579) );
INVx2_ASAP7_75t_L g580 ( .A(n_464), .Y(n_580) );
NOR2xp67_ASAP7_75t_L g581 ( .A(n_479), .B(n_448), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_479), .B(n_448), .Y(n_582) );
NOR2xp33_ASAP7_75t_R g583 ( .A(n_479), .B(n_356), .Y(n_583) );
NOR2xp33_ASAP7_75t_L g584 ( .A(n_495), .B(n_417), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_477), .Y(n_585) );
AOI22xp5_ASAP7_75t_L g586 ( .A1(n_501), .A2(n_382), .B1(n_408), .B2(n_376), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_497), .B(n_362), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_509), .B(n_291), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_584), .B(n_297), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_584), .B(n_307), .Y(n_590) );
CKINVDCx5p33_ASAP7_75t_R g591 ( .A(n_531), .Y(n_591) );
OAI21xp5_ASAP7_75t_L g592 ( .A1(n_520), .A2(n_317), .B(n_305), .Y(n_592) );
AND2x4_ASAP7_75t_L g593 ( .A(n_560), .B(n_376), .Y(n_593) );
BUFx6f_ASAP7_75t_L g594 ( .A(n_506), .Y(n_594) );
INVx4_ASAP7_75t_L g595 ( .A(n_506), .Y(n_595) );
AOI21xp33_ASAP7_75t_L g596 ( .A1(n_501), .A2(n_408), .B(n_382), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_507), .Y(n_597) );
OAI21xp33_ASAP7_75t_L g598 ( .A1(n_512), .A2(n_323), .B(n_308), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_510), .Y(n_599) );
BUFx4f_ASAP7_75t_L g600 ( .A(n_501), .Y(n_600) );
CKINVDCx5p33_ASAP7_75t_R g601 ( .A(n_499), .Y(n_601) );
AND2x2_ASAP7_75t_SL g602 ( .A(n_538), .B(n_368), .Y(n_602) );
NOR2xp33_ASAP7_75t_L g603 ( .A(n_534), .B(n_395), .Y(n_603) );
OR2x6_ASAP7_75t_L g604 ( .A(n_518), .B(n_326), .Y(n_604) );
A2O1A1Ixp33_ASAP7_75t_L g605 ( .A1(n_559), .A2(n_342), .B(n_346), .C(n_338), .Y(n_605) );
INVx2_ASAP7_75t_L g606 ( .A(n_539), .Y(n_606) );
INVx2_ASAP7_75t_L g607 ( .A(n_553), .Y(n_607) );
BUFx12f_ASAP7_75t_L g608 ( .A(n_562), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_585), .Y(n_609) );
BUFx4f_ASAP7_75t_L g610 ( .A(n_519), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_513), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_530), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_514), .B(n_359), .Y(n_613) );
OAI21xp5_ASAP7_75t_L g614 ( .A1(n_558), .A2(n_315), .B(n_304), .Y(n_614) );
O2A1O1Ixp33_ASAP7_75t_L g615 ( .A1(n_527), .A2(n_377), .B(n_378), .C(n_361), .Y(n_615) );
BUFx3_ASAP7_75t_L g616 ( .A(n_498), .Y(n_616) );
CKINVDCx5p33_ASAP7_75t_R g617 ( .A(n_503), .Y(n_617) );
CKINVDCx20_ASAP7_75t_R g618 ( .A(n_560), .Y(n_618) );
OAI22xp5_ASAP7_75t_L g619 ( .A1(n_530), .A2(n_399), .B1(n_405), .B2(n_379), .Y(n_619) );
AOI22xp5_ASAP7_75t_L g620 ( .A1(n_525), .A2(n_358), .B1(n_403), .B2(n_298), .Y(n_620) );
NOR2xp33_ASAP7_75t_L g621 ( .A(n_505), .B(n_410), .Y(n_621) );
O2A1O1Ixp33_ASAP7_75t_L g622 ( .A1(n_527), .A2(n_430), .B(n_433), .C(n_422), .Y(n_622) );
AND2x4_ASAP7_75t_L g623 ( .A(n_525), .B(n_430), .Y(n_623) );
AOI21x1_ASAP7_75t_L g624 ( .A1(n_502), .A2(n_327), .B(n_322), .Y(n_624) );
INVx2_ASAP7_75t_L g625 ( .A(n_554), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_505), .B(n_433), .Y(n_626) );
OA22x2_ASAP7_75t_L g627 ( .A1(n_561), .A2(n_331), .B1(n_332), .B2(n_330), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_555), .Y(n_628) );
AND2x4_ASAP7_75t_L g629 ( .A(n_547), .B(n_333), .Y(n_629) );
AOI21xp5_ASAP7_75t_L g630 ( .A1(n_526), .A2(n_340), .B(n_337), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_557), .Y(n_631) );
INVx2_ASAP7_75t_SL g632 ( .A(n_552), .Y(n_632) );
INVx4_ASAP7_75t_L g633 ( .A(n_506), .Y(n_633) );
CKINVDCx16_ASAP7_75t_R g634 ( .A(n_583), .Y(n_634) );
AOI21xp33_ASAP7_75t_L g635 ( .A1(n_545), .A2(n_383), .B(n_300), .Y(n_635) );
BUFx6f_ASAP7_75t_L g636 ( .A(n_506), .Y(n_636) );
AO22x1_ASAP7_75t_L g637 ( .A1(n_528), .A2(n_306), .B1(n_316), .B2(n_278), .Y(n_637) );
INVx5_ASAP7_75t_L g638 ( .A(n_500), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_544), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_544), .Y(n_640) );
BUFx2_ASAP7_75t_L g641 ( .A(n_583), .Y(n_641) );
AND2x4_ASAP7_75t_SL g642 ( .A(n_556), .B(n_341), .Y(n_642) );
OAI22xp5_ASAP7_75t_L g643 ( .A1(n_515), .A2(n_345), .B1(n_353), .B2(n_344), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_550), .Y(n_644) );
AOI21xp5_ASAP7_75t_L g645 ( .A1(n_526), .A2(n_363), .B(n_354), .Y(n_645) );
BUFx6f_ASAP7_75t_L g646 ( .A(n_500), .Y(n_646) );
BUFx2_ASAP7_75t_L g647 ( .A(n_533), .Y(n_647) );
INVx5_ASAP7_75t_L g648 ( .A(n_500), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_550), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g650 ( .A1(n_505), .A2(n_373), .B1(n_381), .B2(n_372), .Y(n_650) );
O2A1O1Ixp33_ASAP7_75t_SL g651 ( .A1(n_541), .A2(n_388), .B(n_389), .C(n_387), .Y(n_651) );
OA22x2_ASAP7_75t_L g652 ( .A1(n_517), .A2(n_393), .B1(n_394), .B2(n_390), .Y(n_652) );
INVx2_ASAP7_75t_L g653 ( .A(n_542), .Y(n_653) );
A2O1A1Ixp33_ASAP7_75t_L g654 ( .A1(n_564), .A2(n_545), .B(n_548), .C(n_543), .Y(n_654) );
OR2x6_ASAP7_75t_L g655 ( .A(n_536), .B(n_396), .Y(n_655) );
BUFx12f_ASAP7_75t_L g656 ( .A(n_568), .Y(n_656) );
INVxp67_ASAP7_75t_L g657 ( .A(n_549), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_574), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_546), .B(n_318), .Y(n_659) );
BUFx2_ASAP7_75t_L g660 ( .A(n_549), .Y(n_660) );
INVx1_ASAP7_75t_SL g661 ( .A(n_500), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_542), .Y(n_662) );
HB1xp67_ASAP7_75t_L g663 ( .A(n_542), .Y(n_663) );
INVx2_ASAP7_75t_L g664 ( .A(n_567), .Y(n_664) );
INVx2_ASAP7_75t_SL g665 ( .A(n_547), .Y(n_665) );
O2A1O1Ixp33_ASAP7_75t_L g666 ( .A1(n_540), .A2(n_402), .B(n_406), .C(n_398), .Y(n_666) );
INVx4_ASAP7_75t_L g667 ( .A(n_511), .Y(n_667) );
AND2x4_ASAP7_75t_L g668 ( .A(n_516), .B(n_409), .Y(n_668) );
HB1xp67_ASAP7_75t_L g669 ( .A(n_511), .Y(n_669) );
NOR2xp33_ASAP7_75t_L g670 ( .A(n_551), .B(n_336), .Y(n_670) );
BUFx2_ASAP7_75t_L g671 ( .A(n_511), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_504), .B(n_343), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_523), .Y(n_673) );
AOI21xp33_ASAP7_75t_L g674 ( .A1(n_516), .A2(n_365), .B(n_355), .Y(n_674) );
BUFx6f_ASAP7_75t_L g675 ( .A(n_511), .Y(n_675) );
AND2x2_ASAP7_75t_L g676 ( .A(n_551), .B(n_8), .Y(n_676) );
AOI21xp5_ASAP7_75t_L g677 ( .A1(n_540), .A2(n_412), .B(n_411), .Y(n_677) );
OAI22xp5_ASAP7_75t_L g678 ( .A1(n_537), .A2(n_415), .B1(n_375), .B2(n_367), .Y(n_678) );
BUFx3_ASAP7_75t_L g679 ( .A(n_566), .Y(n_679) );
INVx3_ASAP7_75t_L g680 ( .A(n_504), .Y(n_680) );
O2A1O1Ixp33_ASAP7_75t_L g681 ( .A1(n_522), .A2(n_350), .B(n_290), .C(n_364), .Y(n_681) );
INVx2_ASAP7_75t_L g682 ( .A(n_521), .Y(n_682) );
INVx2_ASAP7_75t_SL g683 ( .A(n_551), .Y(n_683) );
NOR2xp33_ASAP7_75t_L g684 ( .A(n_564), .B(n_369), .Y(n_684) );
AND3x1_ASAP7_75t_SL g685 ( .A(n_524), .B(n_8), .C(n_9), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_570), .Y(n_686) );
INVx2_ASAP7_75t_L g687 ( .A(n_529), .Y(n_687) );
NOR2x1_ASAP7_75t_L g688 ( .A(n_532), .B(n_286), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_575), .Y(n_689) );
NOR2xp33_ASAP7_75t_L g690 ( .A(n_532), .B(n_371), .Y(n_690) );
HB1xp67_ASAP7_75t_L g691 ( .A(n_571), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_573), .Y(n_692) );
INVx3_ASAP7_75t_L g693 ( .A(n_565), .Y(n_693) );
A2O1A1Ixp33_ASAP7_75t_L g694 ( .A1(n_535), .A2(n_524), .B(n_578), .C(n_576), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_582), .Y(n_695) );
AOI21xp5_ASAP7_75t_L g696 ( .A1(n_563), .A2(n_301), .B(n_290), .Y(n_696) );
HB1xp67_ASAP7_75t_L g697 ( .A(n_569), .Y(n_697) );
AO21x2_ASAP7_75t_L g698 ( .A1(n_581), .A2(n_351), .B(n_350), .Y(n_698) );
AND2x2_ASAP7_75t_L g699 ( .A(n_535), .B(n_10), .Y(n_699) );
AOI21xp5_ASAP7_75t_L g700 ( .A1(n_572), .A2(n_374), .B(n_391), .Y(n_700) );
AOI22xp5_ASAP7_75t_L g701 ( .A1(n_577), .A2(n_303), .B1(n_392), .B2(n_407), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_579), .Y(n_702) );
BUFx8_ASAP7_75t_L g703 ( .A(n_580), .Y(n_703) );
HB1xp67_ASAP7_75t_L g704 ( .A(n_497), .Y(n_704) );
BUFx10_ASAP7_75t_L g705 ( .A(n_499), .Y(n_705) );
AOI22xp5_ASAP7_75t_L g706 ( .A1(n_501), .A2(n_303), .B1(n_400), .B2(n_348), .Y(n_706) );
AOI22xp33_ASAP7_75t_L g707 ( .A1(n_528), .A2(n_303), .B1(n_348), .B2(n_320), .Y(n_707) );
INVx4_ASAP7_75t_L g708 ( .A(n_506), .Y(n_708) );
BUFx6f_ASAP7_75t_L g709 ( .A(n_506), .Y(n_709) );
BUFx6f_ASAP7_75t_L g710 ( .A(n_506), .Y(n_710) );
INVx2_ASAP7_75t_L g711 ( .A(n_539), .Y(n_711) );
BUFx6f_ASAP7_75t_L g712 ( .A(n_506), .Y(n_712) );
INVx2_ASAP7_75t_L g713 ( .A(n_539), .Y(n_713) );
NAND2x1p5_ASAP7_75t_L g714 ( .A(n_600), .B(n_285), .Y(n_714) );
INVx2_ASAP7_75t_L g715 ( .A(n_628), .Y(n_715) );
AND2x4_ASAP7_75t_L g716 ( .A(n_647), .B(n_11), .Y(n_716) );
AOI21xp33_ASAP7_75t_SL g717 ( .A1(n_602), .A2(n_11), .B(n_12), .Y(n_717) );
OA21x2_ASAP7_75t_L g718 ( .A1(n_592), .A2(n_303), .B(n_285), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_639), .B(n_303), .Y(n_719) );
OAI21x1_ASAP7_75t_SL g720 ( .A1(n_595), .A2(n_303), .B(n_13), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_597), .Y(n_721) );
OAI22xp5_ASAP7_75t_L g722 ( .A1(n_600), .A2(n_348), .B1(n_320), .B2(n_445), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_599), .Y(n_723) );
AOI22xp33_ASAP7_75t_L g724 ( .A1(n_652), .A2(n_643), .B1(n_609), .B2(n_623), .Y(n_724) );
CKINVDCx8_ASAP7_75t_R g725 ( .A(n_591), .Y(n_725) );
CKINVDCx20_ASAP7_75t_R g726 ( .A(n_618), .Y(n_726) );
OAI22xp5_ASAP7_75t_L g727 ( .A1(n_586), .A2(n_348), .B1(n_320), .B2(n_445), .Y(n_727) );
A2O1A1Ixp33_ASAP7_75t_L g728 ( .A1(n_654), .A2(n_320), .B(n_445), .C(n_432), .Y(n_728) );
AOI21xp5_ASAP7_75t_L g729 ( .A1(n_614), .A2(n_445), .B(n_432), .Y(n_729) );
AND2x2_ASAP7_75t_L g730 ( .A(n_704), .B(n_13), .Y(n_730) );
OAI21x1_ASAP7_75t_L g731 ( .A1(n_624), .A2(n_445), .B(n_432), .Y(n_731) );
CKINVDCx14_ASAP7_75t_R g732 ( .A(n_608), .Y(n_732) );
INVx4_ASAP7_75t_L g733 ( .A(n_638), .Y(n_733) );
AOI21x1_ASAP7_75t_L g734 ( .A1(n_696), .A2(n_75), .B(n_73), .Y(n_734) );
OAI21x1_ASAP7_75t_L g735 ( .A1(n_688), .A2(n_79), .B(n_76), .Y(n_735) );
AND2x4_ASAP7_75t_L g736 ( .A(n_612), .B(n_14), .Y(n_736) );
AND2x4_ASAP7_75t_L g737 ( .A(n_595), .B(n_14), .Y(n_737) );
OAI21xp5_ASAP7_75t_L g738 ( .A1(n_673), .A2(n_16), .B(n_17), .Y(n_738) );
NAND2xp5_ASAP7_75t_SL g739 ( .A(n_646), .B(n_89), .Y(n_739) );
OAI21x1_ASAP7_75t_L g740 ( .A1(n_702), .A2(n_92), .B(n_91), .Y(n_740) );
INVx2_ASAP7_75t_L g741 ( .A(n_606), .Y(n_741) );
OAI21x1_ASAP7_75t_L g742 ( .A1(n_614), .A2(n_95), .B(n_94), .Y(n_742) );
INVx1_ASAP7_75t_L g743 ( .A(n_611), .Y(n_743) );
OAI22xp33_ASAP7_75t_L g744 ( .A1(n_586), .A2(n_17), .B1(n_18), .B2(n_19), .Y(n_744) );
INVx2_ASAP7_75t_L g745 ( .A(n_607), .Y(n_745) );
INVx2_ASAP7_75t_L g746 ( .A(n_625), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_640), .B(n_19), .Y(n_747) );
O2A1O1Ixp33_ASAP7_75t_SL g748 ( .A1(n_694), .A2(n_145), .B(n_270), .C(n_267), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_644), .B(n_20), .Y(n_749) );
AOI21xp5_ASAP7_75t_L g750 ( .A1(n_681), .A2(n_99), .B(n_98), .Y(n_750) );
AO31x2_ASAP7_75t_L g751 ( .A1(n_643), .A2(n_21), .A3(n_22), .B(n_23), .Y(n_751) );
INVx3_ASAP7_75t_L g752 ( .A(n_633), .Y(n_752) );
INVx1_ASAP7_75t_L g753 ( .A(n_626), .Y(n_753) );
INVxp67_ASAP7_75t_L g754 ( .A(n_604), .Y(n_754) );
OAI21x1_ASAP7_75t_L g755 ( .A1(n_689), .A2(n_102), .B(n_100), .Y(n_755) );
A2O1A1Ixp33_ASAP7_75t_L g756 ( .A1(n_615), .A2(n_24), .B(n_26), .C(n_27), .Y(n_756) );
INVx1_ASAP7_75t_L g757 ( .A(n_623), .Y(n_757) );
AOI22xp5_ASAP7_75t_L g758 ( .A1(n_587), .A2(n_26), .B1(n_27), .B2(n_28), .Y(n_758) );
NOR2xp33_ASAP7_75t_L g759 ( .A(n_657), .B(n_28), .Y(n_759) );
AOI221xp5_ASAP7_75t_L g760 ( .A1(n_589), .A2(n_29), .B1(n_30), .B2(n_31), .C(n_32), .Y(n_760) );
INVx6_ASAP7_75t_L g761 ( .A(n_703), .Y(n_761) );
OAI21x1_ASAP7_75t_L g762 ( .A1(n_686), .A2(n_158), .B(n_266), .Y(n_762) );
AOI22xp33_ASAP7_75t_SL g763 ( .A1(n_593), .A2(n_31), .B1(n_32), .B2(n_33), .Y(n_763) );
HB1xp67_ASAP7_75t_L g764 ( .A(n_638), .Y(n_764) );
A2O1A1Ixp33_ASAP7_75t_L g765 ( .A1(n_598), .A2(n_33), .B(n_34), .C(n_35), .Y(n_765) );
O2A1O1Ixp33_ASAP7_75t_SL g766 ( .A1(n_706), .A2(n_163), .B(n_265), .C(n_264), .Y(n_766) );
OAI21x1_ASAP7_75t_L g767 ( .A1(n_692), .A2(n_157), .B(n_259), .Y(n_767) );
OA21x2_ASAP7_75t_L g768 ( .A1(n_706), .A2(n_156), .B(n_258), .Y(n_768) );
INVx2_ASAP7_75t_L g769 ( .A(n_711), .Y(n_769) );
OAI21x1_ASAP7_75t_L g770 ( .A1(n_630), .A2(n_154), .B(n_256), .Y(n_770) );
INVx1_ASAP7_75t_L g771 ( .A(n_649), .Y(n_771) );
OAI22xp5_ASAP7_75t_L g772 ( .A1(n_655), .A2(n_35), .B1(n_36), .B2(n_38), .Y(n_772) );
OAI21x1_ASAP7_75t_L g773 ( .A1(n_645), .A2(n_167), .B(n_254), .Y(n_773) );
OAI21x1_ASAP7_75t_L g774 ( .A1(n_664), .A2(n_150), .B(n_253), .Y(n_774) );
INVx1_ASAP7_75t_L g775 ( .A(n_622), .Y(n_775) );
INVx2_ASAP7_75t_L g776 ( .A(n_713), .Y(n_776) );
NOR2xp67_ASAP7_75t_L g777 ( .A(n_656), .B(n_38), .Y(n_777) );
BUFx2_ASAP7_75t_L g778 ( .A(n_604), .Y(n_778) );
OAI21x1_ASAP7_75t_L g779 ( .A1(n_680), .A2(n_147), .B(n_252), .Y(n_779) );
O2A1O1Ixp33_ASAP7_75t_L g780 ( .A1(n_605), .A2(n_39), .B(n_41), .C(n_42), .Y(n_780) );
BUFx12f_ASAP7_75t_L g781 ( .A(n_705), .Y(n_781) );
INVx3_ASAP7_75t_L g782 ( .A(n_633), .Y(n_782) );
AO31x2_ASAP7_75t_L g783 ( .A1(n_677), .A2(n_41), .A3(n_43), .B(n_44), .Y(n_783) );
OAI21x1_ASAP7_75t_L g784 ( .A1(n_680), .A2(n_173), .B(n_247), .Y(n_784) );
OR2x2_ASAP7_75t_L g785 ( .A(n_604), .B(n_45), .Y(n_785) );
INVx2_ASAP7_75t_L g786 ( .A(n_631), .Y(n_786) );
OAI21xp5_ASAP7_75t_L g787 ( .A1(n_695), .A2(n_45), .B(n_46), .Y(n_787) );
OAI21xp5_ASAP7_75t_L g788 ( .A1(n_658), .A2(n_47), .B(n_48), .Y(n_788) );
OAI21x1_ASAP7_75t_L g789 ( .A1(n_682), .A2(n_178), .B(n_243), .Y(n_789) );
INVx2_ASAP7_75t_L g790 ( .A(n_687), .Y(n_790) );
OAI21x1_ASAP7_75t_L g791 ( .A1(n_707), .A2(n_146), .B(n_241), .Y(n_791) );
AO21x2_ASAP7_75t_L g792 ( .A1(n_698), .A2(n_143), .B(n_238), .Y(n_792) );
BUFx8_ASAP7_75t_L g793 ( .A(n_616), .Y(n_793) );
INVx2_ASAP7_75t_L g794 ( .A(n_594), .Y(n_794) );
NOR2xp67_ASAP7_75t_L g795 ( .A(n_601), .B(n_47), .Y(n_795) );
OAI21xp5_ASAP7_75t_L g796 ( .A1(n_666), .A2(n_49), .B(n_51), .Y(n_796) );
OAI21x1_ASAP7_75t_L g797 ( .A1(n_700), .A2(n_179), .B(n_237), .Y(n_797) );
OAI21x1_ASAP7_75t_L g798 ( .A1(n_662), .A2(n_140), .B(n_236), .Y(n_798) );
O2A1O1Ixp33_ASAP7_75t_SL g799 ( .A1(n_661), .A2(n_139), .B(n_235), .C(n_232), .Y(n_799) );
INVx2_ASAP7_75t_L g800 ( .A(n_594), .Y(n_800) );
OR2x6_ASAP7_75t_L g801 ( .A(n_655), .B(n_49), .Y(n_801) );
NOR2xp33_ASAP7_75t_L g802 ( .A(n_620), .B(n_51), .Y(n_802) );
A2O1A1Ixp33_ASAP7_75t_L g803 ( .A1(n_590), .A2(n_52), .B(n_53), .C(n_55), .Y(n_803) );
OAI21x1_ASAP7_75t_L g804 ( .A1(n_653), .A2(n_180), .B(n_228), .Y(n_804) );
CKINVDCx20_ASAP7_75t_R g805 ( .A(n_617), .Y(n_805) );
OAI21xp5_ASAP7_75t_L g806 ( .A1(n_620), .A2(n_52), .B(n_55), .Y(n_806) );
OAI21xp5_ASAP7_75t_L g807 ( .A1(n_668), .A2(n_56), .B(n_57), .Y(n_807) );
NAND3xp33_ASAP7_75t_L g808 ( .A(n_684), .B(n_57), .C(n_58), .Y(n_808) );
INVx2_ASAP7_75t_L g809 ( .A(n_594), .Y(n_809) );
INVx1_ASAP7_75t_L g810 ( .A(n_665), .Y(n_810) );
OAI21x1_ASAP7_75t_L g811 ( .A1(n_693), .A2(n_183), .B(n_225), .Y(n_811) );
A2O1A1Ixp33_ASAP7_75t_L g812 ( .A1(n_613), .A2(n_59), .B(n_61), .C(n_62), .Y(n_812) );
BUFx2_ASAP7_75t_L g813 ( .A(n_655), .Y(n_813) );
OA21x2_ASAP7_75t_L g814 ( .A1(n_588), .A2(n_138), .B(n_224), .Y(n_814) );
AOI22xp33_ASAP7_75t_L g815 ( .A1(n_627), .A2(n_59), .B1(n_61), .B2(n_62), .Y(n_815) );
OR2x6_ASAP7_75t_L g816 ( .A(n_660), .B(n_63), .Y(n_816) );
INVx2_ASAP7_75t_L g817 ( .A(n_636), .Y(n_817) );
BUFx2_ASAP7_75t_L g818 ( .A(n_636), .Y(n_818) );
A2O1A1Ixp33_ASAP7_75t_L g819 ( .A1(n_699), .A2(n_63), .B(n_64), .C(n_65), .Y(n_819) );
AO22x2_ASAP7_75t_L g820 ( .A1(n_683), .A2(n_65), .B1(n_66), .B2(n_67), .Y(n_820) );
BUFx2_ASAP7_75t_L g821 ( .A(n_636), .Y(n_821) );
AO31x2_ASAP7_75t_L g822 ( .A1(n_619), .A2(n_67), .A3(n_68), .B(n_105), .Y(n_822) );
OAI21x1_ASAP7_75t_L g823 ( .A1(n_693), .A2(n_195), .B(n_106), .Y(n_823) );
NAND2xp5_ASAP7_75t_L g824 ( .A(n_668), .B(n_68), .Y(n_824) );
INVx1_ASAP7_75t_L g825 ( .A(n_629), .Y(n_825) );
OAI21x1_ASAP7_75t_L g826 ( .A1(n_669), .A2(n_110), .B(n_112), .Y(n_826) );
OAI21x1_ASAP7_75t_L g827 ( .A1(n_701), .A2(n_113), .B(n_116), .Y(n_827) );
BUFx2_ASAP7_75t_L g828 ( .A(n_709), .Y(n_828) );
AO21x2_ASAP7_75t_L g829 ( .A1(n_698), .A2(n_117), .B(n_119), .Y(n_829) );
OAI21xp5_ASAP7_75t_L g830 ( .A1(n_621), .A2(n_120), .B(n_122), .Y(n_830) );
AOI22xp33_ASAP7_75t_L g831 ( .A1(n_629), .A2(n_124), .B1(n_125), .B2(n_126), .Y(n_831) );
OAI21x1_ASAP7_75t_L g832 ( .A1(n_701), .A2(n_128), .B(n_129), .Y(n_832) );
A2O1A1Ixp33_ASAP7_75t_L g833 ( .A1(n_632), .A2(n_130), .B(n_137), .C(n_188), .Y(n_833) );
INVx1_ASAP7_75t_L g834 ( .A(n_679), .Y(n_834) );
INVx1_ASAP7_75t_L g835 ( .A(n_663), .Y(n_835) );
BUFx3_ASAP7_75t_L g836 ( .A(n_610), .Y(n_836) );
NAND2x1p5_ASAP7_75t_L g837 ( .A(n_638), .B(n_272), .Y(n_837) );
OAI22xp33_ASAP7_75t_L g838 ( .A1(n_596), .A2(n_190), .B1(n_192), .B2(n_193), .Y(n_838) );
OAI21xp5_ASAP7_75t_L g839 ( .A1(n_650), .A2(n_196), .B(n_197), .Y(n_839) );
NAND2xp5_ASAP7_75t_L g840 ( .A(n_642), .B(n_198), .Y(n_840) );
INVx1_ASAP7_75t_L g841 ( .A(n_676), .Y(n_841) );
INVx2_ASAP7_75t_L g842 ( .A(n_709), .Y(n_842) );
INVx1_ASAP7_75t_L g843 ( .A(n_651), .Y(n_843) );
INVx1_ASAP7_75t_L g844 ( .A(n_659), .Y(n_844) );
CKINVDCx11_ASAP7_75t_R g845 ( .A(n_725), .Y(n_845) );
AOI22xp33_ASAP7_75t_SL g846 ( .A1(n_778), .A2(n_634), .B1(n_641), .B2(n_603), .Y(n_846) );
OAI211xp5_ASAP7_75t_L g847 ( .A1(n_717), .A2(n_635), .B(n_670), .C(n_674), .Y(n_847) );
OAI22xp5_ASAP7_75t_L g848 ( .A1(n_801), .A2(n_634), .B1(n_661), .B2(n_648), .Y(n_848) );
OR2x2_ASAP7_75t_L g849 ( .A(n_813), .B(n_637), .Y(n_849) );
INVx1_ASAP7_75t_L g850 ( .A(n_771), .Y(n_850) );
AND2x2_ASAP7_75t_L g851 ( .A(n_801), .B(n_648), .Y(n_851) );
AND2x2_ASAP7_75t_L g852 ( .A(n_801), .B(n_648), .Y(n_852) );
AOI21xp5_ASAP7_75t_L g853 ( .A1(n_729), .A2(n_646), .B(n_675), .Y(n_853) );
AOI22xp33_ASAP7_75t_L g854 ( .A1(n_802), .A2(n_678), .B1(n_690), .B2(n_708), .Y(n_854) );
NAND2xp33_ASAP7_75t_L g855 ( .A(n_714), .B(n_712), .Y(n_855) );
OAI21x1_ASAP7_75t_L g856 ( .A1(n_731), .A2(n_691), .B(n_672), .Y(n_856) );
OAI22xp5_ASAP7_75t_L g857 ( .A1(n_727), .A2(n_724), .B1(n_816), .B2(n_807), .Y(n_857) );
INVx1_ASAP7_75t_L g858 ( .A(n_715), .Y(n_858) );
OAI221xp5_ASAP7_75t_L g859 ( .A1(n_724), .A2(n_708), .B1(n_697), .B2(n_671), .C(n_710), .Y(n_859) );
AOI21xp5_ASAP7_75t_L g860 ( .A1(n_729), .A2(n_675), .B(n_646), .Y(n_860) );
AOI22xp33_ASAP7_75t_L g861 ( .A1(n_802), .A2(n_712), .B1(n_710), .B2(n_667), .Y(n_861) );
INVx2_ASAP7_75t_L g862 ( .A(n_721), .Y(n_862) );
AND2x4_ASAP7_75t_L g863 ( .A(n_754), .B(n_710), .Y(n_863) );
INVx1_ASAP7_75t_L g864 ( .A(n_723), .Y(n_864) );
AOI22xp33_ASAP7_75t_SL g865 ( .A1(n_716), .A2(n_712), .B1(n_685), .B2(n_675), .Y(n_865) );
BUFx6f_ASAP7_75t_L g866 ( .A(n_733), .Y(n_866) );
AND2x2_ASAP7_75t_L g867 ( .A(n_754), .B(n_667), .Y(n_867) );
NAND3xp33_ASAP7_75t_L g868 ( .A(n_728), .B(n_199), .C(n_201), .Y(n_868) );
INVx4_ASAP7_75t_L g869 ( .A(n_761), .Y(n_869) );
OAI22xp5_ASAP7_75t_SL g870 ( .A1(n_726), .A2(n_202), .B1(n_203), .B2(n_204), .Y(n_870) );
AOI21xp33_ASAP7_75t_L g871 ( .A1(n_727), .A2(n_207), .B(n_208), .Y(n_871) );
AOI22xp33_ASAP7_75t_L g872 ( .A1(n_844), .A2(n_209), .B1(n_210), .B2(n_212), .Y(n_872) );
INVx2_ASAP7_75t_L g873 ( .A(n_743), .Y(n_873) );
AOI222xp33_ASAP7_75t_L g874 ( .A1(n_744), .A2(n_213), .B1(n_214), .B2(n_215), .C1(n_216), .C2(n_219), .Y(n_874) );
NAND2xp5_ASAP7_75t_L g875 ( .A(n_753), .B(n_223), .Y(n_875) );
AND2x2_ASAP7_75t_L g876 ( .A(n_730), .B(n_736), .Y(n_876) );
OAI21xp33_ASAP7_75t_L g877 ( .A1(n_806), .A2(n_815), .B(n_796), .Y(n_877) );
AND2x4_ASAP7_75t_L g878 ( .A(n_733), .B(n_752), .Y(n_878) );
OAI321xp33_ASAP7_75t_L g879 ( .A1(n_744), .A2(n_772), .A3(n_806), .B1(n_807), .B2(n_838), .C(n_738), .Y(n_879) );
OAI22xp5_ASAP7_75t_L g880 ( .A1(n_816), .A2(n_736), .B1(n_824), .B2(n_815), .Y(n_880) );
OAI22xp5_ASAP7_75t_L g881 ( .A1(n_816), .A2(n_824), .B1(n_714), .B2(n_775), .Y(n_881) );
INVx1_ASAP7_75t_L g882 ( .A(n_747), .Y(n_882) );
INVx1_ASAP7_75t_L g883 ( .A(n_747), .Y(n_883) );
INVxp67_ASAP7_75t_L g884 ( .A(n_785), .Y(n_884) );
INVx2_ASAP7_75t_L g885 ( .A(n_786), .Y(n_885) );
OAI22xp5_ASAP7_75t_L g886 ( .A1(n_772), .A2(n_820), .B1(n_738), .B2(n_765), .Y(n_886) );
NOR2xp33_ASAP7_75t_L g887 ( .A(n_841), .B(n_825), .Y(n_887) );
OAI222xp33_ASAP7_75t_L g888 ( .A1(n_763), .A2(n_758), .B1(n_737), .B2(n_780), .C1(n_838), .C2(n_749), .Y(n_888) );
AND2x2_ASAP7_75t_L g889 ( .A(n_761), .B(n_763), .Y(n_889) );
AO31x2_ASAP7_75t_L g890 ( .A1(n_765), .A2(n_750), .A3(n_833), .B(n_843), .Y(n_890) );
INVx1_ASAP7_75t_L g891 ( .A(n_749), .Y(n_891) );
AOI22xp33_ASAP7_75t_SL g892 ( .A1(n_761), .A2(n_820), .B1(n_737), .B2(n_788), .Y(n_892) );
AND2x2_ASAP7_75t_L g893 ( .A(n_757), .B(n_834), .Y(n_893) );
AOI22xp33_ASAP7_75t_L g894 ( .A1(n_759), .A2(n_760), .B1(n_835), .B2(n_808), .Y(n_894) );
NAND2xp5_ASAP7_75t_L g895 ( .A(n_759), .B(n_810), .Y(n_895) );
OAI22xp5_ASAP7_75t_L g896 ( .A1(n_820), .A2(n_788), .B1(n_787), .B2(n_819), .Y(n_896) );
AOI22xp33_ASAP7_75t_L g897 ( .A1(n_760), .A2(n_840), .B1(n_793), .B2(n_752), .Y(n_897) );
OAI221xp5_ASAP7_75t_L g898 ( .A1(n_756), .A2(n_819), .B1(n_795), .B2(n_780), .C(n_812), .Y(n_898) );
AOI22xp33_ASAP7_75t_L g899 ( .A1(n_840), .A2(n_793), .B1(n_782), .B2(n_764), .Y(n_899) );
AND2x4_ASAP7_75t_L g900 ( .A(n_782), .B(n_836), .Y(n_900) );
OR2x2_ASAP7_75t_L g901 ( .A(n_764), .B(n_818), .Y(n_901) );
AND2x4_ASAP7_75t_L g902 ( .A(n_821), .B(n_828), .Y(n_902) );
OAI21xp33_ASAP7_75t_L g903 ( .A1(n_756), .A2(n_812), .B(n_803), .Y(n_903) );
INVx1_ASAP7_75t_L g904 ( .A(n_741), .Y(n_904) );
NAND3xp33_ASAP7_75t_L g905 ( .A(n_750), .B(n_803), .C(n_839), .Y(n_905) );
INVx4_ASAP7_75t_L g906 ( .A(n_781), .Y(n_906) );
AND2x2_ASAP7_75t_L g907 ( .A(n_745), .B(n_746), .Y(n_907) );
OAI22xp33_ASAP7_75t_L g908 ( .A1(n_805), .A2(n_777), .B1(n_839), .B2(n_830), .Y(n_908) );
OAI21xp5_ASAP7_75t_L g909 ( .A1(n_719), .A2(n_832), .B(n_827), .Y(n_909) );
AND2x2_ASAP7_75t_L g910 ( .A(n_769), .B(n_776), .Y(n_910) );
BUFx2_ASAP7_75t_L g911 ( .A(n_794), .Y(n_911) );
AOI22xp33_ASAP7_75t_L g912 ( .A1(n_790), .A2(n_719), .B1(n_720), .B2(n_830), .Y(n_912) );
AOI21xp33_ASAP7_75t_L g913 ( .A1(n_718), .A2(n_768), .B(n_829), .Y(n_913) );
OA21x2_ASAP7_75t_L g914 ( .A1(n_742), .A2(n_774), .B(n_789), .Y(n_914) );
HB1xp67_ASAP7_75t_L g915 ( .A(n_800), .Y(n_915) );
OAI22xp5_ASAP7_75t_L g916 ( .A1(n_831), .A2(n_837), .B1(n_768), .B2(n_722), .Y(n_916) );
NOR2xp33_ASAP7_75t_SL g917 ( .A(n_837), .B(n_722), .Y(n_917) );
INVx1_ASAP7_75t_L g918 ( .A(n_751), .Y(n_918) );
OAI22xp5_ASAP7_75t_L g919 ( .A1(n_831), .A2(n_833), .B1(n_718), .B2(n_842), .Y(n_919) );
AND2x2_ASAP7_75t_L g920 ( .A(n_751), .B(n_822), .Y(n_920) );
OR2x2_ASAP7_75t_L g921 ( .A(n_809), .B(n_817), .Y(n_921) );
AOI221xp5_ASAP7_75t_L g922 ( .A1(n_766), .A2(n_732), .B1(n_748), .B2(n_799), .C(n_739), .Y(n_922) );
AND2x2_ASAP7_75t_L g923 ( .A(n_751), .B(n_822), .Y(n_923) );
INVx2_ASAP7_75t_SL g924 ( .A(n_822), .Y(n_924) );
INVx1_ASAP7_75t_L g925 ( .A(n_783), .Y(n_925) );
OAI221xp5_ASAP7_75t_L g926 ( .A1(n_766), .A2(n_814), .B1(n_734), .B2(n_799), .C(n_783), .Y(n_926) );
INVx2_ASAP7_75t_L g927 ( .A(n_783), .Y(n_927) );
OAI22xp5_ASAP7_75t_L g928 ( .A1(n_811), .A2(n_823), .B1(n_826), .B2(n_792), .Y(n_928) );
INVx3_ASAP7_75t_L g929 ( .A(n_735), .Y(n_929) );
OAI22xp5_ASAP7_75t_L g930 ( .A1(n_755), .A2(n_767), .B1(n_762), .B2(n_784), .Y(n_930) );
OAI221xp5_ASAP7_75t_SL g931 ( .A1(n_798), .A2(n_740), .B1(n_779), .B2(n_770), .C(n_773), .Y(n_931) );
AOI21xp5_ASAP7_75t_L g932 ( .A1(n_797), .A2(n_804), .B(n_791), .Y(n_932) );
OAI221xp5_ASAP7_75t_L g933 ( .A1(n_724), .A2(n_538), .B1(n_497), .B2(n_508), .C(n_551), .Y(n_933) );
INVx2_ASAP7_75t_SL g934 ( .A(n_761), .Y(n_934) );
AO31x2_ASAP7_75t_L g935 ( .A1(n_728), .A2(n_729), .A3(n_765), .B(n_750), .Y(n_935) );
AOI22xp33_ASAP7_75t_L g936 ( .A1(n_802), .A2(n_602), .B1(n_508), .B2(n_525), .Y(n_936) );
AOI21xp5_ASAP7_75t_L g937 ( .A1(n_729), .A2(n_481), .B(n_654), .Y(n_937) );
INVx2_ASAP7_75t_L g938 ( .A(n_715), .Y(n_938) );
AO31x2_ASAP7_75t_L g939 ( .A1(n_728), .A2(n_729), .A3(n_765), .B(n_750), .Y(n_939) );
AND2x2_ASAP7_75t_L g940 ( .A(n_813), .B(n_497), .Y(n_940) );
INVx3_ASAP7_75t_L g941 ( .A(n_733), .Y(n_941) );
AND2x2_ASAP7_75t_L g942 ( .A(n_813), .B(n_497), .Y(n_942) );
INVx2_ASAP7_75t_L g943 ( .A(n_715), .Y(n_943) );
INVx2_ASAP7_75t_L g944 ( .A(n_715), .Y(n_944) );
AND2x4_ASAP7_75t_L g945 ( .A(n_754), .B(n_647), .Y(n_945) );
INVx1_ASAP7_75t_L g946 ( .A(n_771), .Y(n_946) );
INVx2_ASAP7_75t_SL g947 ( .A(n_761), .Y(n_947) );
AOI221xp5_ASAP7_75t_L g948 ( .A1(n_844), .A2(n_643), .B1(n_534), .B2(n_744), .C(n_585), .Y(n_948) );
OAI221xp5_ASAP7_75t_L g949 ( .A1(n_724), .A2(n_538), .B1(n_497), .B2(n_508), .C(n_551), .Y(n_949) );
A2O1A1Ixp33_ASAP7_75t_L g950 ( .A1(n_806), .A2(n_600), .B(n_654), .C(n_780), .Y(n_950) );
NOR2xp33_ASAP7_75t_L g951 ( .A(n_754), .B(n_561), .Y(n_951) );
INVx3_ASAP7_75t_L g952 ( .A(n_733), .Y(n_952) );
INVx2_ASAP7_75t_L g953 ( .A(n_715), .Y(n_953) );
NAND4xp25_ASAP7_75t_L g954 ( .A(n_802), .B(n_724), .C(n_815), .D(n_760), .Y(n_954) );
INVx1_ASAP7_75t_L g955 ( .A(n_771), .Y(n_955) );
OAI22xp5_ASAP7_75t_L g956 ( .A1(n_801), .A2(n_600), .B1(n_586), .B2(n_727), .Y(n_956) );
INVx1_ASAP7_75t_L g957 ( .A(n_771), .Y(n_957) );
INVx1_ASAP7_75t_L g958 ( .A(n_771), .Y(n_958) );
INVx2_ASAP7_75t_L g959 ( .A(n_715), .Y(n_959) );
INVx2_ASAP7_75t_L g960 ( .A(n_715), .Y(n_960) );
AOI221xp5_ASAP7_75t_L g961 ( .A1(n_844), .A2(n_643), .B1(n_534), .B2(n_744), .C(n_585), .Y(n_961) );
AOI21xp5_ASAP7_75t_L g962 ( .A1(n_729), .A2(n_481), .B(n_654), .Y(n_962) );
AOI22xp33_ASAP7_75t_SL g963 ( .A1(n_778), .A2(n_602), .B1(n_538), .B2(n_503), .Y(n_963) );
NAND2xp5_ASAP7_75t_L g964 ( .A(n_948), .B(n_961), .Y(n_964) );
HB1xp67_ASAP7_75t_L g965 ( .A(n_940), .Y(n_965) );
HB1xp67_ASAP7_75t_L g966 ( .A(n_942), .Y(n_966) );
HB1xp67_ASAP7_75t_L g967 ( .A(n_901), .Y(n_967) );
AOI22xp33_ASAP7_75t_L g968 ( .A1(n_954), .A2(n_956), .B1(n_880), .B2(n_963), .Y(n_968) );
CKINVDCx5p33_ASAP7_75t_R g969 ( .A(n_845), .Y(n_969) );
AND2x2_ASAP7_75t_L g970 ( .A(n_907), .B(n_910), .Y(n_970) );
NAND2xp5_ASAP7_75t_L g971 ( .A(n_936), .B(n_951), .Y(n_971) );
AND2x2_ASAP7_75t_L g972 ( .A(n_938), .B(n_943), .Y(n_972) );
AND2x4_ASAP7_75t_L g973 ( .A(n_929), .B(n_866), .Y(n_973) );
BUFx6f_ASAP7_75t_L g974 ( .A(n_866), .Y(n_974) );
INVx1_ASAP7_75t_L g975 ( .A(n_925), .Y(n_975) );
AOI211xp5_ASAP7_75t_L g976 ( .A1(n_956), .A2(n_908), .B(n_880), .C(n_857), .Y(n_976) );
AND2x2_ASAP7_75t_L g977 ( .A(n_944), .B(n_953), .Y(n_977) );
INVx1_ASAP7_75t_L g978 ( .A(n_918), .Y(n_978) );
OAI31xp33_ASAP7_75t_L g979 ( .A1(n_857), .A2(n_954), .A3(n_881), .B(n_949), .Y(n_979) );
AND2x2_ASAP7_75t_L g980 ( .A(n_959), .B(n_960), .Y(n_980) );
AND2x2_ASAP7_75t_L g981 ( .A(n_885), .B(n_858), .Y(n_981) );
INVx1_ASAP7_75t_L g982 ( .A(n_927), .Y(n_982) );
INVx1_ASAP7_75t_L g983 ( .A(n_920), .Y(n_983) );
NOR2x1_ASAP7_75t_SL g984 ( .A(n_881), .B(n_848), .Y(n_984) );
INVx1_ASAP7_75t_L g985 ( .A(n_923), .Y(n_985) );
HB1xp67_ASAP7_75t_L g986 ( .A(n_945), .Y(n_986) );
INVx2_ASAP7_75t_SL g987 ( .A(n_866), .Y(n_987) );
AND2x2_ASAP7_75t_L g988 ( .A(n_904), .B(n_862), .Y(n_988) );
AND2x2_ASAP7_75t_L g989 ( .A(n_873), .B(n_882), .Y(n_989) );
AND2x4_ASAP7_75t_L g990 ( .A(n_929), .B(n_878), .Y(n_990) );
AND2x2_ASAP7_75t_L g991 ( .A(n_883), .B(n_891), .Y(n_991) );
OR2x2_ASAP7_75t_L g992 ( .A(n_864), .B(n_886), .Y(n_992) );
AOI22xp33_ASAP7_75t_L g993 ( .A1(n_889), .A2(n_897), .B1(n_892), .B2(n_933), .Y(n_993) );
AND2x2_ASAP7_75t_L g994 ( .A(n_850), .B(n_946), .Y(n_994) );
INVx2_ASAP7_75t_L g995 ( .A(n_856), .Y(n_995) );
INVx2_ASAP7_75t_L g996 ( .A(n_924), .Y(n_996) );
BUFx3_ASAP7_75t_L g997 ( .A(n_878), .Y(n_997) );
AND2x2_ASAP7_75t_L g998 ( .A(n_955), .B(n_957), .Y(n_998) );
AND2x2_ASAP7_75t_L g999 ( .A(n_958), .B(n_893), .Y(n_999) );
INVx1_ASAP7_75t_L g1000 ( .A(n_886), .Y(n_1000) );
OR2x2_ASAP7_75t_L g1001 ( .A(n_896), .B(n_884), .Y(n_1001) );
INVxp67_ASAP7_75t_SL g1002 ( .A(n_848), .Y(n_1002) );
AND2x4_ASAP7_75t_L g1003 ( .A(n_863), .B(n_941), .Y(n_1003) );
INVx1_ASAP7_75t_L g1004 ( .A(n_896), .Y(n_1004) );
HB1xp67_ASAP7_75t_L g1005 ( .A(n_902), .Y(n_1005) );
AND2x2_ASAP7_75t_L g1006 ( .A(n_876), .B(n_863), .Y(n_1006) );
INVx1_ASAP7_75t_L g1007 ( .A(n_921), .Y(n_1007) );
INVx1_ASAP7_75t_L g1008 ( .A(n_915), .Y(n_1008) );
NAND2xp5_ASAP7_75t_L g1009 ( .A(n_887), .B(n_895), .Y(n_1009) );
NAND2xp5_ASAP7_75t_L g1010 ( .A(n_894), .B(n_846), .Y(n_1010) );
BUFx3_ASAP7_75t_L g1011 ( .A(n_941), .Y(n_1011) );
AND2x2_ASAP7_75t_L g1012 ( .A(n_950), .B(n_867), .Y(n_1012) );
INVx2_ASAP7_75t_L g1013 ( .A(n_914), .Y(n_1013) );
NAND2xp5_ASAP7_75t_L g1014 ( .A(n_899), .B(n_851), .Y(n_1014) );
INVx1_ASAP7_75t_L g1015 ( .A(n_877), .Y(n_1015) );
AND2x4_ASAP7_75t_L g1016 ( .A(n_952), .B(n_852), .Y(n_1016) );
INVx1_ASAP7_75t_L g1017 ( .A(n_903), .Y(n_1017) );
INVx1_ASAP7_75t_L g1018 ( .A(n_911), .Y(n_1018) );
AND2x2_ASAP7_75t_L g1019 ( .A(n_952), .B(n_874), .Y(n_1019) );
AND2x4_ASAP7_75t_L g1020 ( .A(n_909), .B(n_860), .Y(n_1020) );
AND2x2_ASAP7_75t_L g1021 ( .A(n_874), .B(n_865), .Y(n_1021) );
AND2x2_ASAP7_75t_L g1022 ( .A(n_912), .B(n_861), .Y(n_1022) );
AND2x2_ASAP7_75t_L g1023 ( .A(n_849), .B(n_890), .Y(n_1023) );
AND2x2_ASAP7_75t_L g1024 ( .A(n_890), .B(n_854), .Y(n_1024) );
AND2x2_ASAP7_75t_L g1025 ( .A(n_890), .B(n_900), .Y(n_1025) );
BUFx2_ASAP7_75t_L g1026 ( .A(n_916), .Y(n_1026) );
OR2x2_ASAP7_75t_L g1027 ( .A(n_898), .B(n_859), .Y(n_1027) );
AND2x2_ASAP7_75t_L g1028 ( .A(n_900), .B(n_935), .Y(n_1028) );
AND2x4_ASAP7_75t_L g1029 ( .A(n_909), .B(n_853), .Y(n_1029) );
AND2x4_ASAP7_75t_L g1030 ( .A(n_868), .B(n_939), .Y(n_1030) );
NOR2x1_ASAP7_75t_L g1031 ( .A(n_855), .B(n_868), .Y(n_1031) );
OR2x2_ASAP7_75t_L g1032 ( .A(n_905), .B(n_869), .Y(n_1032) );
AND2x4_ASAP7_75t_L g1033 ( .A(n_939), .B(n_905), .Y(n_1033) );
AND2x4_ASAP7_75t_L g1034 ( .A(n_939), .B(n_962), .Y(n_1034) );
INVx2_ASAP7_75t_L g1035 ( .A(n_926), .Y(n_1035) );
AND2x4_ASAP7_75t_L g1036 ( .A(n_937), .B(n_932), .Y(n_1036) );
INVx1_ASAP7_75t_L g1037 ( .A(n_928), .Y(n_1037) );
NOR2xp33_ASAP7_75t_L g1038 ( .A(n_869), .B(n_847), .Y(n_1038) );
INVxp67_ASAP7_75t_L g1039 ( .A(n_934), .Y(n_1039) );
CKINVDCx11_ASAP7_75t_R g1040 ( .A(n_906), .Y(n_1040) );
AND2x2_ASAP7_75t_L g1041 ( .A(n_875), .B(n_922), .Y(n_1041) );
INVx1_ASAP7_75t_L g1042 ( .A(n_928), .Y(n_1042) );
INVx1_ASAP7_75t_L g1043 ( .A(n_930), .Y(n_1043) );
INVx1_ASAP7_75t_L g1044 ( .A(n_919), .Y(n_1044) );
OR2x2_ASAP7_75t_L g1045 ( .A(n_947), .B(n_916), .Y(n_1045) );
INVx2_ASAP7_75t_L g1046 ( .A(n_919), .Y(n_1046) );
INVx2_ASAP7_75t_L g1047 ( .A(n_870), .Y(n_1047) );
INVx1_ASAP7_75t_L g1048 ( .A(n_879), .Y(n_1048) );
AND2x2_ASAP7_75t_L g1049 ( .A(n_1023), .B(n_913), .Y(n_1049) );
AO21x2_ASAP7_75t_L g1050 ( .A1(n_995), .A2(n_879), .B(n_888), .Y(n_1050) );
AOI221xp5_ASAP7_75t_L g1051 ( .A1(n_968), .A2(n_871), .B1(n_906), .B2(n_931), .C(n_872), .Y(n_1051) );
AOI211xp5_ASAP7_75t_L g1052 ( .A1(n_1021), .A2(n_871), .B(n_917), .C(n_1047), .Y(n_1052) );
AND2x2_ASAP7_75t_L g1053 ( .A(n_1023), .B(n_917), .Y(n_1053) );
HB1xp67_ASAP7_75t_L g1054 ( .A(n_967), .Y(n_1054) );
AND2x2_ASAP7_75t_L g1055 ( .A(n_983), .B(n_985), .Y(n_1055) );
OAI31xp33_ASAP7_75t_L g1056 ( .A1(n_1021), .A2(n_964), .A3(n_1047), .B(n_1019), .Y(n_1056) );
AND2x2_ASAP7_75t_L g1057 ( .A(n_983), .B(n_985), .Y(n_1057) );
INVx1_ASAP7_75t_L g1058 ( .A(n_978), .Y(n_1058) );
INVx5_ASAP7_75t_L g1059 ( .A(n_974), .Y(n_1059) );
INVxp67_ASAP7_75t_SL g1060 ( .A(n_1008), .Y(n_1060) );
INVx1_ASAP7_75t_L g1061 ( .A(n_978), .Y(n_1061) );
INVx1_ASAP7_75t_L g1062 ( .A(n_975), .Y(n_1062) );
AND2x2_ASAP7_75t_L g1063 ( .A(n_1028), .B(n_1025), .Y(n_1063) );
AND2x4_ASAP7_75t_L g1064 ( .A(n_1028), .B(n_1025), .Y(n_1064) );
AND2x2_ASAP7_75t_L g1065 ( .A(n_1000), .B(n_1004), .Y(n_1065) );
AND2x2_ASAP7_75t_L g1066 ( .A(n_1000), .B(n_1004), .Y(n_1066) );
OAI22xp5_ASAP7_75t_L g1067 ( .A1(n_976), .A2(n_993), .B1(n_1019), .B2(n_1010), .Y(n_1067) );
INVx1_ASAP7_75t_L g1068 ( .A(n_975), .Y(n_1068) );
AND2x2_ASAP7_75t_L g1069 ( .A(n_970), .B(n_976), .Y(n_1069) );
INVx1_ASAP7_75t_L g1070 ( .A(n_982), .Y(n_1070) );
NOR3xp33_ASAP7_75t_L g1071 ( .A(n_1038), .B(n_1039), .C(n_1009), .Y(n_1071) );
AND2x2_ASAP7_75t_L g1072 ( .A(n_970), .B(n_1024), .Y(n_1072) );
HB1xp67_ASAP7_75t_L g1073 ( .A(n_965), .Y(n_1073) );
INVx2_ASAP7_75t_L g1074 ( .A(n_1013), .Y(n_1074) );
AND2x2_ASAP7_75t_L g1075 ( .A(n_1024), .B(n_992), .Y(n_1075) );
INVx1_ASAP7_75t_L g1076 ( .A(n_992), .Y(n_1076) );
AOI22xp33_ASAP7_75t_L g1077 ( .A1(n_979), .A2(n_971), .B1(n_1012), .B2(n_1001), .Y(n_1077) );
INVx2_ASAP7_75t_SL g1078 ( .A(n_974), .Y(n_1078) );
HB1xp67_ASAP7_75t_L g1079 ( .A(n_966), .Y(n_1079) );
AND2x2_ASAP7_75t_L g1080 ( .A(n_999), .B(n_1012), .Y(n_1080) );
AND2x2_ASAP7_75t_L g1081 ( .A(n_999), .B(n_994), .Y(n_1081) );
AOI22xp33_ASAP7_75t_L g1082 ( .A1(n_979), .A2(n_1001), .B1(n_1027), .B2(n_1022), .Y(n_1082) );
AND2x2_ASAP7_75t_L g1083 ( .A(n_994), .B(n_998), .Y(n_1083) );
INVx1_ASAP7_75t_SL g1084 ( .A(n_1040), .Y(n_1084) );
INVx1_ASAP7_75t_L g1085 ( .A(n_996), .Y(n_1085) );
NAND2xp5_ASAP7_75t_L g1086 ( .A(n_991), .B(n_998), .Y(n_1086) );
AOI22xp33_ASAP7_75t_L g1087 ( .A1(n_1027), .A2(n_1022), .B1(n_1041), .B2(n_1026), .Y(n_1087) );
AND2x2_ASAP7_75t_L g1088 ( .A(n_988), .B(n_1026), .Y(n_1088) );
NAND2xp5_ASAP7_75t_L g1089 ( .A(n_1007), .B(n_989), .Y(n_1089) );
INVx1_ASAP7_75t_L g1090 ( .A(n_1045), .Y(n_1090) );
OAI21xp33_ASAP7_75t_L g1091 ( .A1(n_1048), .A2(n_1002), .B(n_1017), .Y(n_1091) );
AND2x2_ASAP7_75t_L g1092 ( .A(n_1017), .B(n_981), .Y(n_1092) );
AND2x4_ASAP7_75t_L g1093 ( .A(n_990), .B(n_973), .Y(n_1093) );
OAI321xp33_ASAP7_75t_L g1094 ( .A1(n_1032), .A2(n_1014), .A3(n_1041), .B1(n_1015), .B2(n_1044), .C(n_1037), .Y(n_1094) );
INVx1_ASAP7_75t_L g1095 ( .A(n_1032), .Y(n_1095) );
INVx1_ASAP7_75t_L g1096 ( .A(n_1043), .Y(n_1096) );
INVx2_ASAP7_75t_SL g1097 ( .A(n_1011), .Y(n_1097) );
NAND2xp5_ASAP7_75t_L g1098 ( .A(n_981), .B(n_972), .Y(n_1098) );
AOI22xp33_ASAP7_75t_L g1099 ( .A1(n_1006), .A2(n_986), .B1(n_1016), .B2(n_1018), .Y(n_1099) );
BUFx2_ASAP7_75t_L g1100 ( .A(n_990), .Y(n_1100) );
AOI22xp5_ASAP7_75t_L g1101 ( .A1(n_1006), .A2(n_1018), .B1(n_977), .B2(n_980), .Y(n_1101) );
CKINVDCx5p33_ASAP7_75t_R g1102 ( .A(n_1084), .Y(n_1102) );
AND2x2_ASAP7_75t_L g1103 ( .A(n_1072), .B(n_1033), .Y(n_1103) );
AND2x2_ASAP7_75t_L g1104 ( .A(n_1072), .B(n_1033), .Y(n_1104) );
AND2x2_ASAP7_75t_L g1105 ( .A(n_1063), .B(n_1033), .Y(n_1105) );
AND2x2_ASAP7_75t_L g1106 ( .A(n_1063), .B(n_1033), .Y(n_1106) );
OR2x2_ASAP7_75t_L g1107 ( .A(n_1088), .B(n_1046), .Y(n_1107) );
AND2x2_ASAP7_75t_L g1108 ( .A(n_1075), .B(n_1034), .Y(n_1108) );
INVx1_ASAP7_75t_L g1109 ( .A(n_1058), .Y(n_1109) );
INVx1_ASAP7_75t_L g1110 ( .A(n_1058), .Y(n_1110) );
AND2x2_ASAP7_75t_L g1111 ( .A(n_1075), .B(n_1034), .Y(n_1111) );
AND2x2_ASAP7_75t_L g1112 ( .A(n_1064), .B(n_1034), .Y(n_1112) );
AND2x4_ASAP7_75t_L g1113 ( .A(n_1093), .B(n_1064), .Y(n_1113) );
AND2x4_ASAP7_75t_L g1114 ( .A(n_1093), .B(n_1029), .Y(n_1114) );
INVx2_ASAP7_75t_L g1115 ( .A(n_1074), .Y(n_1115) );
INVx1_ASAP7_75t_SL g1116 ( .A(n_1081), .Y(n_1116) );
AOI22xp5_ASAP7_75t_L g1117 ( .A1(n_1067), .A2(n_1016), .B1(n_997), .B2(n_1003), .Y(n_1117) );
AND2x2_ASAP7_75t_L g1118 ( .A(n_1064), .B(n_1034), .Y(n_1118) );
NAND2xp5_ASAP7_75t_L g1119 ( .A(n_1083), .B(n_980), .Y(n_1119) );
INVx1_ASAP7_75t_L g1120 ( .A(n_1061), .Y(n_1120) );
NOR2x1_ASAP7_75t_SL g1121 ( .A(n_1097), .B(n_1011), .Y(n_1121) );
AND2x2_ASAP7_75t_L g1122 ( .A(n_1080), .B(n_1042), .Y(n_1122) );
BUFx2_ASAP7_75t_L g1123 ( .A(n_1097), .Y(n_1123) );
INVx1_ASAP7_75t_L g1124 ( .A(n_1062), .Y(n_1124) );
AOI22xp33_ASAP7_75t_L g1125 ( .A1(n_1056), .A2(n_1016), .B1(n_997), .B2(n_1005), .Y(n_1125) );
INVxp67_ASAP7_75t_SL g1126 ( .A(n_1060), .Y(n_1126) );
NOR2xp33_ASAP7_75t_L g1127 ( .A(n_1086), .B(n_969), .Y(n_1127) );
INVx1_ASAP7_75t_L g1128 ( .A(n_1068), .Y(n_1128) );
AND2x2_ASAP7_75t_L g1129 ( .A(n_1080), .B(n_1042), .Y(n_1129) );
OAI221xp5_ASAP7_75t_L g1130 ( .A1(n_1071), .A2(n_997), .B1(n_1011), .B2(n_987), .C(n_1035), .Y(n_1130) );
NAND3xp33_ASAP7_75t_L g1131 ( .A(n_1051), .B(n_1035), .C(n_1036), .Y(n_1131) );
AND2x2_ASAP7_75t_L g1132 ( .A(n_1049), .B(n_984), .Y(n_1132) );
INVx1_ASAP7_75t_L g1133 ( .A(n_1070), .Y(n_1133) );
INVx1_ASAP7_75t_L g1134 ( .A(n_1070), .Y(n_1134) );
AND2x2_ASAP7_75t_L g1135 ( .A(n_1049), .B(n_984), .Y(n_1135) );
AND2x2_ASAP7_75t_L g1136 ( .A(n_1088), .B(n_1036), .Y(n_1136) );
OR2x6_ASAP7_75t_L g1137 ( .A(n_1100), .B(n_990), .Y(n_1137) );
AND2x4_ASAP7_75t_L g1138 ( .A(n_1055), .B(n_1029), .Y(n_1138) );
INVxp67_ASAP7_75t_L g1139 ( .A(n_1073), .Y(n_1139) );
AND2x4_ASAP7_75t_L g1140 ( .A(n_1057), .B(n_1029), .Y(n_1140) );
AND2x2_ASAP7_75t_L g1141 ( .A(n_1057), .B(n_1030), .Y(n_1141) );
AND2x4_ASAP7_75t_L g1142 ( .A(n_1095), .B(n_1020), .Y(n_1142) );
AND2x2_ASAP7_75t_L g1143 ( .A(n_1065), .B(n_1030), .Y(n_1143) );
OAI21xp33_ASAP7_75t_L g1144 ( .A1(n_1116), .A2(n_1091), .B(n_1082), .Y(n_1144) );
AND2x2_ASAP7_75t_L g1145 ( .A(n_1103), .B(n_1053), .Y(n_1145) );
NAND2xp5_ASAP7_75t_L g1146 ( .A(n_1122), .B(n_1054), .Y(n_1146) );
OR2x2_ASAP7_75t_L g1147 ( .A(n_1119), .B(n_1079), .Y(n_1147) );
INVx1_ASAP7_75t_L g1148 ( .A(n_1109), .Y(n_1148) );
AND2x2_ASAP7_75t_L g1149 ( .A(n_1103), .B(n_1053), .Y(n_1149) );
BUFx3_ASAP7_75t_L g1150 ( .A(n_1123), .Y(n_1150) );
AND2x2_ASAP7_75t_L g1151 ( .A(n_1104), .B(n_1090), .Y(n_1151) );
NAND2xp5_ASAP7_75t_L g1152 ( .A(n_1122), .B(n_1092), .Y(n_1152) );
AOI22xp5_ASAP7_75t_L g1153 ( .A1(n_1125), .A2(n_1069), .B1(n_1077), .B2(n_1087), .Y(n_1153) );
INVx1_ASAP7_75t_L g1154 ( .A(n_1109), .Y(n_1154) );
INVx1_ASAP7_75t_L g1155 ( .A(n_1110), .Y(n_1155) );
AND2x2_ASAP7_75t_L g1156 ( .A(n_1104), .B(n_1090), .Y(n_1156) );
AND2x2_ASAP7_75t_L g1157 ( .A(n_1143), .B(n_1066), .Y(n_1157) );
INVx1_ASAP7_75t_L g1158 ( .A(n_1110), .Y(n_1158) );
NAND2xp5_ASAP7_75t_L g1159 ( .A(n_1129), .B(n_1069), .Y(n_1159) );
INVx2_ASAP7_75t_L g1160 ( .A(n_1115), .Y(n_1160) );
NOR2xp33_ASAP7_75t_L g1161 ( .A(n_1139), .B(n_1094), .Y(n_1161) );
AND2x2_ASAP7_75t_L g1162 ( .A(n_1143), .B(n_1065), .Y(n_1162) );
NAND2xp33_ASAP7_75t_SL g1163 ( .A(n_1123), .B(n_1100), .Y(n_1163) );
NOR2xp33_ASAP7_75t_L g1164 ( .A(n_1117), .B(n_1089), .Y(n_1164) );
NAND2xp5_ASAP7_75t_L g1165 ( .A(n_1126), .B(n_1066), .Y(n_1165) );
NAND3xp33_ASAP7_75t_L g1166 ( .A(n_1131), .B(n_1052), .C(n_1091), .Y(n_1166) );
NAND2xp5_ASAP7_75t_L g1167 ( .A(n_1133), .B(n_1101), .Y(n_1167) );
AOI21xp5_ASAP7_75t_L g1168 ( .A1(n_1121), .A2(n_1031), .B(n_1078), .Y(n_1168) );
AOI22xp5_ASAP7_75t_L g1169 ( .A1(n_1130), .A2(n_1101), .B1(n_1099), .B2(n_1016), .Y(n_1169) );
NAND2xp5_ASAP7_75t_L g1170 ( .A(n_1133), .B(n_1076), .Y(n_1170) );
AND2x2_ASAP7_75t_L g1171 ( .A(n_1108), .B(n_1076), .Y(n_1171) );
INVx1_ASAP7_75t_L g1172 ( .A(n_1120), .Y(n_1172) );
NAND2xp5_ASAP7_75t_L g1173 ( .A(n_1134), .B(n_1098), .Y(n_1173) );
AND2x2_ASAP7_75t_L g1174 ( .A(n_1108), .B(n_1096), .Y(n_1174) );
OR2x2_ASAP7_75t_L g1175 ( .A(n_1107), .B(n_1085), .Y(n_1175) );
AOI22xp5_ASAP7_75t_L g1176 ( .A1(n_1153), .A2(n_1132), .B1(n_1135), .B2(n_1140), .Y(n_1176) );
INVx1_ASAP7_75t_L g1177 ( .A(n_1148), .Y(n_1177) );
AOI221xp5_ASAP7_75t_L g1178 ( .A1(n_1161), .A2(n_1111), .B1(n_1106), .B2(n_1105), .C(n_1132), .Y(n_1178) );
XNOR2x1_ASAP7_75t_L g1179 ( .A(n_1147), .B(n_1102), .Y(n_1179) );
AND2x2_ASAP7_75t_L g1180 ( .A(n_1157), .B(n_1113), .Y(n_1180) );
INVx1_ASAP7_75t_L g1181 ( .A(n_1154), .Y(n_1181) );
NAND2xp5_ASAP7_75t_L g1182 ( .A(n_1171), .B(n_1111), .Y(n_1182) );
AOI22xp33_ASAP7_75t_L g1183 ( .A1(n_1166), .A2(n_1127), .B1(n_1140), .B2(n_1138), .Y(n_1183) );
INVx1_ASAP7_75t_L g1184 ( .A(n_1155), .Y(n_1184) );
NOR2xp33_ASAP7_75t_L g1185 ( .A(n_1161), .B(n_1135), .Y(n_1185) );
AOI22xp5_ASAP7_75t_L g1186 ( .A1(n_1164), .A2(n_1140), .B1(n_1138), .B2(n_1136), .Y(n_1186) );
AOI22xp33_ASAP7_75t_L g1187 ( .A1(n_1144), .A2(n_1140), .B1(n_1138), .B2(n_1142), .Y(n_1187) );
OAI221xp5_ASAP7_75t_SL g1188 ( .A1(n_1169), .A2(n_1164), .B1(n_1159), .B2(n_1146), .C(n_1167), .Y(n_1188) );
NAND2xp5_ASAP7_75t_L g1189 ( .A(n_1174), .B(n_1141), .Y(n_1189) );
INVx1_ASAP7_75t_L g1190 ( .A(n_1158), .Y(n_1190) );
INVx1_ASAP7_75t_L g1191 ( .A(n_1172), .Y(n_1191) );
AOI31xp33_ASAP7_75t_L g1192 ( .A1(n_1163), .A2(n_1113), .A3(n_1118), .B(n_1112), .Y(n_1192) );
NOR2xp67_ASAP7_75t_SL g1193 ( .A(n_1150), .B(n_1059), .Y(n_1193) );
INVxp67_ASAP7_75t_L g1194 ( .A(n_1165), .Y(n_1194) );
NOR2xp33_ASAP7_75t_L g1195 ( .A(n_1152), .B(n_1112), .Y(n_1195) );
BUFx2_ASAP7_75t_L g1196 ( .A(n_1163), .Y(n_1196) );
INVx2_ASAP7_75t_L g1197 ( .A(n_1160), .Y(n_1197) );
INVx1_ASAP7_75t_SL g1198 ( .A(n_1175), .Y(n_1198) );
NAND2xp5_ASAP7_75t_L g1199 ( .A(n_1185), .B(n_1157), .Y(n_1199) );
INVx1_ASAP7_75t_L g1200 ( .A(n_1197), .Y(n_1200) );
INVx2_ASAP7_75t_L g1201 ( .A(n_1197), .Y(n_1201) );
INVx2_ASAP7_75t_L g1202 ( .A(n_1177), .Y(n_1202) );
INVx1_ASAP7_75t_L g1203 ( .A(n_1181), .Y(n_1203) );
INVx3_ASAP7_75t_L g1204 ( .A(n_1196), .Y(n_1204) );
INVx1_ASAP7_75t_SL g1205 ( .A(n_1179), .Y(n_1205) );
INVx1_ASAP7_75t_L g1206 ( .A(n_1184), .Y(n_1206) );
NOR3xp33_ASAP7_75t_L g1207 ( .A(n_1188), .B(n_1170), .C(n_1173), .Y(n_1207) );
OAI22xp5_ASAP7_75t_L g1208 ( .A1(n_1192), .A2(n_1137), .B1(n_1149), .B2(n_1145), .Y(n_1208) );
AND2x2_ASAP7_75t_L g1209 ( .A(n_1180), .B(n_1145), .Y(n_1209) );
INVx1_ASAP7_75t_L g1210 ( .A(n_1190), .Y(n_1210) );
INVx1_ASAP7_75t_L g1211 ( .A(n_1191), .Y(n_1211) );
NAND2xp5_ASAP7_75t_L g1212 ( .A(n_1198), .B(n_1162), .Y(n_1212) );
AND2x2_ASAP7_75t_L g1213 ( .A(n_1194), .B(n_1149), .Y(n_1213) );
NAND2xp5_ASAP7_75t_L g1214 ( .A(n_1178), .B(n_1162), .Y(n_1214) );
OR2x2_ASAP7_75t_L g1215 ( .A(n_1212), .B(n_1189), .Y(n_1215) );
AOI22xp5_ASAP7_75t_L g1216 ( .A1(n_1205), .A2(n_1183), .B1(n_1176), .B2(n_1187), .Y(n_1216) );
OAI22xp33_ASAP7_75t_SL g1217 ( .A1(n_1204), .A2(n_1186), .B1(n_1182), .B2(n_1195), .Y(n_1217) );
OAI21xp33_ASAP7_75t_SL g1218 ( .A1(n_1204), .A2(n_1187), .B(n_1183), .Y(n_1218) );
NAND2xp5_ASAP7_75t_L g1219 ( .A(n_1207), .B(n_1174), .Y(n_1219) );
AOI22xp5_ASAP7_75t_L g1220 ( .A1(n_1214), .A2(n_1195), .B1(n_1118), .B2(n_1151), .Y(n_1220) );
AOI22xp5_ASAP7_75t_L g1221 ( .A1(n_1208), .A2(n_1156), .B1(n_1151), .B2(n_1136), .Y(n_1221) );
OAI21xp5_ASAP7_75t_L g1222 ( .A1(n_1204), .A2(n_1168), .B(n_1193), .Y(n_1222) );
AOI322xp5_ASAP7_75t_L g1223 ( .A1(n_1218), .A2(n_1213), .A3(n_1199), .B1(n_1209), .B2(n_1211), .C1(n_1203), .C2(n_1210), .Y(n_1223) );
INVx1_ASAP7_75t_L g1224 ( .A(n_1215), .Y(n_1224) );
AOI221xp5_ASAP7_75t_L g1225 ( .A1(n_1217), .A2(n_1206), .B1(n_1211), .B2(n_1203), .C(n_1202), .Y(n_1225) );
AOI221xp5_ASAP7_75t_L g1226 ( .A1(n_1217), .A2(n_1202), .B1(n_1200), .B2(n_1201), .C(n_1138), .Y(n_1226) );
AOI221xp5_ASAP7_75t_L g1227 ( .A1(n_1219), .A2(n_1216), .B1(n_1222), .B2(n_1220), .C(n_1221), .Y(n_1227) );
INVx2_ASAP7_75t_L g1228 ( .A(n_1224), .Y(n_1228) );
INVx1_ASAP7_75t_L g1229 ( .A(n_1227), .Y(n_1229) );
NOR4xp25_ASAP7_75t_L g1230 ( .A(n_1229), .B(n_1225), .C(n_1226), .D(n_1223), .Y(n_1230) );
INVx4_ASAP7_75t_L g1231 ( .A(n_1228), .Y(n_1231) );
INVx1_ASAP7_75t_L g1232 ( .A(n_1231), .Y(n_1232) );
NAND2xp5_ASAP7_75t_L g1233 ( .A(n_1232), .B(n_1230), .Y(n_1233) );
INVxp67_ASAP7_75t_SL g1234 ( .A(n_1233), .Y(n_1234) );
AOI22xp5_ASAP7_75t_L g1235 ( .A1(n_1234), .A2(n_1050), .B1(n_1114), .B2(n_1142), .Y(n_1235) );
INVx4_ASAP7_75t_L g1236 ( .A(n_1235), .Y(n_1236) );
AOI211xp5_ASAP7_75t_L g1237 ( .A1(n_1236), .A2(n_1175), .B(n_1128), .C(n_1124), .Y(n_1237) );
endmodule