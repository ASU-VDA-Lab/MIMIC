module fake_netlist_5_195_n_1925 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_173, n_25, n_53, n_160, n_188, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1925);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_173;
input n_25;
input n_53;
input n_160;
input n_188;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1925;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_798;
wire n_196;
wire n_350;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_290;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_759;
wire n_1892;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_1916;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_433;
wire n_368;
wire n_604;
wire n_314;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_448;
wire n_259;
wire n_1851;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_1874;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1692;
wire n_1596;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_1902;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1875;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_584;
wire n_681;
wire n_336;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_1904;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1726;
wire n_665;
wire n_1835;
wire n_1584;
wire n_1440;
wire n_421;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1689;
wire n_1524;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1898;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVx1_ASAP7_75t_SL g189 ( 
.A(n_48),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_37),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_115),
.Y(n_191)
);

BUFx10_ASAP7_75t_L g192 ( 
.A(n_59),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_14),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_170),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_179),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_48),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_22),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_144),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_160),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_172),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_42),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_150),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_50),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_41),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_38),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_110),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_109),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g208 ( 
.A(n_21),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_41),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_9),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_125),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_3),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_8),
.Y(n_213)
);

CKINVDCx14_ASAP7_75t_R g214 ( 
.A(n_145),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_152),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_25),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_138),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_116),
.Y(n_218)
);

INVx2_ASAP7_75t_SL g219 ( 
.A(n_52),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_148),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_72),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_53),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_154),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_143),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_173),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_96),
.Y(n_226)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_39),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_120),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_9),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_86),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_90),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_178),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_186),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_84),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_76),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_94),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_169),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_6),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_40),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_66),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_77),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_158),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_10),
.Y(n_243)
);

INVx2_ASAP7_75t_SL g244 ( 
.A(n_140),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_18),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_67),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_3),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_44),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_187),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_126),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_49),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_56),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_161),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_49),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_38),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_73),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_24),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_52),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_129),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_176),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_25),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_108),
.Y(n_262)
);

INVx2_ASAP7_75t_SL g263 ( 
.A(n_89),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_83),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g265 ( 
.A(n_168),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_146),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_63),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_102),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_100),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_39),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_91),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_117),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_153),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_60),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_45),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_151),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_12),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_11),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_23),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_123),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_82),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_147),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_98),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_156),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_142),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_64),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_133),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_35),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_1),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_29),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_15),
.Y(n_291)
);

BUFx10_ASAP7_75t_L g292 ( 
.A(n_132),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_124),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_62),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_149),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_127),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_112),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_136),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_1),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_139),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_19),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_85),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_17),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_6),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_159),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_35),
.Y(n_306)
);

BUFx10_ASAP7_75t_L g307 ( 
.A(n_79),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_58),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_29),
.Y(n_309)
);

BUFx2_ASAP7_75t_L g310 ( 
.A(n_65),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_46),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_69),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_10),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_177),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_65),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_4),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_11),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_4),
.Y(n_318)
);

INVx1_ASAP7_75t_SL g319 ( 
.A(n_16),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_0),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_141),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_47),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_7),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_114),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_106),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_68),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_121),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_88),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_45),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_182),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_24),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_128),
.Y(n_332)
);

BUFx10_ASAP7_75t_L g333 ( 
.A(n_60),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_8),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_67),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_14),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_16),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_188),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_2),
.Y(n_339)
);

BUFx10_ASAP7_75t_L g340 ( 
.A(n_12),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_37),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_162),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_23),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_103),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_19),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_50),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_17),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_61),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_104),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_63),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_59),
.Y(n_351)
);

INVx1_ASAP7_75t_SL g352 ( 
.A(n_171),
.Y(n_352)
);

BUFx2_ASAP7_75t_L g353 ( 
.A(n_32),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_42),
.Y(n_354)
);

INVx2_ASAP7_75t_SL g355 ( 
.A(n_166),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_80),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_33),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_33),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_27),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_22),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_54),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_180),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_118),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_2),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_165),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_21),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_54),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_87),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_28),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_66),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_134),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_163),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_155),
.Y(n_373)
);

INVx1_ASAP7_75t_SL g374 ( 
.A(n_74),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_122),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_28),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_7),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_113),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_68),
.Y(n_379)
);

BUFx2_ASAP7_75t_L g380 ( 
.A(n_208),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_229),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_191),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_191),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_195),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_198),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_195),
.Y(n_386)
);

CKINVDCx16_ASAP7_75t_R g387 ( 
.A(n_229),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_190),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_208),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_200),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_193),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_220),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_196),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_200),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_244),
.B(n_0),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_201),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_202),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_310),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_202),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_310),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_221),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_221),
.Y(n_402)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_197),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_215),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_234),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_205),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_235),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_260),
.Y(n_408)
);

INVxp33_ASAP7_75t_L g409 ( 
.A(n_353),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_265),
.B(n_5),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_194),
.Y(n_411)
);

BUFx6f_ASAP7_75t_SL g412 ( 
.A(n_307),
.Y(n_412)
);

INVxp67_ASAP7_75t_SL g413 ( 
.A(n_227),
.Y(n_413)
);

HB1xp67_ASAP7_75t_L g414 ( 
.A(n_353),
.Y(n_414)
);

OR2x2_ASAP7_75t_L g415 ( 
.A(n_203),
.B(n_5),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_325),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_209),
.Y(n_417)
);

BUFx2_ASAP7_75t_L g418 ( 
.A(n_213),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_244),
.B(n_13),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_235),
.Y(n_420)
);

CKINVDCx16_ASAP7_75t_R g421 ( 
.A(n_226),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_216),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_263),
.B(n_13),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_222),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_363),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_238),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_239),
.Y(n_427)
);

CKINVDCx16_ASAP7_75t_R g428 ( 
.A(n_226),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_230),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_237),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_245),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_230),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_251),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_237),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_242),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_242),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_214),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_252),
.Y(n_438)
);

INVxp33_ASAP7_75t_SL g439 ( 
.A(n_254),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_249),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_255),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_258),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_249),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_199),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_270),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_268),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_275),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_268),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_277),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_271),
.Y(n_450)
);

BUFx3_ASAP7_75t_L g451 ( 
.A(n_228),
.Y(n_451)
);

INVxp67_ASAP7_75t_L g452 ( 
.A(n_340),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_278),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_271),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_286),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_289),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_285),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_206),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_207),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_285),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_293),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_291),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_299),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_293),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_301),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_295),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_295),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_298),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_227),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_303),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_263),
.B(n_15),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_298),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_302),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_306),
.Y(n_474)
);

BUFx6f_ASAP7_75t_L g475 ( 
.A(n_404),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_413),
.B(n_227),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_403),
.Y(n_477)
);

INVx3_ASAP7_75t_L g478 ( 
.A(n_404),
.Y(n_478)
);

AND2x4_ASAP7_75t_L g479 ( 
.A(n_469),
.B(n_228),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_403),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_404),
.Y(n_481)
);

OA21x2_ASAP7_75t_L g482 ( 
.A1(n_469),
.A2(n_315),
.B(n_279),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_404),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_411),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_403),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_404),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_382),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_383),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_384),
.Y(n_489)
);

AND2x4_ASAP7_75t_L g490 ( 
.A(n_386),
.B(n_355),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_390),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_394),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_397),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_399),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_401),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_419),
.B(n_197),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g497 ( 
.A(n_402),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_471),
.B(n_197),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_407),
.Y(n_499)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_420),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_430),
.B(n_197),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_434),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_435),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_436),
.B(n_197),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_429),
.B(n_243),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_395),
.B(n_355),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_440),
.B(n_359),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_443),
.Y(n_508)
);

HB1xp67_ASAP7_75t_L g509 ( 
.A(n_381),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_446),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_448),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_432),
.A2(n_257),
.B1(n_326),
.B2(n_248),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_450),
.Y(n_513)
);

INVx3_ASAP7_75t_L g514 ( 
.A(n_454),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_457),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_460),
.B(n_359),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_461),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_464),
.Y(n_518)
);

INVx3_ASAP7_75t_L g519 ( 
.A(n_466),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_467),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_468),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_472),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_473),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_451),
.B(n_359),
.Y(n_524)
);

BUFx3_ASAP7_75t_L g525 ( 
.A(n_451),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_423),
.B(n_359),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_410),
.B(n_359),
.Y(n_527)
);

AND2x4_ASAP7_75t_L g528 ( 
.A(n_415),
.B(n_256),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_415),
.Y(n_529)
);

AND2x4_ASAP7_75t_L g530 ( 
.A(n_418),
.B(n_256),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_412),
.Y(n_531)
);

AND2x4_ASAP7_75t_L g532 ( 
.A(n_389),
.B(n_269),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_412),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_412),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_388),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g536 ( 
.A(n_398),
.B(n_302),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_400),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_380),
.B(n_321),
.Y(n_538)
);

AND2x4_ASAP7_75t_L g539 ( 
.A(n_452),
.B(n_269),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g540 ( 
.A(n_388),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_391),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_414),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_391),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_393),
.B(n_211),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_393),
.Y(n_545)
);

INVxp33_ASAP7_75t_L g546 ( 
.A(n_409),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_396),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_396),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_406),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_406),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_417),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_417),
.B(n_218),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_439),
.B(n_262),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_422),
.B(n_321),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_482),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_487),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_487),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_482),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_482),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_484),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_540),
.B(n_421),
.Y(n_561)
);

AND2x2_ASAP7_75t_L g562 ( 
.A(n_529),
.B(n_422),
.Y(n_562)
);

AOI22xp33_ASAP7_75t_L g563 ( 
.A1(n_528),
.A2(n_219),
.B1(n_315),
.B2(n_279),
.Y(n_563)
);

AO22x2_ASAP7_75t_L g564 ( 
.A1(n_538),
.A2(n_219),
.B1(n_203),
.B2(n_210),
.Y(n_564)
);

BUFx4f_ASAP7_75t_L g565 ( 
.A(n_540),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_482),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_482),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_482),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_493),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_544),
.B(n_428),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_475),
.Y(n_571)
);

INVx4_ASAP7_75t_L g572 ( 
.A(n_497),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_506),
.B(n_424),
.Y(n_573)
);

BUFx3_ASAP7_75t_L g574 ( 
.A(n_525),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_506),
.B(n_424),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_475),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_540),
.B(n_437),
.Y(n_577)
);

OR2x6_ASAP7_75t_L g578 ( 
.A(n_531),
.B(n_328),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_529),
.B(n_426),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_528),
.B(n_426),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_487),
.Y(n_581)
);

OR2x6_ASAP7_75t_L g582 ( 
.A(n_531),
.B(n_328),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_487),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_493),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_529),
.B(n_524),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_493),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_502),
.Y(n_587)
);

INVx6_ASAP7_75t_L g588 ( 
.A(n_479),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_540),
.B(n_427),
.Y(n_589)
);

BUFx2_ASAP7_75t_L g590 ( 
.A(n_525),
.Y(n_590)
);

OR2x6_ASAP7_75t_L g591 ( 
.A(n_531),
.B(n_338),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_475),
.Y(n_592)
);

AOI22xp33_ASAP7_75t_L g593 ( 
.A1(n_528),
.A2(n_347),
.B1(n_354),
.B2(n_343),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_SL g594 ( 
.A(n_546),
.B(n_387),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_540),
.B(n_427),
.Y(n_595)
);

INVx3_ASAP7_75t_L g596 ( 
.A(n_475),
.Y(n_596)
);

OR2x6_ASAP7_75t_L g597 ( 
.A(n_531),
.B(n_338),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_502),
.Y(n_598)
);

INVx1_ASAP7_75t_SL g599 ( 
.A(n_546),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_494),
.Y(n_600)
);

INVx5_ASAP7_75t_L g601 ( 
.A(n_475),
.Y(n_601)
);

AOI22xp33_ASAP7_75t_L g602 ( 
.A1(n_528),
.A2(n_357),
.B1(n_354),
.B2(n_343),
.Y(n_602)
);

OR2x2_ASAP7_75t_L g603 ( 
.A(n_529),
.B(n_381),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_528),
.B(n_431),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_540),
.B(n_431),
.Y(n_605)
);

INVx1_ASAP7_75t_SL g606 ( 
.A(n_505),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_502),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_494),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_494),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_540),
.B(n_433),
.Y(n_610)
);

BUFx2_ASAP7_75t_L g611 ( 
.A(n_525),
.Y(n_611)
);

OR2x6_ASAP7_75t_L g612 ( 
.A(n_535),
.B(n_342),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_544),
.B(n_444),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_528),
.B(n_433),
.Y(n_614)
);

BUFx4f_ASAP7_75t_L g615 ( 
.A(n_540),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_476),
.B(n_438),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_540),
.B(n_438),
.Y(n_617)
);

AND2x2_ASAP7_75t_L g618 ( 
.A(n_524),
.B(n_441),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_524),
.B(n_441),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_502),
.Y(n_620)
);

NAND3xp33_ASAP7_75t_L g621 ( 
.A(n_496),
.B(n_356),
.C(n_342),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_495),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_503),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_503),
.Y(n_624)
);

NAND2xp33_ASAP7_75t_L g625 ( 
.A(n_535),
.B(n_442),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_503),
.Y(n_626)
);

BUFx8_ASAP7_75t_SL g627 ( 
.A(n_541),
.Y(n_627)
);

AND2x4_ASAP7_75t_L g628 ( 
.A(n_479),
.B(n_490),
.Y(n_628)
);

INVx3_ASAP7_75t_L g629 ( 
.A(n_475),
.Y(n_629)
);

NAND2xp33_ASAP7_75t_L g630 ( 
.A(n_535),
.B(n_474),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_535),
.B(n_442),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_543),
.B(n_445),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_543),
.B(n_445),
.Y(n_633)
);

BUFx6f_ASAP7_75t_L g634 ( 
.A(n_475),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_552),
.B(n_458),
.Y(n_635)
);

AND2x6_ASAP7_75t_L g636 ( 
.A(n_533),
.B(n_280),
.Y(n_636)
);

INVx3_ASAP7_75t_L g637 ( 
.A(n_475),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_503),
.Y(n_638)
);

INVx4_ASAP7_75t_L g639 ( 
.A(n_497),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_495),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_510),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_543),
.B(n_447),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_543),
.B(n_447),
.Y(n_643)
);

INVx3_ASAP7_75t_L g644 ( 
.A(n_475),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_510),
.Y(n_645)
);

BUFx3_ASAP7_75t_L g646 ( 
.A(n_479),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_495),
.Y(n_647)
);

INVx3_ASAP7_75t_L g648 ( 
.A(n_481),
.Y(n_648)
);

INVx2_ASAP7_75t_SL g649 ( 
.A(n_554),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_510),
.Y(n_650)
);

AND2x6_ASAP7_75t_L g651 ( 
.A(n_533),
.B(n_280),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_476),
.B(n_449),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_490),
.B(n_449),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_510),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_511),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_511),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_511),
.Y(n_657)
);

AND2x6_ASAP7_75t_L g658 ( 
.A(n_533),
.B(n_534),
.Y(n_658)
);

BUFx10_ASAP7_75t_L g659 ( 
.A(n_553),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_499),
.Y(n_660)
);

INVx3_ASAP7_75t_L g661 ( 
.A(n_481),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_511),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_515),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_545),
.B(n_453),
.Y(n_664)
);

INVx5_ASAP7_75t_L g665 ( 
.A(n_481),
.Y(n_665)
);

BUFx2_ASAP7_75t_L g666 ( 
.A(n_509),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_515),
.Y(n_667)
);

BUFx3_ASAP7_75t_L g668 ( 
.A(n_479),
.Y(n_668)
);

INVx4_ASAP7_75t_L g669 ( 
.A(n_497),
.Y(n_669)
);

BUFx3_ASAP7_75t_L g670 ( 
.A(n_479),
.Y(n_670)
);

INVx1_ASAP7_75t_SL g671 ( 
.A(n_505),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_545),
.B(n_453),
.Y(n_672)
);

INVx3_ASAP7_75t_L g673 ( 
.A(n_481),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_541),
.B(n_459),
.Y(n_674)
);

BUFx2_ASAP7_75t_L g675 ( 
.A(n_509),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_490),
.B(n_530),
.Y(n_676)
);

AOI22xp5_ASAP7_75t_L g677 ( 
.A1(n_553),
.A2(n_323),
.B1(n_274),
.B2(n_267),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_496),
.B(n_455),
.Y(n_678)
);

BUFx3_ASAP7_75t_L g679 ( 
.A(n_479),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_499),
.Y(n_680)
);

AOI22xp33_ASAP7_75t_SL g681 ( 
.A1(n_512),
.A2(n_392),
.B1(n_408),
.B2(n_416),
.Y(n_681)
);

BUFx4f_ASAP7_75t_L g682 ( 
.A(n_497),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_508),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_515),
.Y(n_684)
);

OR2x6_ASAP7_75t_L g685 ( 
.A(n_545),
.B(n_356),
.Y(n_685)
);

INVx2_ASAP7_75t_SL g686 ( 
.A(n_554),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_545),
.B(n_455),
.Y(n_687)
);

NAND2xp33_ASAP7_75t_SL g688 ( 
.A(n_548),
.B(n_456),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_515),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_548),
.B(n_456),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_548),
.B(n_462),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_498),
.B(n_462),
.Y(n_692)
);

AND2x4_ASAP7_75t_L g693 ( 
.A(n_490),
.B(n_368),
.Y(n_693)
);

AOI22xp33_ASAP7_75t_L g694 ( 
.A1(n_498),
.A2(n_347),
.B1(n_357),
.B2(n_334),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_547),
.B(n_463),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_508),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_517),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_508),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_547),
.B(n_463),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_513),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_513),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_513),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_517),
.Y(n_703)
);

BUFx3_ASAP7_75t_L g704 ( 
.A(n_488),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_585),
.B(n_547),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_616),
.B(n_547),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_585),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_652),
.B(n_550),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_565),
.B(n_615),
.Y(n_709)
);

INVxp67_ASAP7_75t_L g710 ( 
.A(n_599),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_565),
.B(n_615),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_565),
.B(n_550),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_678),
.B(n_550),
.Y(n_713)
);

AOI22xp33_ASAP7_75t_L g714 ( 
.A1(n_621),
.A2(n_536),
.B1(n_527),
.B2(n_532),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_692),
.B(n_550),
.Y(n_715)
);

INVx8_ASAP7_75t_L g716 ( 
.A(n_658),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_676),
.B(n_526),
.Y(n_717)
);

A2O1A1Ixp33_ASAP7_75t_L g718 ( 
.A1(n_649),
.A2(n_554),
.B(n_527),
.C(n_526),
.Y(n_718)
);

INVxp67_ASAP7_75t_L g719 ( 
.A(n_666),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_646),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_704),
.B(n_530),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_573),
.B(n_549),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_646),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_704),
.B(n_530),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_575),
.B(n_549),
.Y(n_725)
);

OAI22xp5_ASAP7_75t_L g726 ( 
.A1(n_649),
.A2(n_686),
.B1(n_580),
.B2(n_614),
.Y(n_726)
);

INVx2_ASAP7_75t_SL g727 ( 
.A(n_603),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_704),
.B(n_530),
.Y(n_728)
);

NAND2xp33_ASAP7_75t_L g729 ( 
.A(n_636),
.B(n_549),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_556),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_569),
.B(n_530),
.Y(n_731)
);

CKINVDCx20_ASAP7_75t_R g732 ( 
.A(n_560),
.Y(n_732)
);

INVx3_ASAP7_75t_L g733 ( 
.A(n_646),
.Y(n_733)
);

AOI22xp33_ASAP7_75t_L g734 ( 
.A1(n_621),
.A2(n_536),
.B1(n_532),
.B2(n_490),
.Y(n_734)
);

NAND2xp33_ASAP7_75t_L g735 ( 
.A(n_636),
.B(n_551),
.Y(n_735)
);

OR2x2_ASAP7_75t_L g736 ( 
.A(n_603),
.B(n_542),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_615),
.B(n_551),
.Y(n_737)
);

AOI22xp5_ASAP7_75t_L g738 ( 
.A1(n_686),
.A2(n_551),
.B1(n_405),
.B2(n_425),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_604),
.B(n_537),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_569),
.B(n_500),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_628),
.B(n_215),
.Y(n_741)
);

O2A1O1Ixp33_ASAP7_75t_L g742 ( 
.A1(n_555),
.A2(n_489),
.B(n_492),
.C(n_491),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_584),
.B(n_500),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_567),
.Y(n_744)
);

OR2x2_ASAP7_75t_L g745 ( 
.A(n_606),
.B(n_542),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_628),
.B(n_215),
.Y(n_746)
);

BUFx6f_ASAP7_75t_L g747 ( 
.A(n_668),
.Y(n_747)
);

INVx4_ASAP7_75t_L g748 ( 
.A(n_574),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_557),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_584),
.B(n_500),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_586),
.B(n_500),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_586),
.B(n_500),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_600),
.B(n_514),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_628),
.B(n_562),
.Y(n_754)
);

BUFx6f_ASAP7_75t_L g755 ( 
.A(n_668),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_600),
.B(n_514),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_608),
.B(n_514),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_608),
.B(n_514),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_668),
.Y(n_759)
);

INVxp33_ASAP7_75t_L g760 ( 
.A(n_594),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_628),
.B(n_215),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_609),
.B(n_514),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_609),
.B(n_519),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_560),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_562),
.B(n_215),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_567),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_579),
.B(n_217),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_581),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_622),
.B(n_519),
.Y(n_769)
);

OAI22xp33_ASAP7_75t_L g770 ( 
.A1(n_612),
.A2(n_537),
.B1(n_542),
.B2(n_470),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_579),
.B(n_217),
.Y(n_771)
);

AND2x2_ASAP7_75t_L g772 ( 
.A(n_618),
.B(n_619),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_690),
.B(n_691),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_618),
.B(n_537),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_622),
.B(n_519),
.Y(n_775)
);

BUFx12f_ASAP7_75t_L g776 ( 
.A(n_666),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_670),
.Y(n_777)
);

AOI22xp33_ASAP7_75t_L g778 ( 
.A1(n_555),
.A2(n_536),
.B1(n_532),
.B2(n_490),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_670),
.Y(n_779)
);

AND2x4_ASAP7_75t_L g780 ( 
.A(n_590),
.B(n_532),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_670),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_581),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_679),
.B(n_217),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_583),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_L g785 ( 
.A(n_570),
.B(n_465),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_SL g786 ( 
.A(n_674),
.B(n_385),
.Y(n_786)
);

BUFx6f_ASAP7_75t_SL g787 ( 
.A(n_659),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_640),
.B(n_519),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_583),
.Y(n_789)
);

BUFx6f_ASAP7_75t_L g790 ( 
.A(n_679),
.Y(n_790)
);

AND2x4_ASAP7_75t_L g791 ( 
.A(n_590),
.B(n_532),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_640),
.B(n_519),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_567),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_679),
.B(n_217),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_647),
.B(n_497),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_568),
.B(n_217),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_587),
.Y(n_797)
);

INVx4_ASAP7_75t_L g798 ( 
.A(n_574),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_568),
.Y(n_799)
);

BUFx3_ASAP7_75t_L g800 ( 
.A(n_574),
.Y(n_800)
);

AND2x2_ASAP7_75t_L g801 ( 
.A(n_675),
.B(n_538),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_587),
.Y(n_802)
);

AOI22xp5_ASAP7_75t_L g803 ( 
.A1(n_613),
.A2(n_538),
.B1(n_534),
.B2(n_532),
.Y(n_803)
);

BUFx6f_ASAP7_75t_L g804 ( 
.A(n_588),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_660),
.Y(n_805)
);

BUFx2_ASAP7_75t_L g806 ( 
.A(n_675),
.Y(n_806)
);

OAI22xp5_ASAP7_75t_L g807 ( 
.A1(n_612),
.A2(n_534),
.B1(n_344),
.B2(n_372),
.Y(n_807)
);

INVxp67_ASAP7_75t_SL g808 ( 
.A(n_568),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_660),
.B(n_497),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_SL g810 ( 
.A(n_653),
.B(n_276),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_631),
.B(n_632),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_680),
.B(n_683),
.Y(n_812)
);

NAND2xp33_ASAP7_75t_L g813 ( 
.A(n_636),
.B(n_223),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_598),
.Y(n_814)
);

AOI22xp5_ASAP7_75t_L g815 ( 
.A1(n_635),
.A2(n_539),
.B1(n_465),
.B2(n_374),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_653),
.B(n_276),
.Y(n_816)
);

OAI22xp5_ASAP7_75t_L g817 ( 
.A1(n_612),
.A2(n_344),
.B1(n_372),
.B2(n_373),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_683),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_633),
.B(n_642),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_696),
.Y(n_820)
);

BUFx2_ASAP7_75t_L g821 ( 
.A(n_688),
.Y(n_821)
);

BUFx6f_ASAP7_75t_L g822 ( 
.A(n_588),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_696),
.Y(n_823)
);

INVxp67_ASAP7_75t_L g824 ( 
.A(n_643),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_698),
.Y(n_825)
);

BUFx6f_ASAP7_75t_L g826 ( 
.A(n_588),
.Y(n_826)
);

INVx8_ASAP7_75t_L g827 ( 
.A(n_658),
.Y(n_827)
);

NOR2xp67_ASAP7_75t_SL g828 ( 
.A(n_558),
.B(n_559),
.Y(n_828)
);

NAND2xp33_ASAP7_75t_L g829 ( 
.A(n_636),
.B(n_224),
.Y(n_829)
);

OR2x2_ASAP7_75t_L g830 ( 
.A(n_671),
.B(n_505),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_700),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_L g832 ( 
.A(n_664),
.B(n_539),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_589),
.B(n_276),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_700),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_SL g835 ( 
.A(n_659),
.B(n_512),
.Y(n_835)
);

INVx2_ASAP7_75t_SL g836 ( 
.A(n_693),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_701),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_595),
.B(n_276),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_672),
.B(n_539),
.Y(n_839)
);

HB1xp67_ASAP7_75t_L g840 ( 
.A(n_611),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_701),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_SL g842 ( 
.A(n_659),
.B(n_307),
.Y(n_842)
);

AOI22xp33_ASAP7_75t_L g843 ( 
.A1(n_558),
.A2(n_290),
.B1(n_370),
.B2(n_210),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_598),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_702),
.B(n_517),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_702),
.B(n_517),
.Y(n_846)
);

AOI22xp33_ASAP7_75t_L g847 ( 
.A1(n_559),
.A2(n_290),
.B1(n_370),
.B2(n_240),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_566),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_566),
.B(n_518),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_588),
.Y(n_850)
);

BUFx6f_ASAP7_75t_L g851 ( 
.A(n_634),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_693),
.B(n_612),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_687),
.B(n_539),
.Y(n_853)
);

BUFx8_ASAP7_75t_L g854 ( 
.A(n_611),
.Y(n_854)
);

INVxp67_ASAP7_75t_L g855 ( 
.A(n_695),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_L g856 ( 
.A(n_699),
.B(n_539),
.Y(n_856)
);

AO22x2_ASAP7_75t_L g857 ( 
.A1(n_693),
.A2(n_368),
.B1(n_240),
.B2(n_246),
.Y(n_857)
);

INVx2_ASAP7_75t_SL g858 ( 
.A(n_693),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_607),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_605),
.B(n_276),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_620),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_612),
.B(n_518),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_659),
.B(n_488),
.Y(n_863)
);

INVx1_ASAP7_75t_SL g864 ( 
.A(n_627),
.Y(n_864)
);

A2O1A1Ixp33_ASAP7_75t_L g865 ( 
.A1(n_706),
.A2(n_630),
.B(n_625),
.C(n_610),
.Y(n_865)
);

CKINVDCx8_ASAP7_75t_R g866 ( 
.A(n_764),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_706),
.B(n_617),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_708),
.B(n_722),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_708),
.B(n_685),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_709),
.A2(n_682),
.B(n_639),
.Y(n_870)
);

OAI21xp5_ASAP7_75t_L g871 ( 
.A1(n_796),
.A2(n_682),
.B(n_561),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_709),
.A2(n_682),
.B(n_639),
.Y(n_872)
);

OAI22x1_ASAP7_75t_L g873 ( 
.A1(n_773),
.A2(n_677),
.B1(n_738),
.B2(n_806),
.Y(n_873)
);

OAI21xp5_ASAP7_75t_L g874 ( 
.A1(n_796),
.A2(n_685),
.B(n_658),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_722),
.B(n_685),
.Y(n_875)
);

CKINVDCx6p67_ASAP7_75t_R g876 ( 
.A(n_732),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_725),
.B(n_685),
.Y(n_877)
);

OAI21xp33_ASAP7_75t_L g878 ( 
.A1(n_785),
.A2(n_677),
.B(n_694),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_820),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_725),
.B(n_685),
.Y(n_880)
);

AO21x1_ASAP7_75t_L g881 ( 
.A1(n_773),
.A2(n_577),
.B(n_378),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_L g882 ( 
.A(n_713),
.B(n_578),
.Y(n_882)
);

NOR3xp33_ASAP7_75t_L g883 ( 
.A(n_785),
.B(n_770),
.C(n_772),
.Y(n_883)
);

AOI22xp5_ASAP7_75t_L g884 ( 
.A1(n_811),
.A2(n_658),
.B1(n_578),
.B2(n_591),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_715),
.B(n_658),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_808),
.B(n_658),
.Y(n_886)
);

NOR2x1_ASAP7_75t_L g887 ( 
.A(n_863),
.B(n_578),
.Y(n_887)
);

HB1xp67_ASAP7_75t_L g888 ( 
.A(n_840),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_711),
.A2(n_639),
.B(n_572),
.Y(n_889)
);

INVxp67_ASAP7_75t_L g890 ( 
.A(n_801),
.Y(n_890)
);

INVx3_ASAP7_75t_L g891 ( 
.A(n_747),
.Y(n_891)
);

AOI22xp5_ASAP7_75t_L g892 ( 
.A1(n_811),
.A2(n_819),
.B1(n_726),
.B2(n_754),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_711),
.A2(n_639),
.B(n_572),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_717),
.A2(n_705),
.B(n_849),
.Y(n_894)
);

O2A1O1Ixp33_ASAP7_75t_L g895 ( 
.A1(n_718),
.A2(n_582),
.B(n_591),
.C(n_578),
.Y(n_895)
);

AO21x1_ASAP7_75t_L g896 ( 
.A1(n_737),
.A2(n_378),
.B(n_373),
.Y(n_896)
);

INVx1_ASAP7_75t_SL g897 ( 
.A(n_745),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_739),
.B(n_658),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_739),
.B(n_564),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_712),
.A2(n_669),
.B(n_572),
.Y(n_900)
);

CKINVDCx20_ASAP7_75t_R g901 ( 
.A(n_854),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_774),
.B(n_681),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_SL g903 ( 
.A(n_819),
.B(n_634),
.Y(n_903)
);

NOR2x1_ASAP7_75t_L g904 ( 
.A(n_800),
.B(n_578),
.Y(n_904)
);

A2O1A1Ixp33_ASAP7_75t_L g905 ( 
.A1(n_832),
.A2(n_563),
.B(n_602),
.C(n_593),
.Y(n_905)
);

OAI22xp5_ASAP7_75t_L g906 ( 
.A1(n_778),
.A2(n_591),
.B1(n_597),
.B2(n_582),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_823),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_721),
.A2(n_669),
.B(n_634),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_823),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_724),
.A2(n_669),
.B(n_634),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_707),
.B(n_564),
.Y(n_911)
);

A2O1A1Ixp33_ASAP7_75t_L g912 ( 
.A1(n_832),
.A2(n_623),
.B(n_624),
.C(n_620),
.Y(n_912)
);

INVx3_ASAP7_75t_L g913 ( 
.A(n_747),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_744),
.B(n_564),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_728),
.A2(n_634),
.B(n_592),
.Y(n_915)
);

O2A1O1Ixp33_ASAP7_75t_SL g916 ( 
.A1(n_737),
.A2(n_592),
.B(n_571),
.C(n_352),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_SL g917 ( 
.A(n_747),
.B(n_755),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_744),
.B(n_564),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_766),
.B(n_636),
.Y(n_919)
);

AND2x2_ASAP7_75t_L g920 ( 
.A(n_727),
.B(n_489),
.Y(n_920)
);

OAI21xp5_ASAP7_75t_L g921 ( 
.A1(n_766),
.A2(n_571),
.B(n_623),
.Y(n_921)
);

O2A1O1Ixp33_ASAP7_75t_L g922 ( 
.A1(n_754),
.A2(n_591),
.B(n_597),
.C(n_582),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_793),
.B(n_636),
.Y(n_923)
);

OAI21xp33_ASAP7_75t_SL g924 ( 
.A1(n_778),
.A2(n_591),
.B(n_582),
.Y(n_924)
);

A2O1A1Ixp33_ASAP7_75t_L g925 ( 
.A1(n_839),
.A2(n_703),
.B(n_697),
.C(n_689),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_793),
.B(n_636),
.Y(n_926)
);

AOI22xp5_ASAP7_75t_L g927 ( 
.A1(n_839),
.A2(n_597),
.B1(n_651),
.B2(n_689),
.Y(n_927)
);

NOR2xp33_ASAP7_75t_L g928 ( 
.A(n_824),
.B(n_597),
.Y(n_928)
);

INVx3_ASAP7_75t_L g929 ( 
.A(n_747),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_SL g930 ( 
.A(n_755),
.B(n_576),
.Y(n_930)
);

O2A1O1Ixp33_ASAP7_75t_SL g931 ( 
.A1(n_833),
.A2(n_703),
.B(n_697),
.C(n_684),
.Y(n_931)
);

BUFx6f_ASAP7_75t_L g932 ( 
.A(n_851),
.Y(n_932)
);

AOI21xp33_ASAP7_75t_L g933 ( 
.A1(n_815),
.A2(n_204),
.B(n_189),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_L g934 ( 
.A(n_855),
.B(n_212),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_719),
.B(n_319),
.Y(n_935)
);

INVx3_ASAP7_75t_L g936 ( 
.A(n_755),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_799),
.B(n_651),
.Y(n_937)
);

INVxp67_ASAP7_75t_L g938 ( 
.A(n_736),
.Y(n_938)
);

AND2x4_ASAP7_75t_L g939 ( 
.A(n_780),
.B(n_791),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_SL g940 ( 
.A(n_780),
.B(n_491),
.Y(n_940)
);

OAI21xp5_ASAP7_75t_L g941 ( 
.A1(n_799),
.A2(n_626),
.B(n_624),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_805),
.Y(n_942)
);

OAI22xp5_ASAP7_75t_L g943 ( 
.A1(n_803),
.A2(n_684),
.B1(n_626),
.B2(n_667),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_848),
.B(n_651),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_848),
.B(n_651),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_710),
.B(n_492),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_714),
.B(n_818),
.Y(n_947)
);

INVx2_ASAP7_75t_SL g948 ( 
.A(n_776),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_714),
.B(n_651),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_825),
.Y(n_950)
);

NOR2x1p5_ASAP7_75t_L g951 ( 
.A(n_830),
.B(n_309),
.Y(n_951)
);

NOR2xp67_ASAP7_75t_L g952 ( 
.A(n_853),
.B(n_520),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_731),
.A2(n_665),
.B(n_601),
.Y(n_953)
);

INVx2_ASAP7_75t_SL g954 ( 
.A(n_854),
.Y(n_954)
);

BUFx3_ASAP7_75t_L g955 ( 
.A(n_791),
.Y(n_955)
);

OAI22xp5_ASAP7_75t_L g956 ( 
.A1(n_853),
.A2(n_650),
.B1(n_667),
.B2(n_663),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_L g957 ( 
.A(n_760),
.B(n_520),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_831),
.B(n_651),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_834),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_837),
.B(n_651),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_SL g961 ( 
.A(n_755),
.B(n_576),
.Y(n_961)
);

OAI21xp5_ASAP7_75t_L g962 ( 
.A1(n_740),
.A2(n_641),
.B(n_638),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_841),
.B(n_673),
.Y(n_963)
);

CKINVDCx14_ASAP7_75t_R g964 ( 
.A(n_821),
.Y(n_964)
);

OAI21xp33_ASAP7_75t_L g965 ( 
.A1(n_842),
.A2(n_835),
.B(n_786),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_852),
.A2(n_665),
.B(n_601),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_856),
.B(n_673),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_720),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_723),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_861),
.Y(n_970)
);

OAI21xp5_ASAP7_75t_L g971 ( 
.A1(n_743),
.A2(n_641),
.B(n_638),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_851),
.A2(n_665),
.B(n_601),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_851),
.A2(n_673),
.B(n_596),
.Y(n_973)
);

AOI22xp33_ASAP7_75t_L g974 ( 
.A1(n_843),
.A2(n_847),
.B1(n_857),
.B2(n_817),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_759),
.Y(n_975)
);

NOR2x1_ASAP7_75t_L g976 ( 
.A(n_800),
.B(n_645),
.Y(n_976)
);

OAI21xp5_ASAP7_75t_L g977 ( 
.A1(n_750),
.A2(n_752),
.B(n_751),
.Y(n_977)
);

OAI22xp5_ASAP7_75t_L g978 ( 
.A1(n_856),
.A2(n_650),
.B1(n_663),
.B2(n_662),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_734),
.B(n_673),
.Y(n_979)
);

OAI21xp5_ASAP7_75t_L g980 ( 
.A1(n_753),
.A2(n_654),
.B(n_645),
.Y(n_980)
);

BUFx4f_ASAP7_75t_L g981 ( 
.A(n_790),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_734),
.B(n_576),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_812),
.B(n_576),
.Y(n_983)
);

OAI21xp5_ASAP7_75t_L g984 ( 
.A1(n_756),
.A2(n_655),
.B(n_654),
.Y(n_984)
);

NOR2xp33_ASAP7_75t_L g985 ( 
.A(n_777),
.B(n_311),
.Y(n_985)
);

OAI22xp5_ASAP7_75t_L g986 ( 
.A1(n_836),
.A2(n_662),
.B1(n_655),
.B2(n_657),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_779),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_765),
.B(n_596),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_729),
.A2(n_629),
.B(n_596),
.Y(n_989)
);

BUFx6f_ASAP7_75t_L g990 ( 
.A(n_790),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_857),
.B(n_340),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_767),
.B(n_771),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_767),
.B(n_661),
.Y(n_993)
);

AO21x1_ASAP7_75t_L g994 ( 
.A1(n_833),
.A2(n_657),
.B(n_656),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_735),
.A2(n_637),
.B(n_629),
.Y(n_995)
);

AOI21x1_ASAP7_75t_L g996 ( 
.A1(n_828),
.A2(n_656),
.B(n_486),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_771),
.B(n_661),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_733),
.B(n_661),
.Y(n_998)
);

OAI21xp33_ASAP7_75t_L g999 ( 
.A1(n_843),
.A2(n_316),
.B(n_313),
.Y(n_999)
);

OAI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_757),
.A2(n_762),
.B(n_758),
.Y(n_1000)
);

OAI22xp5_ASAP7_75t_L g1001 ( 
.A1(n_858),
.A2(n_661),
.B1(n_648),
.B2(n_644),
.Y(n_1001)
);

AND2x4_ASAP7_75t_L g1002 ( 
.A(n_790),
.B(n_246),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_781),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_733),
.B(n_648),
.Y(n_1004)
);

INVxp67_ASAP7_75t_L g1005 ( 
.A(n_810),
.Y(n_1005)
);

INVx4_ASAP7_75t_L g1006 ( 
.A(n_790),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_741),
.A2(n_648),
.B(n_637),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_741),
.A2(n_648),
.B(n_637),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_SL g1009 ( 
.A(n_804),
.B(n_629),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_847),
.B(n_629),
.Y(n_1010)
);

NOR3xp33_ASAP7_75t_L g1011 ( 
.A(n_810),
.B(n_504),
.C(n_501),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_859),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_SL g1013 ( 
.A(n_804),
.B(n_637),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_L g1014 ( 
.A(n_816),
.B(n_320),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_742),
.B(n_644),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_748),
.B(n_644),
.Y(n_1016)
);

OAI21xp33_ASAP7_75t_L g1017 ( 
.A1(n_816),
.A2(n_329),
.B(n_322),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_845),
.Y(n_1018)
);

AND2x2_ASAP7_75t_L g1019 ( 
.A(n_857),
.B(n_340),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_746),
.A2(n_644),
.B(n_481),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_SL g1021 ( 
.A(n_804),
.B(n_225),
.Y(n_1021)
);

OR2x6_ASAP7_75t_L g1022 ( 
.A(n_716),
.B(n_247),
.Y(n_1022)
);

OAI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_763),
.A2(n_486),
.B(n_483),
.Y(n_1023)
);

O2A1O1Ixp33_ASAP7_75t_L g1024 ( 
.A1(n_746),
.A2(n_516),
.B(n_507),
.C(n_504),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_748),
.B(n_521),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_804),
.B(n_231),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_SL g1027 ( 
.A(n_822),
.B(n_232),
.Y(n_1027)
);

NOR2x1_ASAP7_75t_L g1028 ( 
.A(n_798),
.B(n_850),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_SL g1029 ( 
.A(n_822),
.B(n_233),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_SL g1030 ( 
.A(n_822),
.B(n_236),
.Y(n_1030)
);

AND2x2_ASAP7_75t_SL g1031 ( 
.A(n_798),
.B(n_247),
.Y(n_1031)
);

OAI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_769),
.A2(n_483),
.B(n_521),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_775),
.B(n_521),
.Y(n_1033)
);

AOI22xp5_ASAP7_75t_L g1034 ( 
.A1(n_838),
.A2(n_281),
.B1(n_375),
.B2(n_371),
.Y(n_1034)
);

NOR2xp33_ASAP7_75t_SL g1035 ( 
.A(n_864),
.B(n_307),
.Y(n_1035)
);

NAND2x1_ASAP7_75t_L g1036 ( 
.A(n_730),
.B(n_481),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_788),
.B(n_521),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_761),
.A2(n_481),
.B(n_478),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_792),
.B(n_522),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_716),
.A2(n_481),
.B(n_478),
.Y(n_1040)
);

AOI22xp33_ASAP7_75t_L g1041 ( 
.A1(n_838),
.A2(n_860),
.B1(n_862),
.B2(n_288),
.Y(n_1041)
);

AO21x1_ASAP7_75t_L g1042 ( 
.A1(n_860),
.A2(n_360),
.B(n_288),
.Y(n_1042)
);

AND2x2_ASAP7_75t_L g1043 ( 
.A(n_783),
.B(n_192),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_868),
.B(n_846),
.Y(n_1044)
);

HB1xp67_ASAP7_75t_L g1045 ( 
.A(n_888),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_SL g1046 ( 
.A(n_939),
.B(n_822),
.Y(n_1046)
);

OAI21xp33_ASAP7_75t_L g1047 ( 
.A1(n_934),
.A2(n_335),
.B(n_331),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_1018),
.B(n_749),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_867),
.B(n_826),
.Y(n_1049)
);

O2A1O1Ixp33_ASAP7_75t_L g1050 ( 
.A1(n_878),
.A2(n_807),
.B(n_794),
.C(n_783),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_886),
.A2(n_827),
.B(n_716),
.Y(n_1051)
);

AOI22xp5_ASAP7_75t_L g1052 ( 
.A1(n_965),
.A2(n_787),
.B1(n_826),
.B2(n_829),
.Y(n_1052)
);

NOR2xp33_ASAP7_75t_SL g1053 ( 
.A(n_866),
.B(n_787),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_879),
.Y(n_1054)
);

BUFx2_ASAP7_75t_L g1055 ( 
.A(n_888),
.Y(n_1055)
);

BUFx6f_ASAP7_75t_L g1056 ( 
.A(n_932),
.Y(n_1056)
);

OR2x2_ASAP7_75t_L g1057 ( 
.A(n_897),
.B(n_794),
.Y(n_1057)
);

OAI22xp5_ASAP7_75t_L g1058 ( 
.A1(n_974),
.A2(n_892),
.B1(n_875),
.B2(n_880),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_877),
.B(n_826),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_894),
.A2(n_827),
.B(n_813),
.Y(n_1060)
);

NOR2xp33_ASAP7_75t_SL g1061 ( 
.A(n_1031),
.B(n_827),
.Y(n_1061)
);

AOI22xp5_ASAP7_75t_L g1062 ( 
.A1(n_883),
.A2(n_826),
.B1(n_327),
.B2(n_324),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_967),
.A2(n_809),
.B(n_795),
.Y(n_1063)
);

INVx3_ASAP7_75t_L g1064 ( 
.A(n_990),
.Y(n_1064)
);

BUFx6f_ASAP7_75t_L g1065 ( 
.A(n_932),
.Y(n_1065)
);

AOI22xp5_ASAP7_75t_L g1066 ( 
.A1(n_902),
.A2(n_273),
.B1(n_365),
.B2(n_362),
.Y(n_1066)
);

AND2x2_ASAP7_75t_L g1067 ( 
.A(n_946),
.B(n_192),
.Y(n_1067)
);

NOR2xp33_ASAP7_75t_R g1068 ( 
.A(n_964),
.B(n_241),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_SL g1069 ( 
.A(n_939),
.B(n_768),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_907),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_885),
.A2(n_844),
.B(n_814),
.Y(n_1071)
);

OR2x2_ASAP7_75t_L g1072 ( 
.A(n_890),
.B(n_782),
.Y(n_1072)
);

O2A1O1Ixp33_ASAP7_75t_L g1073 ( 
.A1(n_865),
.A2(n_360),
.B(n_261),
.C(n_294),
.Y(n_1073)
);

OAI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_924),
.A2(n_802),
.B(n_797),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_909),
.Y(n_1075)
);

O2A1O1Ixp33_ASAP7_75t_L g1076 ( 
.A1(n_933),
.A2(n_261),
.B(n_294),
.C(n_304),
.Y(n_1076)
);

OAI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_974),
.A2(n_304),
.B1(n_308),
.B2(n_317),
.Y(n_1077)
);

OAI22xp5_ASAP7_75t_L g1078 ( 
.A1(n_947),
.A2(n_361),
.B1(n_317),
.B2(n_318),
.Y(n_1078)
);

OAI22xp5_ASAP7_75t_L g1079 ( 
.A1(n_899),
.A2(n_361),
.B1(n_318),
.B2(n_334),
.Y(n_1079)
);

AO32x1_ASAP7_75t_L g1080 ( 
.A1(n_943),
.A2(n_308),
.A3(n_784),
.B1(n_789),
.B2(n_522),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_970),
.Y(n_1081)
);

A2O1A1Ixp33_ASAP7_75t_SL g1082 ( 
.A1(n_882),
.A2(n_523),
.B(n_522),
.C(n_516),
.Y(n_1082)
);

BUFx6f_ASAP7_75t_L g1083 ( 
.A(n_932),
.Y(n_1083)
);

A2O1A1Ixp33_ASAP7_75t_L g1084 ( 
.A1(n_928),
.A2(n_1014),
.B(n_882),
.C(n_895),
.Y(n_1084)
);

INVxp67_ASAP7_75t_L g1085 ( 
.A(n_934),
.Y(n_1085)
);

INVx4_ASAP7_75t_L g1086 ( 
.A(n_981),
.Y(n_1086)
);

AND2x2_ASAP7_75t_L g1087 ( 
.A(n_938),
.B(n_192),
.Y(n_1087)
);

NOR2xp33_ASAP7_75t_L g1088 ( 
.A(n_938),
.B(n_336),
.Y(n_1088)
);

OAI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_949),
.A2(n_523),
.B(n_522),
.Y(n_1089)
);

OR2x2_ASAP7_75t_L g1090 ( 
.A(n_935),
.B(n_957),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_1012),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_942),
.Y(n_1092)
);

CKINVDCx14_ASAP7_75t_R g1093 ( 
.A(n_876),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_908),
.A2(n_478),
.B(n_483),
.Y(n_1094)
);

OAI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_905),
.A2(n_337),
.B1(n_339),
.B2(n_341),
.Y(n_1095)
);

O2A1O1Ixp33_ASAP7_75t_L g1096 ( 
.A1(n_957),
.A2(n_523),
.B(n_485),
.C(n_480),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_869),
.B(n_523),
.Y(n_1097)
);

OAI22xp5_ASAP7_75t_SL g1098 ( 
.A1(n_901),
.A2(n_358),
.B1(n_345),
.B2(n_346),
.Y(n_1098)
);

OAI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_979),
.A2(n_485),
.B(n_480),
.Y(n_1099)
);

AO22x1_ASAP7_75t_L g1100 ( 
.A1(n_991),
.A2(n_364),
.B1(n_348),
.B2(n_350),
.Y(n_1100)
);

OAI22xp5_ASAP7_75t_L g1101 ( 
.A1(n_1031),
.A2(n_351),
.B1(n_366),
.B2(n_367),
.Y(n_1101)
);

BUFx2_ASAP7_75t_L g1102 ( 
.A(n_1002),
.Y(n_1102)
);

HB1xp67_ASAP7_75t_L g1103 ( 
.A(n_1002),
.Y(n_1103)
);

AND2x2_ASAP7_75t_L g1104 ( 
.A(n_920),
.B(n_192),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_SL g1105 ( 
.A(n_955),
.B(n_250),
.Y(n_1105)
);

A2O1A1Ixp33_ASAP7_75t_L g1106 ( 
.A1(n_928),
.A2(n_253),
.B(n_259),
.C(n_264),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_SL g1107 ( 
.A(n_981),
.B(n_266),
.Y(n_1107)
);

HB1xp67_ASAP7_75t_L g1108 ( 
.A(n_873),
.Y(n_1108)
);

INVx2_ASAP7_75t_SL g1109 ( 
.A(n_951),
.Y(n_1109)
);

AND2x2_ASAP7_75t_SL g1110 ( 
.A(n_1019),
.B(n_307),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_910),
.A2(n_898),
.B(n_874),
.Y(n_1111)
);

AOI21xp33_ASAP7_75t_L g1112 ( 
.A1(n_1014),
.A2(n_369),
.B(n_376),
.Y(n_1112)
);

BUFx6f_ASAP7_75t_L g1113 ( 
.A(n_932),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_983),
.A2(n_478),
.B(n_483),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_950),
.B(n_477),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_959),
.B(n_477),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_SL g1117 ( 
.A(n_990),
.B(n_272),
.Y(n_1117)
);

BUFx6f_ASAP7_75t_SL g1118 ( 
.A(n_954),
.Y(n_1118)
);

BUFx6f_ASAP7_75t_L g1119 ( 
.A(n_990),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_968),
.Y(n_1120)
);

O2A1O1Ixp33_ASAP7_75t_L g1121 ( 
.A1(n_1005),
.A2(n_485),
.B(n_480),
.C(n_477),
.Y(n_1121)
);

OAI22xp5_ASAP7_75t_L g1122 ( 
.A1(n_911),
.A2(n_377),
.B1(n_379),
.B2(n_312),
.Y(n_1122)
);

BUFx6f_ASAP7_75t_L g1123 ( 
.A(n_990),
.Y(n_1123)
);

BUFx6f_ASAP7_75t_L g1124 ( 
.A(n_891),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_987),
.Y(n_1125)
);

INVx4_ASAP7_75t_L g1126 ( 
.A(n_1006),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_1005),
.B(n_282),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_SL g1128 ( 
.A(n_887),
.B(n_283),
.Y(n_1128)
);

BUFx2_ASAP7_75t_L g1129 ( 
.A(n_1022),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_969),
.B(n_284),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_975),
.B(n_287),
.Y(n_1131)
);

AOI22xp33_ASAP7_75t_L g1132 ( 
.A1(n_881),
.A2(n_292),
.B1(n_349),
.B2(n_305),
.Y(n_1132)
);

BUFx4f_ASAP7_75t_L g1133 ( 
.A(n_948),
.Y(n_1133)
);

OAI22xp5_ASAP7_75t_SL g1134 ( 
.A1(n_935),
.A2(n_314),
.B1(n_296),
.B2(n_297),
.Y(n_1134)
);

AO21x1_ASAP7_75t_L g1135 ( 
.A1(n_903),
.A2(n_871),
.B(n_922),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_1016),
.A2(n_478),
.B(n_332),
.Y(n_1136)
);

BUFx2_ASAP7_75t_L g1137 ( 
.A(n_1022),
.Y(n_1137)
);

AOI21x1_ASAP7_75t_L g1138 ( 
.A1(n_903),
.A2(n_300),
.B(n_330),
.Y(n_1138)
);

AO32x1_ASAP7_75t_L g1139 ( 
.A1(n_956),
.A2(n_292),
.A3(n_333),
.B1(n_26),
.B2(n_27),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1003),
.Y(n_1140)
);

BUFx6f_ASAP7_75t_L g1141 ( 
.A(n_913),
.Y(n_1141)
);

BUFx12f_ASAP7_75t_L g1142 ( 
.A(n_1022),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_913),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_985),
.B(n_292),
.Y(n_1144)
);

INVx3_ASAP7_75t_L g1145 ( 
.A(n_1006),
.Y(n_1145)
);

OAI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_982),
.A2(n_925),
.B(n_912),
.Y(n_1146)
);

O2A1O1Ixp5_ASAP7_75t_L g1147 ( 
.A1(n_896),
.A2(n_78),
.B(n_185),
.C(n_184),
.Y(n_1147)
);

INVx2_ASAP7_75t_SL g1148 ( 
.A(n_1043),
.Y(n_1148)
);

NAND3xp33_ASAP7_75t_SL g1149 ( 
.A(n_1035),
.B(n_999),
.C(n_1017),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_998),
.A2(n_75),
.B(n_183),
.Y(n_1150)
);

AO22x1_ASAP7_75t_L g1151 ( 
.A1(n_904),
.A2(n_333),
.B1(n_20),
.B2(n_26),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_952),
.B(n_333),
.Y(n_1152)
);

BUFx6f_ASAP7_75t_L g1153 ( 
.A(n_929),
.Y(n_1153)
);

O2A1O1Ixp33_ASAP7_75t_L g1154 ( 
.A1(n_940),
.A2(n_333),
.B(n_20),
.C(n_30),
.Y(n_1154)
);

OAI22xp5_ASAP7_75t_L g1155 ( 
.A1(n_884),
.A2(n_18),
.B1(n_30),
.B2(n_31),
.Y(n_1155)
);

OAI22xp5_ASAP7_75t_L g1156 ( 
.A1(n_1010),
.A2(n_31),
.B1(n_32),
.B2(n_34),
.Y(n_1156)
);

OAI22xp5_ASAP7_75t_L g1157 ( 
.A1(n_914),
.A2(n_34),
.B1(n_36),
.B2(n_40),
.Y(n_1157)
);

AO21x2_ASAP7_75t_L g1158 ( 
.A1(n_916),
.A2(n_92),
.B(n_175),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_936),
.B(n_36),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_936),
.B(n_43),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_918),
.Y(n_1161)
);

AOI22x1_ASAP7_75t_L g1162 ( 
.A1(n_915),
.A2(n_81),
.B1(n_174),
.B2(n_167),
.Y(n_1162)
);

BUFx2_ASAP7_75t_L g1163 ( 
.A(n_1042),
.Y(n_1163)
);

BUFx6f_ASAP7_75t_L g1164 ( 
.A(n_917),
.Y(n_1164)
);

A2O1A1Ixp33_ASAP7_75t_L g1165 ( 
.A1(n_992),
.A2(n_43),
.B(n_44),
.C(n_46),
.Y(n_1165)
);

INVx2_ASAP7_75t_SL g1166 ( 
.A(n_1021),
.Y(n_1166)
);

AOI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_1021),
.A2(n_95),
.B1(n_164),
.B2(n_157),
.Y(n_1167)
);

NOR3xp33_ASAP7_75t_SL g1168 ( 
.A(n_1026),
.B(n_47),
.C(n_51),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1011),
.B(n_51),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_SL g1170 ( 
.A(n_906),
.B(n_93),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1011),
.B(n_53),
.Y(n_1171)
);

BUFx2_ASAP7_75t_L g1172 ( 
.A(n_976),
.Y(n_1172)
);

A2O1A1Ixp33_ASAP7_75t_L g1173 ( 
.A1(n_927),
.A2(n_960),
.B(n_958),
.C(n_1041),
.Y(n_1173)
);

AND2x2_ASAP7_75t_L g1174 ( 
.A(n_1041),
.B(n_55),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_963),
.Y(n_1175)
);

BUFx6f_ASAP7_75t_L g1176 ( 
.A(n_917),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_996),
.Y(n_1177)
);

OAI22x1_ASAP7_75t_L g1178 ( 
.A1(n_1026),
.A2(n_1027),
.B1(n_1030),
.B2(n_1029),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1004),
.A2(n_97),
.B(n_137),
.Y(n_1179)
);

OR2x2_ASAP7_75t_L g1180 ( 
.A(n_1027),
.B(n_55),
.Y(n_1180)
);

HB1xp67_ASAP7_75t_L g1181 ( 
.A(n_1029),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_SL g1182 ( 
.A(n_1034),
.B(n_1030),
.Y(n_1182)
);

OA22x2_ASAP7_75t_L g1183 ( 
.A1(n_1015),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.Y(n_1183)
);

O2A1O1Ixp33_ASAP7_75t_L g1184 ( 
.A1(n_1024),
.A2(n_57),
.B(n_61),
.C(n_62),
.Y(n_1184)
);

O2A1O1Ixp33_ASAP7_75t_L g1185 ( 
.A1(n_1001),
.A2(n_64),
.B(n_70),
.C(n_71),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_930),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_977),
.B(n_99),
.Y(n_1187)
);

AOI22xp33_ASAP7_75t_L g1188 ( 
.A1(n_1028),
.A2(n_101),
.B1(n_105),
.B2(n_107),
.Y(n_1188)
);

BUFx2_ASAP7_75t_L g1189 ( 
.A(n_1025),
.Y(n_1189)
);

O2A1O1Ixp33_ASAP7_75t_L g1190 ( 
.A1(n_986),
.A2(n_111),
.B(n_119),
.C(n_130),
.Y(n_1190)
);

A2O1A1Ixp33_ASAP7_75t_L g1191 ( 
.A1(n_1000),
.A2(n_131),
.B(n_135),
.C(n_181),
.Y(n_1191)
);

O2A1O1Ixp33_ASAP7_75t_L g1192 ( 
.A1(n_931),
.A2(n_1039),
.B(n_1037),
.C(n_1033),
.Y(n_1192)
);

INVx2_ASAP7_75t_L g1193 ( 
.A(n_930),
.Y(n_1193)
);

AOI21x1_ASAP7_75t_L g1194 ( 
.A1(n_1187),
.A2(n_994),
.B(n_978),
.Y(n_1194)
);

NOR2xp33_ASAP7_75t_L g1195 ( 
.A(n_1090),
.B(n_1013),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1048),
.Y(n_1196)
);

AOI21x1_ASAP7_75t_L g1197 ( 
.A1(n_1138),
.A2(n_870),
.B(n_872),
.Y(n_1197)
);

AO31x2_ASAP7_75t_L g1198 ( 
.A1(n_1135),
.A2(n_889),
.A3(n_893),
.B(n_900),
.Y(n_1198)
);

BUFx3_ASAP7_75t_L g1199 ( 
.A(n_1055),
.Y(n_1199)
);

AND2x2_ASAP7_75t_L g1200 ( 
.A(n_1104),
.B(n_961),
.Y(n_1200)
);

A2O1A1Ixp33_ASAP7_75t_L g1201 ( 
.A1(n_1084),
.A2(n_1073),
.B(n_1144),
.C(n_1050),
.Y(n_1201)
);

NAND3xp33_ASAP7_75t_L g1202 ( 
.A(n_1112),
.B(n_1032),
.C(n_1023),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1060),
.A2(n_945),
.B(n_944),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_1091),
.Y(n_1204)
);

AO21x2_ASAP7_75t_L g1205 ( 
.A1(n_1082),
.A2(n_921),
.B(n_980),
.Y(n_1205)
);

AO32x2_ASAP7_75t_L g1206 ( 
.A1(n_1058),
.A2(n_984),
.A3(n_971),
.B1(n_962),
.B2(n_941),
.Y(n_1206)
);

A2O1A1Ixp33_ASAP7_75t_L g1207 ( 
.A1(n_1058),
.A2(n_1008),
.B(n_1007),
.C(n_989),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1111),
.A2(n_919),
.B(n_923),
.Y(n_1208)
);

AO21x2_ASAP7_75t_L g1209 ( 
.A1(n_1146),
.A2(n_995),
.B(n_966),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_1072),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1048),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1044),
.A2(n_926),
.B(n_937),
.Y(n_1212)
);

NOR2xp33_ASAP7_75t_L g1213 ( 
.A(n_1085),
.B(n_1009),
.Y(n_1213)
);

NAND3xp33_ASAP7_75t_L g1214 ( 
.A(n_1108),
.B(n_1013),
.C(n_997),
.Y(n_1214)
);

AOI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1044),
.A2(n_988),
.B(n_993),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_1092),
.Y(n_1216)
);

BUFx6f_ASAP7_75t_L g1217 ( 
.A(n_1056),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1061),
.A2(n_1040),
.B(n_973),
.Y(n_1218)
);

BUFx3_ASAP7_75t_L g1219 ( 
.A(n_1045),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1061),
.A2(n_1051),
.B(n_1063),
.Y(n_1220)
);

AO32x2_ASAP7_75t_L g1221 ( 
.A1(n_1079),
.A2(n_1036),
.A3(n_1020),
.B1(n_1038),
.B2(n_953),
.Y(n_1221)
);

AOI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1097),
.A2(n_972),
.B(n_1192),
.Y(n_1222)
);

CKINVDCx11_ASAP7_75t_R g1223 ( 
.A(n_1142),
.Y(n_1223)
);

O2A1O1Ixp5_ASAP7_75t_L g1224 ( 
.A1(n_1170),
.A2(n_1182),
.B(n_1171),
.C(n_1169),
.Y(n_1224)
);

AOI221x1_ASAP7_75t_L g1225 ( 
.A1(n_1155),
.A2(n_1156),
.B1(n_1157),
.B2(n_1178),
.C(n_1078),
.Y(n_1225)
);

O2A1O1Ixp33_ASAP7_75t_SL g1226 ( 
.A1(n_1191),
.A2(n_1106),
.B(n_1173),
.C(n_1165),
.Y(n_1226)
);

BUFx12f_ASAP7_75t_L g1227 ( 
.A(n_1109),
.Y(n_1227)
);

OR2x2_ASAP7_75t_L g1228 ( 
.A(n_1057),
.B(n_1102),
.Y(n_1228)
);

OA21x2_ASAP7_75t_L g1229 ( 
.A1(n_1146),
.A2(n_1099),
.B(n_1089),
.Y(n_1229)
);

AO31x2_ASAP7_75t_L g1230 ( 
.A1(n_1097),
.A2(n_1078),
.A3(n_1079),
.B(n_1163),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1059),
.A2(n_1049),
.B(n_1074),
.Y(n_1231)
);

INVx3_ASAP7_75t_L g1232 ( 
.A(n_1124),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_1093),
.Y(n_1233)
);

OAI21x1_ASAP7_75t_L g1234 ( 
.A1(n_1074),
.A2(n_1114),
.B(n_1089),
.Y(n_1234)
);

AO31x2_ASAP7_75t_L g1235 ( 
.A1(n_1077),
.A2(n_1177),
.A3(n_1155),
.B(n_1156),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_1068),
.Y(n_1236)
);

OR2x2_ASAP7_75t_L g1237 ( 
.A(n_1148),
.B(n_1067),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1175),
.A2(n_1128),
.B(n_1189),
.Y(n_1238)
);

OR2x6_ASAP7_75t_L g1239 ( 
.A(n_1086),
.B(n_1129),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_SL g1240 ( 
.A(n_1110),
.B(n_1053),
.Y(n_1240)
);

O2A1O1Ixp33_ASAP7_75t_L g1241 ( 
.A1(n_1184),
.A2(n_1076),
.B(n_1149),
.C(n_1101),
.Y(n_1241)
);

AO31x2_ASAP7_75t_L g1242 ( 
.A1(n_1077),
.A2(n_1157),
.A3(n_1122),
.B(n_1161),
.Y(n_1242)
);

OAI21xp5_ASAP7_75t_SL g1243 ( 
.A1(n_1066),
.A2(n_1101),
.B(n_1047),
.Y(n_1243)
);

AOI221xp5_ASAP7_75t_SL g1244 ( 
.A1(n_1095),
.A2(n_1122),
.B1(n_1154),
.B2(n_1134),
.C(n_1088),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1103),
.B(n_1181),
.Y(n_1245)
);

OR2x2_ASAP7_75t_L g1246 ( 
.A(n_1087),
.B(n_1152),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1120),
.B(n_1140),
.Y(n_1247)
);

INVx2_ASAP7_75t_SL g1248 ( 
.A(n_1133),
.Y(n_1248)
);

BUFx4f_ASAP7_75t_L g1249 ( 
.A(n_1119),
.Y(n_1249)
);

AOI221xp5_ASAP7_75t_L g1250 ( 
.A1(n_1095),
.A2(n_1100),
.B1(n_1098),
.B2(n_1174),
.C(n_1168),
.Y(n_1250)
);

O2A1O1Ixp33_ASAP7_75t_L g1251 ( 
.A1(n_1180),
.A2(n_1185),
.B(n_1166),
.C(n_1127),
.Y(n_1251)
);

AOI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1046),
.A2(n_1069),
.B(n_1052),
.Y(n_1252)
);

INVx3_ASAP7_75t_L g1253 ( 
.A(n_1124),
.Y(n_1253)
);

BUFx6f_ASAP7_75t_L g1254 ( 
.A(n_1056),
.Y(n_1254)
);

AND2x2_ASAP7_75t_SL g1255 ( 
.A(n_1053),
.B(n_1086),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1054),
.Y(n_1256)
);

INVx5_ASAP7_75t_L g1257 ( 
.A(n_1119),
.Y(n_1257)
);

OAI21x1_ASAP7_75t_L g1258 ( 
.A1(n_1186),
.A2(n_1193),
.B(n_1162),
.Y(n_1258)
);

AND2x2_ASAP7_75t_L g1259 ( 
.A(n_1125),
.B(n_1137),
.Y(n_1259)
);

A2O1A1Ixp33_ASAP7_75t_L g1260 ( 
.A1(n_1190),
.A2(n_1167),
.B(n_1062),
.C(n_1132),
.Y(n_1260)
);

AOI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_1136),
.A2(n_1080),
.B(n_1117),
.Y(n_1261)
);

AOI31xp67_ASAP7_75t_L g1262 ( 
.A1(n_1183),
.A2(n_1080),
.A3(n_1159),
.B(n_1160),
.Y(n_1262)
);

AO31x2_ASAP7_75t_L g1263 ( 
.A1(n_1080),
.A2(n_1070),
.A3(n_1075),
.B(n_1150),
.Y(n_1263)
);

BUFx6f_ASAP7_75t_L g1264 ( 
.A(n_1056),
.Y(n_1264)
);

OAI21xp33_ASAP7_75t_SL g1265 ( 
.A1(n_1183),
.A2(n_1131),
.B(n_1130),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1107),
.A2(n_1179),
.B(n_1145),
.Y(n_1266)
);

NAND2x1p5_ASAP7_75t_L g1267 ( 
.A(n_1126),
.B(n_1145),
.Y(n_1267)
);

OR2x6_ASAP7_75t_L g1268 ( 
.A(n_1126),
.B(n_1151),
.Y(n_1268)
);

A2O1A1Ixp33_ASAP7_75t_L g1269 ( 
.A1(n_1096),
.A2(n_1121),
.B(n_1147),
.C(n_1172),
.Y(n_1269)
);

NOR2xp33_ASAP7_75t_L g1270 ( 
.A(n_1105),
.B(n_1176),
.Y(n_1270)
);

BUFx4f_ASAP7_75t_SL g1271 ( 
.A(n_1119),
.Y(n_1271)
);

OAI21x1_ASAP7_75t_L g1272 ( 
.A1(n_1115),
.A2(n_1116),
.B(n_1064),
.Y(n_1272)
);

NOR2xp33_ASAP7_75t_SL g1273 ( 
.A(n_1133),
.B(n_1118),
.Y(n_1273)
);

AOI221x1_ASAP7_75t_L g1274 ( 
.A1(n_1164),
.A2(n_1176),
.B1(n_1139),
.B2(n_1064),
.C(n_1143),
.Y(n_1274)
);

OAI21x1_ASAP7_75t_L g1275 ( 
.A1(n_1081),
.A2(n_1188),
.B(n_1176),
.Y(n_1275)
);

BUFx3_ASAP7_75t_L g1276 ( 
.A(n_1124),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1164),
.Y(n_1277)
);

AO31x2_ASAP7_75t_L g1278 ( 
.A1(n_1158),
.A2(n_1139),
.A3(n_1123),
.B(n_1113),
.Y(n_1278)
);

AOI21xp33_ASAP7_75t_L g1279 ( 
.A1(n_1141),
.A2(n_1153),
.B(n_1123),
.Y(n_1279)
);

OAI21xp5_ASAP7_75t_L g1280 ( 
.A1(n_1158),
.A2(n_1141),
.B(n_1153),
.Y(n_1280)
);

AO21x2_ASAP7_75t_L g1281 ( 
.A1(n_1123),
.A2(n_1065),
.B(n_1083),
.Y(n_1281)
);

BUFx10_ASAP7_75t_L g1282 ( 
.A(n_1118),
.Y(n_1282)
);

O2A1O1Ixp33_ASAP7_75t_L g1283 ( 
.A1(n_1065),
.A2(n_1083),
.B(n_1113),
.C(n_773),
.Y(n_1283)
);

AND2x6_ASAP7_75t_L g1284 ( 
.A(n_1174),
.B(n_887),
.Y(n_1284)
);

AOI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1060),
.A2(n_615),
.B(n_565),
.Y(n_1285)
);

AND2x4_ASAP7_75t_L g1286 ( 
.A(n_1102),
.B(n_955),
.Y(n_1286)
);

AOI21xp5_ASAP7_75t_L g1287 ( 
.A1(n_1060),
.A2(n_615),
.B(n_565),
.Y(n_1287)
);

AND2x2_ASAP7_75t_L g1288 ( 
.A(n_1104),
.B(n_902),
.Y(n_1288)
);

BUFx2_ASAP7_75t_L g1289 ( 
.A(n_1055),
.Y(n_1289)
);

OAI22xp5_ASAP7_75t_L g1290 ( 
.A1(n_1090),
.A2(n_868),
.B1(n_773),
.B2(n_875),
.Y(n_1290)
);

OR2x2_ASAP7_75t_L g1291 ( 
.A(n_1090),
.B(n_599),
.Y(n_1291)
);

CKINVDCx11_ASAP7_75t_R g1292 ( 
.A(n_1142),
.Y(n_1292)
);

OAI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1084),
.A2(n_868),
.B(n_867),
.Y(n_1293)
);

AO31x2_ASAP7_75t_L g1294 ( 
.A1(n_1135),
.A2(n_1058),
.A3(n_1084),
.B(n_881),
.Y(n_1294)
);

AOI221x1_ASAP7_75t_L g1295 ( 
.A1(n_1155),
.A2(n_883),
.B1(n_868),
.B2(n_1084),
.C(n_1058),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1090),
.B(n_868),
.Y(n_1296)
);

AO31x2_ASAP7_75t_L g1297 ( 
.A1(n_1135),
.A2(n_1058),
.A3(n_1084),
.B(n_881),
.Y(n_1297)
);

AOI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1060),
.A2(n_615),
.B(n_565),
.Y(n_1298)
);

AO31x2_ASAP7_75t_L g1299 ( 
.A1(n_1135),
.A2(n_1058),
.A3(n_1084),
.B(n_881),
.Y(n_1299)
);

OAI21x1_ASAP7_75t_L g1300 ( 
.A1(n_1060),
.A2(n_1071),
.B(n_1094),
.Y(n_1300)
);

AOI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1060),
.A2(n_615),
.B(n_565),
.Y(n_1301)
);

OAI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1084),
.A2(n_868),
.B(n_867),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1090),
.B(n_868),
.Y(n_1303)
);

NOR2xp67_ASAP7_75t_L g1304 ( 
.A(n_1166),
.B(n_710),
.Y(n_1304)
);

A2O1A1Ixp33_ASAP7_75t_L g1305 ( 
.A1(n_1084),
.A2(n_868),
.B(n_965),
.C(n_878),
.Y(n_1305)
);

OAI21x1_ASAP7_75t_L g1306 ( 
.A1(n_1060),
.A2(n_1071),
.B(n_1094),
.Y(n_1306)
);

BUFx6f_ASAP7_75t_L g1307 ( 
.A(n_1056),
.Y(n_1307)
);

AOI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1060),
.A2(n_615),
.B(n_565),
.Y(n_1308)
);

AND2x4_ASAP7_75t_L g1309 ( 
.A(n_1102),
.B(n_955),
.Y(n_1309)
);

OAI21xp5_ASAP7_75t_L g1310 ( 
.A1(n_1084),
.A2(n_868),
.B(n_867),
.Y(n_1310)
);

OAI21x1_ASAP7_75t_L g1311 ( 
.A1(n_1060),
.A2(n_1071),
.B(n_1094),
.Y(n_1311)
);

AO32x2_ASAP7_75t_L g1312 ( 
.A1(n_1058),
.A2(n_1079),
.A3(n_1155),
.B1(n_1078),
.B2(n_1156),
.Y(n_1312)
);

INVx3_ASAP7_75t_L g1313 ( 
.A(n_1124),
.Y(n_1313)
);

AO31x2_ASAP7_75t_L g1314 ( 
.A1(n_1135),
.A2(n_1058),
.A3(n_1084),
.B(n_881),
.Y(n_1314)
);

NOR2xp67_ASAP7_75t_L g1315 ( 
.A(n_1166),
.B(n_710),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1090),
.B(n_868),
.Y(n_1316)
);

OAI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_1084),
.A2(n_868),
.B(n_867),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1090),
.B(n_868),
.Y(n_1318)
);

NAND2x1p5_ASAP7_75t_L g1319 ( 
.A(n_1086),
.B(n_981),
.Y(n_1319)
);

OAI22xp33_ASAP7_75t_L g1320 ( 
.A1(n_1090),
.A2(n_786),
.B1(n_835),
.B2(n_842),
.Y(n_1320)
);

OR2x2_ASAP7_75t_L g1321 ( 
.A(n_1090),
.B(n_599),
.Y(n_1321)
);

BUFx3_ASAP7_75t_L g1322 ( 
.A(n_1055),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1090),
.B(n_868),
.Y(n_1323)
);

AO31x2_ASAP7_75t_L g1324 ( 
.A1(n_1135),
.A2(n_1058),
.A3(n_1084),
.B(n_881),
.Y(n_1324)
);

AOI221x1_ASAP7_75t_L g1325 ( 
.A1(n_1155),
.A2(n_883),
.B1(n_868),
.B2(n_1084),
.C(n_1058),
.Y(n_1325)
);

OAI21x1_ASAP7_75t_L g1326 ( 
.A1(n_1060),
.A2(n_1071),
.B(n_1094),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1090),
.B(n_868),
.Y(n_1327)
);

OA21x2_ASAP7_75t_L g1328 ( 
.A1(n_1146),
.A2(n_1084),
.B(n_1135),
.Y(n_1328)
);

A2O1A1Ixp33_ASAP7_75t_L g1329 ( 
.A1(n_1084),
.A2(n_868),
.B(n_965),
.C(n_878),
.Y(n_1329)
);

OAI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1084),
.A2(n_868),
.B(n_867),
.Y(n_1330)
);

BUFx10_ASAP7_75t_L g1331 ( 
.A(n_1118),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1090),
.B(n_868),
.Y(n_1332)
);

AOI21xp5_ASAP7_75t_L g1333 ( 
.A1(n_1060),
.A2(n_615),
.B(n_565),
.Y(n_1333)
);

O2A1O1Ixp33_ASAP7_75t_L g1334 ( 
.A1(n_1144),
.A2(n_773),
.B(n_965),
.C(n_785),
.Y(n_1334)
);

AOI21xp5_ASAP7_75t_L g1335 ( 
.A1(n_1060),
.A2(n_615),
.B(n_565),
.Y(n_1335)
);

BUFx6f_ASAP7_75t_L g1336 ( 
.A(n_1056),
.Y(n_1336)
);

AND2x4_ASAP7_75t_L g1337 ( 
.A(n_1102),
.B(n_955),
.Y(n_1337)
);

A2O1A1Ixp33_ASAP7_75t_L g1338 ( 
.A1(n_1084),
.A2(n_868),
.B(n_965),
.C(n_878),
.Y(n_1338)
);

AO31x2_ASAP7_75t_L g1339 ( 
.A1(n_1135),
.A2(n_1058),
.A3(n_1084),
.B(n_881),
.Y(n_1339)
);

CKINVDCx11_ASAP7_75t_R g1340 ( 
.A(n_1142),
.Y(n_1340)
);

BUFx4_ASAP7_75t_SL g1341 ( 
.A(n_1055),
.Y(n_1341)
);

OR2x6_ASAP7_75t_L g1342 ( 
.A(n_1086),
.B(n_776),
.Y(n_1342)
);

AOI21xp5_ASAP7_75t_L g1343 ( 
.A1(n_1060),
.A2(n_615),
.B(n_565),
.Y(n_1343)
);

AOI22xp5_ASAP7_75t_L g1344 ( 
.A1(n_1110),
.A2(n_786),
.B1(n_764),
.B2(n_674),
.Y(n_1344)
);

AOI21xp5_ASAP7_75t_L g1345 ( 
.A1(n_1060),
.A2(n_615),
.B(n_565),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1048),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1090),
.B(n_868),
.Y(n_1347)
);

AOI22xp33_ASAP7_75t_L g1348 ( 
.A1(n_1250),
.A2(n_1320),
.B1(n_1288),
.B2(n_1284),
.Y(n_1348)
);

AOI22xp33_ASAP7_75t_SL g1349 ( 
.A1(n_1328),
.A2(n_1229),
.B1(n_1310),
.B2(n_1330),
.Y(n_1349)
);

BUFx6f_ASAP7_75t_L g1350 ( 
.A(n_1249),
.Y(n_1350)
);

AOI22xp33_ASAP7_75t_L g1351 ( 
.A1(n_1284),
.A2(n_1344),
.B1(n_1240),
.B2(n_1246),
.Y(n_1351)
);

BUFx6f_ASAP7_75t_L g1352 ( 
.A(n_1249),
.Y(n_1352)
);

AOI22xp33_ASAP7_75t_L g1353 ( 
.A1(n_1284),
.A2(n_1302),
.B1(n_1293),
.B2(n_1317),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1247),
.Y(n_1354)
);

AOI22xp5_ASAP7_75t_L g1355 ( 
.A1(n_1243),
.A2(n_1270),
.B1(n_1304),
.B2(n_1315),
.Y(n_1355)
);

AND2x4_ASAP7_75t_L g1356 ( 
.A(n_1239),
.B(n_1286),
.Y(n_1356)
);

BUFx3_ASAP7_75t_L g1357 ( 
.A(n_1199),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_1204),
.Y(n_1358)
);

OAI22xp33_ASAP7_75t_L g1359 ( 
.A1(n_1225),
.A2(n_1347),
.B1(n_1296),
.B2(n_1303),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1259),
.B(n_1210),
.Y(n_1360)
);

AOI22xp5_ASAP7_75t_L g1361 ( 
.A1(n_1244),
.A2(n_1265),
.B1(n_1255),
.B2(n_1284),
.Y(n_1361)
);

BUFx2_ASAP7_75t_L g1362 ( 
.A(n_1322),
.Y(n_1362)
);

CKINVDCx11_ASAP7_75t_R g1363 ( 
.A(n_1223),
.Y(n_1363)
);

BUFx3_ASAP7_75t_L g1364 ( 
.A(n_1289),
.Y(n_1364)
);

INVx1_ASAP7_75t_SL g1365 ( 
.A(n_1291),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1256),
.Y(n_1366)
);

CKINVDCx20_ASAP7_75t_R g1367 ( 
.A(n_1236),
.Y(n_1367)
);

INVx1_ASAP7_75t_SL g1368 ( 
.A(n_1321),
.Y(n_1368)
);

OAI22xp5_ASAP7_75t_L g1369 ( 
.A1(n_1316),
.A2(n_1318),
.B1(n_1323),
.B2(n_1327),
.Y(n_1369)
);

CKINVDCx20_ASAP7_75t_R g1370 ( 
.A(n_1233),
.Y(n_1370)
);

BUFx2_ASAP7_75t_SL g1371 ( 
.A(n_1248),
.Y(n_1371)
);

INVx1_ASAP7_75t_SL g1372 ( 
.A(n_1341),
.Y(n_1372)
);

BUFx3_ASAP7_75t_L g1373 ( 
.A(n_1219),
.Y(n_1373)
);

BUFx6f_ASAP7_75t_L g1374 ( 
.A(n_1257),
.Y(n_1374)
);

CKINVDCx11_ASAP7_75t_R g1375 ( 
.A(n_1292),
.Y(n_1375)
);

OAI22xp5_ASAP7_75t_L g1376 ( 
.A1(n_1332),
.A2(n_1338),
.B1(n_1329),
.B2(n_1305),
.Y(n_1376)
);

AOI22xp33_ASAP7_75t_L g1377 ( 
.A1(n_1200),
.A2(n_1268),
.B1(n_1290),
.B2(n_1202),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1196),
.Y(n_1378)
);

INVx3_ASAP7_75t_SL g1379 ( 
.A(n_1342),
.Y(n_1379)
);

OAI22xp33_ASAP7_75t_L g1380 ( 
.A1(n_1295),
.A2(n_1325),
.B1(n_1268),
.B2(n_1228),
.Y(n_1380)
);

OAI22xp33_ASAP7_75t_L g1381 ( 
.A1(n_1237),
.A2(n_1346),
.B1(n_1211),
.B2(n_1196),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1211),
.Y(n_1382)
);

BUFx2_ASAP7_75t_L g1383 ( 
.A(n_1286),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_1277),
.Y(n_1384)
);

CKINVDCx11_ASAP7_75t_R g1385 ( 
.A(n_1340),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1245),
.Y(n_1386)
);

BUFx4f_ASAP7_75t_SL g1387 ( 
.A(n_1227),
.Y(n_1387)
);

OAI22xp5_ASAP7_75t_SL g1388 ( 
.A1(n_1342),
.A2(n_1239),
.B1(n_1309),
.B2(n_1337),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_1232),
.Y(n_1389)
);

AOI22xp33_ASAP7_75t_L g1390 ( 
.A1(n_1195),
.A2(n_1328),
.B1(n_1238),
.B2(n_1252),
.Y(n_1390)
);

INVx5_ASAP7_75t_L g1391 ( 
.A(n_1257),
.Y(n_1391)
);

AOI22xp33_ASAP7_75t_L g1392 ( 
.A1(n_1214),
.A2(n_1337),
.B1(n_1309),
.B2(n_1213),
.Y(n_1392)
);

AOI22xp33_ASAP7_75t_L g1393 ( 
.A1(n_1209),
.A2(n_1231),
.B1(n_1275),
.B2(n_1215),
.Y(n_1393)
);

AOI22xp33_ASAP7_75t_SL g1394 ( 
.A1(n_1273),
.A2(n_1312),
.B1(n_1334),
.B2(n_1241),
.Y(n_1394)
);

BUFx6f_ASAP7_75t_L g1395 ( 
.A(n_1217),
.Y(n_1395)
);

AOI22xp33_ASAP7_75t_L g1396 ( 
.A1(n_1319),
.A2(n_1261),
.B1(n_1212),
.B2(n_1266),
.Y(n_1396)
);

CKINVDCx11_ASAP7_75t_R g1397 ( 
.A(n_1282),
.Y(n_1397)
);

BUFx3_ASAP7_75t_L g1398 ( 
.A(n_1331),
.Y(n_1398)
);

BUFx3_ASAP7_75t_L g1399 ( 
.A(n_1331),
.Y(n_1399)
);

CKINVDCx20_ASAP7_75t_R g1400 ( 
.A(n_1271),
.Y(n_1400)
);

AOI22xp33_ASAP7_75t_L g1401 ( 
.A1(n_1276),
.A2(n_1313),
.B1(n_1253),
.B2(n_1205),
.Y(n_1401)
);

INVx5_ASAP7_75t_L g1402 ( 
.A(n_1217),
.Y(n_1402)
);

BUFx6f_ASAP7_75t_L g1403 ( 
.A(n_1217),
.Y(n_1403)
);

AOI22xp33_ASAP7_75t_L g1404 ( 
.A1(n_1253),
.A2(n_1313),
.B1(n_1208),
.B2(n_1280),
.Y(n_1404)
);

CKINVDCx11_ASAP7_75t_R g1405 ( 
.A(n_1254),
.Y(n_1405)
);

AOI22xp33_ASAP7_75t_L g1406 ( 
.A1(n_1272),
.A2(n_1234),
.B1(n_1203),
.B2(n_1220),
.Y(n_1406)
);

AOI22xp33_ASAP7_75t_L g1407 ( 
.A1(n_1222),
.A2(n_1279),
.B1(n_1336),
.B2(n_1264),
.Y(n_1407)
);

OAI22xp5_ASAP7_75t_L g1408 ( 
.A1(n_1201),
.A2(n_1260),
.B1(n_1312),
.B2(n_1269),
.Y(n_1408)
);

AOI22xp33_ASAP7_75t_L g1409 ( 
.A1(n_1254),
.A2(n_1264),
.B1(n_1307),
.B2(n_1336),
.Y(n_1409)
);

OAI22xp33_ASAP7_75t_L g1410 ( 
.A1(n_1274),
.A2(n_1312),
.B1(n_1267),
.B2(n_1224),
.Y(n_1410)
);

AOI22xp33_ASAP7_75t_L g1411 ( 
.A1(n_1258),
.A2(n_1226),
.B1(n_1242),
.B2(n_1218),
.Y(n_1411)
);

INVx6_ASAP7_75t_L g1412 ( 
.A(n_1254),
.Y(n_1412)
);

AOI22xp33_ASAP7_75t_L g1413 ( 
.A1(n_1242),
.A2(n_1264),
.B1(n_1336),
.B2(n_1307),
.Y(n_1413)
);

CKINVDCx20_ASAP7_75t_R g1414 ( 
.A(n_1307),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1283),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1281),
.Y(n_1416)
);

AOI22xp33_ASAP7_75t_L g1417 ( 
.A1(n_1242),
.A2(n_1235),
.B1(n_1251),
.B2(n_1335),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1235),
.Y(n_1418)
);

AOI22xp33_ASAP7_75t_L g1419 ( 
.A1(n_1300),
.A2(n_1306),
.B1(n_1311),
.B2(n_1326),
.Y(n_1419)
);

OAI22xp33_ASAP7_75t_L g1420 ( 
.A1(n_1194),
.A2(n_1235),
.B1(n_1343),
.B2(n_1333),
.Y(n_1420)
);

OAI22xp5_ASAP7_75t_L g1421 ( 
.A1(n_1207),
.A2(n_1345),
.B1(n_1308),
.B2(n_1285),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1230),
.Y(n_1422)
);

CKINVDCx11_ASAP7_75t_R g1423 ( 
.A(n_1262),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1230),
.Y(n_1424)
);

CKINVDCx20_ASAP7_75t_R g1425 ( 
.A(n_1287),
.Y(n_1425)
);

CKINVDCx20_ASAP7_75t_R g1426 ( 
.A(n_1298),
.Y(n_1426)
);

OAI22xp5_ASAP7_75t_L g1427 ( 
.A1(n_1301),
.A2(n_1206),
.B1(n_1230),
.B2(n_1197),
.Y(n_1427)
);

OAI22xp33_ASAP7_75t_SL g1428 ( 
.A1(n_1294),
.A2(n_1297),
.B1(n_1324),
.B2(n_1314),
.Y(n_1428)
);

CKINVDCx20_ASAP7_75t_R g1429 ( 
.A(n_1294),
.Y(n_1429)
);

AOI22xp33_ASAP7_75t_L g1430 ( 
.A1(n_1294),
.A2(n_1297),
.B1(n_1324),
.B2(n_1314),
.Y(n_1430)
);

CKINVDCx11_ASAP7_75t_R g1431 ( 
.A(n_1297),
.Y(n_1431)
);

CKINVDCx11_ASAP7_75t_R g1432 ( 
.A(n_1299),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1263),
.Y(n_1433)
);

AOI22xp33_ASAP7_75t_L g1434 ( 
.A1(n_1299),
.A2(n_1314),
.B1(n_1324),
.B2(n_1339),
.Y(n_1434)
);

CKINVDCx20_ASAP7_75t_R g1435 ( 
.A(n_1299),
.Y(n_1435)
);

OAI22xp33_ASAP7_75t_L g1436 ( 
.A1(n_1339),
.A2(n_1206),
.B1(n_1278),
.B2(n_1221),
.Y(n_1436)
);

INVx4_ASAP7_75t_L g1437 ( 
.A(n_1221),
.Y(n_1437)
);

AOI22xp33_ASAP7_75t_L g1438 ( 
.A1(n_1206),
.A2(n_965),
.B1(n_1250),
.B2(n_878),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1221),
.Y(n_1439)
);

INVx4_ASAP7_75t_L g1440 ( 
.A(n_1198),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1198),
.Y(n_1441)
);

BUFx8_ASAP7_75t_L g1442 ( 
.A(n_1227),
.Y(n_1442)
);

NAND2x1p5_ASAP7_75t_L g1443 ( 
.A(n_1257),
.B(n_981),
.Y(n_1443)
);

OA22x2_ASAP7_75t_L g1444 ( 
.A1(n_1344),
.A2(n_965),
.B1(n_677),
.B2(n_1243),
.Y(n_1444)
);

CKINVDCx6p67_ASAP7_75t_R g1445 ( 
.A(n_1342),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1247),
.Y(n_1446)
);

BUFx8_ASAP7_75t_L g1447 ( 
.A(n_1227),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1196),
.B(n_868),
.Y(n_1448)
);

INVx6_ASAP7_75t_L g1449 ( 
.A(n_1257),
.Y(n_1449)
);

OAI21xp5_ASAP7_75t_SL g1450 ( 
.A1(n_1344),
.A2(n_677),
.B(n_681),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1216),
.Y(n_1451)
);

BUFx10_ASAP7_75t_L g1452 ( 
.A(n_1233),
.Y(n_1452)
);

INVx1_ASAP7_75t_SL g1453 ( 
.A(n_1289),
.Y(n_1453)
);

CKINVDCx20_ASAP7_75t_R g1454 ( 
.A(n_1236),
.Y(n_1454)
);

AOI22xp33_ASAP7_75t_L g1455 ( 
.A1(n_1250),
.A2(n_965),
.B1(n_878),
.B2(n_1110),
.Y(n_1455)
);

CKINVDCx16_ASAP7_75t_R g1456 ( 
.A(n_1273),
.Y(n_1456)
);

OAI21xp33_ASAP7_75t_SL g1457 ( 
.A1(n_1250),
.A2(n_868),
.B(n_974),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1247),
.Y(n_1458)
);

BUFx10_ASAP7_75t_L g1459 ( 
.A(n_1233),
.Y(n_1459)
);

CKINVDCx11_ASAP7_75t_R g1460 ( 
.A(n_1223),
.Y(n_1460)
);

CKINVDCx5p33_ASAP7_75t_R g1461 ( 
.A(n_1341),
.Y(n_1461)
);

NAND2x1p5_ASAP7_75t_L g1462 ( 
.A(n_1257),
.B(n_981),
.Y(n_1462)
);

INVx6_ASAP7_75t_L g1463 ( 
.A(n_1257),
.Y(n_1463)
);

AOI22xp33_ASAP7_75t_L g1464 ( 
.A1(n_1250),
.A2(n_965),
.B1(n_878),
.B2(n_1110),
.Y(n_1464)
);

AOI21xp33_ASAP7_75t_L g1465 ( 
.A1(n_1241),
.A2(n_868),
.B(n_1334),
.Y(n_1465)
);

BUFx10_ASAP7_75t_L g1466 ( 
.A(n_1233),
.Y(n_1466)
);

AOI22xp33_ASAP7_75t_SL g1467 ( 
.A1(n_1328),
.A2(n_1110),
.B1(n_786),
.B2(n_835),
.Y(n_1467)
);

CKINVDCx11_ASAP7_75t_R g1468 ( 
.A(n_1223),
.Y(n_1468)
);

AND2x4_ASAP7_75t_L g1469 ( 
.A(n_1239),
.B(n_1286),
.Y(n_1469)
);

AOI22xp33_ASAP7_75t_L g1470 ( 
.A1(n_1250),
.A2(n_965),
.B1(n_878),
.B2(n_1110),
.Y(n_1470)
);

AOI22xp33_ASAP7_75t_L g1471 ( 
.A1(n_1250),
.A2(n_965),
.B1(n_878),
.B2(n_1110),
.Y(n_1471)
);

AOI22xp33_ASAP7_75t_SL g1472 ( 
.A1(n_1328),
.A2(n_1110),
.B1(n_786),
.B2(n_835),
.Y(n_1472)
);

BUFx4f_ASAP7_75t_L g1473 ( 
.A(n_1255),
.Y(n_1473)
);

NAND2x1p5_ASAP7_75t_L g1474 ( 
.A(n_1257),
.B(n_981),
.Y(n_1474)
);

BUFx10_ASAP7_75t_L g1475 ( 
.A(n_1233),
.Y(n_1475)
);

AOI22xp33_ASAP7_75t_L g1476 ( 
.A1(n_1250),
.A2(n_965),
.B1(n_1110),
.B2(n_878),
.Y(n_1476)
);

AOI22xp33_ASAP7_75t_L g1477 ( 
.A1(n_1250),
.A2(n_965),
.B1(n_1110),
.B2(n_878),
.Y(n_1477)
);

CKINVDCx20_ASAP7_75t_R g1478 ( 
.A(n_1236),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1247),
.Y(n_1479)
);

BUFx10_ASAP7_75t_L g1480 ( 
.A(n_1233),
.Y(n_1480)
);

INVx3_ASAP7_75t_L g1481 ( 
.A(n_1232),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1247),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1247),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1247),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1418),
.Y(n_1485)
);

HB1xp67_ASAP7_75t_L g1486 ( 
.A(n_1386),
.Y(n_1486)
);

OR2x2_ASAP7_75t_L g1487 ( 
.A(n_1422),
.B(n_1424),
.Y(n_1487)
);

BUFx12f_ASAP7_75t_L g1488 ( 
.A(n_1363),
.Y(n_1488)
);

OA21x2_ASAP7_75t_L g1489 ( 
.A1(n_1433),
.A2(n_1411),
.B(n_1430),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1441),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1378),
.Y(n_1491)
);

INVx2_ASAP7_75t_L g1492 ( 
.A(n_1382),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1369),
.B(n_1359),
.Y(n_1493)
);

HB1xp67_ASAP7_75t_L g1494 ( 
.A(n_1365),
.Y(n_1494)
);

AND2x4_ASAP7_75t_L g1495 ( 
.A(n_1366),
.B(n_1384),
.Y(n_1495)
);

BUFx2_ASAP7_75t_L g1496 ( 
.A(n_1416),
.Y(n_1496)
);

INVx2_ASAP7_75t_SL g1497 ( 
.A(n_1449),
.Y(n_1497)
);

INVx2_ASAP7_75t_SL g1498 ( 
.A(n_1449),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1369),
.B(n_1359),
.Y(n_1499)
);

OAI21x1_ASAP7_75t_L g1500 ( 
.A1(n_1421),
.A2(n_1406),
.B(n_1419),
.Y(n_1500)
);

AND2x4_ASAP7_75t_L g1501 ( 
.A(n_1361),
.B(n_1451),
.Y(n_1501)
);

OAI21x1_ASAP7_75t_L g1502 ( 
.A1(n_1421),
.A2(n_1396),
.B(n_1393),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1360),
.B(n_1354),
.Y(n_1503)
);

HB1xp67_ASAP7_75t_L g1504 ( 
.A(n_1368),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1440),
.Y(n_1505)
);

OAI22xp33_ASAP7_75t_L g1506 ( 
.A1(n_1444),
.A2(n_1450),
.B1(n_1473),
.B2(n_1355),
.Y(n_1506)
);

INVx2_ASAP7_75t_SL g1507 ( 
.A(n_1449),
.Y(n_1507)
);

CKINVDCx11_ASAP7_75t_R g1508 ( 
.A(n_1375),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1394),
.B(n_1429),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1428),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1440),
.Y(n_1511)
);

CKINVDCx11_ASAP7_75t_R g1512 ( 
.A(n_1385),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1435),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1394),
.B(n_1349),
.Y(n_1514)
);

INVx2_ASAP7_75t_L g1515 ( 
.A(n_1358),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1408),
.Y(n_1516)
);

INVx4_ASAP7_75t_L g1517 ( 
.A(n_1391),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1408),
.Y(n_1518)
);

HB1xp67_ASAP7_75t_L g1519 ( 
.A(n_1446),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1439),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1415),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1349),
.B(n_1438),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1413),
.B(n_1431),
.Y(n_1523)
);

NAND2xp33_ASAP7_75t_R g1524 ( 
.A(n_1461),
.B(n_1362),
.Y(n_1524)
);

INVx6_ASAP7_75t_L g1525 ( 
.A(n_1391),
.Y(n_1525)
);

OAI21x1_ASAP7_75t_L g1526 ( 
.A1(n_1427),
.A2(n_1417),
.B(n_1404),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1458),
.Y(n_1527)
);

OAI21x1_ASAP7_75t_L g1528 ( 
.A1(n_1417),
.A2(n_1390),
.B(n_1413),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1479),
.Y(n_1529)
);

INVx3_ASAP7_75t_L g1530 ( 
.A(n_1391),
.Y(n_1530)
);

HB1xp67_ASAP7_75t_L g1531 ( 
.A(n_1482),
.Y(n_1531)
);

OAI21x1_ASAP7_75t_L g1532 ( 
.A1(n_1434),
.A2(n_1353),
.B(n_1376),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1483),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1484),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1437),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1437),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1436),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1436),
.Y(n_1538)
);

INVx2_ASAP7_75t_SL g1539 ( 
.A(n_1463),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1381),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1381),
.Y(n_1541)
);

NOR2xp33_ASAP7_75t_L g1542 ( 
.A(n_1383),
.B(n_1473),
.Y(n_1542)
);

OAI22xp5_ASAP7_75t_L g1543 ( 
.A1(n_1467),
.A2(n_1472),
.B1(n_1477),
.B2(n_1476),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1432),
.B(n_1377),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1420),
.Y(n_1545)
);

OR2x2_ASAP7_75t_L g1546 ( 
.A(n_1380),
.B(n_1376),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1420),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1476),
.B(n_1477),
.Y(n_1548)
);

OR2x2_ASAP7_75t_L g1549 ( 
.A(n_1380),
.B(n_1351),
.Y(n_1549)
);

AOI21x1_ASAP7_75t_L g1550 ( 
.A1(n_1448),
.A2(n_1444),
.B(n_1389),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1423),
.B(n_1348),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1448),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1465),
.B(n_1467),
.Y(n_1553)
);

AOI21x1_ASAP7_75t_L g1554 ( 
.A1(n_1356),
.A2(n_1469),
.B(n_1465),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1410),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1410),
.Y(n_1556)
);

NOR2xp33_ASAP7_75t_L g1557 ( 
.A(n_1364),
.B(n_1453),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1455),
.B(n_1464),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1425),
.Y(n_1559)
);

BUFx6f_ASAP7_75t_L g1560 ( 
.A(n_1374),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1472),
.B(n_1471),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1426),
.Y(n_1562)
);

OAI21xp5_ASAP7_75t_L g1563 ( 
.A1(n_1470),
.A2(n_1457),
.B(n_1392),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1469),
.B(n_1373),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1401),
.Y(n_1565)
);

HB1xp67_ASAP7_75t_L g1566 ( 
.A(n_1481),
.Y(n_1566)
);

OAI21xp5_ASAP7_75t_L g1567 ( 
.A1(n_1407),
.A2(n_1462),
.B(n_1443),
.Y(n_1567)
);

OAI21xp5_ASAP7_75t_L g1568 ( 
.A1(n_1443),
.A2(n_1474),
.B(n_1462),
.Y(n_1568)
);

OR2x2_ASAP7_75t_L g1569 ( 
.A(n_1456),
.B(n_1379),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1481),
.B(n_1395),
.Y(n_1570)
);

OAI21x1_ASAP7_75t_L g1571 ( 
.A1(n_1474),
.A2(n_1409),
.B(n_1388),
.Y(n_1571)
);

OAI21x1_ASAP7_75t_L g1572 ( 
.A1(n_1463),
.A2(n_1402),
.B(n_1445),
.Y(n_1572)
);

INVx2_ASAP7_75t_SL g1573 ( 
.A(n_1374),
.Y(n_1573)
);

NAND2x1p5_ASAP7_75t_L g1574 ( 
.A(n_1374),
.B(n_1399),
.Y(n_1574)
);

OAI21x1_ASAP7_75t_L g1575 ( 
.A1(n_1379),
.A2(n_1412),
.B(n_1371),
.Y(n_1575)
);

CKINVDCx16_ASAP7_75t_R g1576 ( 
.A(n_1400),
.Y(n_1576)
);

OAI21x1_ASAP7_75t_L g1577 ( 
.A1(n_1412),
.A2(n_1405),
.B(n_1403),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1395),
.Y(n_1578)
);

OR2x2_ASAP7_75t_L g1579 ( 
.A(n_1357),
.B(n_1398),
.Y(n_1579)
);

BUFx3_ASAP7_75t_L g1580 ( 
.A(n_1414),
.Y(n_1580)
);

INVx6_ASAP7_75t_SL g1581 ( 
.A(n_1452),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1350),
.Y(n_1582)
);

OR2x2_ASAP7_75t_L g1583 ( 
.A(n_1372),
.B(n_1350),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1352),
.B(n_1480),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1352),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1452),
.B(n_1459),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1397),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1459),
.Y(n_1588)
);

INVxp67_ASAP7_75t_SL g1589 ( 
.A(n_1442),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1466),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1466),
.Y(n_1591)
);

BUFx12f_ASAP7_75t_L g1592 ( 
.A(n_1508),
.Y(n_1592)
);

AND2x4_ASAP7_75t_L g1593 ( 
.A(n_1575),
.B(n_1370),
.Y(n_1593)
);

AND2x4_ASAP7_75t_L g1594 ( 
.A(n_1575),
.B(n_1478),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1559),
.B(n_1475),
.Y(n_1595)
);

NOR2x1_ASAP7_75t_SL g1596 ( 
.A(n_1546),
.B(n_1468),
.Y(n_1596)
);

OA21x2_ASAP7_75t_L g1597 ( 
.A1(n_1526),
.A2(n_1475),
.B(n_1387),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1540),
.B(n_1442),
.Y(n_1598)
);

NAND3xp33_ASAP7_75t_L g1599 ( 
.A(n_1563),
.B(n_1447),
.C(n_1460),
.Y(n_1599)
);

A2O1A1Ixp33_ASAP7_75t_L g1600 ( 
.A1(n_1543),
.A2(n_1367),
.B(n_1454),
.C(n_1387),
.Y(n_1600)
);

O2A1O1Ixp33_ASAP7_75t_SL g1601 ( 
.A1(n_1506),
.A2(n_1447),
.B(n_1548),
.C(n_1558),
.Y(n_1601)
);

OAI21xp5_ASAP7_75t_L g1602 ( 
.A1(n_1493),
.A2(n_1499),
.B(n_1546),
.Y(n_1602)
);

AOI221xp5_ASAP7_75t_L g1603 ( 
.A1(n_1561),
.A2(n_1553),
.B1(n_1551),
.B2(n_1516),
.C(n_1518),
.Y(n_1603)
);

OAI21x1_ASAP7_75t_L g1604 ( 
.A1(n_1500),
.A2(n_1502),
.B(n_1554),
.Y(n_1604)
);

NOR2x1_ASAP7_75t_L g1605 ( 
.A(n_1590),
.B(n_1588),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1513),
.B(n_1562),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1495),
.Y(n_1607)
);

A2O1A1Ixp33_ASAP7_75t_L g1608 ( 
.A1(n_1549),
.A2(n_1561),
.B(n_1551),
.C(n_1532),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1513),
.B(n_1562),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1540),
.B(n_1541),
.Y(n_1610)
);

OR2x2_ASAP7_75t_L g1611 ( 
.A(n_1510),
.B(n_1494),
.Y(n_1611)
);

INVxp67_ASAP7_75t_L g1612 ( 
.A(n_1519),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1544),
.B(n_1523),
.Y(n_1613)
);

OR2x6_ASAP7_75t_L g1614 ( 
.A(n_1528),
.B(n_1532),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1541),
.B(n_1516),
.Y(n_1615)
);

OAI211xp5_ASAP7_75t_L g1616 ( 
.A1(n_1549),
.A2(n_1553),
.B(n_1509),
.C(n_1514),
.Y(n_1616)
);

NOR2xp33_ASAP7_75t_L g1617 ( 
.A(n_1557),
.B(n_1576),
.Y(n_1617)
);

AO32x2_ASAP7_75t_L g1618 ( 
.A1(n_1497),
.A2(n_1507),
.A3(n_1498),
.B1(n_1539),
.B2(n_1510),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1518),
.B(n_1552),
.Y(n_1619)
);

NAND2x1_ASAP7_75t_L g1620 ( 
.A(n_1525),
.B(n_1521),
.Y(n_1620)
);

AND2x4_ASAP7_75t_L g1621 ( 
.A(n_1491),
.B(n_1492),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1523),
.B(n_1486),
.Y(n_1622)
);

OR2x2_ASAP7_75t_L g1623 ( 
.A(n_1504),
.B(n_1531),
.Y(n_1623)
);

AND2x4_ASAP7_75t_L g1624 ( 
.A(n_1495),
.B(n_1577),
.Y(n_1624)
);

OAI22xp5_ASAP7_75t_SL g1625 ( 
.A1(n_1587),
.A2(n_1569),
.B1(n_1589),
.B2(n_1488),
.Y(n_1625)
);

OAI22xp5_ASAP7_75t_L g1626 ( 
.A1(n_1514),
.A2(n_1503),
.B1(n_1522),
.B2(n_1555),
.Y(n_1626)
);

OA21x2_ASAP7_75t_L g1627 ( 
.A1(n_1528),
.A2(n_1547),
.B(n_1545),
.Y(n_1627)
);

OAI21xp5_ASAP7_75t_L g1628 ( 
.A1(n_1554),
.A2(n_1567),
.B(n_1550),
.Y(n_1628)
);

NOR2xp33_ASAP7_75t_L g1629 ( 
.A(n_1564),
.B(n_1583),
.Y(n_1629)
);

NOR2xp33_ASAP7_75t_L g1630 ( 
.A(n_1583),
.B(n_1580),
.Y(n_1630)
);

A2O1A1Ixp33_ASAP7_75t_L g1631 ( 
.A1(n_1542),
.A2(n_1571),
.B(n_1556),
.C(n_1547),
.Y(n_1631)
);

AO32x2_ASAP7_75t_L g1632 ( 
.A1(n_1497),
.A2(n_1507),
.A3(n_1498),
.B1(n_1539),
.B2(n_1537),
.Y(n_1632)
);

O2A1O1Ixp33_ASAP7_75t_SL g1633 ( 
.A1(n_1587),
.A2(n_1586),
.B(n_1590),
.C(n_1569),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1485),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1485),
.Y(n_1635)
);

NOR2xp33_ASAP7_75t_L g1636 ( 
.A(n_1580),
.B(n_1579),
.Y(n_1636)
);

INVx1_ASAP7_75t_SL g1637 ( 
.A(n_1566),
.Y(n_1637)
);

NOR2xp33_ASAP7_75t_L g1638 ( 
.A(n_1579),
.B(n_1588),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1487),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1501),
.B(n_1570),
.Y(n_1640)
);

OR2x6_ASAP7_75t_L g1641 ( 
.A(n_1572),
.B(n_1525),
.Y(n_1641)
);

OAI21xp5_ASAP7_75t_L g1642 ( 
.A1(n_1550),
.A2(n_1565),
.B(n_1571),
.Y(n_1642)
);

INVx1_ASAP7_75t_SL g1643 ( 
.A(n_1496),
.Y(n_1643)
);

AOI21xp33_ASAP7_75t_L g1644 ( 
.A1(n_1565),
.A2(n_1533),
.B(n_1529),
.Y(n_1644)
);

O2A1O1Ixp33_ASAP7_75t_L g1645 ( 
.A1(n_1527),
.A2(n_1534),
.B(n_1568),
.C(n_1591),
.Y(n_1645)
);

AO32x2_ASAP7_75t_L g1646 ( 
.A1(n_1537),
.A2(n_1538),
.A3(n_1517),
.B1(n_1573),
.B2(n_1536),
.Y(n_1646)
);

AOI221xp5_ASAP7_75t_L g1647 ( 
.A1(n_1538),
.A2(n_1591),
.B1(n_1515),
.B2(n_1535),
.C(n_1536),
.Y(n_1647)
);

NOR2xp67_ASAP7_75t_SL g1648 ( 
.A(n_1488),
.B(n_1525),
.Y(n_1648)
);

OA21x2_ASAP7_75t_L g1649 ( 
.A1(n_1490),
.A2(n_1511),
.B(n_1505),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1634),
.Y(n_1650)
);

OR2x2_ASAP7_75t_L g1651 ( 
.A(n_1627),
.B(n_1535),
.Y(n_1651)
);

HB1xp67_ASAP7_75t_L g1652 ( 
.A(n_1649),
.Y(n_1652)
);

AOI21xp33_ASAP7_75t_L g1653 ( 
.A1(n_1616),
.A2(n_1489),
.B(n_1490),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1635),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1614),
.B(n_1489),
.Y(n_1655)
);

AND2x4_ASAP7_75t_SL g1656 ( 
.A(n_1641),
.B(n_1517),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1614),
.B(n_1627),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1614),
.B(n_1489),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1646),
.B(n_1489),
.Y(n_1659)
);

BUFx3_ASAP7_75t_L g1660 ( 
.A(n_1641),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1646),
.B(n_1604),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1646),
.B(n_1520),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1621),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1612),
.B(n_1639),
.Y(n_1664)
);

BUFx2_ASAP7_75t_L g1665 ( 
.A(n_1618),
.Y(n_1665)
);

NOR2x1p5_ASAP7_75t_L g1666 ( 
.A(n_1599),
.B(n_1530),
.Y(n_1666)
);

HB1xp67_ASAP7_75t_L g1667 ( 
.A(n_1643),
.Y(n_1667)
);

CKINVDCx5p33_ASAP7_75t_R g1668 ( 
.A(n_1592),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1632),
.Y(n_1669)
);

INVx4_ASAP7_75t_L g1670 ( 
.A(n_1593),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1632),
.Y(n_1671)
);

BUFx2_ASAP7_75t_L g1672 ( 
.A(n_1618),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1632),
.Y(n_1673)
);

BUFx2_ASAP7_75t_L g1674 ( 
.A(n_1618),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1619),
.Y(n_1675)
);

HB1xp67_ASAP7_75t_L g1676 ( 
.A(n_1643),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1655),
.B(n_1597),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1675),
.B(n_1611),
.Y(n_1678)
);

AOI22xp33_ASAP7_75t_L g1679 ( 
.A1(n_1653),
.A2(n_1602),
.B1(n_1603),
.B2(n_1606),
.Y(n_1679)
);

OAI22xp5_ASAP7_75t_L g1680 ( 
.A1(n_1665),
.A2(n_1616),
.B1(n_1603),
.B2(n_1608),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1650),
.Y(n_1681)
);

NOR2xp33_ASAP7_75t_L g1682 ( 
.A(n_1664),
.B(n_1633),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1655),
.B(n_1597),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1655),
.B(n_1628),
.Y(n_1684)
);

BUFx2_ASAP7_75t_L g1685 ( 
.A(n_1660),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1658),
.B(n_1628),
.Y(n_1686)
);

NOR3xp33_ASAP7_75t_L g1687 ( 
.A(n_1653),
.B(n_1600),
.C(n_1601),
.Y(n_1687)
);

OAI221xp5_ASAP7_75t_SL g1688 ( 
.A1(n_1665),
.A2(n_1631),
.B1(n_1645),
.B2(n_1613),
.C(n_1647),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1652),
.Y(n_1689)
);

OAI221xp5_ASAP7_75t_L g1690 ( 
.A1(n_1668),
.A2(n_1602),
.B1(n_1598),
.B2(n_1642),
.C(n_1626),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1658),
.B(n_1642),
.Y(n_1691)
);

OAI211xp5_ASAP7_75t_L g1692 ( 
.A1(n_1665),
.A2(n_1645),
.B(n_1626),
.C(n_1598),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1658),
.B(n_1659),
.Y(n_1693)
);

NAND3xp33_ASAP7_75t_L g1694 ( 
.A(n_1661),
.B(n_1605),
.C(n_1647),
.Y(n_1694)
);

OAI31xp33_ASAP7_75t_SL g1695 ( 
.A1(n_1657),
.A2(n_1593),
.A3(n_1594),
.B(n_1630),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1661),
.B(n_1607),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1652),
.Y(n_1697)
);

OAI221xp5_ASAP7_75t_L g1698 ( 
.A1(n_1668),
.A2(n_1625),
.B1(n_1638),
.B2(n_1636),
.C(n_1648),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1654),
.Y(n_1699)
);

OAI22xp5_ASAP7_75t_L g1700 ( 
.A1(n_1672),
.A2(n_1623),
.B1(n_1609),
.B2(n_1610),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1662),
.Y(n_1701)
);

NOR2xp33_ASAP7_75t_L g1702 ( 
.A(n_1664),
.B(n_1663),
.Y(n_1702)
);

OR2x2_ASAP7_75t_L g1703 ( 
.A(n_1674),
.B(n_1637),
.Y(n_1703)
);

BUFx2_ASAP7_75t_L g1704 ( 
.A(n_1660),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1674),
.B(n_1622),
.Y(n_1705)
);

OAI22xp5_ASAP7_75t_L g1706 ( 
.A1(n_1674),
.A2(n_1629),
.B1(n_1615),
.B2(n_1594),
.Y(n_1706)
);

AND2x4_ASAP7_75t_L g1707 ( 
.A(n_1660),
.B(n_1656),
.Y(n_1707)
);

INVxp67_ASAP7_75t_L g1708 ( 
.A(n_1667),
.Y(n_1708)
);

BUFx3_ASAP7_75t_L g1709 ( 
.A(n_1676),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1657),
.B(n_1640),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1657),
.B(n_1624),
.Y(n_1711)
);

AOI221xp5_ASAP7_75t_L g1712 ( 
.A1(n_1669),
.A2(n_1644),
.B1(n_1615),
.B2(n_1619),
.C(n_1595),
.Y(n_1712)
);

HB1xp67_ASAP7_75t_L g1713 ( 
.A(n_1667),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_1662),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1693),
.B(n_1669),
.Y(n_1715)
);

INVx2_ASAP7_75t_L g1716 ( 
.A(n_1689),
.Y(n_1716)
);

BUFx2_ASAP7_75t_L g1717 ( 
.A(n_1707),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1681),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1681),
.Y(n_1719)
);

INVx2_ASAP7_75t_L g1720 ( 
.A(n_1689),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1693),
.B(n_1671),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1689),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1678),
.B(n_1671),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1697),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1697),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_1701),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1693),
.B(n_1673),
.Y(n_1727)
);

HB1xp67_ASAP7_75t_L g1728 ( 
.A(n_1713),
.Y(n_1728)
);

INVx2_ASAP7_75t_SL g1729 ( 
.A(n_1709),
.Y(n_1729)
);

INVx3_ASAP7_75t_L g1730 ( 
.A(n_1714),
.Y(n_1730)
);

BUFx3_ASAP7_75t_L g1731 ( 
.A(n_1704),
.Y(n_1731)
);

OR2x2_ASAP7_75t_L g1732 ( 
.A(n_1703),
.B(n_1651),
.Y(n_1732)
);

OR2x6_ASAP7_75t_L g1733 ( 
.A(n_1694),
.B(n_1620),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1696),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1699),
.Y(n_1735)
);

INVx3_ASAP7_75t_R g1736 ( 
.A(n_1685),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1699),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1678),
.B(n_1675),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1717),
.B(n_1684),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1730),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1738),
.B(n_1682),
.Y(n_1741)
);

NOR3x1_ASAP7_75t_L g1742 ( 
.A(n_1717),
.B(n_1692),
.C(n_1690),
.Y(n_1742)
);

AOI22xp33_ASAP7_75t_L g1743 ( 
.A1(n_1733),
.A2(n_1687),
.B1(n_1680),
.B2(n_1690),
.Y(n_1743)
);

HB1xp67_ASAP7_75t_L g1744 ( 
.A(n_1731),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1735),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1738),
.B(n_1682),
.Y(n_1746)
);

INVx4_ASAP7_75t_L g1747 ( 
.A(n_1731),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1735),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1717),
.B(n_1684),
.Y(n_1749)
);

OR2x2_ASAP7_75t_L g1750 ( 
.A(n_1723),
.B(n_1703),
.Y(n_1750)
);

OAI31xp33_ASAP7_75t_SL g1751 ( 
.A1(n_1736),
.A2(n_1692),
.A3(n_1680),
.B(n_1694),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_1730),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1735),
.Y(n_1753)
);

OR2x2_ASAP7_75t_L g1754 ( 
.A(n_1723),
.B(n_1703),
.Y(n_1754)
);

INVxp67_ASAP7_75t_SL g1755 ( 
.A(n_1728),
.Y(n_1755)
);

INVx2_ASAP7_75t_L g1756 ( 
.A(n_1730),
.Y(n_1756)
);

OR2x2_ASAP7_75t_L g1757 ( 
.A(n_1732),
.B(n_1700),
.Y(n_1757)
);

OR2x2_ASAP7_75t_L g1758 ( 
.A(n_1732),
.B(n_1700),
.Y(n_1758)
);

OR2x2_ASAP7_75t_L g1759 ( 
.A(n_1732),
.B(n_1708),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1728),
.B(n_1705),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1715),
.B(n_1684),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1737),
.Y(n_1762)
);

INVx2_ASAP7_75t_L g1763 ( 
.A(n_1730),
.Y(n_1763)
);

AOI22xp5_ASAP7_75t_L g1764 ( 
.A1(n_1733),
.A2(n_1687),
.B1(n_1679),
.B2(n_1666),
.Y(n_1764)
);

HB1xp67_ASAP7_75t_L g1765 ( 
.A(n_1731),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1737),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1737),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1715),
.B(n_1686),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1718),
.B(n_1705),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1718),
.Y(n_1770)
);

INVx2_ASAP7_75t_L g1771 ( 
.A(n_1730),
.Y(n_1771)
);

AOI22xp33_ASAP7_75t_L g1772 ( 
.A1(n_1733),
.A2(n_1666),
.B1(n_1670),
.B2(n_1679),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1730),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1718),
.B(n_1705),
.Y(n_1774)
);

OR2x2_ASAP7_75t_L g1775 ( 
.A(n_1733),
.B(n_1708),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1715),
.B(n_1686),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1721),
.B(n_1686),
.Y(n_1777)
);

INVx2_ASAP7_75t_L g1778 ( 
.A(n_1726),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1719),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1719),
.Y(n_1780)
);

CKINVDCx16_ASAP7_75t_R g1781 ( 
.A(n_1731),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1721),
.B(n_1711),
.Y(n_1782)
);

INVxp67_ASAP7_75t_L g1783 ( 
.A(n_1729),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1719),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1745),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1746),
.B(n_1691),
.Y(n_1786)
);

NOR2xp33_ASAP7_75t_L g1787 ( 
.A(n_1741),
.B(n_1512),
.Y(n_1787)
);

NOR2x1_ASAP7_75t_L g1788 ( 
.A(n_1747),
.B(n_1733),
.Y(n_1788)
);

OR2x2_ASAP7_75t_L g1789 ( 
.A(n_1741),
.B(n_1706),
.Y(n_1789)
);

INVx2_ASAP7_75t_L g1790 ( 
.A(n_1747),
.Y(n_1790)
);

BUFx2_ASAP7_75t_L g1791 ( 
.A(n_1783),
.Y(n_1791)
);

AND2x4_ASAP7_75t_L g1792 ( 
.A(n_1747),
.B(n_1729),
.Y(n_1792)
);

OAI21x1_ASAP7_75t_L g1793 ( 
.A1(n_1740),
.A2(n_1756),
.B(n_1752),
.Y(n_1793)
);

INVx1_ASAP7_75t_SL g1794 ( 
.A(n_1781),
.Y(n_1794)
);

OAI211xp5_ASAP7_75t_L g1795 ( 
.A1(n_1751),
.A2(n_1688),
.B(n_1712),
.C(n_1695),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1781),
.B(n_1733),
.Y(n_1796)
);

INVx1_ASAP7_75t_SL g1797 ( 
.A(n_1744),
.Y(n_1797)
);

OR2x2_ASAP7_75t_L g1798 ( 
.A(n_1760),
.B(n_1706),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1745),
.Y(n_1799)
);

OR2x2_ASAP7_75t_L g1800 ( 
.A(n_1760),
.B(n_1688),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1739),
.B(n_1733),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1739),
.B(n_1729),
.Y(n_1802)
);

INVx2_ASAP7_75t_SL g1803 ( 
.A(n_1765),
.Y(n_1803)
);

OAI21xp33_ASAP7_75t_L g1804 ( 
.A1(n_1751),
.A2(n_1695),
.B(n_1683),
.Y(n_1804)
);

OR2x2_ASAP7_75t_L g1805 ( 
.A(n_1757),
.B(n_1734),
.Y(n_1805)
);

OR2x2_ASAP7_75t_L g1806 ( 
.A(n_1757),
.B(n_1734),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1748),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_1743),
.B(n_1691),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1748),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1742),
.B(n_1691),
.Y(n_1810)
);

OR2x2_ASAP7_75t_L g1811 ( 
.A(n_1758),
.B(n_1734),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1753),
.Y(n_1812)
);

NAND2xp33_ASAP7_75t_L g1813 ( 
.A(n_1764),
.B(n_1713),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1753),
.Y(n_1814)
);

AND2x4_ASAP7_75t_L g1815 ( 
.A(n_1747),
.B(n_1782),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1762),
.Y(n_1816)
);

OR2x2_ASAP7_75t_L g1817 ( 
.A(n_1758),
.B(n_1734),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1742),
.B(n_1702),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1764),
.B(n_1702),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1755),
.B(n_1710),
.Y(n_1820)
);

INVx2_ASAP7_75t_SL g1821 ( 
.A(n_1749),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1785),
.Y(n_1822)
);

INVx2_ASAP7_75t_L g1823 ( 
.A(n_1821),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1799),
.Y(n_1824)
);

AOI22xp5_ASAP7_75t_L g1825 ( 
.A1(n_1795),
.A2(n_1772),
.B1(n_1749),
.B2(n_1683),
.Y(n_1825)
);

AOI221x1_ASAP7_75t_L g1826 ( 
.A1(n_1804),
.A2(n_1762),
.B1(n_1767),
.B2(n_1766),
.C(n_1779),
.Y(n_1826)
);

NOR2xp33_ASAP7_75t_L g1827 ( 
.A(n_1787),
.B(n_1794),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_L g1828 ( 
.A(n_1818),
.B(n_1782),
.Y(n_1828)
);

XOR2x2_ASAP7_75t_L g1829 ( 
.A(n_1787),
.B(n_1596),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1807),
.Y(n_1830)
);

AOI22xp5_ASAP7_75t_L g1831 ( 
.A1(n_1813),
.A2(n_1810),
.B1(n_1819),
.B2(n_1808),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1796),
.B(n_1761),
.Y(n_1832)
);

OAI32xp33_ASAP7_75t_L g1833 ( 
.A1(n_1800),
.A2(n_1775),
.A3(n_1759),
.B1(n_1754),
.B2(n_1750),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1809),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1812),
.Y(n_1835)
);

AND2x2_ASAP7_75t_L g1836 ( 
.A(n_1802),
.B(n_1761),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1814),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1797),
.B(n_1791),
.Y(n_1838)
);

AOI21xp5_ASAP7_75t_L g1839 ( 
.A1(n_1813),
.A2(n_1698),
.B(n_1775),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1816),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1803),
.B(n_1790),
.Y(n_1841)
);

INVx1_ASAP7_75t_SL g1842 ( 
.A(n_1802),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1803),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1821),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1790),
.Y(n_1845)
);

OAI21xp33_ASAP7_75t_L g1846 ( 
.A1(n_1789),
.A2(n_1759),
.B(n_1683),
.Y(n_1846)
);

AOI221xp5_ASAP7_75t_L g1847 ( 
.A1(n_1796),
.A2(n_1712),
.B1(n_1767),
.B2(n_1766),
.C(n_1779),
.Y(n_1847)
);

NAND2xp33_ASAP7_75t_L g1848 ( 
.A(n_1788),
.B(n_1798),
.Y(n_1848)
);

NOR2xp67_ASAP7_75t_L g1849 ( 
.A(n_1815),
.B(n_1750),
.Y(n_1849)
);

INVx1_ASAP7_75t_SL g1850 ( 
.A(n_1842),
.Y(n_1850)
);

INVx2_ASAP7_75t_L g1851 ( 
.A(n_1836),
.Y(n_1851)
);

AOI22xp5_ASAP7_75t_L g1852 ( 
.A1(n_1831),
.A2(n_1815),
.B1(n_1801),
.B2(n_1820),
.Y(n_1852)
);

INVx2_ASAP7_75t_L g1853 ( 
.A(n_1836),
.Y(n_1853)
);

OAI221xp5_ASAP7_75t_L g1854 ( 
.A1(n_1825),
.A2(n_1801),
.B1(n_1698),
.B2(n_1811),
.C(n_1806),
.Y(n_1854)
);

AOI322xp5_ASAP7_75t_L g1855 ( 
.A1(n_1827),
.A2(n_1786),
.A3(n_1768),
.B1(n_1776),
.B2(n_1777),
.C1(n_1815),
.C2(n_1727),
.Y(n_1855)
);

INVx2_ASAP7_75t_L g1856 ( 
.A(n_1823),
.Y(n_1856)
);

AOI21xp33_ASAP7_75t_L g1857 ( 
.A1(n_1827),
.A2(n_1792),
.B(n_1805),
.Y(n_1857)
);

OR2x2_ASAP7_75t_L g1858 ( 
.A(n_1828),
.B(n_1817),
.Y(n_1858)
);

INVx3_ASAP7_75t_L g1859 ( 
.A(n_1823),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1822),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1824),
.Y(n_1861)
);

AOI22xp5_ASAP7_75t_L g1862 ( 
.A1(n_1849),
.A2(n_1792),
.B1(n_1677),
.B2(n_1707),
.Y(n_1862)
);

OAI321xp33_ASAP7_75t_L g1863 ( 
.A1(n_1839),
.A2(n_1754),
.A3(n_1774),
.B1(n_1769),
.B2(n_1704),
.C(n_1770),
.Y(n_1863)
);

INVx1_ASAP7_75t_SL g1864 ( 
.A(n_1838),
.Y(n_1864)
);

OR2x2_ASAP7_75t_L g1865 ( 
.A(n_1843),
.B(n_1769),
.Y(n_1865)
);

AOI222xp33_ASAP7_75t_L g1866 ( 
.A1(n_1848),
.A2(n_1792),
.B1(n_1768),
.B2(n_1777),
.C1(n_1776),
.C2(n_1774),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1830),
.Y(n_1867)
);

INVx2_ASAP7_75t_SL g1868 ( 
.A(n_1844),
.Y(n_1868)
);

INVx3_ASAP7_75t_L g1869 ( 
.A(n_1832),
.Y(n_1869)
);

AOI21xp33_ASAP7_75t_L g1870 ( 
.A1(n_1848),
.A2(n_1780),
.B(n_1770),
.Y(n_1870)
);

AOI322xp5_ASAP7_75t_L g1871 ( 
.A1(n_1864),
.A2(n_1846),
.A3(n_1847),
.B1(n_1835),
.B2(n_1834),
.C1(n_1840),
.C2(n_1837),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1851),
.Y(n_1872)
);

INVxp67_ASAP7_75t_L g1873 ( 
.A(n_1869),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1851),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1869),
.B(n_1841),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_L g1876 ( 
.A(n_1869),
.B(n_1850),
.Y(n_1876)
);

AOI332xp33_ASAP7_75t_L g1877 ( 
.A1(n_1860),
.A2(n_1845),
.A3(n_1826),
.B1(n_1833),
.B2(n_1778),
.B3(n_1780),
.C1(n_1784),
.C2(n_1829),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1853),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_SL g1879 ( 
.A(n_1863),
.B(n_1829),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1853),
.Y(n_1880)
);

INVxp33_ASAP7_75t_SL g1881 ( 
.A(n_1852),
.Y(n_1881)
);

OAI211xp5_ASAP7_75t_L g1882 ( 
.A1(n_1870),
.A2(n_1736),
.B(n_1704),
.C(n_1617),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1873),
.B(n_1868),
.Y(n_1883)
);

OAI221xp5_ASAP7_75t_SL g1884 ( 
.A1(n_1871),
.A2(n_1882),
.B1(n_1877),
.B2(n_1876),
.C(n_1875),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1881),
.B(n_1868),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1872),
.Y(n_1886)
);

NOR2xp33_ASAP7_75t_L g1887 ( 
.A(n_1879),
.B(n_1857),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1874),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1878),
.B(n_1856),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_SL g1890 ( 
.A(n_1879),
.B(n_1866),
.Y(n_1890)
);

OAI21xp33_ASAP7_75t_L g1891 ( 
.A1(n_1880),
.A2(n_1855),
.B(n_1854),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1872),
.Y(n_1892)
);

AO22x2_ASAP7_75t_L g1893 ( 
.A1(n_1890),
.A2(n_1856),
.B1(n_1859),
.B2(n_1867),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1889),
.Y(n_1894)
);

AOI221xp5_ASAP7_75t_L g1895 ( 
.A1(n_1884),
.A2(n_1861),
.B1(n_1859),
.B2(n_1858),
.C(n_1865),
.Y(n_1895)
);

NAND3xp33_ASAP7_75t_SL g1896 ( 
.A(n_1887),
.B(n_1862),
.C(n_1859),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1885),
.B(n_1721),
.Y(n_1897)
);

NAND4xp25_ASAP7_75t_L g1898 ( 
.A(n_1891),
.B(n_1524),
.C(n_1584),
.D(n_1670),
.Y(n_1898)
);

OAI322xp33_ASAP7_75t_L g1899 ( 
.A1(n_1897),
.A2(n_1883),
.A3(n_1894),
.B1(n_1886),
.B2(n_1888),
.C1(n_1892),
.C2(n_1884),
.Y(n_1899)
);

AOI321xp33_ASAP7_75t_L g1900 ( 
.A1(n_1895),
.A2(n_1584),
.A3(n_1677),
.B1(n_1778),
.B2(n_1585),
.C(n_1582),
.Y(n_1900)
);

NAND3xp33_ASAP7_75t_SL g1901 ( 
.A(n_1893),
.B(n_1574),
.C(n_1581),
.Y(n_1901)
);

AOI221xp5_ASAP7_75t_L g1902 ( 
.A1(n_1896),
.A2(n_1784),
.B1(n_1778),
.B2(n_1756),
.C(n_1752),
.Y(n_1902)
);

AOI211xp5_ASAP7_75t_L g1903 ( 
.A1(n_1898),
.A2(n_1581),
.B(n_1793),
.C(n_1736),
.Y(n_1903)
);

AOI211xp5_ASAP7_75t_L g1904 ( 
.A1(n_1896),
.A2(n_1581),
.B(n_1793),
.C(n_1677),
.Y(n_1904)
);

OR3x2_ASAP7_75t_L g1905 ( 
.A(n_1899),
.B(n_1582),
.C(n_1578),
.Y(n_1905)
);

NOR2x1_ASAP7_75t_L g1906 ( 
.A(n_1901),
.B(n_1716),
.Y(n_1906)
);

NAND4xp75_ASAP7_75t_L g1907 ( 
.A(n_1902),
.B(n_1773),
.C(n_1771),
.D(n_1763),
.Y(n_1907)
);

INVx2_ASAP7_75t_L g1908 ( 
.A(n_1904),
.Y(n_1908)
);

NAND2x1p5_ASAP7_75t_L g1909 ( 
.A(n_1900),
.B(n_1560),
.Y(n_1909)
);

OR2x2_ASAP7_75t_L g1910 ( 
.A(n_1909),
.B(n_1740),
.Y(n_1910)
);

OAI21xp33_ASAP7_75t_L g1911 ( 
.A1(n_1908),
.A2(n_1903),
.B(n_1773),
.Y(n_1911)
);

NAND3xp33_ASAP7_75t_L g1912 ( 
.A(n_1906),
.B(n_1773),
.C(n_1771),
.Y(n_1912)
);

AOI22xp5_ASAP7_75t_L g1913 ( 
.A1(n_1911),
.A2(n_1905),
.B1(n_1907),
.B2(n_1771),
.Y(n_1913)
);

AOI22xp5_ASAP7_75t_SL g1914 ( 
.A1(n_1913),
.A2(n_1910),
.B1(n_1709),
.B2(n_1574),
.Y(n_1914)
);

OAI22xp5_ASAP7_75t_L g1915 ( 
.A1(n_1914),
.A2(n_1912),
.B1(n_1752),
.B2(n_1763),
.Y(n_1915)
);

AOI22xp5_ASAP7_75t_L g1916 ( 
.A1(n_1914),
.A2(n_1763),
.B1(n_1756),
.B2(n_1740),
.Y(n_1916)
);

AOI22x1_ASAP7_75t_L g1917 ( 
.A1(n_1915),
.A2(n_1574),
.B1(n_1722),
.B2(n_1724),
.Y(n_1917)
);

XOR2x2_ASAP7_75t_L g1918 ( 
.A(n_1916),
.B(n_1573),
.Y(n_1918)
);

OAI21xp5_ASAP7_75t_SL g1919 ( 
.A1(n_1918),
.A2(n_1716),
.B(n_1724),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1917),
.Y(n_1920)
);

AOI21xp5_ASAP7_75t_L g1921 ( 
.A1(n_1920),
.A2(n_1725),
.B(n_1716),
.Y(n_1921)
);

HB1xp67_ASAP7_75t_L g1922 ( 
.A(n_1921),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1922),
.Y(n_1923)
);

OAI221xp5_ASAP7_75t_R g1924 ( 
.A1(n_1923),
.A2(n_1919),
.B1(n_1716),
.B2(n_1722),
.C(n_1724),
.Y(n_1924)
);

AOI211xp5_ASAP7_75t_L g1925 ( 
.A1(n_1924),
.A2(n_1560),
.B(n_1722),
.C(n_1720),
.Y(n_1925)
);


endmodule