module fake_jpeg_15438_n_242 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_242);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_242;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx3_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVxp33_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx4f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_40),
.Y(n_46)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx3_ASAP7_75t_SL g47 ( 
.A(n_37),
.Y(n_47)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_0),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_37),
.A2(n_20),
.B1(n_22),
.B2(n_18),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_48),
.A2(n_49),
.B1(n_33),
.B2(n_31),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_38),
.A2(n_22),
.B1(n_19),
.B2(n_21),
.Y(n_49)
);

NAND2xp33_ASAP7_75t_SL g51 ( 
.A(n_44),
.B(n_25),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_51),
.A2(n_31),
.B(n_27),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_39),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_59),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_43),
.A2(n_28),
.B1(n_21),
.B2(n_18),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_55),
.Y(n_95)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_35),
.Y(n_59)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_60),
.B(n_65),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_25),
.C(n_17),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_62),
.B(n_27),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_41),
.B(n_24),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_36),
.B(n_26),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_66),
.B(n_67),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_68),
.A2(n_81),
.B1(n_47),
.B2(n_85),
.Y(n_109)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_69),
.Y(n_105)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_72),
.B(n_73),
.Y(n_102)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

AOI21xp33_ASAP7_75t_L g74 ( 
.A1(n_46),
.A2(n_24),
.B(n_26),
.Y(n_74)
);

A2O1A1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_74),
.A2(n_92),
.B(n_17),
.C(n_23),
.Y(n_113)
);

INVx13_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_75),
.B(n_78),
.Y(n_110)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_76),
.Y(n_120)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_77),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_67),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_66),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_79),
.B(n_80),
.Y(n_118)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_82),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_83),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_104)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_85),
.Y(n_123)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_57),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_86),
.B(n_89),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_50),
.B(n_63),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_100),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_61),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_90),
.B(n_91),
.Y(n_108)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_64),
.A2(n_45),
.B1(n_42),
.B2(n_33),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_93),
.A2(n_96),
.B1(n_99),
.B2(n_5),
.Y(n_121)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_60),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_L g119 ( 
.A1(n_94),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_58),
.A2(n_45),
.B1(n_42),
.B2(n_32),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_62),
.Y(n_97)
);

NOR3xp33_ASAP7_75t_SL g125 ( 
.A(n_97),
.B(n_12),
.C(n_15),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_58),
.B(n_32),
.Y(n_98)
);

BUFx24_ASAP7_75t_SL g111 ( 
.A(n_98),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_50),
.A2(n_30),
.B1(n_1),
.B2(n_2),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_63),
.B(n_25),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_83),
.B(n_59),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_101),
.B(n_112),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_104),
.B(n_68),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_97),
.A2(n_47),
.B1(n_61),
.B2(n_4),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_107),
.A2(n_93),
.B(n_91),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_109),
.B(n_121),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_84),
.B(n_17),
.Y(n_112)
);

NOR2x1_ASAP7_75t_R g148 ( 
.A(n_113),
.B(n_125),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_100),
.B(n_23),
.C(n_34),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_115),
.B(n_117),
.C(n_99),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_75),
.B(n_34),
.C(n_11),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_119),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_83),
.B(n_6),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_122),
.B(n_124),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_92),
.B(n_6),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_127),
.B(n_134),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_105),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_128),
.B(n_129),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_71),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_105),
.Y(n_130)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_130),
.Y(n_157)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_116),
.Y(n_132)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_132),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_120),
.B(n_108),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_133),
.B(n_144),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_103),
.B(n_88),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_136),
.B(n_140),
.Y(n_161)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_137),
.Y(n_167)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_106),
.Y(n_138)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_138),
.Y(n_170)
);

NOR2x1_ASAP7_75t_L g139 ( 
.A(n_113),
.B(n_82),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_139),
.A2(n_149),
.B1(n_124),
.B2(n_95),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_103),
.B(n_87),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_107),
.Y(n_142)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_142),
.Y(n_172)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_121),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_143),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_110),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_101),
.B(n_96),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_145),
.B(n_86),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_118),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_146),
.B(n_147),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_120),
.B(n_77),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_119),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_150),
.Y(n_169)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_114),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_151),
.B(n_128),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_152),
.A2(n_131),
.B1(n_126),
.B2(n_127),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_139),
.A2(n_95),
.B(n_114),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_153),
.A2(n_159),
.B(n_158),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_142),
.A2(n_125),
.B1(n_117),
.B2(n_104),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_155),
.A2(n_154),
.B1(n_170),
.B2(n_172),
.Y(n_185)
);

A2O1A1O1Ixp25_ASAP7_75t_L g156 ( 
.A1(n_148),
.A2(n_122),
.B(n_111),
.C(n_112),
.D(n_115),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_156),
.A2(n_158),
.B(n_135),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_144),
.A2(n_123),
.B(n_70),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_143),
.A2(n_123),
.B(n_69),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_163),
.B(n_145),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_164),
.B(n_173),
.Y(n_181)
);

OA21x2_ASAP7_75t_L g168 ( 
.A1(n_149),
.A2(n_81),
.B(n_76),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_168),
.B(n_141),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_140),
.B(n_94),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_166),
.B(n_126),
.C(n_136),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_174),
.B(n_179),
.C(n_182),
.Y(n_193)
);

O2A1O1Ixp33_ASAP7_75t_L g202 ( 
.A1(n_175),
.A2(n_186),
.B(n_159),
.C(n_165),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_176),
.A2(n_185),
.B1(n_167),
.B2(n_160),
.Y(n_204)
);

NOR3xp33_ASAP7_75t_SL g177 ( 
.A(n_156),
.B(n_148),
.C(n_135),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_177),
.B(n_155),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_164),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_178),
.B(n_180),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_157),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_166),
.B(n_163),
.C(n_161),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_183),
.B(n_187),
.C(n_188),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_162),
.B(n_138),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_184),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_161),
.B(n_134),
.C(n_137),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_173),
.B(n_132),
.C(n_130),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_157),
.Y(n_189)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_189),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_170),
.B(n_151),
.Y(n_190)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_190),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g191 ( 
.A(n_168),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_191),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_191),
.A2(n_172),
.B1(n_169),
.B2(n_168),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_192),
.A2(n_198),
.B1(n_185),
.B2(n_186),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_183),
.B(n_153),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_195),
.B(n_197),
.C(n_205),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_179),
.B(n_174),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_200),
.B(n_204),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_202),
.A2(n_160),
.B(n_7),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_187),
.B(n_171),
.C(n_167),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_199),
.B(n_176),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_206),
.B(n_210),
.C(n_215),
.Y(n_221)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_207),
.Y(n_217)
);

NOR3xp33_ASAP7_75t_L g208 ( 
.A(n_200),
.B(n_177),
.C(n_181),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_208),
.B(n_212),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_204),
.B(n_188),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_211),
.A2(n_214),
.B1(n_9),
.B2(n_12),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_196),
.B(n_90),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_194),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_213),
.B(n_192),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_203),
.A2(n_6),
.B(n_7),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_199),
.B(n_11),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_208),
.B(n_201),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_218),
.B(n_220),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_222),
.B(n_14),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_216),
.B(n_205),
.C(n_193),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_223),
.B(n_224),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_216),
.B(n_193),
.C(n_197),
.Y(n_224)
);

AOI21x1_ASAP7_75t_L g225 ( 
.A1(n_218),
.A2(n_209),
.B(n_202),
.Y(n_225)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_225),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_221),
.B(n_210),
.C(n_195),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_226),
.B(n_230),
.Y(n_234)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_228),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_219),
.A2(n_217),
.B(n_209),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_227),
.B(n_15),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_231),
.B(n_16),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_234),
.A2(n_229),
.B(n_226),
.Y(n_235)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_235),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_236),
.B(n_237),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_232),
.B(n_16),
.C(n_9),
.Y(n_237)
);

BUFx24_ASAP7_75t_SL g240 ( 
.A(n_239),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_240),
.B(n_238),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_241),
.B(n_233),
.Y(n_242)
);


endmodule