module fake_aes_3998_n_685 (n_44, n_81, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_51, n_39, n_685);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_685;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_529;
wire n_455;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_420;
wire n_342;
wire n_423;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_409;
wire n_363;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_684;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g87 ( .A(n_9), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_17), .Y(n_88) );
CKINVDCx5p33_ASAP7_75t_R g89 ( .A(n_82), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_56), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_47), .Y(n_91) );
BUFx2_ASAP7_75t_L g92 ( .A(n_22), .Y(n_92) );
CKINVDCx20_ASAP7_75t_R g93 ( .A(n_5), .Y(n_93) );
CKINVDCx14_ASAP7_75t_R g94 ( .A(n_86), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_75), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_3), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_77), .Y(n_97) );
BUFx3_ASAP7_75t_L g98 ( .A(n_1), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_61), .Y(n_99) );
INVx2_ASAP7_75t_L g100 ( .A(n_45), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_34), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_30), .Y(n_102) );
INVx2_ASAP7_75t_L g103 ( .A(n_81), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_72), .Y(n_104) );
BUFx3_ASAP7_75t_L g105 ( .A(n_48), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_10), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_53), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_62), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g109 ( .A(n_2), .Y(n_109) );
INVxp67_ASAP7_75t_SL g110 ( .A(n_20), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_26), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_69), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g113 ( .A(n_78), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_23), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_0), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_38), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_73), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_50), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_6), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_41), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_15), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_3), .Y(n_122) );
AND2x4_ASAP7_75t_L g123 ( .A(n_92), .B(n_0), .Y(n_123) );
BUFx6f_ASAP7_75t_L g124 ( .A(n_105), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_98), .Y(n_125) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_105), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_113), .Y(n_127) );
OA21x2_ASAP7_75t_L g128 ( .A1(n_100), .A2(n_44), .B(n_84), .Y(n_128) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_100), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_98), .Y(n_130) );
AOI22xp5_ASAP7_75t_L g131 ( .A1(n_115), .A2(n_1), .B1(n_2), .B2(n_4), .Y(n_131) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_103), .Y(n_132) );
OAI22x1_ASAP7_75t_L g133 ( .A1(n_115), .A2(n_4), .B1(n_5), .B2(n_6), .Y(n_133) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_103), .Y(n_134) );
BUFx8_ASAP7_75t_L g135 ( .A(n_92), .Y(n_135) );
AND2x2_ASAP7_75t_L g136 ( .A(n_94), .B(n_7), .Y(n_136) );
INVx3_ASAP7_75t_L g137 ( .A(n_87), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_88), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_90), .Y(n_139) );
BUFx3_ASAP7_75t_L g140 ( .A(n_116), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_91), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_116), .Y(n_142) );
BUFx2_ASAP7_75t_L g143 ( .A(n_119), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_119), .B(n_7), .Y(n_144) );
AOI22xp33_ASAP7_75t_L g145 ( .A1(n_123), .A2(n_122), .B1(n_106), .B2(n_96), .Y(n_145) );
NOR2xp33_ASAP7_75t_SL g146 ( .A(n_135), .B(n_89), .Y(n_146) );
NAND2xp5_ASAP7_75t_SL g147 ( .A(n_135), .B(n_89), .Y(n_147) );
OAI22xp5_ASAP7_75t_L g148 ( .A1(n_143), .A2(n_121), .B1(n_93), .B2(n_109), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_129), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_129), .Y(n_150) );
INVx4_ASAP7_75t_L g151 ( .A(n_123), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_143), .B(n_121), .Y(n_152) );
NAND2xp33_ASAP7_75t_L g153 ( .A(n_138), .B(n_99), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_129), .Y(n_154) );
OAI22xp33_ASAP7_75t_SL g155 ( .A1(n_123), .A2(n_120), .B1(n_118), .B2(n_99), .Y(n_155) );
OAI22xp33_ASAP7_75t_L g156 ( .A1(n_131), .A2(n_120), .B1(n_118), .B2(n_107), .Y(n_156) );
BUFx3_ASAP7_75t_L g157 ( .A(n_124), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_129), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_129), .Y(n_159) );
BUFx4f_ASAP7_75t_L g160 ( .A(n_123), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_129), .Y(n_161) );
CKINVDCx5p33_ASAP7_75t_R g162 ( .A(n_135), .Y(n_162) );
CKINVDCx11_ASAP7_75t_R g163 ( .A(n_135), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_132), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_132), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_132), .Y(n_166) );
NAND2xp5_ASAP7_75t_SL g167 ( .A(n_138), .B(n_107), .Y(n_167) );
NAND2xp5_ASAP7_75t_SL g168 ( .A(n_139), .B(n_108), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_132), .Y(n_169) );
NAND2xp33_ASAP7_75t_SL g170 ( .A(n_136), .B(n_108), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_139), .B(n_111), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_132), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_141), .B(n_111), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_141), .B(n_112), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_125), .B(n_112), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_132), .Y(n_176) );
INVx4_ASAP7_75t_L g177 ( .A(n_128), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_134), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_134), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_151), .B(n_136), .Y(n_180) );
NAND2xp5_ASAP7_75t_SL g181 ( .A(n_160), .B(n_144), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g182 ( .A1(n_160), .A2(n_128), .B(n_125), .Y(n_182) );
AOI22xp33_ASAP7_75t_L g183 ( .A1(n_160), .A2(n_140), .B1(n_137), .B2(n_130), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_151), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_171), .B(n_137), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g186 ( .A(n_152), .B(n_137), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_151), .Y(n_187) );
BUFx6f_ASAP7_75t_L g188 ( .A(n_157), .Y(n_188) );
CKINVDCx6p67_ASAP7_75t_R g189 ( .A(n_163), .Y(n_189) );
AOI22xp33_ASAP7_75t_L g190 ( .A1(n_151), .A2(n_140), .B1(n_130), .B2(n_133), .Y(n_190) );
NOR2xp33_ASAP7_75t_SL g191 ( .A(n_146), .B(n_110), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_173), .B(n_142), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_157), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_157), .Y(n_194) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_155), .B(n_95), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_174), .B(n_142), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_175), .B(n_97), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g198 ( .A(n_167), .B(n_127), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_168), .B(n_101), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_145), .B(n_102), .Y(n_200) );
INVx3_ASAP7_75t_L g201 ( .A(n_177), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_153), .B(n_104), .Y(n_202) );
AOI22xp33_ASAP7_75t_L g203 ( .A1(n_155), .A2(n_133), .B1(n_126), .B2(n_124), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_149), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_170), .B(n_114), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_149), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_177), .Y(n_207) );
AOI22xp5_ASAP7_75t_L g208 ( .A1(n_146), .A2(n_117), .B1(n_134), .B2(n_128), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_147), .B(n_124), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_162), .B(n_124), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_162), .B(n_124), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_177), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g213 ( .A(n_156), .B(n_128), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_177), .B(n_126), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_148), .B(n_126), .Y(n_215) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_154), .B(n_126), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_179), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_154), .B(n_126), .Y(n_218) );
INVx2_ASAP7_75t_SL g219 ( .A(n_179), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_179), .Y(n_220) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_191), .B(n_124), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_180), .B(n_186), .Y(n_222) );
INVxp67_ASAP7_75t_L g223 ( .A(n_180), .Y(n_223) );
INVx4_ASAP7_75t_L g224 ( .A(n_189), .Y(n_224) );
OAI22xp5_ASAP7_75t_SL g225 ( .A1(n_190), .A2(n_8), .B1(n_9), .B2(n_10), .Y(n_225) );
AO21x1_ASAP7_75t_L g226 ( .A1(n_182), .A2(n_164), .B(n_176), .Y(n_226) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_191), .B(n_126), .Y(n_227) );
BUFx12f_ASAP7_75t_L g228 ( .A(n_189), .Y(n_228) );
AOI22xp33_ASAP7_75t_L g229 ( .A1(n_213), .A2(n_134), .B1(n_176), .B2(n_164), .Y(n_229) );
OAI22xp5_ASAP7_75t_L g230 ( .A1(n_203), .A2(n_183), .B1(n_200), .B2(n_185), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_205), .B(n_8), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_195), .B(n_134), .Y(n_232) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_207), .B(n_134), .Y(n_233) );
INVx4_ASAP7_75t_L g234 ( .A(n_188), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_184), .Y(n_235) );
NOR2x1_ASAP7_75t_L g236 ( .A(n_198), .B(n_158), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_207), .A2(n_178), .B(n_158), .Y(n_237) );
AOI221xp5_ASAP7_75t_L g238 ( .A1(n_197), .A2(n_159), .B1(n_178), .B2(n_169), .C(n_166), .Y(n_238) );
NOR2x1_ASAP7_75t_R g239 ( .A(n_215), .B(n_11), .Y(n_239) );
AO21x1_ASAP7_75t_L g240 ( .A1(n_208), .A2(n_159), .B(n_169), .Y(n_240) );
OAI22xp5_ASAP7_75t_L g241 ( .A1(n_192), .A2(n_172), .B1(n_166), .B2(n_165), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_212), .A2(n_172), .B(n_165), .Y(n_242) );
NOR2xp33_ASAP7_75t_SL g243 ( .A(n_212), .B(n_161), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_196), .B(n_11), .Y(n_244) );
INVx2_ASAP7_75t_L g245 ( .A(n_201), .Y(n_245) );
AND2x2_ASAP7_75t_L g246 ( .A(n_199), .B(n_12), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_202), .B(n_12), .Y(n_247) );
AOI21xp5_ASAP7_75t_L g248 ( .A1(n_214), .A2(n_161), .B(n_150), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_181), .B(n_13), .Y(n_249) );
NAND2xp5_ASAP7_75t_SL g250 ( .A(n_201), .B(n_150), .Y(n_250) );
AOI21xp5_ASAP7_75t_L g251 ( .A1(n_201), .A2(n_54), .B(n_83), .Y(n_251) );
AND2x2_ASAP7_75t_L g252 ( .A(n_184), .B(n_13), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_187), .B(n_14), .Y(n_253) );
INVx3_ASAP7_75t_L g254 ( .A(n_234), .Y(n_254) );
AO21x2_ASAP7_75t_L g255 ( .A1(n_240), .A2(n_208), .B(n_209), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_223), .B(n_187), .Y(n_256) );
NAND3xp33_ASAP7_75t_SL g257 ( .A(n_231), .B(n_244), .C(n_247), .Y(n_257) );
OAI21x1_ASAP7_75t_L g258 ( .A1(n_226), .A2(n_218), .B(n_210), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_222), .B(n_211), .Y(n_259) );
AOI22xp5_ASAP7_75t_L g260 ( .A1(n_231), .A2(n_193), .B1(n_194), .B2(n_217), .Y(n_260) );
OA21x2_ASAP7_75t_L g261 ( .A1(n_229), .A2(n_216), .B(n_220), .Y(n_261) );
AOI21xp5_ASAP7_75t_L g262 ( .A1(n_250), .A2(n_193), .B(n_194), .Y(n_262) );
AOI21xp5_ASAP7_75t_L g263 ( .A1(n_250), .A2(n_219), .B(n_220), .Y(n_263) );
NOR2x1_ASAP7_75t_SL g264 ( .A(n_228), .B(n_188), .Y(n_264) );
AND2x4_ASAP7_75t_L g265 ( .A(n_235), .B(n_188), .Y(n_265) );
AOI22xp5_ASAP7_75t_L g266 ( .A1(n_225), .A2(n_217), .B1(n_188), .B2(n_206), .Y(n_266) );
AOI21xp5_ASAP7_75t_L g267 ( .A1(n_237), .A2(n_219), .B(n_206), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_252), .Y(n_268) );
BUFx2_ASAP7_75t_L g269 ( .A(n_228), .Y(n_269) );
OR2x2_ASAP7_75t_L g270 ( .A(n_224), .B(n_188), .Y(n_270) );
AOI21xp5_ASAP7_75t_L g271 ( .A1(n_242), .A2(n_204), .B(n_55), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_253), .Y(n_272) );
AOI21x1_ASAP7_75t_SL g273 ( .A1(n_249), .A2(n_57), .B(n_85), .Y(n_273) );
OAI22xp5_ASAP7_75t_L g274 ( .A1(n_230), .A2(n_204), .B1(n_15), .B2(n_16), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_268), .B(n_246), .Y(n_275) );
NAND2x1p5_ASAP7_75t_L g276 ( .A(n_254), .B(n_234), .Y(n_276) );
AOI21xp5_ASAP7_75t_L g277 ( .A1(n_257), .A2(n_221), .B(n_227), .Y(n_277) );
OAI21xp5_ASAP7_75t_L g278 ( .A1(n_259), .A2(n_229), .B(n_233), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_256), .B(n_239), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_272), .B(n_236), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_265), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_258), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_258), .Y(n_283) );
OAI21x1_ASAP7_75t_L g284 ( .A1(n_273), .A2(n_221), .B(n_227), .Y(n_284) );
INVx6_ASAP7_75t_L g285 ( .A(n_270), .Y(n_285) );
AO21x2_ASAP7_75t_L g286 ( .A1(n_255), .A2(n_232), .B(n_251), .Y(n_286) );
OAI21x1_ASAP7_75t_L g287 ( .A1(n_271), .A2(n_248), .B(n_233), .Y(n_287) );
OAI21x1_ASAP7_75t_L g288 ( .A1(n_261), .A2(n_241), .B(n_245), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_261), .Y(n_289) );
AOI22xp5_ASAP7_75t_L g290 ( .A1(n_266), .A2(n_238), .B1(n_245), .B2(n_243), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_265), .Y(n_291) );
OR2x2_ASAP7_75t_L g292 ( .A(n_270), .B(n_14), .Y(n_292) );
OR2x2_ASAP7_75t_L g293 ( .A(n_254), .B(n_16), .Y(n_293) );
AOI21x1_ASAP7_75t_L g294 ( .A1(n_274), .A2(n_18), .B(n_19), .Y(n_294) );
AO21x2_ASAP7_75t_L g295 ( .A1(n_255), .A2(n_21), .B(n_24), .Y(n_295) );
OR2x2_ASAP7_75t_L g296 ( .A(n_254), .B(n_265), .Y(n_296) );
OAI21xp5_ASAP7_75t_L g297 ( .A1(n_260), .A2(n_25), .B(n_27), .Y(n_297) );
INVx3_ASAP7_75t_L g298 ( .A(n_276), .Y(n_298) );
AND2x2_ASAP7_75t_L g299 ( .A(n_281), .B(n_255), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_293), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_293), .Y(n_301) );
AND2x4_ASAP7_75t_L g302 ( .A(n_281), .B(n_264), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_289), .Y(n_303) );
BUFx3_ASAP7_75t_L g304 ( .A(n_276), .Y(n_304) );
AND2x4_ASAP7_75t_L g305 ( .A(n_291), .B(n_264), .Y(n_305) );
AO21x2_ASAP7_75t_L g306 ( .A1(n_282), .A2(n_262), .B(n_267), .Y(n_306) );
AOI22xp33_ASAP7_75t_L g307 ( .A1(n_279), .A2(n_261), .B1(n_269), .B2(n_263), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_291), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_289), .Y(n_309) );
AND2x4_ASAP7_75t_L g310 ( .A(n_282), .B(n_28), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_289), .Y(n_311) );
INVxp67_ASAP7_75t_L g312 ( .A(n_292), .Y(n_312) );
INVx3_ASAP7_75t_L g313 ( .A(n_276), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_282), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_283), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_283), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_283), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_288), .Y(n_318) );
OAI21x1_ASAP7_75t_L g319 ( .A1(n_284), .A2(n_29), .B(n_31), .Y(n_319) );
BUFx3_ASAP7_75t_L g320 ( .A(n_285), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_292), .Y(n_321) );
HB1xp67_ASAP7_75t_L g322 ( .A(n_285), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_288), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_296), .Y(n_324) );
INVx2_ASAP7_75t_SL g325 ( .A(n_285), .Y(n_325) );
BUFx2_ASAP7_75t_L g326 ( .A(n_285), .Y(n_326) );
OA21x2_ASAP7_75t_L g327 ( .A1(n_284), .A2(n_32), .B(n_33), .Y(n_327) );
OA21x2_ASAP7_75t_L g328 ( .A1(n_277), .A2(n_35), .B(n_36), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_295), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_296), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_295), .Y(n_331) );
INVxp67_ASAP7_75t_SL g332 ( .A(n_297), .Y(n_332) );
AND2x4_ASAP7_75t_L g333 ( .A(n_286), .B(n_37), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_295), .B(n_286), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_280), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_303), .Y(n_336) );
BUFx2_ASAP7_75t_L g337 ( .A(n_304), .Y(n_337) );
AND2x2_ASAP7_75t_L g338 ( .A(n_299), .B(n_286), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_311), .Y(n_339) );
INVx3_ASAP7_75t_L g340 ( .A(n_310), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_303), .Y(n_341) );
CKINVDCx5p33_ASAP7_75t_R g342 ( .A(n_304), .Y(n_342) );
NAND2x1_ASAP7_75t_L g343 ( .A(n_310), .B(n_290), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_311), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_303), .Y(n_345) );
INVx3_ASAP7_75t_L g346 ( .A(n_310), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_299), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_303), .Y(n_348) );
OR2x2_ASAP7_75t_L g349 ( .A(n_321), .B(n_275), .Y(n_349) );
OR2x2_ASAP7_75t_L g350 ( .A(n_321), .B(n_278), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_299), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_316), .Y(n_352) );
AND2x2_ASAP7_75t_L g353 ( .A(n_324), .B(n_294), .Y(n_353) );
BUFx2_ASAP7_75t_L g354 ( .A(n_304), .Y(n_354) );
INVx3_ASAP7_75t_L g355 ( .A(n_310), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_316), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_324), .B(n_294), .Y(n_357) );
BUFx3_ASAP7_75t_L g358 ( .A(n_298), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_330), .B(n_290), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_335), .B(n_287), .Y(n_360) );
INVx5_ASAP7_75t_SL g361 ( .A(n_302), .Y(n_361) );
OR2x2_ASAP7_75t_L g362 ( .A(n_312), .B(n_287), .Y(n_362) );
INVx2_ASAP7_75t_SL g363 ( .A(n_298), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_330), .B(n_308), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_308), .B(n_39), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_309), .B(n_40), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_317), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_317), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_309), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_312), .B(n_80), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_309), .Y(n_371) );
BUFx2_ASAP7_75t_L g372 ( .A(n_298), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_300), .B(n_42), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_314), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_300), .B(n_79), .Y(n_375) );
BUFx3_ASAP7_75t_L g376 ( .A(n_298), .Y(n_376) );
HB1xp67_ASAP7_75t_L g377 ( .A(n_322), .Y(n_377) );
INVx3_ASAP7_75t_L g378 ( .A(n_310), .Y(n_378) );
INVx1_ASAP7_75t_SL g379 ( .A(n_313), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_314), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_301), .B(n_43), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_314), .Y(n_382) );
OR2x2_ASAP7_75t_L g383 ( .A(n_301), .B(n_46), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_314), .Y(n_384) );
HB1xp67_ASAP7_75t_L g385 ( .A(n_322), .Y(n_385) );
INVx4_ASAP7_75t_L g386 ( .A(n_313), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_315), .Y(n_387) );
INVxp67_ASAP7_75t_L g388 ( .A(n_326), .Y(n_388) );
OAI22xp5_ASAP7_75t_L g389 ( .A1(n_313), .A2(n_49), .B1(n_51), .B2(n_52), .Y(n_389) );
BUFx3_ASAP7_75t_L g390 ( .A(n_313), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_315), .Y(n_391) );
NOR2x1_ASAP7_75t_L g392 ( .A(n_302), .B(n_58), .Y(n_392) );
BUFx3_ASAP7_75t_L g393 ( .A(n_326), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_315), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_315), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_334), .B(n_59), .Y(n_396) );
AND2x2_ASAP7_75t_L g397 ( .A(n_347), .B(n_334), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_339), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_347), .B(n_334), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_336), .Y(n_400) );
OR2x2_ASAP7_75t_L g401 ( .A(n_351), .B(n_326), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_339), .Y(n_402) );
INVx4_ASAP7_75t_L g403 ( .A(n_386), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_364), .B(n_325), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_344), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_351), .B(n_329), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_344), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_336), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_364), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_338), .B(n_329), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_349), .B(n_325), .Y(n_411) );
INVx4_ASAP7_75t_L g412 ( .A(n_386), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_352), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_341), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_338), .B(n_329), .Y(n_415) );
BUFx3_ASAP7_75t_L g416 ( .A(n_342), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_352), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_341), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_369), .B(n_329), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_369), .B(n_331), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_345), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_356), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_371), .B(n_331), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_345), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_371), .B(n_331), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_348), .Y(n_426) );
OR2x2_ASAP7_75t_L g427 ( .A(n_362), .B(n_307), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_348), .B(n_333), .Y(n_428) );
INVxp33_ASAP7_75t_L g429 ( .A(n_337), .Y(n_429) );
INVx1_ASAP7_75t_SL g430 ( .A(n_337), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_374), .Y(n_431) );
OR2x2_ASAP7_75t_L g432 ( .A(n_362), .B(n_307), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_356), .B(n_333), .Y(n_433) );
INVx2_ASAP7_75t_SL g434 ( .A(n_354), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_367), .B(n_333), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_349), .B(n_325), .Y(n_436) );
HB1xp67_ASAP7_75t_L g437 ( .A(n_377), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_368), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_368), .B(n_333), .Y(n_439) );
HB1xp67_ASAP7_75t_L g440 ( .A(n_385), .Y(n_440) );
OR2x2_ASAP7_75t_L g441 ( .A(n_360), .B(n_318), .Y(n_441) );
AND2x4_ASAP7_75t_L g442 ( .A(n_386), .B(n_333), .Y(n_442) );
INVx3_ASAP7_75t_L g443 ( .A(n_386), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_380), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_359), .B(n_302), .Y(n_445) );
NAND2xp5_ASAP7_75t_SL g446 ( .A(n_392), .B(n_302), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_374), .Y(n_447) );
BUFx2_ASAP7_75t_L g448 ( .A(n_354), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_380), .Y(n_449) );
INVx4_ASAP7_75t_L g450 ( .A(n_358), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_384), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_384), .B(n_323), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_387), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_359), .B(n_302), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_387), .B(n_318), .Y(n_455) );
BUFx3_ASAP7_75t_L g456 ( .A(n_372), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_382), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_391), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_382), .Y(n_459) );
OR2x2_ASAP7_75t_L g460 ( .A(n_350), .B(n_318), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_350), .Y(n_461) );
INVxp67_ASAP7_75t_SL g462 ( .A(n_394), .Y(n_462) );
NAND3xp33_ASAP7_75t_L g463 ( .A(n_370), .B(n_305), .C(n_320), .Y(n_463) );
INVx2_ASAP7_75t_SL g464 ( .A(n_390), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_388), .B(n_305), .Y(n_465) );
OR2x2_ASAP7_75t_L g466 ( .A(n_394), .B(n_323), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_383), .Y(n_467) );
OR2x2_ASAP7_75t_L g468 ( .A(n_395), .B(n_323), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_395), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_353), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_353), .B(n_306), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_393), .B(n_320), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_357), .B(n_306), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_357), .B(n_306), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_383), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_365), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_396), .B(n_306), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_340), .B(n_332), .Y(n_478) );
INVx1_ASAP7_75t_SL g479 ( .A(n_430), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_437), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_440), .Y(n_481) );
OR2x2_ASAP7_75t_L g482 ( .A(n_409), .B(n_361), .Y(n_482) );
OR2x2_ASAP7_75t_L g483 ( .A(n_461), .B(n_361), .Y(n_483) );
INVxp67_ASAP7_75t_SL g484 ( .A(n_462), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_398), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_402), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_405), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_397), .B(n_393), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_407), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_397), .B(n_361), .Y(n_490) );
NAND2x1_ASAP7_75t_SL g491 ( .A(n_403), .B(n_392), .Y(n_491) );
AND3x2_ASAP7_75t_L g492 ( .A(n_448), .B(n_373), .C(n_381), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_399), .B(n_343), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_399), .B(n_343), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_413), .B(n_379), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_417), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_422), .B(n_340), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_438), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_470), .B(n_340), .Y(n_499) );
HB1xp67_ASAP7_75t_L g500 ( .A(n_434), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_445), .B(n_454), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_400), .Y(n_502) );
AND2x4_ASAP7_75t_L g503 ( .A(n_403), .B(n_390), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_470), .B(n_340), .Y(n_504) );
OR2x2_ASAP7_75t_L g505 ( .A(n_404), .B(n_361), .Y(n_505) );
INVx1_ASAP7_75t_SL g506 ( .A(n_416), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_444), .B(n_346), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_449), .B(n_346), .Y(n_508) );
NAND2x1p5_ASAP7_75t_L g509 ( .A(n_403), .B(n_358), .Y(n_509) );
OR2x2_ASAP7_75t_L g510 ( .A(n_401), .B(n_390), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_411), .Y(n_511) );
NAND2x1p5_ASAP7_75t_L g512 ( .A(n_412), .B(n_376), .Y(n_512) );
OR2x2_ASAP7_75t_L g513 ( .A(n_401), .B(n_346), .Y(n_513) );
BUFx2_ASAP7_75t_L g514 ( .A(n_412), .Y(n_514) );
NOR2xp67_ASAP7_75t_L g515 ( .A(n_412), .B(n_378), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_472), .B(n_363), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_436), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_451), .B(n_355), .Y(n_518) );
AND2x2_ASAP7_75t_SL g519 ( .A(n_442), .B(n_378), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_453), .B(n_355), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_400), .Y(n_521) );
INVx2_ASAP7_75t_L g522 ( .A(n_408), .Y(n_522) );
BUFx3_ASAP7_75t_L g523 ( .A(n_450), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_410), .B(n_355), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_458), .Y(n_525) );
INVx2_ASAP7_75t_SL g526 ( .A(n_450), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_460), .Y(n_527) );
HB1xp67_ASAP7_75t_L g528 ( .A(n_456), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_406), .B(n_378), .Y(n_529) );
NOR2xp33_ASAP7_75t_L g530 ( .A(n_465), .B(n_320), .Y(n_530) );
NOR2x1p5_ASAP7_75t_L g531 ( .A(n_443), .B(n_375), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_410), .B(n_366), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_415), .B(n_366), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_415), .B(n_381), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_460), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_450), .B(n_373), .Y(n_536) );
INVx2_ASAP7_75t_L g537 ( .A(n_414), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_406), .B(n_471), .Y(n_538) );
AND2x4_ASAP7_75t_L g539 ( .A(n_442), .B(n_319), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_429), .B(n_327), .Y(n_540) );
AND2x4_ASAP7_75t_L g541 ( .A(n_442), .B(n_319), .Y(n_541) );
NOR2xp33_ASAP7_75t_L g542 ( .A(n_476), .B(n_389), .Y(n_542) );
NOR2xp33_ASAP7_75t_L g543 ( .A(n_467), .B(n_60), .Y(n_543) );
NAND4xp25_ASAP7_75t_L g544 ( .A(n_463), .B(n_427), .C(n_432), .D(n_446), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_475), .Y(n_545) );
HB1xp67_ASAP7_75t_L g546 ( .A(n_456), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_418), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_471), .B(n_328), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_429), .B(n_327), .Y(n_549) );
OR2x2_ASAP7_75t_L g550 ( .A(n_427), .B(n_327), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_418), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_433), .B(n_327), .Y(n_552) );
INVx2_ASAP7_75t_L g553 ( .A(n_421), .Y(n_553) );
INVxp67_ASAP7_75t_L g554 ( .A(n_464), .Y(n_554) );
INVx2_ASAP7_75t_L g555 ( .A(n_421), .Y(n_555) );
INVxp67_ASAP7_75t_SL g556 ( .A(n_424), .Y(n_556) );
INVx2_ASAP7_75t_L g557 ( .A(n_424), .Y(n_557) );
HB1xp67_ASAP7_75t_L g558 ( .A(n_484), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_480), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_479), .B(n_435), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_479), .B(n_435), .Y(n_561) );
NAND3xp33_ASAP7_75t_L g562 ( .A(n_544), .B(n_432), .C(n_446), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_481), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_485), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_486), .Y(n_565) );
INVx2_ASAP7_75t_L g566 ( .A(n_514), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_487), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_527), .B(n_473), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_489), .Y(n_569) );
INVx2_ASAP7_75t_SL g570 ( .A(n_506), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_496), .Y(n_571) );
HB1xp67_ASAP7_75t_L g572 ( .A(n_500), .Y(n_572) );
OR2x2_ASAP7_75t_L g573 ( .A(n_538), .B(n_441), .Y(n_573) );
OR2x2_ASAP7_75t_L g574 ( .A(n_538), .B(n_488), .Y(n_574) );
INVx2_ASAP7_75t_L g575 ( .A(n_523), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_535), .B(n_473), .Y(n_576) );
AOI311xp33_ASAP7_75t_L g577 ( .A1(n_511), .A2(n_477), .A3(n_474), .B(n_439), .C(n_478), .Y(n_577) );
NOR2xp33_ASAP7_75t_L g578 ( .A(n_517), .B(n_474), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_490), .B(n_478), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_545), .B(n_419), .Y(n_580) );
OR2x2_ASAP7_75t_L g581 ( .A(n_488), .B(n_441), .Y(n_581) );
OAI21xp33_ASAP7_75t_L g582 ( .A1(n_544), .A2(n_428), .B(n_419), .Y(n_582) );
OR2x2_ASAP7_75t_L g583 ( .A(n_529), .B(n_469), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_501), .B(n_428), .Y(n_584) );
OAI31xp33_ASAP7_75t_L g585 ( .A1(n_531), .A2(n_452), .A3(n_455), .B(n_425), .Y(n_585) );
OAI21xp5_ASAP7_75t_L g586 ( .A1(n_491), .A2(n_328), .B(n_319), .Y(n_586) );
INVx2_ASAP7_75t_L g587 ( .A(n_526), .Y(n_587) );
INVx1_ASAP7_75t_SL g588 ( .A(n_528), .Y(n_588) );
INVxp33_ASAP7_75t_SL g589 ( .A(n_546), .Y(n_589) );
AOI21xp5_ASAP7_75t_L g590 ( .A1(n_515), .A2(n_469), .B(n_426), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g591 ( .A(n_554), .B(n_447), .Y(n_591) );
OAI221xp5_ASAP7_75t_L g592 ( .A1(n_542), .A2(n_431), .B1(n_426), .B2(n_459), .C(n_457), .Y(n_592) );
OR2x2_ASAP7_75t_L g593 ( .A(n_529), .B(n_447), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_498), .Y(n_594) );
INVx1_ASAP7_75t_SL g595 ( .A(n_503), .Y(n_595) );
AND2x2_ASAP7_75t_L g596 ( .A(n_524), .B(n_420), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_525), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_551), .B(n_423), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_495), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_516), .B(n_455), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_532), .B(n_452), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_495), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_502), .B(n_431), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_497), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_533), .B(n_468), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_507), .Y(n_606) );
AOI22xp5_ASAP7_75t_L g607 ( .A1(n_530), .A2(n_328), .B1(n_466), .B2(n_468), .Y(n_607) );
INVx2_ASAP7_75t_L g608 ( .A(n_521), .Y(n_608) );
INVx2_ASAP7_75t_SL g609 ( .A(n_503), .Y(n_609) );
INVx3_ASAP7_75t_L g610 ( .A(n_509), .Y(n_610) );
NAND2xp5_ASAP7_75t_SL g611 ( .A(n_519), .B(n_466), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_508), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_508), .Y(n_613) );
INVx2_ASAP7_75t_L g614 ( .A(n_522), .Y(n_614) );
OAI22xp33_ASAP7_75t_L g615 ( .A1(n_610), .A2(n_512), .B1(n_509), .B2(n_505), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_604), .B(n_518), .Y(n_616) );
INVx1_ASAP7_75t_SL g617 ( .A(n_588), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_558), .Y(n_618) );
INVx2_ASAP7_75t_L g619 ( .A(n_588), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_599), .Y(n_620) );
INVx1_ASAP7_75t_SL g621 ( .A(n_589), .Y(n_621) );
AOI222xp33_ASAP7_75t_L g622 ( .A1(n_562), .A2(n_548), .B1(n_493), .B2(n_494), .C1(n_536), .C2(n_540), .Y(n_622) );
AOI21xp5_ASAP7_75t_L g623 ( .A1(n_585), .A2(n_512), .B(n_556), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_602), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_606), .B(n_520), .Y(n_625) );
OAI221xp5_ASAP7_75t_L g626 ( .A1(n_577), .A2(n_493), .B1(n_550), .B2(n_548), .C(n_482), .Y(n_626) );
OAI22xp33_ASAP7_75t_L g627 ( .A1(n_610), .A2(n_483), .B1(n_510), .B2(n_513), .Y(n_627) );
OAI21xp33_ASAP7_75t_L g628 ( .A1(n_582), .A2(n_499), .B(n_504), .Y(n_628) );
OR2x2_ASAP7_75t_L g629 ( .A(n_573), .B(n_499), .Y(n_629) );
OAI21xp5_ASAP7_75t_L g630 ( .A1(n_585), .A2(n_543), .B(n_549), .Y(n_630) );
NAND2x1_ASAP7_75t_L g631 ( .A(n_609), .B(n_539), .Y(n_631) );
INVx2_ASAP7_75t_L g632 ( .A(n_572), .Y(n_632) );
OAI22xp33_ASAP7_75t_L g633 ( .A1(n_595), .A2(n_492), .B1(n_539), .B2(n_541), .Y(n_633) );
AOI22xp5_ASAP7_75t_L g634 ( .A1(n_578), .A2(n_541), .B1(n_534), .B2(n_552), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_581), .Y(n_635) );
INVx2_ASAP7_75t_L g636 ( .A(n_583), .Y(n_636) );
NAND2xp5_ASAP7_75t_SL g637 ( .A(n_570), .B(n_557), .Y(n_637) );
AOI21xp5_ASAP7_75t_L g638 ( .A1(n_611), .A2(n_555), .B(n_553), .Y(n_638) );
OAI21xp33_ASAP7_75t_L g639 ( .A1(n_568), .A2(n_547), .B(n_537), .Y(n_639) );
AO21x1_ASAP7_75t_L g640 ( .A1(n_590), .A2(n_328), .B(n_63), .Y(n_640) );
XNOR2x2_ASAP7_75t_L g641 ( .A(n_595), .B(n_592), .Y(n_641) );
OAI221xp5_ASAP7_75t_L g642 ( .A1(n_607), .A2(n_328), .B1(n_64), .B2(n_65), .C(n_66), .Y(n_642) );
OAI221xp5_ASAP7_75t_L g643 ( .A1(n_621), .A2(n_566), .B1(n_563), .B2(n_559), .C(n_575), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_618), .Y(n_644) );
OAI211xp5_ASAP7_75t_SL g645 ( .A1(n_621), .A2(n_587), .B(n_564), .C(n_565), .Y(n_645) );
AOI31xp33_ASAP7_75t_L g646 ( .A1(n_623), .A2(n_586), .A3(n_574), .B(n_561), .Y(n_646) );
AOI22xp5_ASAP7_75t_L g647 ( .A1(n_622), .A2(n_613), .B1(n_612), .B2(n_576), .Y(n_647) );
OAI32xp33_ASAP7_75t_L g648 ( .A1(n_617), .A2(n_576), .A3(n_568), .B1(n_580), .B2(n_593), .Y(n_648) );
OAI322xp33_ASAP7_75t_L g649 ( .A1(n_641), .A2(n_580), .A3(n_594), .B1(n_567), .B2(n_569), .C1(n_571), .C2(n_597), .Y(n_649) );
HB1xp67_ASAP7_75t_L g650 ( .A(n_617), .Y(n_650) );
AOI21xp33_ASAP7_75t_SL g651 ( .A1(n_633), .A2(n_591), .B(n_586), .Y(n_651) );
AOI211xp5_ASAP7_75t_L g652 ( .A1(n_615), .A2(n_560), .B(n_579), .C(n_598), .Y(n_652) );
AOI21xp33_ASAP7_75t_L g653 ( .A1(n_622), .A2(n_603), .B(n_598), .Y(n_653) );
AOI322xp5_ASAP7_75t_L g654 ( .A1(n_628), .A2(n_601), .A3(n_605), .B1(n_584), .B2(n_596), .C1(n_600), .C2(n_614), .Y(n_654) );
AOI221xp5_ASAP7_75t_L g655 ( .A1(n_626), .A2(n_608), .B1(n_68), .B2(n_70), .C(n_71), .Y(n_655) );
AOI22xp5_ASAP7_75t_L g656 ( .A1(n_630), .A2(n_67), .B1(n_74), .B2(n_76), .Y(n_656) );
OAI21xp33_ASAP7_75t_SL g657 ( .A1(n_637), .A2(n_634), .B(n_619), .Y(n_657) );
OAI21xp5_ASAP7_75t_L g658 ( .A1(n_631), .A2(n_632), .B(n_638), .Y(n_658) );
OAI211xp5_ASAP7_75t_SL g659 ( .A1(n_639), .A2(n_642), .B(n_620), .C(n_624), .Y(n_659) );
NOR2xp33_ASAP7_75t_L g660 ( .A(n_635), .B(n_616), .Y(n_660) );
OAI221xp5_ASAP7_75t_L g661 ( .A1(n_625), .A2(n_629), .B1(n_636), .B2(n_627), .C(n_640), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_618), .Y(n_662) );
INVxp67_ASAP7_75t_L g663 ( .A(n_621), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_618), .Y(n_664) );
OAI221xp5_ASAP7_75t_L g665 ( .A1(n_628), .A2(n_621), .B1(n_630), .B2(n_577), .C(n_585), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_618), .Y(n_666) );
OAI22xp5_ASAP7_75t_L g667 ( .A1(n_665), .A2(n_652), .B1(n_646), .B2(n_647), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_650), .Y(n_668) );
NOR2xp33_ASAP7_75t_L g669 ( .A(n_663), .B(n_657), .Y(n_669) );
AOI211x1_ASAP7_75t_SL g670 ( .A1(n_659), .A2(n_658), .B(n_645), .C(n_653), .Y(n_670) );
O2A1O1Ixp33_ASAP7_75t_L g671 ( .A1(n_649), .A2(n_661), .B(n_651), .C(n_643), .Y(n_671) );
INVxp33_ASAP7_75t_SL g672 ( .A(n_669), .Y(n_672) );
NOR2x1_ASAP7_75t_L g673 ( .A(n_671), .B(n_667), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_670), .B(n_654), .Y(n_674) );
INVx2_ASAP7_75t_L g675 ( .A(n_673), .Y(n_675) );
AND3x4_ASAP7_75t_L g676 ( .A(n_672), .B(n_655), .C(n_668), .Y(n_676) );
INVx2_ASAP7_75t_L g677 ( .A(n_675), .Y(n_677) );
AND2x2_ASAP7_75t_SL g678 ( .A(n_676), .B(n_674), .Y(n_678) );
INVx3_ASAP7_75t_L g679 ( .A(n_677), .Y(n_679) );
XNOR2x1_ASAP7_75t_L g680 ( .A(n_678), .B(n_656), .Y(n_680) );
INVxp67_ASAP7_75t_SL g681 ( .A(n_679), .Y(n_681) );
OA22x2_ASAP7_75t_L g682 ( .A1(n_681), .A2(n_679), .B1(n_680), .B2(n_644), .Y(n_682) );
OR2x6_ASAP7_75t_L g683 ( .A(n_682), .B(n_666), .Y(n_683) );
AOI21xp5_ASAP7_75t_L g684 ( .A1(n_683), .A2(n_643), .B(n_648), .Y(n_684) );
AOI22xp33_ASAP7_75t_SL g685 ( .A1(n_684), .A2(n_664), .B1(n_662), .B2(n_660), .Y(n_685) );
endmodule