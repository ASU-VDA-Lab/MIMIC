module real_jpeg_1002_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_288;
wire n_249;
wire n_176;
wire n_166;
wire n_292;
wire n_221;
wire n_215;
wire n_286;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_271;
wire n_281;
wire n_131;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_293;
wire n_48;
wire n_164;
wire n_184;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_290;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_285;
wire n_172;
wire n_45;
wire n_211;
wire n_268;
wire n_42;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_258;
wire n_195;
wire n_110;
wire n_205;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_279;
wire n_59;
wire n_169;
wire n_128;
wire n_295;
wire n_244;
wire n_179;
wire n_167;
wire n_202;
wire n_133;
wire n_213;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_273;
wire n_89;
wire n_16;

INVx2_ASAP7_75t_L g73 ( 
.A(n_0),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_1),
.Y(n_97)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_2),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_3),
.A2(n_21),
.B1(n_22),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_3),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_3),
.A2(n_51),
.B1(n_60),
.B2(n_61),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_3),
.A2(n_33),
.B1(n_34),
.B2(n_51),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_3),
.A2(n_51),
.B1(n_70),
.B2(n_71),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_3),
.B(n_29),
.C(n_34),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_3),
.B(n_32),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_3),
.B(n_57),
.C(n_61),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_3),
.B(n_97),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_3),
.B(n_68),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_3),
.B(n_69),
.C(n_71),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_3),
.B(n_63),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_4),
.A2(n_21),
.B1(n_22),
.B2(n_49),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g49 ( 
.A(n_4),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_4),
.A2(n_49),
.B1(n_60),
.B2(n_61),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_4),
.A2(n_33),
.B1(n_34),
.B2(n_49),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_4),
.A2(n_49),
.B1(n_70),
.B2(n_71),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_5),
.A2(n_21),
.B1(n_22),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_5),
.Y(n_40)
);

OAI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_5),
.A2(n_33),
.B1(n_34),
.B2(n_40),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_5),
.A2(n_40),
.B1(n_70),
.B2(n_71),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_5),
.A2(n_40),
.B1(n_60),
.B2(n_61),
.Y(n_115)
);

BUFx4f_ASAP7_75t_L g57 ( 
.A(n_6),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g20 ( 
.A1(n_7),
.A2(n_21),
.B1(n_22),
.B2(n_25),
.Y(n_20)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_7),
.A2(n_25),
.B1(n_33),
.B2(n_34),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_7),
.A2(n_25),
.B1(n_60),
.B2(n_61),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_7),
.A2(n_25),
.B1(n_70),
.B2(n_71),
.Y(n_100)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g69 ( 
.A(n_9),
.Y(n_69)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_SL g294 ( 
.A(n_12),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_12),
.B(n_296),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_13),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_294),
.B(n_295),
.Y(n_14)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_42),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_41),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_38),
.Y(n_17)
);

OR2x2_ASAP7_75t_L g41 ( 
.A(n_18),
.B(n_38),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_26),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_20),
.A2(n_27),
.B1(n_37),
.B2(n_39),
.Y(n_38)
);

O2A1O1Ixp33_ASAP7_75t_L g28 ( 
.A1(n_21),
.A2(n_29),
.B(n_31),
.C(n_32),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_21),
.B(n_29),
.Y(n_31)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_22),
.B(n_158),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_26),
.B(n_50),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_37),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_28),
.A2(n_32),
.B1(n_47),
.B2(n_50),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_28),
.B(n_50),
.Y(n_81)
);

AO22x1_ASAP7_75t_SL g32 ( 
.A1(n_29),
.A2(n_33),
.B1(n_34),
.B2(n_36),
.Y(n_32)
);

INVx2_ASAP7_75t_SL g36 ( 
.A(n_29),
.Y(n_36)
);

BUFx4f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_33),
.A2(n_34),
.B1(n_57),
.B2(n_58),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_34),
.B(n_212),
.Y(n_211)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_37),
.A2(n_39),
.B(n_81),
.Y(n_80)
);

OA21x2_ASAP7_75t_L g130 ( 
.A1(n_37),
.A2(n_48),
.B(n_81),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_38),
.B(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_38),
.B(n_44),
.Y(n_293)
);

AO21x1_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_82),
.B(n_293),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_78),
.C(n_80),
.Y(n_44)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_45),
.B(n_290),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_52),
.C(n_65),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_46),
.A2(n_103),
.B1(n_107),
.B2(n_108),
.Y(n_102)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_46),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_46),
.A2(n_108),
.B1(n_145),
.B2(n_163),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_46),
.B(n_145),
.C(n_155),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_46),
.A2(n_108),
.B1(n_280),
.B2(n_281),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_52),
.A2(n_65),
.B1(n_267),
.B2(n_282),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_52),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_54),
.B1(n_63),
.B2(n_64),
.Y(n_52)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_53),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_54),
.A2(n_63),
.B1(n_104),
.B2(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_55),
.B(n_59),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_55),
.B(n_106),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_55),
.A2(n_59),
.B(n_106),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_56),
.B(n_59),
.Y(n_55)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_57),
.Y(n_58)
);

AOI22x1_ASAP7_75t_L g59 ( 
.A1(n_57),
.A2(n_58),
.B1(n_60),
.B2(n_61),
.Y(n_59)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_59),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_59),
.A2(n_269),
.B(n_270),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_60),
.A2(n_61),
.B1(n_69),
.B2(n_74),
.Y(n_76)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_61),
.B(n_229),
.Y(n_228)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

AO21x1_ASAP7_75t_L g103 ( 
.A1(n_63),
.A2(n_104),
.B(n_105),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_79),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_65),
.A2(n_267),
.B1(n_268),
.B2(n_271),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_65),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_65),
.B(n_130),
.C(n_268),
.Y(n_283)
);

AND2x2_ASAP7_75t_SL g65 ( 
.A(n_66),
.B(n_77),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_75),
.Y(n_66)
);

OA22x2_ASAP7_75t_L g91 ( 
.A1(n_67),
.A2(n_75),
.B1(n_92),
.B2(n_93),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_67),
.A2(n_115),
.B(n_116),
.Y(n_114)
);

OA22x2_ASAP7_75t_L g127 ( 
.A1(n_67),
.A2(n_75),
.B1(n_92),
.B2(n_93),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_67),
.A2(n_75),
.B(n_93),
.Y(n_171)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_68),
.B(n_76),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_68),
.A2(n_77),
.B1(n_118),
.B2(n_144),
.Y(n_143)
);

AO22x1_ASAP7_75t_SL g68 ( 
.A1(n_69),
.A2(n_70),
.B1(n_71),
.B2(n_74),
.Y(n_68)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_69),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_70),
.B(n_97),
.Y(n_96)
);

INVx3_ASAP7_75t_SL g70 ( 
.A(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_71),
.B(n_222),
.Y(n_221)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_75),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_78),
.B(n_80),
.Y(n_290)
);

OAI21x1_ASAP7_75t_SL g82 ( 
.A1(n_83),
.A2(n_288),
.B(n_292),
.Y(n_82)
);

AOI21x1_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_259),
.B(n_285),
.Y(n_83)
);

OAI21x1_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_149),
.B(n_258),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_131),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_86),
.B(n_131),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_109),
.C(n_120),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_87),
.B(n_109),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_89),
.B1(n_101),
.B2(n_102),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_88),
.B(n_103),
.C(n_108),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_94),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_90),
.A2(n_91),
.B1(n_94),
.B2(n_195),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_90),
.A2(n_91),
.B1(n_236),
.B2(n_237),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_90),
.A2(n_91),
.B1(n_209),
.B2(n_249),
.Y(n_248)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_91),
.B(n_204),
.C(n_209),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_91),
.B(n_160),
.C(n_236),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_93),
.Y(n_117)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_94),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_98),
.B1(n_99),
.B2(n_100),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_95),
.B(n_99),
.Y(n_112)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_96),
.B(n_125),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_96),
.A2(n_97),
.B1(n_125),
.B2(n_161),
.Y(n_160)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_97),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_98),
.A2(n_99),
.B(n_124),
.Y(n_123)
);

OA21x2_ASAP7_75t_L g180 ( 
.A1(n_99),
.A2(n_124),
.B(n_181),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_100),
.B(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_103),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_103),
.B(n_129),
.C(n_171),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_103),
.A2(n_107),
.B1(n_171),
.B2(n_176),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_103),
.A2(n_107),
.B1(n_126),
.B2(n_127),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_103),
.B(n_126),
.C(n_244),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_105),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_106),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_113),
.B1(n_114),
.B2(n_119),
.Y(n_109)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_110),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_110),
.B(n_114),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_110),
.A2(n_119),
.B1(n_139),
.B2(n_140),
.Y(n_138)
);

INVxp33_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_112),
.B(n_125),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_115),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_118),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_119),
.A2(n_135),
.B(n_140),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_120),
.B(n_256),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_128),
.C(n_129),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_121),
.A2(n_122),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_126),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_123),
.A2(n_126),
.B1(n_127),
.B2(n_168),
.Y(n_167)
);

CKINVDCx14_ASAP7_75t_R g168 ( 
.A(n_123),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_126),
.A2(n_127),
.B1(n_228),
.B2(n_230),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_126),
.B(n_230),
.Y(n_238)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_128),
.A2(n_129),
.B1(n_130),
.B2(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_128),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_129),
.A2(n_130),
.B1(n_174),
.B2(n_175),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_129),
.A2(n_130),
.B1(n_265),
.B2(n_266),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_129),
.A2(n_130),
.B1(n_278),
.B2(n_279),
.Y(n_277)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_130),
.B(n_279),
.C(n_283),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_148),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_133),
.A2(n_134),
.B1(n_141),
.B2(n_142),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_134),
.B(n_141),
.C(n_148),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_136),
.B1(n_137),
.B2(n_138),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_139),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_145),
.B(n_147),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_143),
.B(n_145),
.Y(n_147)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_145),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_145),
.B(n_179),
.C(n_180),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_145),
.A2(n_163),
.B1(n_205),
.B2(n_208),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_147),
.A2(n_263),
.B1(n_264),
.B2(n_272),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_147),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_253),
.B(n_257),
.Y(n_149)
);

OAI211xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_182),
.B(n_196),
.C(n_197),
.Y(n_150)
);

OR2x2_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_172),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_152),
.B(n_172),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_154),
.B1(n_164),
.B2(n_165),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_153),
.B(n_167),
.C(n_169),
.Y(n_184)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_155),
.B(n_162),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_159),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_156),
.A2(n_157),
.B1(n_159),
.B2(n_160),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_159),
.A2(n_160),
.B1(n_234),
.B2(n_235),
.Y(n_233)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_160),
.B(n_224),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_160),
.B(n_224),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_161),
.Y(n_181)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_167),
.B1(n_169),
.B2(n_170),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_171),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_177),
.C(n_178),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_173),
.B(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_177),
.B(n_178),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_179),
.A2(n_180),
.B1(n_206),
.B2(n_207),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_179),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_180),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_180),
.B(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

NAND3xp33_ASAP7_75t_SL g197 ( 
.A(n_183),
.B(n_198),
.C(n_199),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

OR2x2_ASAP7_75t_L g196 ( 
.A(n_184),
.B(n_185),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_186),
.B(n_188),
.C(n_194),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_188),
.A2(n_189),
.B1(n_193),
.B2(n_194),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

OAI21x1_ASAP7_75t_SL g199 ( 
.A1(n_200),
.A2(n_215),
.B(n_252),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_201),
.B(n_203),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_201),
.B(n_203),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_204),
.B(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_205),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_207),
.B(n_227),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_207),
.B(n_227),
.Y(n_231)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_209),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_213),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_210),
.A2(n_211),
.B1(n_213),
.B2(n_214),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_216),
.A2(n_246),
.B(n_251),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_217),
.A2(n_240),
.B(n_245),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_232),
.B(n_239),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_226),
.B(n_231),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_223),
.B(n_225),
.Y(n_219)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_228),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_233),
.B(n_238),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_233),
.B(n_238),
.Y(n_239)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_236),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_241),
.B(n_242),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_247),
.B(n_250),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_247),
.B(n_250),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_254),
.B(n_255),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_275),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_261),
.B(n_274),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_261),
.B(n_274),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_273),
.Y(n_261)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_264),
.B(n_272),
.C(n_273),
.Y(n_284)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

CKINVDCx14_ASAP7_75t_R g271 ( 
.A(n_268),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_275),
.A2(n_286),
.B(n_287),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_276),
.B(n_284),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_276),
.B(n_284),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_283),
.Y(n_276)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_291),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_289),
.B(n_291),
.Y(n_292)
);


endmodule