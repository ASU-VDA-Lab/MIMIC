module fake_jpeg_20190_n_289 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_289);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_289;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx4f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_18),
.B(n_25),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_31),
.Y(n_61)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_20),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_18),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx4_ASAP7_75t_SL g45 ( 
.A(n_31),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_45),
.Y(n_48)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_39),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_47),
.B(n_56),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_33),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_51),
.B(n_57),
.Y(n_76)
);

CKINVDCx9p33_ASAP7_75t_R g55 ( 
.A(n_39),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g80 ( 
.A(n_55),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_33),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_34),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_58),
.B(n_60),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_42),
.A2(n_40),
.B1(n_41),
.B2(n_31),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_59),
.A2(n_63),
.B1(n_67),
.B2(n_71),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_42),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_61),
.B(n_69),
.Y(n_94)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_40),
.A2(n_27),
.B1(n_23),
.B2(n_25),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_65),
.Y(n_108)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

AOI21xp33_ASAP7_75t_L g67 ( 
.A1(n_45),
.A2(n_34),
.B(n_23),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_45),
.B(n_28),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_40),
.A2(n_27),
.B1(n_24),
.B2(n_28),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_36),
.B(n_21),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_72),
.A2(n_29),
.B1(n_26),
.B2(n_20),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_45),
.B(n_35),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_73),
.Y(n_111)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_51),
.A2(n_41),
.B1(n_27),
.B2(n_44),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_77),
.A2(n_110),
.B1(n_30),
.B2(n_22),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_79),
.B(n_102),
.Y(n_114)
);

INVx13_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

BUFx4f_ASAP7_75t_SL g112 ( 
.A(n_81),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_72),
.A2(n_38),
.B(n_41),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_82),
.A2(n_103),
.B(n_106),
.Y(n_127)
);

OAI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_61),
.A2(n_36),
.B1(n_44),
.B2(n_37),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_87),
.A2(n_88),
.B1(n_101),
.B2(n_104),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_L g88 ( 
.A1(n_53),
.A2(n_44),
.B1(n_37),
.B2(n_46),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_66),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_89),
.B(n_90),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_50),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_91),
.Y(n_113)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_53),
.Y(n_92)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_92),
.Y(n_129)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_70),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_95),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_49),
.A2(n_29),
.B1(n_26),
.B2(n_35),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_96),
.Y(n_131)
);

BUFx2_ASAP7_75t_SL g97 ( 
.A(n_48),
.Y(n_97)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_97),
.Y(n_122)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_62),
.Y(n_98)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_98),
.Y(n_126)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_70),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_99),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_L g101 ( 
.A1(n_49),
.A2(n_44),
.B1(n_37),
.B2(n_38),
.Y(n_101)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_68),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_61),
.B(n_37),
.Y(n_103)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_64),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_107),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_75),
.B(n_30),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_64),
.Y(n_107)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_74),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_109),
.B(n_65),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_75),
.A2(n_19),
.B1(n_22),
.B2(n_21),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_111),
.A2(n_68),
.B1(n_19),
.B2(n_48),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_116),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_108),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_117),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_119),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_82),
.B(n_65),
.C(n_54),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_120),
.B(n_101),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_76),
.B(n_54),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_123),
.B(n_124),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_76),
.B(n_52),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_91),
.B(n_52),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_125),
.B(n_135),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_128),
.B(n_88),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_94),
.B(n_30),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_130),
.A2(n_139),
.B(n_80),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_79),
.A2(n_22),
.B1(n_21),
.B2(n_19),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_132),
.A2(n_136),
.B1(n_131),
.B2(n_80),
.Y(n_156)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_84),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_134),
.B(n_86),
.Y(n_143)
);

AO22x2_ASAP7_75t_L g135 ( 
.A1(n_93),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_81),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_103),
.B(n_1),
.Y(n_137)
);

AND2x2_ASAP7_75t_SL g162 ( 
.A(n_137),
.B(n_106),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_103),
.B(n_3),
.Y(n_139)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_126),
.Y(n_140)
);

INVx13_ASAP7_75t_L g177 ( 
.A(n_140),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_129),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_142),
.B(n_145),
.Y(n_172)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_143),
.Y(n_171)
);

O2A1O1Ixp33_ASAP7_75t_L g144 ( 
.A1(n_114),
.A2(n_85),
.B(n_92),
.C(n_78),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_144),
.A2(n_161),
.B(n_163),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_115),
.B(n_111),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_146),
.B(n_169),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_147),
.A2(n_156),
.B1(n_139),
.B2(n_122),
.Y(n_187)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_125),
.Y(n_148)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_148),
.Y(n_173)
);

OA21x2_ASAP7_75t_L g149 ( 
.A1(n_131),
.A2(n_85),
.B(n_109),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_149),
.B(n_157),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g150 ( 
.A(n_113),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_150),
.B(n_151),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_121),
.B(n_100),
.Y(n_151)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_126),
.Y(n_152)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_152),
.Y(n_196)
);

NAND3xp33_ASAP7_75t_L g153 ( 
.A(n_137),
.B(n_16),
.C(n_14),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_153),
.B(n_160),
.Y(n_185)
);

BUFx24_ASAP7_75t_SL g154 ( 
.A(n_130),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_154),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_112),
.B(n_83),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_117),
.Y(n_158)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_158),
.Y(n_186)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_134),
.Y(n_159)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_159),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_112),
.B(n_102),
.Y(n_160)
);

O2A1O1Ixp33_ASAP7_75t_L g161 ( 
.A1(n_132),
.A2(n_99),
.B(n_95),
.C(n_84),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_162),
.B(n_124),
.Y(n_182)
);

HAxp5_ASAP7_75t_SL g163 ( 
.A(n_127),
.B(n_106),
.CON(n_163),
.SN(n_163)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_112),
.B(n_98),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_165),
.B(n_166),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_118),
.B(n_83),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_169),
.B(n_127),
.C(n_120),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_170),
.B(n_183),
.C(n_141),
.Y(n_206)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_148),
.Y(n_174)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_174),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_146),
.B(n_123),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g214 ( 
.A(n_175),
.B(n_194),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_163),
.B(n_133),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_178),
.A2(n_187),
.B(n_189),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_162),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_180),
.B(n_142),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_182),
.B(n_188),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_164),
.B(n_130),
.C(n_139),
.Y(n_183)
);

OR2x2_ASAP7_75t_L g184 ( 
.A(n_168),
.B(n_136),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_184),
.A2(n_147),
.B(n_135),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_164),
.B(n_168),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_155),
.A2(n_149),
.B(n_147),
.Y(n_189)
);

AND2x6_ASAP7_75t_L g193 ( 
.A(n_149),
.B(n_135),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_193),
.B(n_133),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_162),
.B(n_156),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_191),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_197),
.B(n_202),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_198),
.A2(n_205),
.B1(n_217),
.B2(n_219),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_187),
.B(n_157),
.Y(n_200)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_200),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_176),
.B(n_170),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_201),
.B(n_204),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_172),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_203),
.B(n_211),
.Y(n_226)
);

A2O1A1O1Ixp25_ASAP7_75t_L g204 ( 
.A1(n_190),
.A2(n_144),
.B(n_155),
.C(n_135),
.D(n_161),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_206),
.B(n_194),
.C(n_175),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_179),
.A2(n_141),
.B(n_138),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_207),
.B(n_208),
.Y(n_235)
);

XOR2x2_ASAP7_75t_L g208 ( 
.A(n_176),
.B(n_150),
.Y(n_208)
);

OAI31xp33_ASAP7_75t_SL g209 ( 
.A1(n_193),
.A2(n_122),
.A3(n_152),
.B(n_159),
.Y(n_209)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_209),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_179),
.A2(n_158),
.B(n_140),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_178),
.A2(n_167),
.B(n_105),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_212),
.B(n_216),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_171),
.B(n_167),
.Y(n_215)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_215),
.Y(n_231)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_195),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_188),
.B(n_86),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_189),
.A2(n_108),
.B(n_5),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_218),
.B(n_4),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_174),
.B(n_4),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_200),
.A2(n_178),
.B1(n_173),
.B2(n_184),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_220),
.A2(n_204),
.B1(n_213),
.B2(n_210),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_200),
.A2(n_197),
.B1(n_199),
.B2(n_209),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_221),
.B(n_233),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_222),
.B(n_224),
.C(n_206),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_201),
.B(n_182),
.C(n_183),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_207),
.B(n_192),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_228),
.B(n_219),
.Y(n_239)
);

OA22x2_ASAP7_75t_L g233 ( 
.A1(n_211),
.A2(n_190),
.B1(n_180),
.B2(n_196),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_205),
.A2(n_185),
.B1(n_186),
.B2(n_196),
.Y(n_234)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_234),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_236),
.B(n_237),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_214),
.B(n_181),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_238),
.B(n_240),
.Y(n_261)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_239),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_224),
.B(n_214),
.C(n_208),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g241 ( 
.A(n_231),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_241),
.B(n_244),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_222),
.B(n_217),
.C(n_212),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_243),
.Y(n_254)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_225),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_227),
.B(n_213),
.C(n_210),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_245),
.Y(n_256)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_230),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_246),
.A2(n_248),
.B1(n_250),
.B2(n_232),
.Y(n_255)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_220),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_223),
.A2(n_218),
.B(n_216),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_251),
.A2(n_226),
.B(n_229),
.Y(n_253)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_253),
.Y(n_266)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_255),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_245),
.B(n_233),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_257),
.Y(n_265)
);

INVxp33_ASAP7_75t_L g258 ( 
.A(n_249),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_258),
.B(n_260),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_242),
.A2(n_227),
.B1(n_233),
.B2(n_235),
.Y(n_260)
);

A2O1A1Ixp33_ASAP7_75t_SL g262 ( 
.A1(n_249),
.A2(n_235),
.B(n_236),
.C(n_177),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_262),
.B(n_243),
.C(n_248),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_264),
.B(n_262),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_261),
.B(n_238),
.C(n_240),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_267),
.B(n_268),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_256),
.B(n_237),
.C(n_247),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_257),
.B(n_247),
.C(n_251),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_270),
.B(n_259),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_271),
.B(n_274),
.Y(n_280)
);

NOR2xp67_ASAP7_75t_R g273 ( 
.A(n_266),
.B(n_252),
.Y(n_273)
);

NAND3xp33_ASAP7_75t_L g277 ( 
.A(n_273),
.B(n_269),
.C(n_263),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_265),
.A2(n_259),
.B(n_241),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_265),
.A2(n_254),
.B(n_262),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_275),
.B(n_276),
.Y(n_278)
);

A2O1A1Ixp33_ASAP7_75t_L g282 ( 
.A1(n_277),
.A2(n_5),
.B(n_6),
.C(n_7),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_272),
.A2(n_177),
.B1(n_16),
.B2(n_7),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_279),
.B(n_8),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_278),
.A2(n_280),
.B(n_6),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_281),
.B(n_282),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_283),
.B(n_8),
.C(n_9),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_285),
.A2(n_9),
.B(n_10),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_286),
.A2(n_284),
.B1(n_10),
.B2(n_12),
.Y(n_287)
);

AO21x2_ASAP7_75t_L g288 ( 
.A1(n_287),
.A2(n_9),
.B(n_10),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_288),
.B(n_13),
.Y(n_289)
);


endmodule