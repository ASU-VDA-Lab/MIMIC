module fake_jpeg_27187_n_262 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_262);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_262;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_107;
wire n_39;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_9),
.B(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_24),
.B(n_11),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_28),
.B(n_29),
.Y(n_44)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

HB1xp67_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_22),
.B(n_0),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_26),
.C(n_22),
.Y(n_42)
);

BUFx10_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_34),
.Y(n_59)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_45),
.B(n_34),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_35),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_34),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_47),
.A2(n_33),
.B1(n_16),
.B2(n_32),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_48),
.A2(n_46),
.B1(n_37),
.B2(n_41),
.Y(n_71)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_57),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_47),
.A2(n_33),
.B1(n_16),
.B2(n_32),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_52),
.A2(n_46),
.B1(n_37),
.B2(n_41),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_43),
.A2(n_16),
.B1(n_25),
.B2(n_18),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_30),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_55),
.B(n_56),
.Y(n_78)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_38),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_62),
.Y(n_76)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_30),
.Y(n_62)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_45),
.B(n_29),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_64),
.A2(n_29),
.B1(n_13),
.B2(n_20),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_66),
.Y(n_99)
);

INVx2_ASAP7_75t_SL g68 ( 
.A(n_54),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_68),
.B(n_54),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_71),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_59),
.A2(n_45),
.B1(n_42),
.B2(n_46),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_73),
.A2(n_75),
.B1(n_77),
.B2(n_64),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_63),
.A2(n_42),
.B1(n_44),
.B2(n_38),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_51),
.A2(n_43),
.B1(n_41),
.B2(n_38),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_49),
.A2(n_43),
.B1(n_14),
.B2(n_25),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_79),
.A2(n_26),
.B(n_57),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_81),
.B(n_14),
.Y(n_97)
);

AND2x6_ASAP7_75t_L g83 ( 
.A(n_73),
.B(n_52),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_83),
.A2(n_81),
.B(n_57),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_78),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_85),
.Y(n_113)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_91),
.Y(n_103)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_88),
.A2(n_65),
.B(n_74),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_89),
.A2(n_67),
.B1(n_69),
.B2(n_71),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_80),
.A2(n_50),
.B1(n_61),
.B2(n_58),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_90),
.A2(n_82),
.B1(n_72),
.B2(n_49),
.Y(n_116)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_78),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_70),
.B(n_62),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_92),
.B(n_93),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_70),
.B(n_55),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_76),
.B(n_31),
.C(n_54),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_94),
.B(n_98),
.Y(n_104)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_96),
.Y(n_109)
);

INVx13_ASAP7_75t_L g96 ( 
.A(n_66),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_97),
.B(n_100),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_76),
.B(n_75),
.C(n_67),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_67),
.B(n_31),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_101),
.A2(n_107),
.B1(n_117),
.B2(n_40),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_89),
.A2(n_82),
.B1(n_72),
.B2(n_50),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_102),
.A2(n_118),
.B1(n_91),
.B2(n_68),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_86),
.A2(n_83),
.B1(n_98),
.B2(n_95),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_106),
.A2(n_116),
.B1(n_84),
.B2(n_94),
.Y(n_126)
);

OAI22xp33_ASAP7_75t_L g107 ( 
.A1(n_84),
.A2(n_61),
.B1(n_68),
.B2(n_56),
.Y(n_107)
);

NAND2xp33_ASAP7_75t_SL g130 ( 
.A(n_108),
.B(n_98),
.Y(n_130)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_112),
.B(n_40),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_88),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_114),
.B(n_119),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_85),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_115),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_84),
.A2(n_82),
.B1(n_65),
.B2(n_56),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_92),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_103),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_120),
.B(n_123),
.Y(n_142)
);

NAND3xp33_ASAP7_75t_L g121 ( 
.A(n_111),
.B(n_100),
.C(n_93),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_121),
.B(n_135),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_122),
.B(n_126),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_109),
.Y(n_123)
);

AOI22x1_ASAP7_75t_L g124 ( 
.A1(n_108),
.A2(n_83),
.B1(n_84),
.B2(n_90),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_124),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g125 ( 
.A(n_110),
.Y(n_125)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_125),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_119),
.B(n_99),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_127),
.B(n_129),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_113),
.A2(n_96),
.B1(n_99),
.B2(n_49),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_128),
.A2(n_130),
.B(n_102),
.Y(n_152)
);

INVx13_ASAP7_75t_L g129 ( 
.A(n_109),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_106),
.A2(n_97),
.B1(n_58),
.B2(n_96),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_132),
.B(n_133),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_117),
.A2(n_74),
.B1(n_38),
.B2(n_66),
.Y(n_133)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_111),
.Y(n_135)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_136),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_113),
.B(n_31),
.Y(n_137)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_137),
.Y(n_149)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_103),
.Y(n_138)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_138),
.Y(n_150)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_139),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_101),
.A2(n_14),
.B1(n_20),
.B2(n_13),
.Y(n_140)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_140),
.Y(n_157)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_118),
.Y(n_141)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_141),
.Y(n_159)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_124),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_144),
.B(n_40),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_SL g146 ( 
.A(n_126),
.B(n_104),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_146),
.B(n_162),
.Y(n_170)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_129),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_148),
.B(n_156),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_131),
.B(n_104),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_151),
.B(n_161),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_152),
.A2(n_123),
.B1(n_105),
.B2(n_137),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_120),
.B(n_104),
.C(n_115),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_153),
.B(n_156),
.C(n_15),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_138),
.B(n_132),
.C(n_141),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_124),
.B(n_110),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_133),
.B(n_112),
.Y(n_162)
);

A2O1A1O1Ixp25_ASAP7_75t_L g163 ( 
.A1(n_135),
.A2(n_105),
.B(n_116),
.C(n_17),
.D(n_28),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_163),
.B(n_17),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_165),
.A2(n_169),
.B1(n_183),
.B2(n_148),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_155),
.A2(n_122),
.B1(n_134),
.B2(n_136),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_167),
.A2(n_176),
.B1(n_149),
.B2(n_154),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_164),
.A2(n_13),
.B(n_20),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_168),
.B(n_171),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_144),
.A2(n_40),
.B1(n_26),
.B2(n_25),
.Y(n_169)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_142),
.Y(n_171)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_172),
.Y(n_193)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_173),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_174),
.B(n_161),
.Y(n_192)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_145),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_175),
.B(n_177),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_160),
.A2(n_40),
.B1(n_26),
.B2(n_39),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_157),
.B(n_23),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_150),
.B(n_21),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_178),
.B(n_181),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_179),
.B(n_184),
.C(n_27),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_146),
.B(n_39),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_180),
.B(n_151),
.Y(n_186)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_162),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_163),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_182),
.A2(n_11),
.B(n_12),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_158),
.A2(n_18),
.B1(n_21),
.B2(n_11),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_153),
.B(n_23),
.Y(n_184)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_185),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_186),
.B(n_192),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_179),
.B(n_147),
.C(n_143),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_187),
.B(n_188),
.C(n_190),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_180),
.B(n_170),
.C(n_166),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_170),
.B(n_152),
.C(n_159),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_194),
.A2(n_19),
.B1(n_23),
.B2(n_17),
.Y(n_216)
);

BUFx2_ASAP7_75t_L g197 ( 
.A(n_167),
.Y(n_197)
);

BUFx12_ASAP7_75t_L g202 ( 
.A(n_197),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_166),
.B(n_154),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_198),
.B(n_199),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_174),
.B(n_17),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_200),
.B(n_40),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_201),
.A2(n_168),
.B1(n_176),
.B2(n_18),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_203),
.A2(n_199),
.B1(n_192),
.B2(n_197),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_187),
.B(n_169),
.C(n_15),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_206),
.B(n_207),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_196),
.B(n_15),
.C(n_27),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_193),
.A2(n_21),
.B1(n_8),
.B2(n_9),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_209),
.B(n_195),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_189),
.A2(n_9),
.B(n_12),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_210),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_211),
.B(n_213),
.Y(n_227)
);

A2O1A1Ixp33_ASAP7_75t_SL g212 ( 
.A1(n_190),
.A2(n_27),
.B(n_19),
.C(n_3),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_212),
.A2(n_19),
.B1(n_2),
.B2(n_3),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_188),
.B(n_27),
.C(n_17),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_191),
.B(n_10),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_215),
.B(n_8),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_216),
.A2(n_19),
.B1(n_2),
.B2(n_3),
.Y(n_224)
);

OAI22xp33_ASAP7_75t_L g229 ( 
.A1(n_217),
.A2(n_223),
.B1(n_202),
.B2(n_212),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_214),
.B(n_186),
.C(n_198),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_218),
.B(n_219),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_204),
.B(n_23),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_220),
.B(n_225),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_221),
.B(n_224),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_204),
.B(n_19),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_205),
.A2(n_8),
.B1(n_19),
.B2(n_4),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_226),
.B(n_1),
.Y(n_237)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_229),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_228),
.A2(n_212),
.B(n_202),
.Y(n_230)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_230),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_218),
.A2(n_214),
.B(n_227),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_231),
.A2(n_236),
.B(n_1),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_217),
.A2(n_202),
.B(n_208),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_233),
.A2(n_225),
.B(n_223),
.Y(n_239)
);

XNOR2x1_ASAP7_75t_L g234 ( 
.A(n_220),
.B(n_208),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_234),
.B(n_4),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_222),
.A2(n_19),
.B(n_2),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_237),
.B(n_5),
.Y(n_246)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_239),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_235),
.A2(n_19),
.B(n_4),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_241),
.B(n_243),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_242),
.B(n_232),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_237),
.B(n_1),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_245),
.B(n_5),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_246),
.B(n_7),
.Y(n_251)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_247),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_248),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_244),
.A2(n_238),
.B1(n_6),
.B2(n_7),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_250),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_254),
.B(n_252),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_256),
.B(n_257),
.C(n_243),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_255),
.B(n_240),
.C(n_249),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_258),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_259),
.A2(n_253),
.B(n_251),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_260),
.A2(n_5),
.B(n_6),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_261),
.B(n_5),
.Y(n_262)
);


endmodule