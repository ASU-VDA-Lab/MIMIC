module fake_jpeg_8351_n_168 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_168);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_168;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_1),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_9),
.Y(n_12)
);

INVx8_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_7),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx24_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_14),
.B(n_5),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_25),
.B(n_28),
.Y(n_37)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_14),
.B(n_5),
.Y(n_28)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_29),
.B(n_31),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_31),
.B(n_21),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_34),
.B(n_25),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_19),
.Y(n_36)
);

OR2x4_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_20),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

HB1xp67_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_44),
.Y(n_58)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_28),
.Y(n_46)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_38),
.A2(n_16),
.B1(n_13),
.B2(n_40),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_47),
.A2(n_17),
.B1(n_12),
.B2(n_21),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_49),
.A2(n_36),
.B(n_19),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_15),
.Y(n_50)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_38),
.A2(n_13),
.B1(n_16),
.B2(n_40),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_52),
.A2(n_29),
.B1(n_13),
.B2(n_17),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_53),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_36),
.B(n_15),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_54),
.B(n_55),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_32),
.B(n_15),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_21),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_19),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_L g59 ( 
.A1(n_49),
.A2(n_40),
.B1(n_38),
.B2(n_16),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_59),
.A2(n_61),
.B1(n_62),
.B2(n_67),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_52),
.A2(n_13),
.B1(n_36),
.B2(n_27),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_64),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_SL g64 ( 
.A(n_54),
.B(n_20),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_39),
.Y(n_66)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_33),
.C(n_39),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_47),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_71),
.B(n_43),
.Y(n_80)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_73),
.B(n_75),
.Y(n_96)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_71),
.Y(n_75)
);

CKINVDCx12_ASAP7_75t_R g76 ( 
.A(n_69),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_76),
.B(n_77),
.Y(n_88)
);

CKINVDCx12_ASAP7_75t_R g77 ( 
.A(n_68),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_63),
.A2(n_56),
.B(n_50),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_78),
.A2(n_84),
.B(n_65),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_58),
.B(n_46),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_79),
.B(n_80),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_60),
.A2(n_35),
.B1(n_17),
.B2(n_12),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_81),
.A2(n_12),
.B(n_57),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_82),
.B(n_23),
.Y(n_98)
);

AND2x4_ASAP7_75t_L g84 ( 
.A(n_64),
.B(n_26),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_70),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_68),
.Y(n_92)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_81),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_86),
.B(n_89),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_57),
.C(n_60),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_93),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_79),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_92),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_74),
.B(n_58),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_73),
.A2(n_62),
.B1(n_65),
.B2(n_61),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_94),
.A2(n_72),
.B1(n_75),
.B2(n_83),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_95),
.A2(n_78),
.B(n_84),
.Y(n_109)
);

NOR4xp25_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_5),
.C(n_8),
.D(n_7),
.Y(n_97)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_97),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_98),
.B(n_72),
.Y(n_103)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_99),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_88),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_101),
.B(n_106),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_100),
.C(n_104),
.Y(n_123)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_96),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_107),
.A2(n_112),
.B1(n_114),
.B2(n_18),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_SL g124 ( 
.A(n_109),
.B(n_33),
.Y(n_124)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_90),
.Y(n_110)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_110),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_91),
.B(n_87),
.Y(n_111)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_111),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_89),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_86),
.A2(n_84),
.B1(n_35),
.B2(n_39),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_113),
.A2(n_51),
.B1(n_33),
.B2(n_42),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_95),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_106),
.A2(n_99),
.B1(n_97),
.B2(n_98),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_115),
.A2(n_117),
.B1(n_126),
.B2(n_127),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_102),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_116),
.B(n_120),
.Y(n_129)
);

BUFx2_ASAP7_75t_L g118 ( 
.A(n_110),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_118),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_112),
.A2(n_93),
.B(n_22),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_123),
.B(n_125),
.C(n_104),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_124),
.B(n_108),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_108),
.B(n_48),
.C(n_51),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_100),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_124),
.A2(n_114),
.B(n_105),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_128),
.B(n_132),
.Y(n_144)
);

FAx1_ASAP7_75t_SL g131 ( 
.A(n_123),
.B(n_109),
.CI(n_105),
.CON(n_131),
.SN(n_131)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_131),
.B(n_137),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_133),
.B(n_135),
.C(n_136),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_125),
.B(n_113),
.C(n_48),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_122),
.B(n_45),
.C(n_42),
.Y(n_136)
);

FAx1_ASAP7_75t_SL g137 ( 
.A(n_117),
.B(n_26),
.CI(n_42),
.CON(n_137),
.SN(n_137)
);

NOR2xp67_ASAP7_75t_SL g138 ( 
.A(n_131),
.B(n_118),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_138),
.A2(n_128),
.B(n_131),
.Y(n_146)
);

OR2x2_ASAP7_75t_L g140 ( 
.A(n_129),
.B(n_121),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_140),
.B(n_145),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_133),
.B(n_119),
.C(n_116),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_141),
.B(n_142),
.C(n_11),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_129),
.B(n_136),
.C(n_132),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_134),
.A2(n_30),
.B1(n_27),
.B2(n_23),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_146),
.A2(n_149),
.B(n_151),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_143),
.A2(n_130),
.B(n_135),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_147),
.A2(n_6),
.B(n_10),
.Y(n_155)
);

XNOR2x2_ASAP7_75t_SL g148 ( 
.A(n_143),
.B(n_137),
.Y(n_148)
);

AOI21x1_ASAP7_75t_SL g157 ( 
.A1(n_148),
.A2(n_4),
.B(n_8),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_139),
.A2(n_134),
.B(n_137),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_144),
.A2(n_45),
.B(n_22),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_7),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_153),
.B(n_156),
.C(n_4),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_150),
.B(n_41),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_154),
.A2(n_41),
.B1(n_30),
.B2(n_2),
.Y(n_161)
);

AO21x1_ASAP7_75t_L g162 ( 
.A1(n_155),
.A2(n_0),
.B(n_1),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_150),
.B(n_6),
.Y(n_156)
);

OA21x2_ASAP7_75t_SL g160 ( 
.A1(n_157),
.A2(n_4),
.B(n_1),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_159),
.A2(n_0),
.B1(n_3),
.B2(n_41),
.Y(n_165)
);

OAI321xp33_ASAP7_75t_L g163 ( 
.A1(n_160),
.A2(n_161),
.A3(n_162),
.B1(n_158),
.B2(n_1),
.C(n_2),
.Y(n_163)
);

FAx1_ASAP7_75t_SL g167 ( 
.A(n_163),
.B(n_165),
.CI(n_3),
.CON(n_167),
.SN(n_167)
);

AOI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_162),
.A2(n_41),
.B(n_2),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_164),
.A2(n_0),
.B(n_3),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_166),
.B(n_167),
.Y(n_168)
);


endmodule