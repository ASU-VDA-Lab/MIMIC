module fake_jpeg_28720_n_252 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_252);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_252;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g18 ( 
.A(n_1),
.B(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_14),
.B(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_2),
.B(n_10),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx10_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_32),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_24),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_23),
.B(n_18),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_23),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_45),
.A2(n_24),
.B1(n_34),
.B2(n_25),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_48),
.A2(n_65),
.B1(n_66),
.B2(n_29),
.Y(n_93)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_52),
.B(n_72),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_17),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_54),
.B(n_55),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_18),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_58),
.B(n_64),
.Y(n_92)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_63),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_43),
.B(n_33),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_37),
.A2(n_24),
.B1(n_34),
.B2(n_25),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_37),
.A2(n_23),
.B1(n_33),
.B2(n_34),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_67),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_42),
.B(n_25),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_68),
.B(n_69),
.Y(n_97)
);

CKINVDCx14_ASAP7_75t_R g69 ( 
.A(n_42),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_70),
.Y(n_101)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_43),
.B(n_16),
.Y(n_72)
);

AO22x1_ASAP7_75t_SL g73 ( 
.A1(n_59),
.A2(n_46),
.B1(n_38),
.B2(n_39),
.Y(n_73)
);

OA22x2_ASAP7_75t_SL g111 ( 
.A1(n_73),
.A2(n_39),
.B1(n_57),
.B2(n_35),
.Y(n_111)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_74),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_51),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_75),
.B(n_99),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_L g76 ( 
.A1(n_59),
.A2(n_46),
.B1(n_28),
.B2(n_26),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_76),
.A2(n_93),
.B1(n_95),
.B2(n_104),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_47),
.A2(n_28),
.B1(n_26),
.B2(n_30),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_77),
.A2(n_35),
.B1(n_32),
.B2(n_2),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_78),
.Y(n_125)
);

BUFx6f_ASAP7_75t_SL g79 ( 
.A(n_53),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_79),
.Y(n_113)
);

INVx2_ASAP7_75t_SL g80 ( 
.A(n_47),
.Y(n_80)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_80),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_54),
.A2(n_28),
.B1(n_30),
.B2(n_17),
.Y(n_82)
);

AOI32xp33_ASAP7_75t_L g109 ( 
.A1(n_82),
.A2(n_22),
.A3(n_19),
.B1(n_29),
.B2(n_27),
.Y(n_109)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_83),
.Y(n_119)
);

BUFx12_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_84),
.B(n_91),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_56),
.B(n_27),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_85),
.B(n_22),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_86),
.Y(n_120)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_71),
.Y(n_89)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_89),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_62),
.Y(n_91)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_94),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_50),
.A2(n_29),
.B1(n_19),
.B2(n_21),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_56),
.B(n_30),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_70),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_100),
.B(n_105),
.Y(n_130)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_60),
.Y(n_102)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_102),
.Y(n_126)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_63),
.Y(n_103)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_103),
.Y(n_128)
);

OAI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_50),
.A2(n_46),
.B1(n_35),
.B2(n_32),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_62),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_109),
.B(n_127),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_110),
.B(n_131),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_111),
.A2(n_73),
.B1(n_96),
.B2(n_90),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_88),
.A2(n_57),
.B1(n_22),
.B2(n_27),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_114),
.A2(n_124),
.B1(n_0),
.B2(n_1),
.Y(n_145)
);

OAI21xp33_ASAP7_75t_L g116 ( 
.A1(n_92),
.A2(n_21),
.B(n_19),
.Y(n_116)
);

OAI21xp33_ASAP7_75t_L g155 ( 
.A1(n_116),
.A2(n_4),
.B(n_6),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_99),
.A2(n_76),
.B1(n_87),
.B2(n_97),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_117),
.A2(n_121),
.B1(n_82),
.B2(n_80),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_87),
.A2(n_21),
.B1(n_17),
.B2(n_35),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_106),
.B(n_16),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_85),
.B(n_35),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_129),
.B(n_32),
.Y(n_142)
);

O2A1O1Ixp33_ASAP7_75t_L g131 ( 
.A1(n_73),
.A2(n_35),
.B(n_32),
.C(n_3),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_88),
.B(n_0),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_132),
.B(n_7),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_133),
.A2(n_134),
.B1(n_135),
.B2(n_136),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_108),
.A2(n_90),
.B1(n_96),
.B2(n_101),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_108),
.A2(n_101),
.B1(n_98),
.B2(n_81),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_110),
.A2(n_107),
.B(n_129),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_137),
.A2(n_143),
.B(n_11),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_117),
.A2(n_98),
.B1(n_81),
.B2(n_105),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_138),
.A2(n_139),
.B1(n_154),
.B2(n_115),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_111),
.A2(n_78),
.B1(n_74),
.B2(n_79),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_112),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_140),
.B(n_141),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_130),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_142),
.B(n_147),
.Y(n_163)
);

NAND2x1_ASAP7_75t_SL g143 ( 
.A(n_111),
.B(n_84),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_125),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_144),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_145),
.A2(n_121),
.B1(n_127),
.B2(n_118),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_118),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_146),
.B(n_158),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_114),
.B(n_132),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_119),
.Y(n_148)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_148),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_119),
.B(n_1),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_150),
.B(n_152),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_123),
.B(n_3),
.Y(n_152)
);

A2O1A1Ixp33_ASAP7_75t_L g153 ( 
.A1(n_111),
.A2(n_84),
.B(n_5),
.C(n_6),
.Y(n_153)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_153),
.Y(n_175)
);

OAI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_131),
.A2(n_115),
.B1(n_126),
.B2(n_123),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g180 ( 
.A(n_155),
.Y(n_180)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_126),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_156),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_128),
.B(n_7),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_157),
.B(n_150),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_137),
.B(n_122),
.C(n_128),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_159),
.B(n_168),
.C(n_172),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_160),
.B(n_171),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_162),
.A2(n_139),
.B1(n_136),
.B2(n_135),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_165),
.A2(n_134),
.B1(n_143),
.B2(n_145),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_141),
.B(n_122),
.Y(n_167)
);

CKINVDCx14_ASAP7_75t_R g199 ( 
.A(n_167),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_142),
.B(n_120),
.C(n_125),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_133),
.B(n_147),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_138),
.B(n_120),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_149),
.B(n_8),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_173),
.B(n_176),
.C(n_160),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_154),
.A2(n_113),
.B1(n_9),
.B2(n_11),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_174),
.A2(n_153),
.B(n_144),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_151),
.B(n_8),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_152),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_178),
.B(n_157),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_179),
.A2(n_153),
.B(n_149),
.Y(n_183)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_170),
.Y(n_182)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_182),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_183),
.A2(n_200),
.B(n_173),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_184),
.B(n_186),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_185),
.A2(n_193),
.B1(n_194),
.B2(n_197),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_164),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_170),
.Y(n_187)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_187),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_166),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_188),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_189),
.A2(n_192),
.B1(n_181),
.B2(n_169),
.Y(n_211)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_172),
.Y(n_191)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_191),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_175),
.A2(n_179),
.B1(n_165),
.B2(n_161),
.Y(n_192)
);

NOR3xp33_ASAP7_75t_SL g193 ( 
.A(n_180),
.B(n_151),
.C(n_158),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_175),
.A2(n_143),
.B(n_156),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_196),
.A2(n_174),
.B(n_159),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_181),
.B(n_148),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_198),
.B(n_176),
.Y(n_206)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_168),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_201),
.A2(n_205),
.B(n_209),
.Y(n_221)
);

AOI211xp5_ASAP7_75t_L g202 ( 
.A1(n_183),
.A2(n_171),
.B(n_177),
.C(n_163),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_202),
.A2(n_211),
.B1(n_189),
.B2(n_192),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_196),
.A2(n_163),
.B(n_161),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_206),
.B(n_212),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_190),
.B(n_15),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_190),
.B(n_11),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_213),
.B(n_195),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_214),
.A2(n_193),
.B(n_184),
.Y(n_215)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_215),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_212),
.B(n_200),
.C(n_191),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_216),
.B(n_218),
.Y(n_230)
);

NOR3xp33_ASAP7_75t_L g217 ( 
.A(n_207),
.B(n_186),
.C(n_199),
.Y(n_217)
);

BUFx24_ASAP7_75t_SL g228 ( 
.A(n_217),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_208),
.B(n_195),
.C(n_198),
.Y(n_218)
);

AOI31xp67_ASAP7_75t_L g219 ( 
.A1(n_203),
.A2(n_188),
.A3(n_194),
.B(n_197),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_219),
.A2(n_223),
.B1(n_224),
.B2(n_225),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_204),
.B(n_187),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_220),
.B(n_222),
.Y(n_234)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_210),
.Y(n_223)
);

INVxp33_ASAP7_75t_L g225 ( 
.A(n_211),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_221),
.B(n_209),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_227),
.B(n_12),
.Y(n_240)
);

XOR2x1_ASAP7_75t_SL g231 ( 
.A(n_221),
.B(n_202),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_231),
.A2(n_225),
.B1(n_182),
.B2(n_218),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_224),
.A2(n_185),
.B1(n_201),
.B2(n_205),
.Y(n_232)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_232),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_235),
.B(n_228),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_230),
.B(n_216),
.C(n_226),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_236),
.B(n_240),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_233),
.A2(n_206),
.B1(n_213),
.B2(n_226),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_237),
.A2(n_227),
.B1(n_234),
.B2(n_229),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_231),
.A2(n_222),
.B(n_13),
.Y(n_239)
);

CKINVDCx14_ASAP7_75t_R g241 ( 
.A(n_239),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_242),
.B(n_243),
.Y(n_247)
);

OR2x2_ASAP7_75t_L g245 ( 
.A(n_244),
.B(n_238),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_245),
.A2(n_246),
.B(n_12),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_244),
.A2(n_239),
.B(n_240),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_247),
.B(n_241),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_248),
.A2(n_249),
.B(n_14),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_250),
.B(n_15),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_251),
.B(n_15),
.Y(n_252)
);


endmodule