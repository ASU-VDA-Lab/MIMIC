module fake_jpeg_15481_n_145 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_145);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_145;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_12),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_8),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx4f_ASAP7_75t_SL g28 ( 
.A(n_4),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_37),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_16),
.B(n_0),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_32),
.B(n_25),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_18),
.B(n_0),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_33),
.B(n_26),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_34),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_37),
.A2(n_26),
.B1(n_16),
.B2(n_25),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_39),
.B(n_42),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_33),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_50),
.Y(n_57)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_20),
.Y(n_48)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_30),
.B(n_28),
.C(n_27),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_52),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_30),
.B(n_27),
.Y(n_52)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

O2A1O1Ixp33_ASAP7_75t_L g56 ( 
.A1(n_50),
.A2(n_28),
.B(n_34),
.C(n_14),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_49),
.Y(n_77)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_60),
.B(n_61),
.Y(n_70)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_62),
.B(n_63),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

CKINVDCx14_ASAP7_75t_R g65 ( 
.A(n_39),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_65),
.B(n_23),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_28),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_66),
.B(n_45),
.Y(n_69)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_68),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_69),
.B(n_81),
.Y(n_85)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_72),
.B(n_53),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_58),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_73),
.B(n_77),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_57),
.A2(n_64),
.B1(n_67),
.B2(n_66),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_74),
.A2(n_63),
.B1(n_59),
.B2(n_53),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_64),
.B(n_52),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_75),
.A2(n_49),
.B1(n_46),
.B2(n_15),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_44),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_76),
.B(n_83),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_57),
.A2(n_38),
.B(n_23),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_78),
.B(n_60),
.Y(n_86)
);

AND2x2_ASAP7_75t_SL g83 ( 
.A(n_56),
.B(n_15),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_86),
.B(n_88),
.Y(n_100)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_89),
.Y(n_104)
);

NOR2x1_ASAP7_75t_L g90 ( 
.A(n_83),
.B(n_77),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_90),
.B(n_93),
.Y(n_98)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_84),
.Y(n_91)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_91),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_78),
.Y(n_106)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_84),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_69),
.B(n_55),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_94),
.B(n_95),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_70),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_41),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_96),
.B(n_75),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_102),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_91),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_93),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_103),
.Y(n_112)
);

OA22x2_ASAP7_75t_L g116 ( 
.A1(n_106),
.A2(n_79),
.B1(n_21),
.B2(n_20),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_97),
.A2(n_76),
.B1(n_74),
.B2(n_77),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_107),
.A2(n_109),
.B1(n_87),
.B2(n_80),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_90),
.A2(n_83),
.B(n_73),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_SL g119 ( 
.A(n_108),
.B(n_24),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_92),
.A2(n_80),
.B1(n_72),
.B2(n_79),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_98),
.A2(n_87),
.B1(n_96),
.B2(n_85),
.Y(n_110)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_110),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_111),
.B(n_113),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_104),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_100),
.B(n_86),
.C(n_88),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_114),
.B(n_115),
.C(n_106),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_100),
.B(n_82),
.C(n_71),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_SL g120 ( 
.A(n_116),
.B(n_119),
.Y(n_120)
);

AOI322xp5_ASAP7_75t_L g118 ( 
.A1(n_108),
.A2(n_35),
.A3(n_13),
.B1(n_21),
.B2(n_14),
.C1(n_24),
.C2(n_7),
.Y(n_118)
);

BUFx24_ASAP7_75t_SL g126 ( 
.A(n_118),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_117),
.A2(n_104),
.B1(n_99),
.B2(n_105),
.Y(n_121)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_121),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_122),
.B(n_116),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_116),
.B(n_105),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_123),
.A2(n_112),
.B(n_24),
.Y(n_131)
);

MAJx2_ASAP7_75t_L g125 ( 
.A(n_119),
.B(n_101),
.C(n_10),
.Y(n_125)
);

NOR4xp25_ASAP7_75t_L g133 ( 
.A(n_125),
.B(n_9),
.C(n_11),
.D(n_4),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_124),
.B(n_112),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_128),
.A2(n_127),
.B1(n_126),
.B2(n_120),
.Y(n_134)
);

BUFx24_ASAP7_75t_SL g135 ( 
.A(n_130),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_131),
.A2(n_132),
.B(n_133),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_124),
.A2(n_10),
.B(n_12),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_134),
.A2(n_136),
.B1(n_1),
.B2(n_6),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_129),
.A2(n_13),
.B1(n_3),
.B2(n_5),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_135),
.B(n_130),
.C(n_22),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_138),
.B(n_139),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_137),
.B(n_24),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_140),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_141),
.Y(n_143)
);

NOR3xp33_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_142),
.C(n_22),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_1),
.Y(n_145)
);


endmodule