module fake_jpeg_30184_n_503 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_503);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_503;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

HB1xp67_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_11),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

INVx11_ASAP7_75t_SL g46 ( 
.A(n_14),
.Y(n_46)
);

CKINVDCx5p33_ASAP7_75t_R g47 ( 
.A(n_7),
.Y(n_47)
);

BUFx16f_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

INVx11_ASAP7_75t_L g144 ( 
.A(n_51),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_52),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_53),
.Y(n_138)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_54),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_55),
.Y(n_118)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_56),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_20),
.B(n_7),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_57),
.B(n_89),
.Y(n_123)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_58),
.Y(n_119)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_59),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_7),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_60),
.B(n_88),
.Y(n_113)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_61),
.Y(n_124)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_48),
.Y(n_62)
);

INVx13_ASAP7_75t_L g107 ( 
.A(n_62),
.Y(n_107)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_63),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_64),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_29),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_65),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_66),
.Y(n_161)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_18),
.Y(n_67)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_67),
.Y(n_120)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_68),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_69),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g150 ( 
.A(n_70),
.Y(n_150)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_71),
.Y(n_129)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_18),
.Y(n_72)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_72),
.Y(n_125)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_28),
.Y(n_73)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_73),
.Y(n_134)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_48),
.Y(n_74)
);

INVx5_ASAP7_75t_SL g117 ( 
.A(n_74),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_29),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g156 ( 
.A(n_75),
.Y(n_156)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_76),
.Y(n_147)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

INVx2_ASAP7_75t_SL g143 ( 
.A(n_77),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_38),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g159 ( 
.A(n_78),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_38),
.Y(n_79)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_32),
.Y(n_80)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_80),
.Y(n_133)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_81),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_38),
.Y(n_82)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_82),
.Y(n_137)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_83),
.Y(n_142)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g112 ( 
.A(n_84),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_42),
.Y(n_85)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_85),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_42),
.Y(n_86)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_86),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_42),
.Y(n_87)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_87),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_20),
.B(n_8),
.Y(n_89)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_28),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g127 ( 
.A(n_90),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_19),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g146 ( 
.A(n_91),
.Y(n_146)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_19),
.Y(n_92)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_35),
.Y(n_93)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_93),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_47),
.B(n_6),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_94),
.B(n_27),
.Y(n_102)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_40),
.Y(n_95)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_95),
.Y(n_128)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_19),
.Y(n_96)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_96),
.Y(n_139)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_23),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_97),
.B(n_98),
.Y(n_126)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_23),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_27),
.B(n_6),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_99),
.B(n_100),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_23),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_33),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_101),
.B(n_34),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_102),
.B(n_121),
.Y(n_193)
);

NAND2x1_ASAP7_75t_L g109 ( 
.A(n_62),
.B(n_36),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_109),
.B(n_140),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_53),
.A2(n_36),
.B1(n_26),
.B2(n_39),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_111),
.A2(n_116),
.B1(n_155),
.B2(n_17),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_52),
.A2(n_49),
.B1(n_44),
.B2(n_43),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_83),
.B(n_35),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_55),
.A2(n_64),
.B1(n_65),
.B2(n_66),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_132),
.A2(n_135),
.B1(n_149),
.B2(n_157),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_75),
.A2(n_33),
.B1(n_34),
.B2(n_44),
.Y(n_135)
);

AO22x1_ASAP7_75t_L g136 ( 
.A1(n_70),
.A2(n_36),
.B1(n_30),
.B2(n_17),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_136),
.A2(n_0),
.B(n_1),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_78),
.A2(n_86),
.B1(n_79),
.B2(n_82),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_92),
.A2(n_34),
.B1(n_33),
.B2(n_41),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_152),
.A2(n_85),
.B1(n_17),
.B2(n_50),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_70),
.B(n_43),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_153),
.B(n_107),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_69),
.A2(n_39),
.B1(n_26),
.B2(n_41),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_91),
.A2(n_49),
.B1(n_50),
.B2(n_45),
.Y(n_157)
);

HAxp5_ASAP7_75t_SL g160 ( 
.A(n_90),
.B(n_30),
.CON(n_160),
.SN(n_160)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_160),
.B(n_17),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_161),
.A2(n_100),
.B1(n_96),
.B2(n_87),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_162),
.A2(n_199),
.B1(n_133),
.B2(n_110),
.Y(n_220)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_122),
.Y(n_163)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_163),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_164),
.A2(n_167),
.B1(n_168),
.B2(n_179),
.Y(n_244)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_137),
.Y(n_165)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_165),
.Y(n_223)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_119),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_166),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_130),
.A2(n_63),
.B1(n_51),
.B2(n_26),
.Y(n_167)
);

OAI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_159),
.A2(n_68),
.B1(n_81),
.B2(n_21),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_156),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_169),
.B(n_170),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_156),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_123),
.B(n_16),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_171),
.B(n_174),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_136),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_172),
.B(n_191),
.Y(n_222)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_126),
.Y(n_173)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_173),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_113),
.B(n_16),
.Y(n_174)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_142),
.Y(n_175)
);

INVx8_ASAP7_75t_L g231 ( 
.A(n_175),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_103),
.B(n_45),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_176),
.B(n_190),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_108),
.A2(n_74),
.B1(n_88),
.B2(n_21),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_178),
.A2(n_181),
.B1(n_183),
.B2(n_145),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_152),
.A2(n_41),
.B1(n_39),
.B2(n_26),
.Y(n_179)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_117),
.Y(n_180)
);

INVx13_ASAP7_75t_L g224 ( 
.A(n_180),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_114),
.A2(n_10),
.B1(n_14),
.B2(n_13),
.Y(n_181)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_150),
.Y(n_182)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_182),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_148),
.A2(n_10),
.B1(n_14),
.B2(n_13),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_146),
.Y(n_184)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_184),
.Y(n_251)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_151),
.Y(n_185)
);

INVx6_ASAP7_75t_L g247 ( 
.A(n_185),
.Y(n_247)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_117),
.Y(n_186)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_186),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_104),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_187),
.Y(n_233)
);

INVx5_ASAP7_75t_L g188 ( 
.A(n_144),
.Y(n_188)
);

INVx11_ASAP7_75t_L g249 ( 
.A(n_188),
.Y(n_249)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_158),
.Y(n_189)
);

CKINVDCx14_ASAP7_75t_R g238 ( 
.A(n_189),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_124),
.B(n_129),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_159),
.Y(n_191)
);

INVx8_ASAP7_75t_L g192 ( 
.A(n_105),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_192),
.Y(n_241)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_138),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_194),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_196),
.B(n_202),
.Y(n_229)
);

OA22x2_ASAP7_75t_L g214 ( 
.A1(n_197),
.A2(n_211),
.B1(n_161),
.B2(n_133),
.Y(n_214)
);

OR2x2_ASAP7_75t_L g227 ( 
.A(n_198),
.B(n_208),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_155),
.A2(n_111),
.B1(n_134),
.B2(n_106),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_146),
.B(n_17),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_200),
.B(n_209),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_120),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_201),
.Y(n_239)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_105),
.Y(n_202)
);

BUFx2_ASAP7_75t_L g203 ( 
.A(n_110),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_203),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_115),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_204),
.A2(n_210),
.B1(n_39),
.B2(n_2),
.Y(n_250)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_112),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_205),
.B(n_206),
.Y(n_248)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_106),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_128),
.B(n_109),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_207),
.B(n_41),
.Y(n_246)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_127),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_127),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_160),
.A2(n_41),
.B1(n_39),
.B2(n_26),
.Y(n_210)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_154),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_212),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_214),
.B(n_246),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_172),
.A2(n_115),
.B1(n_118),
.B2(n_141),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_215),
.A2(n_236),
.B1(n_178),
.B2(n_180),
.Y(n_263)
);

NOR2x1_ASAP7_75t_L g217 ( 
.A(n_198),
.B(n_107),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_217),
.B(n_211),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_220),
.A2(n_228),
.B1(n_235),
.B2(n_237),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_195),
.B(n_112),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_225),
.B(n_240),
.C(n_198),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_177),
.A2(n_141),
.B1(n_131),
.B2(n_118),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_L g236 ( 
.A1(n_173),
.A2(n_131),
.B1(n_125),
.B2(n_139),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_177),
.A2(n_143),
.B1(n_147),
.B2(n_144),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_195),
.B(n_143),
.C(n_154),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_250),
.A2(n_182),
.B1(n_204),
.B2(n_194),
.Y(n_278)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_218),
.Y(n_252)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_252),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_253),
.B(n_258),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_254),
.B(n_244),
.Y(n_305)
);

BUFx2_ASAP7_75t_L g255 ( 
.A(n_241),
.Y(n_255)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_255),
.Y(n_310)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_218),
.Y(n_256)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_256),
.Y(n_288)
);

A2O1A1Ixp33_ASAP7_75t_SL g257 ( 
.A1(n_214),
.A2(n_199),
.B(n_167),
.C(n_164),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_257),
.A2(n_266),
.B(n_282),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_225),
.B(n_195),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_L g259 ( 
.A1(n_237),
.A2(n_163),
.B1(n_203),
.B2(n_184),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_L g298 ( 
.A1(n_259),
.A2(n_263),
.B1(n_238),
.B2(n_245),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_216),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_260),
.B(n_262),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_243),
.B(n_176),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_261),
.B(n_264),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_216),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_243),
.B(n_171),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_247),
.Y(n_265)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_265),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_222),
.A2(n_186),
.B(n_181),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_247),
.Y(n_267)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_267),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_248),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_268),
.B(n_277),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_226),
.B(n_190),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_269),
.B(n_274),
.Y(n_301)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_241),
.Y(n_270)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_270),
.Y(n_309)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_251),
.Y(n_271)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_271),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_226),
.B(n_200),
.Y(n_274)
);

OA22x2_ASAP7_75t_SL g275 ( 
.A1(n_222),
.A2(n_179),
.B1(n_185),
.B2(n_165),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_275),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_235),
.A2(n_189),
.B1(n_209),
.B2(n_208),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_276),
.A2(n_278),
.B1(n_280),
.B2(n_238),
.Y(n_312)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_247),
.Y(n_277)
);

INVx2_ASAP7_75t_SL g279 ( 
.A(n_245),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_279),
.B(n_285),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_228),
.A2(n_220),
.B1(n_221),
.B2(n_214),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_230),
.B(n_174),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_281),
.B(n_284),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_227),
.A2(n_214),
.B(n_240),
.Y(n_282)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_232),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_283),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_230),
.B(n_193),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_251),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_284),
.B(n_221),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_292),
.B(n_252),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_260),
.B(n_227),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_295),
.B(n_297),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_261),
.B(n_227),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_L g341 ( 
.A1(n_298),
.A2(n_234),
.B1(n_255),
.B2(n_242),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_281),
.B(n_274),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_300),
.B(n_302),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_269),
.B(n_229),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_258),
.B(n_214),
.C(n_246),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_303),
.B(n_183),
.C(n_212),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_264),
.B(n_229),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_304),
.B(n_279),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_305),
.B(n_314),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_254),
.A2(n_217),
.B(n_244),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_307),
.A2(n_313),
.B(n_270),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_283),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_308),
.B(n_279),
.Y(n_333)
);

MAJx2_ASAP7_75t_L g311 ( 
.A(n_253),
.B(n_217),
.C(n_248),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_311),
.B(n_224),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_312),
.A2(n_277),
.B1(n_267),
.B2(n_265),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_282),
.A2(n_239),
.B(n_233),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_272),
.A2(n_242),
.B1(n_219),
.B2(n_234),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_314),
.A2(n_280),
.B1(n_273),
.B2(n_276),
.Y(n_321)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_310),
.Y(n_318)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_318),
.Y(n_354)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_320),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_321),
.A2(n_322),
.B1(n_323),
.B2(n_324),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_317),
.A2(n_273),
.B1(n_257),
.B2(n_272),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_306),
.A2(n_257),
.B1(n_272),
.B2(n_275),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_306),
.A2(n_257),
.B1(n_275),
.B2(n_266),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_286),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_325),
.B(n_327),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_L g371 ( 
.A1(n_326),
.A2(n_346),
.B(n_337),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_292),
.B(n_256),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_286),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_328),
.A2(n_332),
.B1(n_334),
.B2(n_336),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_307),
.A2(n_257),
.B1(n_263),
.B2(n_285),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_329),
.A2(n_339),
.B1(n_297),
.B2(n_312),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_293),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_331),
.Y(n_360)
);

HB1xp67_ASAP7_75t_L g332 ( 
.A(n_310),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g355 ( 
.A1(n_333),
.A2(n_337),
.B(n_293),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_287),
.B(n_213),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_296),
.B(n_271),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_335),
.B(n_311),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_287),
.B(n_213),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_313),
.B(n_241),
.Y(n_337)
);

AND2x2_ASAP7_75t_SL g338 ( 
.A(n_305),
.B(n_231),
.Y(n_338)
);

FAx1_ASAP7_75t_SL g358 ( 
.A(n_338),
.B(n_343),
.CI(n_289),
.CON(n_358),
.SN(n_358)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_303),
.A2(n_302),
.B1(n_305),
.B2(n_304),
.Y(n_339)
);

NAND3xp33_ASAP7_75t_L g340 ( 
.A(n_295),
.B(n_219),
.C(n_232),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_SL g370 ( 
.A1(n_340),
.A2(n_294),
.B(n_202),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_341),
.A2(n_347),
.B1(n_294),
.B2(n_299),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_315),
.B(n_224),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_342),
.A2(n_345),
.B1(n_231),
.B2(n_223),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_344),
.B(n_301),
.C(n_300),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_315),
.B(n_224),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_348),
.B(n_296),
.Y(n_350)
);

OA21x2_ASAP7_75t_L g349 ( 
.A1(n_346),
.A2(n_305),
.B(n_289),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g391 ( 
.A1(n_349),
.A2(n_355),
.B(n_325),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_350),
.B(n_353),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_352),
.B(n_374),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_335),
.B(n_311),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_357),
.B(n_367),
.Y(n_392)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_358),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_359),
.A2(n_318),
.B1(n_249),
.B2(n_3),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_362),
.B(n_365),
.C(n_366),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_321),
.A2(n_316),
.B1(n_288),
.B2(n_308),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_363),
.A2(n_364),
.B1(n_372),
.B2(n_373),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_322),
.A2(n_316),
.B1(n_288),
.B2(n_290),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_348),
.B(n_301),
.C(n_291),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_339),
.B(n_291),
.C(n_309),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_330),
.B(n_309),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_SL g368 ( 
.A(n_319),
.B(n_290),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_368),
.B(n_369),
.C(n_378),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_330),
.B(n_299),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_370),
.B(n_376),
.Y(n_384)
);

AOI21xp5_ASAP7_75t_L g385 ( 
.A1(n_371),
.A2(n_331),
.B(n_327),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_329),
.A2(n_231),
.B1(n_188),
.B2(n_223),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_326),
.A2(n_324),
.B1(n_323),
.B2(n_338),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_326),
.A2(n_206),
.B1(n_249),
.B2(n_192),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_375),
.B(n_333),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_SL g376 ( 
.A1(n_337),
.A2(n_175),
.B(n_249),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_344),
.B(n_343),
.C(n_319),
.Y(n_378)
);

BUFx24_ASAP7_75t_SL g379 ( 
.A(n_377),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_379),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_385),
.B(n_352),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_386),
.B(n_391),
.Y(n_421)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_361),
.Y(n_387)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_387),
.Y(n_412)
);

AND2x2_ASAP7_75t_SL g388 ( 
.A(n_358),
.B(n_338),
.Y(n_388)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_388),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_350),
.B(n_338),
.C(n_320),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_389),
.B(n_390),
.C(n_9),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_353),
.B(n_347),
.C(n_328),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_393),
.A2(n_372),
.B1(n_375),
.B2(n_351),
.Y(n_411)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_358),
.Y(n_394)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_394),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_360),
.B(n_356),
.Y(n_395)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_395),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_367),
.B(n_1),
.Y(n_396)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_396),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_362),
.B(n_6),
.Y(n_397)
);

CKINVDCx16_ASAP7_75t_R g409 ( 
.A(n_397),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_369),
.B(n_363),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_398),
.B(n_399),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_364),
.B(n_2),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_355),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_400),
.B(n_401),
.Y(n_422)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_354),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_373),
.Y(n_402)
);

CKINVDCx16_ASAP7_75t_R g413 ( 
.A(n_402),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_SL g404 ( 
.A(n_378),
.B(n_9),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g423 ( 
.A1(n_404),
.A2(n_385),
.B1(n_387),
.B2(n_383),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_SL g408 ( 
.A(n_388),
.B(n_349),
.C(n_371),
.Y(n_408)
);

NOR2xp67_ASAP7_75t_L g437 ( 
.A(n_408),
.B(n_406),
.Y(n_437)
);

XOR2x1_ASAP7_75t_L g439 ( 
.A(n_410),
.B(n_405),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_411),
.A2(n_414),
.B1(n_405),
.B2(n_410),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_402),
.A2(n_351),
.B1(n_366),
.B2(n_349),
.Y(n_414)
);

FAx1_ASAP7_75t_SL g416 ( 
.A(n_388),
.B(n_368),
.CI(n_357),
.CON(n_416),
.SN(n_416)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_416),
.B(n_423),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_SL g418 ( 
.A(n_389),
.B(n_365),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_418),
.B(n_419),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_403),
.B(n_359),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_381),
.A2(n_9),
.B1(n_11),
.B2(n_10),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_425),
.A2(n_420),
.B1(n_415),
.B2(n_417),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_426),
.B(n_390),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_380),
.B(n_2),
.C(n_3),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_427),
.B(n_396),
.C(n_380),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_428),
.B(n_435),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_412),
.B(n_395),
.Y(n_430)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_430),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_424),
.B(n_404),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_432),
.B(n_440),
.Y(n_447)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_422),
.Y(n_433)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_433),
.Y(n_458)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_422),
.Y(n_434)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_434),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_426),
.B(n_382),
.C(n_403),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_436),
.B(n_418),
.C(n_392),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_437),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_409),
.B(n_400),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_438),
.B(n_441),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_439),
.B(n_444),
.Y(n_446)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_415),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_419),
.B(n_382),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_442),
.A2(n_413),
.B1(n_391),
.B2(n_383),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_443),
.B(n_445),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_414),
.B(n_392),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_417),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_448),
.B(n_441),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_450),
.A2(n_454),
.B1(n_459),
.B2(n_416),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_442),
.A2(n_394),
.B1(n_408),
.B2(n_406),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_436),
.B(n_421),
.C(n_398),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_455),
.B(n_456),
.C(n_446),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_444),
.B(n_421),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_456),
.B(n_431),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_429),
.A2(n_439),
.B1(n_386),
.B2(n_407),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_428),
.A2(n_411),
.B1(n_421),
.B2(n_384),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_461),
.A2(n_420),
.B1(n_431),
.B2(n_393),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_462),
.B(n_467),
.Y(n_485)
);

OR2x2_ASAP7_75t_L g463 ( 
.A(n_449),
.B(n_416),
.Y(n_463)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_463),
.Y(n_484)
);

OAI22xp33_ASAP7_75t_L g464 ( 
.A1(n_449),
.A2(n_399),
.B1(n_407),
.B2(n_401),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_464),
.B(n_465),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_SL g465 ( 
.A(n_452),
.B(n_435),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_466),
.B(n_468),
.Y(n_476)
);

CKINVDCx16_ASAP7_75t_R g469 ( 
.A(n_447),
.Y(n_469)
);

CKINVDCx16_ASAP7_75t_R g477 ( 
.A(n_469),
.Y(n_477)
);

AOI21xp5_ASAP7_75t_L g482 ( 
.A1(n_470),
.A2(n_471),
.B(n_472),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_447),
.B(n_427),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_451),
.B(n_5),
.Y(n_472)
);

OAI21xp5_ASAP7_75t_SL g473 ( 
.A1(n_458),
.A2(n_10),
.B(n_11),
.Y(n_473)
);

AO22x1_ASAP7_75t_L g480 ( 
.A1(n_473),
.A2(n_454),
.B1(n_450),
.B2(n_459),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_457),
.B(n_12),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_474),
.A2(n_475),
.B1(n_460),
.B2(n_461),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_453),
.B(n_4),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_466),
.B(n_446),
.C(n_455),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_478),
.B(n_479),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g490 ( 
.A1(n_480),
.A2(n_464),
.B1(n_3),
.B2(n_4),
.Y(n_490)
);

OA21x2_ASAP7_75t_L g483 ( 
.A1(n_462),
.A2(n_448),
.B(n_3),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_SL g487 ( 
.A(n_483),
.B(n_473),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_476),
.B(n_468),
.C(n_463),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_486),
.B(n_489),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_487),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_476),
.B(n_467),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_490),
.Y(n_492)
);

INVxp67_ASAP7_75t_L g491 ( 
.A(n_478),
.Y(n_491)
);

O2A1O1Ixp33_ASAP7_75t_SL g495 ( 
.A1(n_491),
.A2(n_480),
.B(n_483),
.C(n_481),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_495),
.B(n_483),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_493),
.B(n_491),
.C(n_488),
.Y(n_496)
);

AOI21x1_ASAP7_75t_L g498 ( 
.A1(n_496),
.A2(n_497),
.B(n_489),
.Y(n_498)
);

INVxp67_ASAP7_75t_L g499 ( 
.A(n_498),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_499),
.B(n_492),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_500),
.B(n_477),
.C(n_482),
.Y(n_501)
);

OAI21xp33_ASAP7_75t_SL g502 ( 
.A1(n_501),
.A2(n_494),
.B(n_484),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_502),
.A2(n_2),
.B1(n_485),
.B2(n_499),
.Y(n_503)
);


endmodule