module real_jpeg_28208_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_215;
wire n_166;
wire n_176;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_139;
wire n_33;
wire n_188;
wire n_65;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_285;
wire n_172;
wire n_45;
wire n_211;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_277;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_187;
wire n_97;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_279;
wire n_59;
wire n_169;
wire n_128;
wire n_167;
wire n_244;
wire n_179;
wire n_216;
wire n_202;
wire n_133;
wire n_213;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_283;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_273;
wire n_96;
wire n_253;
wire n_269;
wire n_89;
wire n_16;

INVx11_ASAP7_75t_L g87 ( 
.A(n_0),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_0),
.B(n_215),
.Y(n_220)
);

INVx5_ASAP7_75t_L g231 ( 
.A(n_0),
.Y(n_231)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_2),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

OAI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_2),
.A2(n_23),
.B1(n_24),
.B2(n_31),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_2),
.A2(n_31),
.B1(n_45),
.B2(n_49),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_2),
.A2(n_31),
.B1(n_51),
.B2(n_53),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_4),
.A2(n_29),
.B1(n_30),
.B2(n_117),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_4),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_4),
.A2(n_23),
.B1(n_24),
.B2(n_117),
.Y(n_143)
);

OAI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_4),
.A2(n_45),
.B1(n_49),
.B2(n_117),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_4),
.A2(n_51),
.B1(n_53),
.B2(n_117),
.Y(n_215)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_6),
.A2(n_23),
.B1(n_24),
.B2(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_6),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_6),
.A2(n_45),
.B1(n_49),
.B2(n_68),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_6),
.A2(n_51),
.B1(n_53),
.B2(n_68),
.Y(n_133)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g36 ( 
.A1(n_8),
.A2(n_29),
.B(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_8),
.B(n_29),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_8),
.A2(n_45),
.B1(n_49),
.B2(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_8),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_8),
.A2(n_51),
.B1(n_53),
.B2(n_57),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_8),
.A2(n_23),
.B1(n_24),
.B2(n_57),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_8),
.B(n_20),
.Y(n_170)
);

AOI21xp33_ASAP7_75t_SL g181 ( 
.A1(n_8),
.A2(n_10),
.B(n_45),
.Y(n_181)
);

AOI21xp33_ASAP7_75t_L g206 ( 
.A1(n_8),
.A2(n_48),
.B(n_51),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_8),
.B(n_64),
.Y(n_210)
);

BUFx24_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_10),
.Y(n_61)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_10),
.Y(n_63)
);

INVx11_ASAP7_75t_SL g52 ( 
.A(n_11),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_125),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_123),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_93),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_15),
.B(n_93),
.Y(n_124)
);

BUFx24_ASAP7_75t_SL g286 ( 
.A(n_15),
.Y(n_286)
);

FAx1_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_72),
.CI(n_80),
.CON(n_15),
.SN(n_15)
);

AOI22xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_38),
.B2(n_39),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_18),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_32),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_19),
.B(n_113),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_27),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_20),
.B(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

A2O1A1Ixp33_ASAP7_75t_L g34 ( 
.A1(n_21),
.A2(n_22),
.B(n_29),
.C(n_35),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_21),
.A2(n_34),
.B(n_36),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_21),
.B(n_116),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_24),
.B2(n_26),
.Y(n_21)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_22),
.B(n_29),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_23),
.B(n_26),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

O2A1O1Ixp33_ASAP7_75t_L g60 ( 
.A1(n_24),
.A2(n_61),
.B(n_62),
.C(n_64),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_24),
.B(n_63),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_24),
.A2(n_156),
.B1(n_157),
.B2(n_158),
.Y(n_155)
);

A2O1A1Ixp33_ASAP7_75t_L g179 ( 
.A1(n_24),
.A2(n_57),
.B(n_180),
.C(n_181),
.Y(n_179)
);

BUFx2_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

CKINVDCx14_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_28),
.B(n_34),
.Y(n_260)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_33),
.B(n_139),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_34),
.B(n_36),
.Y(n_33)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_34),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_35),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_36),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_37),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_40),
.A2(n_41),
.B1(n_58),
.B2(n_59),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_40),
.B(n_138),
.C(n_140),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_40),
.A2(n_41),
.B1(n_140),
.B2(n_141),
.Y(n_164)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_54),
.B(n_55),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_42),
.A2(n_90),
.B(n_91),
.Y(n_89)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_43),
.B(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_43),
.B(n_56),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_43),
.B(n_188),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_50),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_44)
);

INVx4_ASAP7_75t_SL g49 ( 
.A(n_45),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_45),
.A2(n_49),
.B1(n_63),
.B2(n_65),
.Y(n_64)
);

A2O1A1Ixp33_ASAP7_75t_L g205 ( 
.A1(n_45),
.A2(n_47),
.B(n_57),
.C(n_206),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_47),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_47),
.A2(n_48),
.B1(n_51),
.B2(n_53),
.Y(n_50)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_50),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_50),
.B(n_56),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_50),
.B(n_79),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_50),
.B(n_188),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_51),
.Y(n_53)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_53),
.B(n_86),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_53),
.B(n_230),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_54),
.A2(n_78),
.B(n_90),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_54),
.B(n_57),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_57),
.B(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_66),
.B(n_69),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_60),
.B(n_71),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_60),
.B(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_60),
.B(n_143),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_60),
.Y(n_263)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_63),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_64),
.B(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_64),
.B(n_143),
.Y(n_142)
);

INVx6_ASAP7_75t_L g180 ( 
.A(n_65),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_67),
.A2(n_74),
.B(n_75),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_69),
.B(n_106),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_70),
.B(n_153),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_72),
.A2(n_73),
.B(n_76),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_76),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_74),
.B(n_151),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_74),
.A2(n_151),
.B(n_263),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_75),
.B(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_78),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_77),
.B(n_197),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_78),
.B(n_187),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_84),
.B(n_92),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_81),
.A2(n_82),
.B1(n_120),
.B2(n_121),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_89),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_83),
.A2(n_84),
.B1(n_92),
.B2(n_122),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_83),
.A2(n_84),
.B1(n_179),
.B2(n_182),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_83),
.A2(n_84),
.B1(n_89),
.B2(n_277),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_84),
.B(n_179),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_85),
.A2(n_86),
.B(n_88),
.Y(n_84)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_85),
.B(n_88),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_85),
.B(n_215),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_86),
.B(n_88),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_86),
.B(n_102),
.Y(n_134)
);

INVx11_ASAP7_75t_L g160 ( 
.A(n_86),
.Y(n_160)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

CKINVDCx14_ASAP7_75t_R g277 ( 
.A(n_89),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_91),
.B(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_91),
.B(n_197),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_92),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_118),
.C(n_119),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_94),
.A2(n_95),
.B1(n_283),
.B2(n_284),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_105),
.C(n_109),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_96),
.B(n_273),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_104),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_97),
.B(n_104),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_99),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_98),
.B(n_214),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_99),
.A2(n_133),
.B(n_160),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_100),
.B(n_219),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_101),
.B(n_103),
.Y(n_100)
);

INVxp33_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_103),
.A2(n_133),
.B(n_134),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_105),
.A2(n_109),
.B1(n_110),
.B2(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_105),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_107),
.B(n_142),
.Y(n_184)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_108),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_113),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_114),
.B(n_115),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_118),
.B(n_119),
.Y(n_284)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_280),
.B(n_285),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_127),
.A2(n_267),
.B(n_279),
.Y(n_126)
);

O2A1O1Ixp33_ASAP7_75t_SL g127 ( 
.A1(n_128),
.A2(n_173),
.B(n_249),
.C(n_266),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_161),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_129),
.B(n_161),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_144),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_137),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_131),
.B(n_137),
.C(n_144),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_135),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_132),
.B(n_135),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_134),
.B(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_134),
.B(n_214),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_136),
.B(n_187),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_138),
.B(n_164),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_139),
.B(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_145),
.B(n_154),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_147),
.B1(n_148),
.B2(n_149),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_146),
.B(n_149),
.C(n_154),
.Y(n_264)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_152),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_159),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_155),
.B(n_159),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_165),
.C(n_167),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_162),
.A2(n_163),
.B1(n_244),
.B2(n_245),
.Y(n_243)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_165),
.A2(n_166),
.B1(n_167),
.B2(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_167),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.C(n_171),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_168),
.B(n_192),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_169),
.A2(n_170),
.B1(n_171),
.B2(n_193),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_170),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_171),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_172),
.B(n_220),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_174),
.B(n_248),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_241),
.B(n_247),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_199),
.B(n_240),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_189),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_177),
.B(n_189),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_183),
.C(n_185),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_178),
.B(n_238),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_179),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_183),
.A2(n_184),
.B1(n_185),
.B2(n_186),
.Y(n_238)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_186),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_190),
.A2(n_191),
.B1(n_194),
.B2(n_195),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_190),
.B(n_196),
.C(n_198),
.Y(n_242)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_198),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_235),
.B(n_239),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_216),
.B(n_234),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_207),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_202),
.B(n_207),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_203),
.B(n_205),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_203),
.A2(n_204),
.B1(n_205),
.B2(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_205),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_213),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_210),
.B1(n_211),
.B2(n_212),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_209),
.B(n_212),
.C(n_213),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_210),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_212),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_223),
.B(n_233),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_221),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_218),
.B(n_221),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_220),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_224),
.A2(n_227),
.B(n_232),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_225),
.B(n_226),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_236),
.B(n_237),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_242),
.B(n_243),
.Y(n_247)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_250),
.B(n_251),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_252),
.A2(n_253),
.B1(n_264),
.B2(n_265),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_254),
.B(n_255),
.C(n_265),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_256),
.B(n_259),
.C(n_261),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_258),
.A2(n_259),
.B1(n_261),
.B2(n_262),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_264),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_268),
.B(n_269),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_278),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_271),
.A2(n_272),
.B1(n_275),
.B2(n_276),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_271),
.B(n_276),
.C(n_278),
.Y(n_281)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_276),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_281),
.B(n_282),
.Y(n_285)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);


endmodule