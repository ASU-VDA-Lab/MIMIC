module real_aes_7652_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_754;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g532 ( .A1(n_0), .A2(n_178), .B(n_533), .C(n_536), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_1), .B(n_483), .Y(n_537) );
INVx1_ASAP7_75t_L g104 ( .A(n_2), .Y(n_104) );
INVx1_ASAP7_75t_L g190 ( .A(n_3), .Y(n_190) );
NAND2xp5_ASAP7_75t_SL g523 ( .A(n_4), .B(n_150), .Y(n_523) );
AOI21xp5_ASAP7_75t_L g476 ( .A1(n_5), .A2(n_456), .B(n_477), .Y(n_476) );
AO21x2_ASAP7_75t_L g485 ( .A1(n_6), .A2(n_170), .B(n_486), .Y(n_485) );
AOI22xp33_ASAP7_75t_L g198 ( .A1(n_7), .A2(n_35), .B1(n_144), .B2(n_199), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_8), .B(n_170), .Y(n_179) );
AND2x6_ASAP7_75t_L g162 ( .A(n_9), .B(n_163), .Y(n_162) );
A2O1A1Ixp33_ASAP7_75t_L g545 ( .A1(n_10), .A2(n_162), .B(n_461), .C(n_546), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_11), .B(n_110), .Y(n_109) );
NOR2xp33_ASAP7_75t_L g123 ( .A(n_11), .B(n_36), .Y(n_123) );
INVx1_ASAP7_75t_L g140 ( .A(n_12), .Y(n_140) );
INVx1_ASAP7_75t_L g183 ( .A(n_13), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_14), .B(n_148), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g491 ( .A(n_15), .B(n_150), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_16), .B(n_136), .Y(n_254) );
AO32x2_ASAP7_75t_L g196 ( .A1(n_17), .A2(n_135), .A3(n_161), .B1(n_170), .B2(n_197), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_18), .B(n_144), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_19), .B(n_136), .Y(n_192) );
AOI22xp33_ASAP7_75t_L g200 ( .A1(n_20), .A2(n_50), .B1(n_144), .B2(n_199), .Y(n_200) );
AOI22xp33_ASAP7_75t_SL g238 ( .A1(n_21), .A2(n_78), .B1(n_144), .B2(n_148), .Y(n_238) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_22), .B(n_144), .Y(n_211) );
A2O1A1Ixp33_ASAP7_75t_L g509 ( .A1(n_23), .A2(n_161), .B(n_461), .C(n_510), .Y(n_509) );
OAI22xp5_ASAP7_75t_SL g125 ( .A1(n_24), .A2(n_55), .B1(n_126), .B2(n_127), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_24), .Y(n_126) );
A2O1A1Ixp33_ASAP7_75t_L g488 ( .A1(n_25), .A2(n_161), .B(n_461), .C(n_489), .Y(n_488) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_26), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_27), .B(n_165), .Y(n_164) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_28), .A2(n_456), .B(n_530), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_29), .B(n_165), .Y(n_213) );
INVx2_ASAP7_75t_L g146 ( .A(n_30), .Y(n_146) );
A2O1A1Ixp33_ASAP7_75t_L g498 ( .A1(n_31), .A2(n_459), .B(n_469), .C(n_499), .Y(n_498) );
NAND2xp5_ASAP7_75t_SL g143 ( .A(n_32), .B(n_144), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_33), .B(n_165), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_34), .B(n_220), .Y(n_490) );
INVx1_ASAP7_75t_L g110 ( .A(n_36), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_37), .B(n_508), .Y(n_507) );
CKINVDCx20_ASAP7_75t_R g550 ( .A(n_38), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_39), .B(n_150), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_40), .B(n_456), .Y(n_487) );
A2O1A1Ixp33_ASAP7_75t_L g458 ( .A1(n_41), .A2(n_459), .B(n_463), .C(n_469), .Y(n_458) );
NAND2xp5_ASAP7_75t_SL g173 ( .A(n_42), .B(n_144), .Y(n_173) );
INVx1_ASAP7_75t_L g534 ( .A(n_43), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g236 ( .A1(n_44), .A2(n_89), .B1(n_199), .B2(n_237), .Y(n_236) );
INVx1_ASAP7_75t_L g464 ( .A(n_45), .Y(n_464) );
NAND2xp5_ASAP7_75t_SL g176 ( .A(n_46), .B(n_144), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_47), .B(n_144), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_48), .B(n_456), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_49), .B(n_156), .Y(n_177) );
AOI22xp33_ASAP7_75t_SL g252 ( .A1(n_51), .A2(n_56), .B1(n_144), .B2(n_148), .Y(n_252) );
CKINVDCx20_ASAP7_75t_R g515 ( .A(n_52), .Y(n_515) );
NAND2xp5_ASAP7_75t_SL g158 ( .A(n_53), .B(n_144), .Y(n_158) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_54), .B(n_144), .Y(n_217) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_55), .Y(n_127) );
OAI22xp5_ASAP7_75t_SL g444 ( .A1(n_55), .A2(n_127), .B1(n_128), .B2(n_445), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_57), .B(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g163 ( .A(n_58), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_59), .B(n_456), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_60), .B(n_483), .Y(n_482) );
A2O1A1Ixp33_ASAP7_75t_L g479 ( .A1(n_61), .A2(n_156), .B(n_186), .C(n_480), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_62), .B(n_144), .Y(n_191) );
INVx1_ASAP7_75t_L g139 ( .A(n_63), .Y(n_139) );
AOI22xp33_ASAP7_75t_L g100 ( .A1(n_64), .A2(n_101), .B1(n_111), .B2(n_754), .Y(n_100) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_65), .Y(n_116) );
NAND2xp5_ASAP7_75t_SL g501 ( .A(n_66), .B(n_150), .Y(n_501) );
AO32x2_ASAP7_75t_L g234 ( .A1(n_67), .A2(n_161), .A3(n_170), .B1(n_235), .B2(n_239), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_68), .B(n_151), .Y(n_547) );
INVx1_ASAP7_75t_L g154 ( .A(n_69), .Y(n_154) );
INVx1_ASAP7_75t_L g208 ( .A(n_70), .Y(n_208) );
CKINVDCx16_ASAP7_75t_R g531 ( .A(n_71), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_72), .B(n_466), .Y(n_511) );
A2O1A1Ixp33_ASAP7_75t_L g520 ( .A1(n_73), .A2(n_461), .B(n_469), .C(n_521), .Y(n_520) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_74), .B(n_148), .Y(n_209) );
CKINVDCx16_ASAP7_75t_R g478 ( .A(n_75), .Y(n_478) );
INVx1_ASAP7_75t_L g108 ( .A(n_76), .Y(n_108) );
NAND2xp5_ASAP7_75t_SL g512 ( .A(n_77), .B(n_465), .Y(n_512) );
AOI222xp33_ASAP7_75t_L g439 ( .A1(n_79), .A2(n_83), .B1(n_440), .B2(n_747), .C1(n_752), .C2(n_753), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_80), .B(n_199), .Y(n_223) );
CKINVDCx20_ASAP7_75t_R g503 ( .A(n_81), .Y(n_503) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_82), .B(n_148), .Y(n_212) );
INVx1_ASAP7_75t_L g752 ( .A(n_83), .Y(n_752) );
INVx2_ASAP7_75t_L g137 ( .A(n_84), .Y(n_137) );
CKINVDCx20_ASAP7_75t_R g527 ( .A(n_85), .Y(n_527) );
NAND2xp5_ASAP7_75t_SL g548 ( .A(n_86), .B(n_160), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_87), .B(n_148), .Y(n_174) );
INVx2_ASAP7_75t_L g105 ( .A(n_88), .Y(n_105) );
OR2x2_ASAP7_75t_L g120 ( .A(n_88), .B(n_121), .Y(n_120) );
OR2x2_ASAP7_75t_L g443 ( .A(n_88), .B(n_122), .Y(n_443) );
AOI22xp33_ASAP7_75t_L g251 ( .A1(n_90), .A2(n_99), .B1(n_148), .B2(n_149), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_91), .B(n_456), .Y(n_497) );
INVx1_ASAP7_75t_L g500 ( .A(n_92), .Y(n_500) );
INVxp67_ASAP7_75t_L g481 ( .A(n_93), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_94), .B(n_148), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_95), .B(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g522 ( .A(n_96), .Y(n_522) );
INVx1_ASAP7_75t_L g543 ( .A(n_97), .Y(n_543) );
AND2x2_ASAP7_75t_L g471 ( .A(n_98), .B(n_165), .Y(n_471) );
INVx1_ASAP7_75t_SL g101 ( .A(n_102), .Y(n_101) );
INVx1_ASAP7_75t_L g755 ( .A(n_102), .Y(n_755) );
OR2x2_ASAP7_75t_L g102 ( .A(n_103), .B(n_109), .Y(n_102) );
NAND3xp33_ASAP7_75t_SL g103 ( .A(n_104), .B(n_105), .C(n_106), .Y(n_103) );
AND2x2_ASAP7_75t_L g122 ( .A(n_104), .B(n_123), .Y(n_122) );
OR2x2_ASAP7_75t_L g448 ( .A(n_105), .B(n_122), .Y(n_448) );
NOR2x2_ASAP7_75t_L g753 ( .A(n_105), .B(n_121), .Y(n_753) );
OA211x2_ASAP7_75t_L g111 ( .A1(n_106), .A2(n_112), .B(n_117), .C(n_436), .Y(n_111) );
INVx1_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_SL g112 ( .A(n_113), .Y(n_112) );
INVx1_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
INVx1_ASAP7_75t_SL g438 ( .A(n_114), .Y(n_438) );
BUFx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
OAI21xp5_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_124), .B(n_432), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
HB1xp67_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx2_ASAP7_75t_L g435 ( .A(n_120), .Y(n_435) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
XNOR2xp5_ASAP7_75t_L g124 ( .A(n_125), .B(n_128), .Y(n_124) );
INVx1_ASAP7_75t_SL g445 ( .A(n_128), .Y(n_445) );
OR3x1_ASAP7_75t_L g128 ( .A(n_129), .B(n_360), .C(n_409), .Y(n_128) );
NAND5xp2_ASAP7_75t_L g129 ( .A(n_130), .B(n_275), .C(n_303), .D(n_333), .E(n_347), .Y(n_129) );
AOI221xp5_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_193), .B1(n_225), .B2(n_230), .C(n_241), .Y(n_130) );
NOR2xp33_ASAP7_75t_L g131 ( .A(n_132), .B(n_166), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_132), .B(n_227), .Y(n_226) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx2_ASAP7_75t_L g255 ( .A(n_133), .Y(n_255) );
AND2x2_ASAP7_75t_L g263 ( .A(n_133), .B(n_169), .Y(n_263) );
AND2x2_ASAP7_75t_L g286 ( .A(n_133), .B(n_168), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_133), .B(n_180), .Y(n_301) );
OR2x2_ASAP7_75t_L g310 ( .A(n_133), .B(n_248), .Y(n_310) );
HB1xp67_ASAP7_75t_L g313 ( .A(n_133), .Y(n_313) );
AND2x2_ASAP7_75t_L g421 ( .A(n_133), .B(n_248), .Y(n_421) );
OA21x2_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_141), .B(n_164), .Y(n_133) );
OA21x2_ASAP7_75t_L g180 ( .A1(n_134), .A2(n_181), .B(n_192), .Y(n_180) );
INVx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
NOR2xp33_ASAP7_75t_L g549 ( .A(n_135), .B(n_550), .Y(n_549) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_136), .Y(n_170) );
AND2x2_ASAP7_75t_L g136 ( .A(n_137), .B(n_138), .Y(n_136) );
AND2x2_ASAP7_75t_SL g165 ( .A(n_137), .B(n_138), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_139), .B(n_140), .Y(n_138) );
OAI21xp5_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_153), .B(n_161), .Y(n_141) );
AOI21xp5_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_147), .B(n_150), .Y(n_142) );
INVx3_ASAP7_75t_L g207 ( .A(n_144), .Y(n_207) );
HB1xp67_ASAP7_75t_L g524 ( .A(n_144), .Y(n_524) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx1_ASAP7_75t_L g199 ( .A(n_145), .Y(n_199) );
BUFx3_ASAP7_75t_L g237 ( .A(n_145), .Y(n_237) );
AND2x6_ASAP7_75t_L g461 ( .A(n_145), .B(n_462), .Y(n_461) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx1_ASAP7_75t_L g149 ( .A(n_146), .Y(n_149) );
INVx1_ASAP7_75t_L g157 ( .A(n_146), .Y(n_157) );
INVx2_ASAP7_75t_L g184 ( .A(n_148), .Y(n_184) );
INVx3_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
AOI21xp5_ASAP7_75t_L g172 ( .A1(n_150), .A2(n_173), .B(n_174), .Y(n_172) );
INVx2_ASAP7_75t_L g178 ( .A(n_150), .Y(n_178) );
O2A1O1Ixp5_ASAP7_75t_SL g206 ( .A1(n_150), .A2(n_207), .B(n_208), .C(n_209), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g480 ( .A(n_150), .B(n_481), .Y(n_480) );
INVx5_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
OAI22xp5_ASAP7_75t_SL g235 ( .A1(n_151), .A2(n_160), .B1(n_236), .B2(n_238), .Y(n_235) );
INVx3_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_152), .Y(n_160) );
BUFx6f_ASAP7_75t_L g188 ( .A(n_152), .Y(n_188) );
INVx1_ASAP7_75t_L g220 ( .A(n_152), .Y(n_220) );
AND2x2_ASAP7_75t_L g457 ( .A(n_152), .B(n_157), .Y(n_457) );
INVx1_ASAP7_75t_L g462 ( .A(n_152), .Y(n_462) );
O2A1O1Ixp5_ASAP7_75t_L g153 ( .A1(n_154), .A2(n_155), .B(n_158), .C(n_159), .Y(n_153) );
O2A1O1Ixp33_ASAP7_75t_L g189 ( .A1(n_155), .A2(n_178), .B(n_190), .C(n_191), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_155), .A2(n_511), .B(n_512), .Y(n_510) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_159), .A2(n_222), .B(n_223), .Y(n_221) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
OAI22xp5_ASAP7_75t_L g197 ( .A1(n_160), .A2(n_178), .B1(n_198), .B2(n_200), .Y(n_197) );
OAI22xp5_ASAP7_75t_L g250 ( .A1(n_160), .A2(n_178), .B1(n_251), .B2(n_252), .Y(n_250) );
INVx4_ASAP7_75t_L g535 ( .A(n_160), .Y(n_535) );
NAND3xp33_ASAP7_75t_L g274 ( .A(n_161), .B(n_249), .C(n_250), .Y(n_274) );
BUFx3_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
OAI21xp5_ASAP7_75t_L g171 ( .A1(n_162), .A2(n_172), .B(n_175), .Y(n_171) );
OAI21xp5_ASAP7_75t_L g181 ( .A1(n_162), .A2(n_182), .B(n_189), .Y(n_181) );
OAI21xp5_ASAP7_75t_L g205 ( .A1(n_162), .A2(n_206), .B(n_210), .Y(n_205) );
OAI21xp5_ASAP7_75t_L g215 ( .A1(n_162), .A2(n_216), .B(n_221), .Y(n_215) );
AND2x4_ASAP7_75t_L g456 ( .A(n_162), .B(n_457), .Y(n_456) );
INVx4_ASAP7_75t_SL g470 ( .A(n_162), .Y(n_470) );
NAND2x1p5_ASAP7_75t_L g544 ( .A(n_162), .B(n_457), .Y(n_544) );
OA21x2_ASAP7_75t_L g204 ( .A1(n_165), .A2(n_205), .B(n_213), .Y(n_204) );
OA21x2_ASAP7_75t_L g214 ( .A1(n_165), .A2(n_215), .B(n_224), .Y(n_214) );
INVx2_ASAP7_75t_L g239 ( .A(n_165), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g454 ( .A1(n_165), .A2(n_455), .B(n_458), .Y(n_454) );
AOI21xp5_ASAP7_75t_L g496 ( .A1(n_165), .A2(n_497), .B(n_498), .Y(n_496) );
INVx1_ASAP7_75t_L g516 ( .A(n_165), .Y(n_516) );
NOR2xp33_ASAP7_75t_L g369 ( .A(n_166), .B(n_313), .Y(n_369) );
INVx2_ASAP7_75t_SL g166 ( .A(n_167), .Y(n_166) );
OAI311xp33_ASAP7_75t_L g311 ( .A1(n_167), .A2(n_312), .A3(n_313), .B1(n_314), .C1(n_329), .Y(n_311) );
AND2x2_ASAP7_75t_L g167 ( .A(n_168), .B(n_180), .Y(n_167) );
AND2x2_ASAP7_75t_L g272 ( .A(n_168), .B(n_273), .Y(n_272) );
INVx2_ASAP7_75t_L g279 ( .A(n_168), .Y(n_279) );
AND2x2_ASAP7_75t_L g400 ( .A(n_168), .B(n_229), .Y(n_400) );
INVx3_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_169), .B(n_229), .Y(n_228) );
AND2x2_ASAP7_75t_L g256 ( .A(n_169), .B(n_180), .Y(n_256) );
AND2x2_ASAP7_75t_L g308 ( .A(n_169), .B(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g322 ( .A(n_169), .B(n_255), .Y(n_322) );
OA21x2_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_171), .B(n_179), .Y(n_169) );
INVx4_ASAP7_75t_L g249 ( .A(n_170), .Y(n_249) );
HB1xp67_ASAP7_75t_L g475 ( .A(n_170), .Y(n_475) );
AOI21xp5_ASAP7_75t_L g486 ( .A1(n_170), .A2(n_487), .B(n_488), .Y(n_486) );
AOI21xp5_ASAP7_75t_L g175 ( .A1(n_176), .A2(n_177), .B(n_178), .Y(n_175) );
INVx2_ASAP7_75t_L g229 ( .A(n_180), .Y(n_229) );
AND2x2_ASAP7_75t_L g271 ( .A(n_180), .B(n_255), .Y(n_271) );
O2A1O1Ixp33_ASAP7_75t_L g182 ( .A1(n_183), .A2(n_184), .B(n_185), .C(n_186), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g489 ( .A1(n_184), .A2(n_490), .B(n_491), .Y(n_489) );
AOI21xp5_ASAP7_75t_L g546 ( .A1(n_184), .A2(n_547), .B(n_548), .Y(n_546) );
O2A1O1Ixp33_ASAP7_75t_L g521 ( .A1(n_186), .A2(n_522), .B(n_523), .C(n_524), .Y(n_521) );
INVx1_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_187), .A2(n_211), .B(n_212), .Y(n_210) );
INVx4_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx2_ASAP7_75t_L g466 ( .A(n_188), .Y(n_466) );
AND2x2_ASAP7_75t_L g193 ( .A(n_194), .B(n_201), .Y(n_193) );
OR2x2_ASAP7_75t_L g366 ( .A(n_194), .B(n_367), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_194), .B(n_372), .Y(n_383) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
NOR2xp33_ASAP7_75t_L g378 ( .A(n_195), .B(n_379), .Y(n_378) );
BUFx2_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
INVx2_ASAP7_75t_L g240 ( .A(n_196), .Y(n_240) );
AND2x2_ASAP7_75t_L g307 ( .A(n_196), .B(n_234), .Y(n_307) );
AND2x2_ASAP7_75t_L g318 ( .A(n_196), .B(n_214), .Y(n_318) );
AND2x2_ASAP7_75t_L g327 ( .A(n_196), .B(n_328), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_201), .B(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_201), .B(n_268), .Y(n_312) );
INVx2_ASAP7_75t_SL g201 ( .A(n_202), .Y(n_201) );
OR2x2_ASAP7_75t_L g299 ( .A(n_202), .B(n_258), .Y(n_299) );
OR2x2_ASAP7_75t_L g202 ( .A(n_203), .B(n_214), .Y(n_202) );
INVx2_ASAP7_75t_L g232 ( .A(n_203), .Y(n_232) );
AND2x2_ASAP7_75t_L g326 ( .A(n_203), .B(n_327), .Y(n_326) );
INVx2_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
INVx2_ASAP7_75t_L g244 ( .A(n_204), .Y(n_244) );
OR2x2_ASAP7_75t_L g343 ( .A(n_204), .B(n_344), .Y(n_343) );
HB1xp67_ASAP7_75t_L g406 ( .A(n_204), .Y(n_406) );
AND2x2_ASAP7_75t_L g245 ( .A(n_214), .B(n_240), .Y(n_245) );
INVx1_ASAP7_75t_L g266 ( .A(n_214), .Y(n_266) );
AND2x2_ASAP7_75t_L g287 ( .A(n_214), .B(n_288), .Y(n_287) );
INVx2_ASAP7_75t_L g328 ( .A(n_214), .Y(n_328) );
INVx1_ASAP7_75t_L g344 ( .A(n_214), .Y(n_344) );
HB1xp67_ASAP7_75t_L g419 ( .A(n_214), .Y(n_419) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_217), .A2(n_218), .B(n_219), .Y(n_216) );
INVx1_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
INVxp67_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_227), .B(n_332), .Y(n_373) );
OAI22xp5_ASAP7_75t_L g375 ( .A1(n_227), .A2(n_317), .B1(n_366), .B2(n_376), .Y(n_375) );
INVx1_ASAP7_75t_SL g227 ( .A(n_228), .Y(n_227) );
OAI211xp5_ASAP7_75t_SL g409 ( .A1(n_228), .A2(n_410), .B(n_412), .C(n_430), .Y(n_409) );
INVx2_ASAP7_75t_L g262 ( .A(n_229), .Y(n_262) );
AND2x2_ASAP7_75t_L g320 ( .A(n_229), .B(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g331 ( .A(n_229), .B(n_332), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_230), .B(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g230 ( .A(n_231), .B(n_233), .Y(n_230) );
AND2x2_ASAP7_75t_L g304 ( .A(n_231), .B(n_268), .Y(n_304) );
BUFx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
AND2x2_ASAP7_75t_L g336 ( .A(n_232), .B(n_327), .Y(n_336) );
AND2x2_ASAP7_75t_L g355 ( .A(n_232), .B(n_269), .Y(n_355) );
AND2x4_ASAP7_75t_L g291 ( .A(n_233), .B(n_265), .Y(n_291) );
AND2x2_ASAP7_75t_L g429 ( .A(n_233), .B(n_405), .Y(n_429) );
AND2x2_ASAP7_75t_L g233 ( .A(n_234), .B(n_240), .Y(n_233) );
BUFx6f_ASAP7_75t_L g258 ( .A(n_234), .Y(n_258) );
INVx1_ASAP7_75t_L g269 ( .A(n_234), .Y(n_269) );
INVx1_ASAP7_75t_L g368 ( .A(n_234), .Y(n_368) );
HB1xp67_ASAP7_75t_L g468 ( .A(n_237), .Y(n_468) );
INVx2_ASAP7_75t_L g536 ( .A(n_237), .Y(n_536) );
INVx1_ASAP7_75t_L g513 ( .A(n_239), .Y(n_513) );
OR2x2_ASAP7_75t_L g259 ( .A(n_240), .B(n_244), .Y(n_259) );
AND2x2_ASAP7_75t_L g268 ( .A(n_240), .B(n_269), .Y(n_268) );
NOR2xp67_ASAP7_75t_L g288 ( .A(n_240), .B(n_289), .Y(n_288) );
OAI221xp5_ASAP7_75t_L g241 ( .A1(n_242), .A2(n_246), .B1(n_257), .B2(n_260), .C(n_264), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
A2O1A1Ixp33_ASAP7_75t_L g264 ( .A1(n_243), .A2(n_265), .B(n_267), .C(n_270), .Y(n_264) );
AND2x2_ASAP7_75t_L g243 ( .A(n_244), .B(n_245), .Y(n_243) );
INVx1_ASAP7_75t_L g289 ( .A(n_244), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_244), .B(n_368), .Y(n_367) );
AND2x2_ASAP7_75t_SL g372 ( .A(n_244), .B(n_266), .Y(n_372) );
HB1xp67_ASAP7_75t_L g379 ( .A(n_244), .Y(n_379) );
AND2x2_ASAP7_75t_L g297 ( .A(n_245), .B(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g334 ( .A(n_245), .B(n_335), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_247), .B(n_256), .Y(n_246) );
INVx2_ASAP7_75t_L g325 ( .A(n_247), .Y(n_325) );
AOI222xp33_ASAP7_75t_L g374 ( .A1(n_247), .A2(n_258), .B1(n_375), .B2(n_377), .C1(n_378), .C2(n_380), .Y(n_374) );
AND2x2_ASAP7_75t_L g431 ( .A(n_247), .B(n_400), .Y(n_431) );
AND2x2_ASAP7_75t_L g247 ( .A(n_248), .B(n_255), .Y(n_247) );
INVx1_ASAP7_75t_L g321 ( .A(n_248), .Y(n_321) );
AO21x1_ASAP7_75t_L g248 ( .A1(n_249), .A2(n_250), .B(n_253), .Y(n_248) );
INVx3_ASAP7_75t_L g483 ( .A(n_249), .Y(n_483) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_249), .B(n_503), .Y(n_502) );
AO21x2_ASAP7_75t_L g518 ( .A1(n_249), .A2(n_519), .B(n_526), .Y(n_518) );
NOR2xp33_ASAP7_75t_L g526 ( .A(n_249), .B(n_527), .Y(n_526) );
AO21x2_ASAP7_75t_L g541 ( .A1(n_249), .A2(n_542), .B(n_549), .Y(n_541) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
AND2x4_ASAP7_75t_L g273 ( .A(n_254), .B(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g359 ( .A(n_256), .B(n_293), .Y(n_359) );
AOI21xp33_ASAP7_75t_L g370 ( .A1(n_257), .A2(n_371), .B(n_373), .Y(n_370) );
OR2x2_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
INVx2_ASAP7_75t_L g298 ( .A(n_258), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_258), .B(n_265), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_258), .B(n_411), .Y(n_410) );
INVx1_ASAP7_75t_SL g260 ( .A(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g261 ( .A(n_262), .B(n_263), .Y(n_261) );
INVx3_ASAP7_75t_L g324 ( .A(n_262), .Y(n_324) );
OR2x2_ASAP7_75t_L g376 ( .A(n_262), .B(n_298), .Y(n_376) );
AND2x2_ASAP7_75t_L g292 ( .A(n_263), .B(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g330 ( .A(n_263), .B(n_331), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_263), .B(n_324), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_263), .B(n_320), .Y(n_346) );
AND2x2_ASAP7_75t_L g350 ( .A(n_263), .B(n_332), .Y(n_350) );
INVxp67_ASAP7_75t_L g282 ( .A(n_265), .Y(n_282) );
BUFx3_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
OAI22xp5_ASAP7_75t_L g339 ( .A1(n_267), .A2(n_340), .B1(n_345), .B2(n_346), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_267), .B(n_372), .Y(n_402) );
INVx1_ASAP7_75t_SL g267 ( .A(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g388 ( .A(n_268), .B(n_379), .Y(n_388) );
AND2x2_ASAP7_75t_L g417 ( .A(n_268), .B(n_418), .Y(n_417) );
AND2x2_ASAP7_75t_L g422 ( .A(n_268), .B(n_372), .Y(n_422) );
INVx1_ASAP7_75t_L g335 ( .A(n_269), .Y(n_335) );
BUFx2_ASAP7_75t_L g341 ( .A(n_269), .Y(n_341) );
INVx1_ASAP7_75t_L g426 ( .A(n_270), .Y(n_426) );
AND2x2_ASAP7_75t_L g270 ( .A(n_271), .B(n_272), .Y(n_270) );
NAND2x1p5_ASAP7_75t_L g277 ( .A(n_271), .B(n_278), .Y(n_277) );
INVx1_ASAP7_75t_L g302 ( .A(n_272), .Y(n_302) );
NOR2x1_ASAP7_75t_L g278 ( .A(n_273), .B(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g285 ( .A(n_273), .B(n_286), .Y(n_285) );
INVx2_ASAP7_75t_L g294 ( .A(n_273), .Y(n_294) );
INVx3_ASAP7_75t_L g332 ( .A(n_273), .Y(n_332) );
OR2x2_ASAP7_75t_L g398 ( .A(n_273), .B(n_399), .Y(n_398) );
AOI211xp5_ASAP7_75t_L g275 ( .A1(n_276), .A2(n_280), .B(n_283), .C(n_295), .Y(n_275) );
AOI221xp5_ASAP7_75t_L g412 ( .A1(n_276), .A2(n_413), .B1(n_420), .B2(n_422), .C(n_423), .Y(n_412) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
NAND2xp5_ASAP7_75t_SL g283 ( .A(n_284), .B(n_290), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_285), .B(n_287), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_286), .B(n_324), .Y(n_338) );
AND2x2_ASAP7_75t_L g380 ( .A(n_286), .B(n_320), .Y(n_380) );
INVx1_ASAP7_75t_SL g393 ( .A(n_287), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_287), .B(n_341), .Y(n_396) );
INVx1_ASAP7_75t_L g414 ( .A(n_288), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_291), .B(n_292), .Y(n_290) );
AOI221xp5_ASAP7_75t_L g381 ( .A1(n_292), .A2(n_382), .B1(n_384), .B2(n_388), .C(n_389), .Y(n_381) );
AND2x2_ASAP7_75t_L g408 ( .A(n_293), .B(n_400), .Y(n_408) );
INVx2_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g392 ( .A(n_294), .Y(n_392) );
AOI21xp33_ASAP7_75t_SL g295 ( .A1(n_296), .A2(n_299), .B(n_300), .Y(n_295) );
INVx1_ASAP7_75t_SL g296 ( .A(n_297), .Y(n_296) );
OR2x2_ASAP7_75t_L g363 ( .A(n_298), .B(n_364), .Y(n_363) );
INVx2_ASAP7_75t_L g349 ( .A(n_299), .Y(n_349) );
INVx1_ASAP7_75t_L g377 ( .A(n_300), .Y(n_377) );
OR2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
O2A1O1Ixp33_ASAP7_75t_L g303 ( .A1(n_304), .A2(n_305), .B(n_308), .C(n_311), .Y(n_303) );
OAI31xp33_ASAP7_75t_L g430 ( .A1(n_304), .A2(n_342), .A3(n_429), .B(n_431), .Y(n_430) );
INVxp67_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g404 ( .A(n_307), .B(n_405), .Y(n_404) );
INVx1_ASAP7_75t_SL g425 ( .A(n_307), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_309), .B(n_324), .Y(n_352) );
INVx1_ASAP7_75t_SL g309 ( .A(n_310), .Y(n_309) );
OR2x2_ASAP7_75t_L g427 ( .A(n_310), .B(n_324), .Y(n_427) );
AOI22xp5_ASAP7_75t_L g314 ( .A1(n_315), .A2(n_319), .B1(n_323), .B2(n_326), .Y(n_314) );
NAND2xp33_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
INVx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_318), .B(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g354 ( .A(n_318), .B(n_355), .Y(n_354) );
AND2x2_ASAP7_75t_L g357 ( .A(n_318), .B(n_341), .Y(n_357) );
AND2x2_ASAP7_75t_L g411 ( .A(n_318), .B(n_406), .Y(n_411) );
AND2x2_ASAP7_75t_L g319 ( .A(n_320), .B(n_322), .Y(n_319) );
INVx1_ASAP7_75t_L g386 ( .A(n_322), .Y(n_386) );
NOR2xp67_ASAP7_75t_L g323 ( .A(n_324), .B(n_325), .Y(n_323) );
OAI32xp33_ASAP7_75t_L g389 ( .A1(n_324), .A2(n_358), .A3(n_390), .B1(n_392), .B2(n_393), .Y(n_389) );
INVx1_ASAP7_75t_L g364 ( .A(n_327), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_327), .B(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g387 ( .A(n_331), .Y(n_387) );
O2A1O1Ixp33_ASAP7_75t_L g333 ( .A1(n_334), .A2(n_336), .B(n_337), .C(n_339), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_335), .B(n_372), .Y(n_371) );
AOI221xp5_ASAP7_75t_L g347 ( .A1(n_336), .A2(n_348), .B1(n_349), .B2(n_350), .C(n_351), .Y(n_347) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_341), .B(n_342), .Y(n_340) );
INVx2_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g348 ( .A(n_346), .Y(n_348) );
OAI22xp5_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_353), .B1(n_356), .B2(n_358), .Y(n_351) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
NAND4xp25_ASAP7_75t_SL g413 ( .A(n_356), .B(n_414), .C(n_415), .D(n_416), .Y(n_413) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_SL g358 ( .A(n_359), .Y(n_358) );
NAND4xp25_ASAP7_75t_SL g360 ( .A(n_361), .B(n_374), .C(n_381), .D(n_394), .Y(n_360) );
O2A1O1Ixp33_ASAP7_75t_L g361 ( .A1(n_362), .A2(n_365), .B(n_369), .C(n_370), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_SL g391 ( .A(n_367), .Y(n_391) );
INVx2_ASAP7_75t_L g415 ( .A(n_372), .Y(n_415) );
OR2x2_ASAP7_75t_L g424 ( .A(n_379), .B(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx2_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
OR2x2_ASAP7_75t_L g385 ( .A(n_386), .B(n_387), .Y(n_385) );
AOI21xp5_ASAP7_75t_L g394 ( .A1(n_395), .A2(n_397), .B(n_401), .Y(n_394) );
INVxp67_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx2_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
AND2x2_ASAP7_75t_L g420 ( .A(n_400), .B(n_421), .Y(n_420) );
AOI21xp33_ASAP7_75t_SL g401 ( .A1(n_402), .A2(n_403), .B(n_407), .Y(n_401) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
CKINVDCx16_ASAP7_75t_R g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
OAI22xp5_ASAP7_75t_L g423 ( .A1(n_424), .A2(n_426), .B1(n_427), .B2(n_428), .Y(n_423) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
NAND3xp33_ASAP7_75t_SL g436 ( .A(n_432), .B(n_437), .C(n_439), .Y(n_436) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVxp67_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
OAI22xp5_ASAP7_75t_L g440 ( .A1(n_441), .A2(n_444), .B1(n_446), .B2(n_449), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g748 ( .A(n_442), .Y(n_748) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g749 ( .A(n_444), .Y(n_749) );
INVx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g750 ( .A(n_447), .Y(n_750) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx4_ASAP7_75t_L g751 ( .A(n_449), .Y(n_751) );
BUFx6f_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
OR5x1_ASAP7_75t_L g450 ( .A(n_451), .B(n_620), .C(n_698), .D(n_722), .E(n_739), .Y(n_450) );
OAI211xp5_ASAP7_75t_SL g451 ( .A1(n_452), .A2(n_492), .B(n_538), .C(n_597), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_453), .B(n_472), .Y(n_452) );
AND2x2_ASAP7_75t_L g551 ( .A(n_453), .B(n_474), .Y(n_551) );
INVx5_ASAP7_75t_SL g579 ( .A(n_453), .Y(n_579) );
AND2x2_ASAP7_75t_L g615 ( .A(n_453), .B(n_600), .Y(n_615) );
OR2x2_ASAP7_75t_L g654 ( .A(n_453), .B(n_473), .Y(n_654) );
OR2x2_ASAP7_75t_L g685 ( .A(n_453), .B(n_576), .Y(n_685) );
NOR2xp33_ASAP7_75t_L g721 ( .A(n_453), .B(n_589), .Y(n_721) );
AND2x2_ASAP7_75t_L g733 ( .A(n_453), .B(n_576), .Y(n_733) );
OR2x6_ASAP7_75t_L g453 ( .A(n_454), .B(n_471), .Y(n_453) );
BUFx2_ASAP7_75t_L g508 ( .A(n_456), .Y(n_508) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
O2A1O1Ixp33_ASAP7_75t_L g477 ( .A1(n_460), .A2(n_470), .B(n_478), .C(n_479), .Y(n_477) );
O2A1O1Ixp33_ASAP7_75t_SL g530 ( .A1(n_460), .A2(n_470), .B(n_531), .C(n_532), .Y(n_530) );
INVx5_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
O2A1O1Ixp33_ASAP7_75t_L g463 ( .A1(n_464), .A2(n_465), .B(n_467), .C(n_468), .Y(n_463) );
O2A1O1Ixp33_ASAP7_75t_L g499 ( .A1(n_465), .A2(n_468), .B(n_500), .C(n_501), .Y(n_499) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
AND2x2_ASAP7_75t_L g732 ( .A(n_472), .B(n_733), .Y(n_732) );
INVx1_ASAP7_75t_SL g472 ( .A(n_473), .Y(n_472) );
OR2x2_ASAP7_75t_L g595 ( .A(n_473), .B(n_596), .Y(n_595) );
OR2x2_ASAP7_75t_L g473 ( .A(n_474), .B(n_484), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_474), .B(n_576), .Y(n_575) );
HB1xp67_ASAP7_75t_L g588 ( .A(n_474), .Y(n_588) );
INVx3_ASAP7_75t_L g603 ( .A(n_474), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_474), .B(n_484), .Y(n_627) );
OR2x2_ASAP7_75t_L g636 ( .A(n_474), .B(n_579), .Y(n_636) );
AND2x2_ASAP7_75t_L g640 ( .A(n_474), .B(n_600), .Y(n_640) );
AND2x2_ASAP7_75t_L g646 ( .A(n_474), .B(n_647), .Y(n_646) );
INVxp67_ASAP7_75t_L g683 ( .A(n_474), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_474), .B(n_541), .Y(n_697) );
OA21x2_ASAP7_75t_L g474 ( .A1(n_475), .A2(n_476), .B(n_482), .Y(n_474) );
OA21x2_ASAP7_75t_L g528 ( .A1(n_483), .A2(n_529), .B(n_537), .Y(n_528) );
OR2x2_ASAP7_75t_L g589 ( .A(n_484), .B(n_541), .Y(n_589) );
AND2x2_ASAP7_75t_L g600 ( .A(n_484), .B(n_576), .Y(n_600) );
AND2x2_ASAP7_75t_L g612 ( .A(n_484), .B(n_603), .Y(n_612) );
NAND2xp5_ASAP7_75t_SL g635 ( .A(n_484), .B(n_541), .Y(n_635) );
INVx1_ASAP7_75t_SL g647 ( .A(n_484), .Y(n_647) );
INVx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
AND2x2_ASAP7_75t_L g540 ( .A(n_485), .B(n_541), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_485), .B(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_494), .B(n_504), .Y(n_493) );
AND2x2_ASAP7_75t_L g560 ( .A(n_494), .B(n_561), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_494), .B(n_517), .Y(n_564) );
AND2x2_ASAP7_75t_L g567 ( .A(n_494), .B(n_568), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_494), .B(n_570), .Y(n_569) );
OR2x2_ASAP7_75t_L g592 ( .A(n_494), .B(n_583), .Y(n_592) );
HB1xp67_ASAP7_75t_L g611 ( .A(n_494), .Y(n_611) );
AND2x2_ASAP7_75t_L g632 ( .A(n_494), .B(n_633), .Y(n_632) );
OR2x2_ASAP7_75t_L g642 ( .A(n_494), .B(n_643), .Y(n_642) );
AND2x2_ASAP7_75t_L g688 ( .A(n_494), .B(n_571), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_494), .B(n_594), .Y(n_715) );
INVx5_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
BUFx2_ASAP7_75t_L g585 ( .A(n_495), .Y(n_585) );
AND2x2_ASAP7_75t_L g651 ( .A(n_495), .B(n_583), .Y(n_651) );
AND2x2_ASAP7_75t_L g735 ( .A(n_495), .B(n_603), .Y(n_735) );
OR2x6_ASAP7_75t_L g495 ( .A(n_496), .B(n_502), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_504), .B(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g724 ( .A(n_504), .Y(n_724) );
AND2x2_ASAP7_75t_L g504 ( .A(n_505), .B(n_517), .Y(n_504) );
AND2x2_ASAP7_75t_L g554 ( .A(n_505), .B(n_555), .Y(n_554) );
AND2x4_ASAP7_75t_L g563 ( .A(n_505), .B(n_561), .Y(n_563) );
INVx5_ASAP7_75t_L g571 ( .A(n_505), .Y(n_571) );
AND2x2_ASAP7_75t_L g594 ( .A(n_505), .B(n_528), .Y(n_594) );
HB1xp67_ASAP7_75t_L g631 ( .A(n_505), .Y(n_631) );
OR2x6_ASAP7_75t_L g505 ( .A(n_506), .B(n_514), .Y(n_505) );
AOI21xp5_ASAP7_75t_SL g506 ( .A1(n_507), .A2(n_509), .B(n_513), .Y(n_506) );
NOR2xp33_ASAP7_75t_L g514 ( .A(n_515), .B(n_516), .Y(n_514) );
INVx1_ASAP7_75t_L g672 ( .A(n_517), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_517), .B(n_688), .Y(n_687) );
AND2x2_ASAP7_75t_L g705 ( .A(n_517), .B(n_571), .Y(n_705) );
A2O1A1Ixp33_ASAP7_75t_L g734 ( .A1(n_517), .A2(n_628), .B(n_735), .C(n_736), .Y(n_734) );
AND2x2_ASAP7_75t_L g517 ( .A(n_518), .B(n_528), .Y(n_517) );
BUFx2_ASAP7_75t_L g555 ( .A(n_518), .Y(n_555) );
INVx2_ASAP7_75t_L g559 ( .A(n_518), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_520), .B(n_525), .Y(n_519) );
INVx2_ASAP7_75t_L g561 ( .A(n_528), .Y(n_561) );
AND2x2_ASAP7_75t_L g568 ( .A(n_528), .B(n_559), .Y(n_568) );
AND2x2_ASAP7_75t_L g659 ( .A(n_528), .B(n_571), .Y(n_659) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_534), .B(n_535), .Y(n_533) );
AOI211x1_ASAP7_75t_SL g538 ( .A1(n_539), .A2(n_552), .B(n_565), .C(n_590), .Y(n_538) );
INVx1_ASAP7_75t_L g656 ( .A(n_539), .Y(n_656) );
AND2x2_ASAP7_75t_L g539 ( .A(n_540), .B(n_551), .Y(n_539) );
INVx5_ASAP7_75t_SL g576 ( .A(n_541), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_541), .B(n_646), .Y(n_645) );
AOI311xp33_ASAP7_75t_L g664 ( .A1(n_541), .A2(n_665), .A3(n_667), .B(n_668), .C(n_674), .Y(n_664) );
A2O1A1Ixp33_ASAP7_75t_L g699 ( .A1(n_541), .A2(n_612), .B(n_700), .C(n_703), .Y(n_699) );
OAI21xp5_ASAP7_75t_L g542 ( .A1(n_543), .A2(n_544), .B(n_545), .Y(n_542) );
INVxp67_ASAP7_75t_L g619 ( .A(n_551), .Y(n_619) );
NAND4xp25_ASAP7_75t_SL g552 ( .A(n_553), .B(n_556), .C(n_562), .D(n_564), .Y(n_552) );
NOR2xp33_ASAP7_75t_L g617 ( .A(n_553), .B(n_618), .Y(n_617) );
INVx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g610 ( .A(n_554), .B(n_611), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_557), .B(n_560), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_557), .B(n_563), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_557), .B(n_570), .Y(n_690) );
BUFx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_558), .B(n_571), .Y(n_708) );
HB1xp67_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx2_ASAP7_75t_L g583 ( .A(n_559), .Y(n_583) );
INVxp67_ASAP7_75t_L g618 ( .A(n_560), .Y(n_618) );
AND2x4_ASAP7_75t_L g570 ( .A(n_561), .B(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g644 ( .A(n_561), .B(n_583), .Y(n_644) );
INVx1_ASAP7_75t_L g671 ( .A(n_561), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_561), .B(n_658), .Y(n_718) );
NOR2xp33_ASAP7_75t_L g652 ( .A(n_562), .B(n_632), .Y(n_652) );
INVx1_ASAP7_75t_SL g562 ( .A(n_563), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_563), .B(n_585), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_563), .B(n_632), .Y(n_731) );
INVx1_ASAP7_75t_L g742 ( .A(n_564), .Y(n_742) );
A2O1A1Ixp33_ASAP7_75t_L g565 ( .A1(n_566), .A2(n_569), .B(n_572), .C(n_580), .Y(n_565) );
INVx1_ASAP7_75t_SL g566 ( .A(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g584 ( .A(n_568), .B(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_L g622 ( .A(n_568), .B(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g604 ( .A(n_569), .Y(n_604) );
AND2x2_ASAP7_75t_L g581 ( .A(n_570), .B(n_582), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_570), .B(n_632), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_570), .B(n_651), .Y(n_675) );
OR2x2_ASAP7_75t_L g591 ( .A(n_571), .B(n_592), .Y(n_591) );
INVx2_ASAP7_75t_L g623 ( .A(n_571), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_571), .B(n_583), .Y(n_638) );
AND2x2_ASAP7_75t_L g695 ( .A(n_571), .B(n_651), .Y(n_695) );
HB1xp67_ASAP7_75t_L g702 ( .A(n_571), .Y(n_702) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
AOI221xp5_ASAP7_75t_L g706 ( .A1(n_573), .A2(n_585), .B1(n_707), .B2(n_709), .C(n_712), .Y(n_706) );
AND2x2_ASAP7_75t_L g573 ( .A(n_574), .B(n_577), .Y(n_573) );
INVx1_ASAP7_75t_SL g574 ( .A(n_575), .Y(n_574) );
OR2x2_ASAP7_75t_L g596 ( .A(n_576), .B(n_579), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_576), .B(n_646), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_576), .B(n_603), .Y(n_711) );
INVx1_ASAP7_75t_SL g577 ( .A(n_578), .Y(n_577) );
OR2x2_ASAP7_75t_L g696 ( .A(n_578), .B(n_697), .Y(n_696) );
OR2x2_ASAP7_75t_L g710 ( .A(n_578), .B(n_711), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_579), .B(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g607 ( .A(n_579), .B(n_600), .Y(n_607) );
AND2x2_ASAP7_75t_L g677 ( .A(n_579), .B(n_678), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_579), .B(n_626), .Y(n_723) );
NOR2xp33_ASAP7_75t_L g726 ( .A(n_579), .B(n_727), .Y(n_726) );
OAI21xp5_ASAP7_75t_SL g580 ( .A1(n_581), .A2(n_584), .B(n_586), .Y(n_580) );
INVx2_ASAP7_75t_L g613 ( .A(n_581), .Y(n_613) );
HB1xp67_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g633 ( .A(n_583), .Y(n_633) );
OR2x2_ASAP7_75t_L g637 ( .A(n_585), .B(n_638), .Y(n_637) );
OR2x2_ASAP7_75t_L g740 ( .A(n_585), .B(n_708), .Y(n_740) );
INVx1_ASAP7_75t_SL g586 ( .A(n_587), .Y(n_586) );
OR2x2_ASAP7_75t_L g587 ( .A(n_588), .B(n_589), .Y(n_587) );
AOI21xp33_ASAP7_75t_SL g590 ( .A1(n_591), .A2(n_593), .B(n_595), .Y(n_590) );
INVx1_ASAP7_75t_L g744 ( .A(n_591), .Y(n_744) );
INVx2_ASAP7_75t_SL g658 ( .A(n_592), .Y(n_658) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
A2O1A1Ixp33_ASAP7_75t_L g739 ( .A1(n_595), .A2(n_676), .B(n_740), .C(n_741), .Y(n_739) );
OAI322xp33_ASAP7_75t_SL g608 ( .A1(n_596), .A2(n_609), .A3(n_612), .B1(n_613), .B2(n_614), .C1(n_616), .C2(n_619), .Y(n_608) );
INVx2_ASAP7_75t_L g628 ( .A(n_596), .Y(n_628) );
AOI221xp5_ASAP7_75t_L g597 ( .A1(n_598), .A2(n_604), .B1(n_605), .B2(n_607), .C(n_608), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
OAI22xp33_ASAP7_75t_SL g674 ( .A1(n_599), .A2(n_675), .B1(n_676), .B2(n_679), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_600), .B(n_601), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_600), .B(n_603), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_600), .B(n_738), .Y(n_737) );
INVx2_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
OR2x2_ASAP7_75t_L g673 ( .A(n_602), .B(n_635), .Y(n_673) );
INVx1_ASAP7_75t_L g663 ( .A(n_603), .Y(n_663) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
AOI21xp5_ASAP7_75t_L g716 ( .A1(n_607), .A2(n_717), .B(n_719), .Y(n_716) );
AOI21xp33_ASAP7_75t_L g641 ( .A1(n_609), .A2(n_642), .B(n_645), .Y(n_641) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
NOR2xp67_ASAP7_75t_SL g670 ( .A(n_611), .B(n_671), .Y(n_670) );
NOR2xp33_ASAP7_75t_L g703 ( .A(n_611), .B(n_704), .Y(n_703) );
INVx1_ASAP7_75t_SL g727 ( .A(n_612), .Y(n_727) );
INVx1_ASAP7_75t_SL g614 ( .A(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
NAND4xp25_ASAP7_75t_L g620 ( .A(n_621), .B(n_648), .C(n_664), .D(n_680), .Y(n_620) );
AOI211xp5_ASAP7_75t_L g621 ( .A1(n_622), .A2(n_624), .B(n_629), .C(n_641), .Y(n_621) );
INVx1_ASAP7_75t_L g713 ( .A(n_622), .Y(n_713) );
AND2x2_ASAP7_75t_L g661 ( .A(n_623), .B(n_644), .Y(n_661) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_626), .B(n_628), .Y(n_625) );
INVx1_ASAP7_75t_SL g626 ( .A(n_627), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_628), .B(n_663), .Y(n_662) );
OAI22xp33_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_634), .B1(n_637), .B2(n_639), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_631), .B(n_632), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_631), .B(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g679 ( .A(n_632), .Y(n_679) );
O2A1O1Ixp33_ASAP7_75t_L g693 ( .A1(n_632), .A2(n_671), .B(n_694), .C(n_696), .Y(n_693) );
OR2x2_ASAP7_75t_L g634 ( .A(n_635), .B(n_636), .Y(n_634) );
INVx1_ASAP7_75t_L g678 ( .A(n_635), .Y(n_678) );
INVx1_ASAP7_75t_L g738 ( .A(n_636), .Y(n_738) );
NAND2xp33_ASAP7_75t_SL g728 ( .A(n_637), .B(n_729), .Y(n_728) );
INVx1_ASAP7_75t_SL g639 ( .A(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx2_ASAP7_75t_L g667 ( .A(n_646), .Y(n_667) );
O2A1O1Ixp33_ASAP7_75t_L g648 ( .A1(n_649), .A2(n_652), .B(n_653), .C(n_655), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
OAI22xp5_ASAP7_75t_L g655 ( .A1(n_656), .A2(n_657), .B1(n_660), .B2(n_662), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_658), .B(n_659), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_658), .B(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_663), .B(n_684), .Y(n_746) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
AOI21xp33_ASAP7_75t_SL g668 ( .A1(n_669), .A2(n_672), .B(n_673), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_SL g676 ( .A(n_677), .Y(n_676) );
AOI221xp5_ASAP7_75t_L g680 ( .A1(n_681), .A2(n_686), .B1(n_689), .B2(n_691), .C(n_693), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_683), .B(n_684), .Y(n_682) );
INVx1_ASAP7_75t_SL g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVxp67_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
OAI22xp5_ASAP7_75t_L g712 ( .A1(n_696), .A2(n_713), .B1(n_714), .B2(n_715), .Y(n_712) );
NAND3xp33_ASAP7_75t_SL g698 ( .A(n_699), .B(n_706), .C(n_716), .Y(n_698) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_SL g704 ( .A(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
CKINVDCx16_ASAP7_75t_R g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVxp67_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
OAI211xp5_ASAP7_75t_L g722 ( .A1(n_723), .A2(n_724), .B(n_725), .C(n_734), .Y(n_722) );
INVx1_ASAP7_75t_L g743 ( .A(n_723), .Y(n_743) );
AOI22xp33_ASAP7_75t_L g725 ( .A1(n_726), .A2(n_728), .B1(n_730), .B2(n_732), .Y(n_725) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
AOI22xp5_ASAP7_75t_L g741 ( .A1(n_742), .A2(n_743), .B1(n_744), .B2(n_745), .Y(n_741) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
OAI22x1_ASAP7_75t_SL g747 ( .A1(n_748), .A2(n_749), .B1(n_750), .B2(n_751), .Y(n_747) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
endmodule