module fake_jpeg_27148_n_336 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_336);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_336;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_15),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx6f_ASAP7_75t_SL g29 ( 
.A(n_15),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx4f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_21),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_45),
.Y(n_60)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

HB1xp67_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_28),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_0),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_16),
.B(n_14),
.Y(n_46)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_28),
.Y(n_53)
);

CKINVDCx14_ASAP7_75t_R g80 ( 
.A(n_48),
.Y(n_80)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_49),
.Y(n_67)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_52),
.B(n_53),
.Y(n_79)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_55),
.B(n_62),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_56),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_39),
.A2(n_19),
.B1(n_29),
.B2(n_32),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_58),
.A2(n_19),
.B1(n_22),
.B2(n_26),
.Y(n_87)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

BUFx4f_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_64),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_37),
.B(n_16),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_65),
.B(n_31),
.Y(n_83)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx2_ASAP7_75t_SL g76 ( 
.A(n_66),
.Y(n_76)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_69),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_53),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_70),
.B(n_71),
.Y(n_108)
);

OAI211xp5_ASAP7_75t_L g71 ( 
.A1(n_60),
.A2(n_18),
.B(n_17),
.C(n_20),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_54),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_72),
.B(n_74),
.Y(n_124)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_75),
.Y(n_107)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_77),
.B(n_84),
.Y(n_136)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_78),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_60),
.A2(n_19),
.B1(n_17),
.B2(n_18),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_82),
.A2(n_88),
.B1(n_96),
.B2(n_106),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_83),
.B(n_91),
.Y(n_110)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_47),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_85),
.B(n_86),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_53),
.B(n_20),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_87),
.A2(n_102),
.B1(n_35),
.B2(n_33),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_52),
.A2(n_31),
.B1(n_22),
.B2(n_26),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_55),
.B(n_31),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_89),
.A2(n_92),
.B(n_94),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_90),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_47),
.B(n_44),
.C(n_41),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_64),
.B(n_31),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_62),
.A2(n_24),
.B1(n_34),
.B2(n_16),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_93),
.A2(n_35),
.B1(n_33),
.B2(n_25),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_64),
.B(n_28),
.Y(n_94)
);

CKINVDCx14_ASAP7_75t_R g95 ( 
.A(n_57),
.Y(n_95)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_95),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_51),
.A2(n_30),
.B1(n_34),
.B2(n_24),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_51),
.Y(n_97)
);

INVx1_ASAP7_75t_SL g116 ( 
.A(n_97),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_61),
.B(n_16),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_98),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_61),
.Y(n_99)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_99),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_57),
.B(n_23),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_100),
.B(n_101),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_59),
.B(n_30),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_66),
.A2(n_25),
.B1(n_24),
.B2(n_12),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_59),
.Y(n_103)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_103),
.Y(n_125)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_54),
.Y(n_105)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_105),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_52),
.A2(n_34),
.B1(n_23),
.B2(n_28),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_82),
.A2(n_25),
.B1(n_23),
.B2(n_28),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_109),
.A2(n_113),
.B1(n_96),
.B2(n_94),
.Y(n_139)
);

OA22x2_ASAP7_75t_L g113 ( 
.A1(n_85),
.A2(n_44),
.B1(n_41),
.B2(n_40),
.Y(n_113)
);

A2O1A1Ixp33_ASAP7_75t_L g114 ( 
.A1(n_79),
.A2(n_25),
.B(n_23),
.C(n_10),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_114),
.A2(n_89),
.B(n_97),
.Y(n_149)
);

BUFx2_ASAP7_75t_L g115 ( 
.A(n_73),
.Y(n_115)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_115),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_81),
.B(n_23),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_126),
.B(n_129),
.Y(n_140)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_100),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_127),
.B(n_128),
.Y(n_155)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_92),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_81),
.B(n_40),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_92),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_130),
.B(n_133),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_132),
.Y(n_167)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_101),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_135),
.A2(n_104),
.B1(n_80),
.B2(n_91),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_133),
.B(n_79),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_137),
.B(n_150),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_139),
.A2(n_76),
.B1(n_121),
.B2(n_120),
.Y(n_199)
);

AND2x4_ASAP7_75t_L g141 ( 
.A(n_123),
.B(n_94),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_141),
.A2(n_142),
.B(n_161),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_110),
.A2(n_77),
.B(n_67),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_136),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_143),
.B(n_144),
.Y(n_176)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_115),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_118),
.B(n_72),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_145),
.B(n_160),
.Y(n_177)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_119),
.Y(n_146)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_146),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_147),
.A2(n_158),
.B1(n_165),
.B2(n_116),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_110),
.A2(n_74),
.B1(n_89),
.B2(n_88),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_148),
.A2(n_156),
.B1(n_127),
.B2(n_130),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_149),
.A2(n_131),
.B(n_122),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_108),
.B(n_104),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_115),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_151),
.Y(n_168)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_119),
.Y(n_152)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_152),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_117),
.B(n_83),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_153),
.B(n_159),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_120),
.Y(n_154)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_154),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_110),
.A2(n_84),
.B1(n_68),
.B2(n_69),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_123),
.B(n_106),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_157),
.B(n_113),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_112),
.A2(n_68),
.B1(n_103),
.B2(n_75),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_117),
.B(n_99),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_124),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_128),
.A2(n_67),
.B(n_1),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_111),
.B(n_105),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_162),
.B(n_166),
.Y(n_195)
);

MAJx2_ASAP7_75t_L g163 ( 
.A(n_126),
.B(n_25),
.C(n_35),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_163),
.B(n_114),
.C(n_111),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_112),
.A2(n_78),
.B1(n_76),
.B2(n_73),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_113),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_151),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_172),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_141),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_174),
.B(n_175),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_147),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_142),
.B(n_129),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_178),
.B(n_193),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_180),
.A2(n_11),
.B1(n_10),
.B2(n_3),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_161),
.A2(n_141),
.B(n_166),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_181),
.A2(n_190),
.B(n_191),
.Y(n_222)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_159),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_182),
.B(n_185),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_183),
.B(n_14),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_139),
.A2(n_156),
.B1(n_148),
.B2(n_165),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_184),
.A2(n_192),
.B1(n_199),
.B2(n_160),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_153),
.B(n_125),
.Y(n_185)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_158),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_187),
.B(n_189),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_154),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_188),
.B(n_200),
.Y(n_202)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_140),
.Y(n_189)
);

NOR2x1_ASAP7_75t_R g190 ( 
.A(n_141),
.B(n_149),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_140),
.A2(n_113),
.B1(n_125),
.B2(n_122),
.Y(n_192)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_155),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_194),
.B(n_201),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_196),
.A2(n_197),
.B(n_198),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_157),
.A2(n_116),
.B(n_1),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_164),
.A2(n_0),
.B(n_1),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_146),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_152),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_203),
.A2(n_230),
.B1(n_183),
.B2(n_198),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_178),
.B(n_163),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_205),
.B(n_225),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_187),
.A2(n_167),
.B1(n_143),
.B2(n_144),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_206),
.A2(n_174),
.B1(n_172),
.B2(n_168),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_181),
.A2(n_137),
.B(n_167),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_207),
.A2(n_208),
.B(n_209),
.Y(n_241)
);

O2A1O1Ixp33_ASAP7_75t_L g208 ( 
.A1(n_195),
.A2(n_138),
.B(n_134),
.C(n_107),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_179),
.A2(n_134),
.B(n_138),
.Y(n_209)
);

CKINVDCx14_ASAP7_75t_R g210 ( 
.A(n_177),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_210),
.B(n_216),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_184),
.A2(n_175),
.B1(n_192),
.B2(n_182),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_211),
.A2(n_219),
.B1(n_191),
.B2(n_186),
.Y(n_231)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_176),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_212),
.B(n_214),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_193),
.B(n_107),
.C(n_73),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_213),
.B(n_229),
.C(n_204),
.Y(n_252)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_169),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_194),
.B(n_121),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_170),
.B(n_107),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_217),
.Y(n_234)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_169),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_218),
.B(n_226),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_180),
.A2(n_76),
.B1(n_33),
.B2(n_15),
.Y(n_219)
);

XNOR2x1_ASAP7_75t_L g225 ( 
.A(n_190),
.B(n_14),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_185),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_189),
.B(n_168),
.Y(n_228)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_228),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_231),
.A2(n_242),
.B1(n_208),
.B2(n_206),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_233),
.A2(n_250),
.B1(n_171),
.B2(n_173),
.Y(n_263)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_228),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_235),
.B(n_240),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_223),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_237),
.B(n_245),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_212),
.B(n_170),
.Y(n_238)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_238),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_239),
.A2(n_247),
.B(n_249),
.Y(n_275)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_202),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_211),
.A2(n_203),
.B1(n_220),
.B2(n_226),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_230),
.A2(n_219),
.B1(n_220),
.B2(n_224),
.Y(n_243)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_243),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_227),
.B(n_205),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_244),
.B(n_252),
.Y(n_273)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_221),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_221),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_246),
.B(n_215),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_225),
.A2(n_179),
.B1(n_196),
.B2(n_197),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_222),
.A2(n_209),
.B(n_223),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_214),
.A2(n_188),
.B1(n_186),
.B2(n_201),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_213),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_254),
.Y(n_267)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_255),
.Y(n_277)
);

NAND2xp67_ASAP7_75t_SL g257 ( 
.A(n_249),
.B(n_207),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_257),
.A2(n_258),
.B1(n_269),
.B2(n_233),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_238),
.B(n_218),
.Y(n_259)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_259),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_252),
.B(n_227),
.C(n_222),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_260),
.B(n_261),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_244),
.B(n_215),
.C(n_204),
.Y(n_261)
);

INVxp33_ASAP7_75t_SL g262 ( 
.A(n_237),
.Y(n_262)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_262),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_263),
.A2(n_242),
.B1(n_235),
.B2(n_232),
.Y(n_284)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_234),
.Y(n_265)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_265),
.Y(n_280)
);

NOR3xp33_ASAP7_75t_SL g268 ( 
.A(n_248),
.B(n_229),
.C(n_171),
.Y(n_268)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_268),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_231),
.A2(n_173),
.B1(n_2),
.B2(n_3),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_241),
.A2(n_1),
.B(n_2),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_270),
.A2(n_253),
.B1(n_4),
.B2(n_5),
.Y(n_291)
);

BUFx2_ASAP7_75t_L g272 ( 
.A(n_234),
.Y(n_272)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_272),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_SL g274 ( 
.A(n_236),
.B(n_2),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_274),
.B(n_236),
.Y(n_281)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_276),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_281),
.B(n_288),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_284),
.A2(n_285),
.B1(n_287),
.B2(n_289),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_263),
.A2(n_232),
.B1(n_246),
.B2(n_245),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_264),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_286),
.B(n_290),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_271),
.A2(n_241),
.B1(n_240),
.B2(n_250),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_273),
.B(n_251),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_257),
.A2(n_253),
.B1(n_247),
.B2(n_251),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_266),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_291),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_288),
.B(n_267),
.C(n_273),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_295),
.B(n_297),
.C(n_302),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_282),
.B(n_275),
.C(n_261),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_282),
.B(n_289),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_298),
.B(n_304),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_279),
.B(n_280),
.Y(n_299)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_299),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_285),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_301),
.B(n_281),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_287),
.B(n_275),
.C(n_260),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_SL g303 ( 
.A1(n_292),
.A2(n_265),
.B1(n_256),
.B2(n_270),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_303),
.A2(n_272),
.B1(n_4),
.B2(n_5),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_284),
.B(n_266),
.C(n_258),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_283),
.A2(n_277),
.B(n_278),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_306),
.B(n_269),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_308),
.B(n_310),
.Y(n_321)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_299),
.Y(n_310)
);

OR2x2_ASAP7_75t_L g320 ( 
.A(n_311),
.B(n_293),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_297),
.B(n_274),
.Y(n_313)
);

BUFx24_ASAP7_75t_SL g322 ( 
.A(n_313),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_306),
.B(n_268),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_314),
.A2(n_296),
.B1(n_304),
.B2(n_302),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_315),
.A2(n_316),
.B1(n_6),
.B2(n_7),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_294),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_316)
);

NOR2xp67_ASAP7_75t_L g317 ( 
.A(n_312),
.B(n_305),
.Y(n_317)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_317),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_318),
.B(n_319),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_315),
.A2(n_295),
.B1(n_300),
.B2(n_298),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_320),
.B(n_323),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_321),
.B(n_312),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_326),
.A2(n_328),
.B(n_320),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_322),
.B(n_313),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_324),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_329),
.A2(n_330),
.B(n_307),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_325),
.Y(n_332)
);

OAI321xp33_ASAP7_75t_L g333 ( 
.A1(n_332),
.A2(n_327),
.A3(n_309),
.B1(n_308),
.B2(n_293),
.C(n_9),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_333),
.A2(n_6),
.B(n_7),
.Y(n_334)
);

O2A1O1Ixp33_ASAP7_75t_SL g335 ( 
.A1(n_334),
.A2(n_6),
.B(n_8),
.C(n_9),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_8),
.Y(n_336)
);


endmodule