module fake_jpeg_12075_n_645 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_645);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_645;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_6),
.B(n_0),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_8),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_10),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_6),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

BUFx8_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_16),
.Y(n_51)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_10),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_3),
.A2(n_12),
.B(n_15),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_0),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_5),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_11),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_7),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_60),
.Y(n_145)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_61),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_62),
.Y(n_148)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_63),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_64),
.Y(n_152)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_65),
.Y(n_160)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_66),
.Y(n_153)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_67),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_31),
.Y(n_68)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_68),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_19),
.B(n_8),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_69),
.B(n_93),
.Y(n_140)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_70),
.Y(n_130)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_71),
.Y(n_150)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_28),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g125 ( 
.A(n_72),
.Y(n_125)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_73),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_74),
.Y(n_178)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

INVx5_ASAP7_75t_L g188 ( 
.A(n_75),
.Y(n_188)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_36),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g132 ( 
.A(n_76),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_77),
.Y(n_184)
);

INVx4_ASAP7_75t_SL g78 ( 
.A(n_44),
.Y(n_78)
);

INVx13_ASAP7_75t_L g169 ( 
.A(n_78),
.Y(n_169)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_79),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_36),
.Y(n_80)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_80),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_81),
.Y(n_196)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

INVx2_ASAP7_75t_SL g126 ( 
.A(n_82),
.Y(n_126)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_83),
.Y(n_146)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_26),
.Y(n_84)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_84),
.Y(n_139)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_26),
.Y(n_85)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_85),
.Y(n_147)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_21),
.Y(n_86)
);

INVx11_ASAP7_75t_L g137 ( 
.A(n_86),
.Y(n_137)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_26),
.Y(n_87)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_87),
.Y(n_155)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_88),
.Y(n_200)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_20),
.Y(n_89)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_89),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_23),
.Y(n_90)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_90),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_22),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_91),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_23),
.Y(n_92)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_92),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_19),
.B(n_8),
.Y(n_93)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_28),
.Y(n_94)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_94),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_38),
.Y(n_95)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_95),
.Y(n_173)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_22),
.Y(n_96)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_96),
.Y(n_171)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_25),
.Y(n_97)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_97),
.Y(n_133)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_21),
.Y(n_98)
);

BUFx10_ASAP7_75t_L g191 ( 
.A(n_98),
.Y(n_191)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_29),
.Y(n_99)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_99),
.Y(n_182)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_21),
.Y(n_100)
);

BUFx2_ASAP7_75t_SL g159 ( 
.A(n_100),
.Y(n_159)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_20),
.Y(n_101)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_101),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_38),
.Y(n_102)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_102),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_55),
.B(n_29),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_103),
.B(n_116),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_38),
.Y(n_104)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_104),
.Y(n_179)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_20),
.Y(n_105)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_105),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_45),
.Y(n_106)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_106),
.Y(n_181)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_45),
.Y(n_107)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_107),
.Y(n_186)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_20),
.Y(n_108)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_108),
.Y(n_199)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_28),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_109),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_45),
.Y(n_110)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_110),
.Y(n_195)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_20),
.Y(n_111)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_111),
.Y(n_203)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_25),
.Y(n_112)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_112),
.Y(n_149)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_24),
.Y(n_113)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_113),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_49),
.Y(n_114)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_114),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_49),
.Y(n_115)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_115),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_49),
.Y(n_116)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_35),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_117),
.B(n_118),
.Y(n_142)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_24),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g119 ( 
.A(n_44),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_119),
.B(n_42),
.Y(n_136)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_24),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_120),
.B(n_121),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_35),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_24),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_122),
.B(n_123),
.Y(n_193)
);

BUFx5_ASAP7_75t_L g123 ( 
.A(n_44),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_63),
.A2(n_47),
.B1(n_35),
.B2(n_24),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_135),
.A2(n_144),
.B1(n_157),
.B2(n_174),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_136),
.Y(n_210)
);

A2O1A1Ixp33_ASAP7_75t_L g141 ( 
.A1(n_103),
.A2(n_55),
.B(n_53),
.C(n_34),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_141),
.B(n_156),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_63),
.B(n_48),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_143),
.B(n_165),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_65),
.A2(n_47),
.B1(n_54),
.B2(n_51),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_91),
.B(n_32),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_90),
.A2(n_47),
.B1(n_32),
.B2(n_54),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_75),
.B(n_43),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_109),
.B(n_59),
.C(n_34),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_167),
.B(n_172),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_83),
.B(n_51),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_75),
.A2(n_42),
.B1(n_53),
.B2(n_59),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_117),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_176),
.B(n_187),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_66),
.A2(n_42),
.B1(n_41),
.B2(n_27),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_180),
.A2(n_57),
.B1(n_102),
.B2(n_95),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_107),
.B(n_48),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_183),
.B(n_189),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_83),
.A2(n_57),
.B(n_30),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_68),
.B(n_43),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_78),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_190),
.B(n_7),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_80),
.B(n_40),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_194),
.B(n_197),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_76),
.B(n_40),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_88),
.B(n_30),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_198),
.B(n_201),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_121),
.B(n_27),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_119),
.B(n_42),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_202),
.B(n_204),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_119),
.B(n_42),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_166),
.Y(n_205)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_205),
.Y(n_286)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_185),
.Y(n_206)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_206),
.Y(n_295)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_133),
.Y(n_208)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_208),
.Y(n_294)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_149),
.Y(n_209)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_209),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_142),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_211),
.B(n_242),
.Y(n_281)
);

BUFx6f_ASAP7_75t_SL g212 ( 
.A(n_191),
.Y(n_212)
);

BUFx24_ASAP7_75t_L g323 ( 
.A(n_212),
.Y(n_323)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_127),
.Y(n_214)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_214),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_193),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_215),
.B(n_272),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_193),
.Y(n_216)
);

CKINVDCx14_ASAP7_75t_R g300 ( 
.A(n_216),
.Y(n_300)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_130),
.Y(n_217)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_217),
.Y(n_318)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_129),
.Y(n_218)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_218),
.Y(n_301)
);

OAI21xp33_ASAP7_75t_L g220 ( 
.A1(n_138),
.A2(n_9),
.B(n_18),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_220),
.B(n_239),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_L g221 ( 
.A1(n_138),
.A2(n_60),
.B1(n_62),
.B2(n_64),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_221),
.A2(n_254),
.B1(n_168),
.B2(n_195),
.Y(n_290)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_188),
.Y(n_224)
);

BUFx2_ASAP7_75t_L g314 ( 
.A(n_224),
.Y(n_314)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_192),
.Y(n_225)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_225),
.Y(n_320)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_188),
.Y(n_227)
);

INVx4_ASAP7_75t_L g285 ( 
.A(n_227),
.Y(n_285)
);

AO22x1_ASAP7_75t_SL g228 ( 
.A1(n_141),
.A2(n_41),
.B1(n_74),
.B2(n_77),
.Y(n_228)
);

AOI22x1_ASAP7_75t_L g308 ( 
.A1(n_228),
.A2(n_164),
.B1(n_162),
.B2(n_160),
.Y(n_308)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_151),
.Y(n_229)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_229),
.Y(n_291)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_199),
.Y(n_230)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_230),
.Y(n_322)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_131),
.Y(n_231)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_231),
.Y(n_331)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_151),
.Y(n_233)
);

INVx5_ASAP7_75t_L g284 ( 
.A(n_233),
.Y(n_284)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_134),
.Y(n_234)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_234),
.Y(n_332)
);

INVx8_ASAP7_75t_L g236 ( 
.A(n_200),
.Y(n_236)
);

INVx5_ASAP7_75t_L g317 ( 
.A(n_236),
.Y(n_317)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_186),
.Y(n_238)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_238),
.Y(n_329)
);

INVx4_ASAP7_75t_SL g239 ( 
.A(n_169),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_135),
.A2(n_116),
.B1(n_115),
.B2(n_114),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_240),
.A2(n_257),
.B1(n_274),
.B2(n_164),
.Y(n_296)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_203),
.Y(n_241)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_241),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_140),
.B(n_0),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_139),
.B(n_147),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_243),
.B(n_245),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_132),
.A2(n_81),
.B1(n_106),
.B2(n_104),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_244),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_142),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_155),
.Y(n_246)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_246),
.Y(n_334)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_124),
.Y(n_247)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_247),
.Y(n_339)
);

INVx4_ASAP7_75t_L g248 ( 
.A(n_200),
.Y(n_248)
);

INVx6_ASAP7_75t_L g313 ( 
.A(n_248),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_249),
.A2(n_152),
.B1(n_159),
.B2(n_13),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_174),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_250),
.B(n_262),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_145),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_251),
.Y(n_293)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_177),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g327 ( 
.A(n_252),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_145),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_253),
.Y(n_328)
);

AOI22xp33_ASAP7_75t_L g254 ( 
.A1(n_161),
.A2(n_110),
.B1(n_92),
.B2(n_52),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_171),
.B(n_10),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_255),
.B(n_258),
.Y(n_303)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_186),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_256),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_180),
.A2(n_52),
.B1(n_37),
.B2(n_7),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_124),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_182),
.B(n_7),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_259),
.B(n_265),
.Y(n_319)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_158),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_260),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_163),
.B(n_0),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_261),
.B(n_273),
.C(n_278),
.Y(n_289)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_170),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_132),
.A2(n_125),
.B1(n_128),
.B2(n_150),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_263),
.A2(n_264),
.B1(n_276),
.B2(n_146),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_125),
.A2(n_52),
.B1(n_37),
.B2(n_12),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_163),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_126),
.B(n_170),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_266),
.B(n_267),
.Y(n_325)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_153),
.Y(n_267)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_153),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_268),
.B(n_269),
.Y(n_287)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_173),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_270),
.B(n_271),
.Y(n_324)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_173),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_175),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_126),
.B(n_1),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_162),
.A2(n_37),
.B1(n_12),
.B2(n_13),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_175),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_275),
.B(n_277),
.Y(n_342)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_177),
.Y(n_276)
);

INVx4_ASAP7_75t_L g277 ( 
.A(n_154),
.Y(n_277)
);

AND2x2_ASAP7_75t_SL g278 ( 
.A(n_128),
.B(n_146),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_169),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_279),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_280),
.Y(n_379)
);

AOI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_250),
.A2(n_154),
.B1(n_168),
.B2(n_179),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_SL g343 ( 
.A1(n_288),
.A2(n_335),
.B1(n_252),
.B2(n_224),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_290),
.B(n_278),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_296),
.A2(n_311),
.B1(n_316),
.B2(n_326),
.Y(n_344)
);

OR2x2_ASAP7_75t_L g298 ( 
.A(n_207),
.B(n_181),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_298),
.B(n_261),
.Y(n_351)
);

MAJx2_ASAP7_75t_L g302 ( 
.A(n_242),
.B(n_191),
.C(n_137),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_302),
.B(n_307),
.C(n_3),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_237),
.A2(n_191),
.B(n_137),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g359 ( 
.A1(n_305),
.A2(n_333),
.B(n_309),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_235),
.B(n_195),
.Y(n_307)
);

OA21x2_ASAP7_75t_L g378 ( 
.A1(n_308),
.A2(n_212),
.B(n_2),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_228),
.A2(n_148),
.B1(n_184),
.B2(n_178),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_310),
.A2(n_321),
.B1(n_278),
.B2(n_251),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_222),
.A2(n_181),
.B1(n_179),
.B2(n_160),
.Y(n_311)
);

XNOR2x2_ASAP7_75t_L g315 ( 
.A(n_226),
.B(n_37),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_315),
.B(n_258),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_240),
.A2(n_196),
.B1(n_184),
.B2(n_178),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_228),
.A2(n_196),
.B1(n_152),
.B2(n_148),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_L g330 ( 
.A1(n_216),
.A2(n_5),
.B1(n_14),
.B2(n_13),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g367 ( 
.A1(n_330),
.A2(n_233),
.B1(n_229),
.B2(n_247),
.Y(n_367)
);

AOI32xp33_ASAP7_75t_L g333 ( 
.A1(n_219),
.A2(n_5),
.A3(n_14),
.B1(n_13),
.B2(n_18),
.Y(n_333)
);

AOI22xp33_ASAP7_75t_SL g335 ( 
.A1(n_236),
.A2(n_268),
.B1(n_267),
.B2(n_248),
.Y(n_335)
);

BUFx24_ASAP7_75t_SL g336 ( 
.A(n_213),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_336),
.B(n_1),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_232),
.A2(n_1),
.B(n_2),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_L g363 ( 
.A1(n_340),
.A2(n_276),
.B(n_241),
.Y(n_363)
);

AOI21xp33_ASAP7_75t_L g341 ( 
.A1(n_223),
.A2(n_14),
.B(n_2),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_SL g358 ( 
.A(n_341),
.B(n_1),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_L g414 ( 
.A1(n_343),
.A2(n_363),
.B(n_291),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_SL g345 ( 
.A(n_307),
.B(n_281),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_345),
.B(n_390),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_303),
.B(n_210),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_346),
.B(n_349),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_347),
.A2(n_352),
.B1(n_354),
.B2(n_356),
.Y(n_394)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_325),
.Y(n_348)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_348),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_306),
.B(n_261),
.Y(n_349)
);

CKINVDCx14_ASAP7_75t_R g425 ( 
.A(n_350),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_SL g417 ( 
.A1(n_351),
.A2(n_377),
.B(n_327),
.Y(n_417)
);

AOI22xp33_ASAP7_75t_L g352 ( 
.A1(n_321),
.A2(n_205),
.B1(n_206),
.B2(n_273),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_286),
.Y(n_353)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_353),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_308),
.A2(n_220),
.B1(n_273),
.B2(n_256),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_286),
.Y(n_355)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_355),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_308),
.A2(n_299),
.B1(n_292),
.B2(n_311),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_296),
.A2(n_218),
.B1(n_214),
.B2(n_238),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_357),
.A2(n_369),
.B1(n_378),
.B2(n_385),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_358),
.B(n_359),
.Y(n_416)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_295),
.Y(n_360)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_360),
.Y(n_401)
);

MAJx2_ASAP7_75t_L g407 ( 
.A(n_361),
.B(n_388),
.C(n_329),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_319),
.B(n_287),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_362),
.B(n_366),
.Y(n_413)
);

BUFx3_ASAP7_75t_L g364 ( 
.A(n_314),
.Y(n_364)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_364),
.Y(n_429)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_295),
.Y(n_365)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_365),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_298),
.B(n_230),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_367),
.B(n_381),
.Y(n_424)
);

INVx1_ASAP7_75t_SL g368 ( 
.A(n_314),
.Y(n_368)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_368),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_316),
.A2(n_253),
.B1(n_225),
.B2(n_271),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_299),
.A2(n_272),
.B1(n_270),
.B2(n_277),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_370),
.A2(n_284),
.B1(n_291),
.B2(n_317),
.Y(n_420)
);

INVx4_ASAP7_75t_L g371 ( 
.A(n_337),
.Y(n_371)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_371),
.Y(n_411)
);

INVx4_ASAP7_75t_SL g372 ( 
.A(n_337),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_372),
.Y(n_393)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_324),
.Y(n_373)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_373),
.Y(n_421)
);

INVx3_ASAP7_75t_L g374 ( 
.A(n_313),
.Y(n_374)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_374),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_340),
.B(n_227),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_375),
.B(n_376),
.Y(n_431)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_297),
.Y(n_376)
);

HAxp5_ASAP7_75t_SL g377 ( 
.A(n_315),
.B(n_239),
.CON(n_377),
.SN(n_377)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_329),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_380),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_342),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_382),
.B(n_383),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_293),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_339),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_384),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_289),
.A2(n_305),
.B1(n_326),
.B2(n_282),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_289),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_386),
.A2(n_317),
.B1(n_285),
.B2(n_284),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_323),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_387),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_302),
.B(n_4),
.C(n_283),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_389),
.B(n_309),
.C(n_334),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_309),
.B(n_4),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_294),
.B(n_4),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_391),
.Y(n_435)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_297),
.Y(n_392)
);

AND2x2_ASAP7_75t_SL g415 ( 
.A(n_392),
.B(n_338),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g438 ( 
.A(n_400),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_345),
.B(n_300),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_405),
.B(n_407),
.C(n_409),
.Y(n_440)
);

AOI32xp33_ASAP7_75t_L g406 ( 
.A1(n_377),
.A2(n_304),
.A3(n_312),
.B1(n_318),
.B2(n_332),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_SL g466 ( 
.A1(n_406),
.A2(n_412),
.B(n_417),
.Y(n_466)
);

O2A1O1Ixp33_ASAP7_75t_L g408 ( 
.A1(n_350),
.A2(n_304),
.B(n_331),
.C(n_323),
.Y(n_408)
);

O2A1O1Ixp33_ASAP7_75t_L g473 ( 
.A1(n_408),
.A2(n_412),
.B(n_417),
.C(n_434),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_388),
.B(n_301),
.C(n_322),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_356),
.A2(n_354),
.B1(n_347),
.B2(n_348),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_410),
.A2(n_420),
.B1(n_430),
.B2(n_378),
.Y(n_441)
);

AO22x1_ASAP7_75t_L g412 ( 
.A1(n_363),
.A2(n_339),
.B1(n_338),
.B2(n_322),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_L g453 ( 
.A1(n_414),
.A2(n_418),
.B(n_426),
.Y(n_453)
);

INVx1_ASAP7_75t_SL g461 ( 
.A(n_415),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_SL g418 ( 
.A1(n_389),
.A2(n_301),
.B(n_320),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_422),
.B(n_357),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_L g423 ( 
.A1(n_385),
.A2(n_375),
.B(n_359),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_L g458 ( 
.A1(n_423),
.A2(n_368),
.B(n_384),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_SL g426 ( 
.A1(n_366),
.A2(n_320),
.B(n_285),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_L g430 ( 
.A1(n_346),
.A2(n_313),
.B1(n_328),
.B2(n_293),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_361),
.B(n_328),
.C(n_323),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_433),
.B(n_370),
.C(n_379),
.Y(n_444)
);

AOI22x1_ASAP7_75t_L g436 ( 
.A1(n_410),
.A2(n_344),
.B1(n_378),
.B2(n_350),
.Y(n_436)
);

OAI22xp33_ASAP7_75t_SL g505 ( 
.A1(n_436),
.A2(n_411),
.B1(n_429),
.B2(n_461),
.Y(n_505)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_398),
.Y(n_437)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_437),
.Y(n_475)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_398),
.Y(n_439)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_439),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_L g485 ( 
.A1(n_441),
.A2(n_451),
.B1(n_393),
.B2(n_396),
.Y(n_485)
);

OAI32xp33_ASAP7_75t_L g442 ( 
.A1(n_425),
.A2(n_349),
.A3(n_373),
.B1(n_390),
.B2(n_358),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_442),
.B(n_447),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_435),
.B(n_382),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_443),
.B(n_448),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_444),
.B(n_470),
.C(n_401),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_445),
.B(n_459),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_SL g446 ( 
.A(n_435),
.B(n_386),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_SL g480 ( 
.A(n_446),
.B(n_463),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_415),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_421),
.B(n_392),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_415),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_449),
.B(n_456),
.Y(n_487)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_399),
.Y(n_450)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_450),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_394),
.A2(n_379),
.B1(n_374),
.B2(n_371),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_395),
.B(n_413),
.Y(n_452)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_452),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_397),
.A2(n_383),
.B1(n_376),
.B2(n_355),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_454),
.A2(n_465),
.B1(n_472),
.B2(n_408),
.Y(n_477)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_399),
.Y(n_455)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_455),
.Y(n_493)
);

A2O1A1Ixp33_ASAP7_75t_L g456 ( 
.A1(n_403),
.A2(n_365),
.B(n_353),
.C(n_360),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_401),
.Y(n_457)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_457),
.Y(n_499)
);

OAI21xp5_ASAP7_75t_SL g488 ( 
.A1(n_458),
.A2(n_393),
.B(n_409),
.Y(n_488)
);

OAI21xp5_ASAP7_75t_L g459 ( 
.A1(n_423),
.A2(n_387),
.B(n_364),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_395),
.B(n_372),
.Y(n_460)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_460),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_421),
.B(n_372),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_462),
.B(n_464),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_SL g463 ( 
.A(n_413),
.B(n_4),
.Y(n_463)
);

CKINVDCx16_ASAP7_75t_R g464 ( 
.A(n_415),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_L g465 ( 
.A1(n_397),
.A2(n_403),
.B1(n_414),
.B2(n_406),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_428),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_467),
.B(n_469),
.Y(n_490)
);

CKINVDCx16_ASAP7_75t_R g468 ( 
.A(n_424),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_468),
.B(n_427),
.Y(n_500)
);

INVx1_ASAP7_75t_SL g469 ( 
.A(n_404),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_419),
.B(n_405),
.C(n_407),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_431),
.B(n_426),
.Y(n_471)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_471),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_L g472 ( 
.A1(n_431),
.A2(n_394),
.B1(n_422),
.B2(n_416),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_473),
.B(n_396),
.Y(n_489)
);

INVxp33_ASAP7_75t_SL g474 ( 
.A(n_433),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_474),
.B(n_432),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_L g516 ( 
.A1(n_477),
.A2(n_481),
.B1(n_464),
.B2(n_453),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_440),
.B(n_419),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_478),
.B(n_491),
.Y(n_523)
);

AOI22x1_ASAP7_75t_SL g481 ( 
.A1(n_465),
.A2(n_412),
.B1(n_407),
.B2(n_418),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_472),
.A2(n_430),
.B1(n_420),
.B2(n_434),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_SL g511 ( 
.A1(n_482),
.A2(n_451),
.B1(n_471),
.B2(n_453),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_SL g515 ( 
.A1(n_485),
.A2(n_497),
.B1(n_505),
.B2(n_489),
.Y(n_515)
);

AOI21xp5_ASAP7_75t_L g527 ( 
.A1(n_488),
.A2(n_496),
.B(n_458),
.Y(n_527)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_489),
.Y(n_510)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_440),
.B(n_400),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_494),
.B(n_438),
.C(n_444),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_SL g495 ( 
.A(n_470),
.B(n_402),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g538 ( 
.A(n_495),
.B(n_498),
.Y(n_538)
);

NAND2x1p5_ASAP7_75t_L g496 ( 
.A(n_466),
.B(n_402),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_441),
.A2(n_432),
.B1(n_411),
.B2(n_427),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_SL g498 ( 
.A(n_452),
.B(n_404),
.Y(n_498)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_500),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_501),
.B(n_503),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_448),
.Y(n_503)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_460),
.Y(n_507)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_507),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_467),
.Y(n_508)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_508),
.Y(n_537)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_462),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_509),
.B(n_463),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_L g550 ( 
.A1(n_511),
.A2(n_516),
.B1(n_521),
.B2(n_486),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_483),
.B(n_456),
.Y(n_513)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_513),
.Y(n_543)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_490),
.Y(n_514)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_514),
.Y(n_564)
);

OAI22xp5_ASAP7_75t_SL g542 ( 
.A1(n_515),
.A2(n_484),
.B1(n_487),
.B2(n_502),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_517),
.B(n_529),
.C(n_536),
.Y(n_547)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_490),
.Y(n_518)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_518),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_483),
.B(n_456),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_519),
.B(n_522),
.Y(n_544)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_479),
.Y(n_520)
);

INVx1_ASAP7_75t_SL g549 ( 
.A(n_520),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_SL g521 ( 
.A1(n_477),
.A2(n_504),
.B1(n_482),
.B2(n_484),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_502),
.B(n_443),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g524 ( 
.A(n_494),
.B(n_466),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g540 ( 
.A(n_524),
.B(n_532),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_508),
.B(n_446),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_525),
.B(n_526),
.Y(n_545)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_479),
.Y(n_526)
);

O2A1O1Ixp33_ASAP7_75t_L g560 ( 
.A1(n_527),
.A2(n_473),
.B(n_496),
.C(n_507),
.Y(n_560)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_493),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_528),
.B(n_531),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_491),
.B(n_459),
.C(n_461),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_480),
.B(n_468),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_530),
.B(n_534),
.Y(n_552)
);

XNOR2xp5_ASAP7_75t_L g532 ( 
.A(n_495),
.B(n_436),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_L g534 ( 
.A1(n_504),
.A2(n_445),
.B1(n_449),
.B2(n_447),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_478),
.B(n_469),
.C(n_436),
.Y(n_536)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_493),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_539),
.B(n_492),
.Y(n_556)
);

XOR2xp5_ASAP7_75t_L g568 ( 
.A(n_542),
.B(n_557),
.Y(n_568)
);

OAI21xp5_ASAP7_75t_SL g546 ( 
.A1(n_527),
.A2(n_489),
.B(n_486),
.Y(n_546)
);

AOI21xp5_ASAP7_75t_L g574 ( 
.A1(n_546),
.A2(n_562),
.B(n_563),
.Y(n_574)
);

OAI22xp5_ASAP7_75t_SL g548 ( 
.A1(n_515),
.A2(n_519),
.B1(n_513),
.B2(n_514),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_548),
.B(n_526),
.Y(n_579)
);

OAI22xp5_ASAP7_75t_SL g572 ( 
.A1(n_550),
.A2(n_533),
.B1(n_539),
.B2(n_528),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_523),
.B(n_501),
.C(n_488),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_551),
.B(n_553),
.Y(n_582)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_523),
.B(n_496),
.C(n_486),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_517),
.B(n_524),
.C(n_529),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g567 ( 
.A(n_554),
.B(n_561),
.C(n_511),
.Y(n_567)
);

XNOR2xp5_ASAP7_75t_L g555 ( 
.A(n_532),
.B(n_481),
.Y(n_555)
);

XNOR2xp5_ASAP7_75t_L g566 ( 
.A(n_555),
.B(n_558),
.Y(n_566)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_556),
.Y(n_573)
);

XOR2xp5_ASAP7_75t_L g557 ( 
.A(n_538),
.B(n_506),
.Y(n_557)
);

XNOR2xp5_ASAP7_75t_L g558 ( 
.A(n_538),
.B(n_498),
.Y(n_558)
);

XNOR2xp5_ASAP7_75t_SL g559 ( 
.A(n_536),
.B(n_487),
.Y(n_559)
);

XOR2xp5_ASAP7_75t_L g569 ( 
.A(n_559),
.B(n_521),
.Y(n_569)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_560),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g561 ( 
.A(n_512),
.B(n_497),
.C(n_454),
.Y(n_561)
);

AOI21xp5_ASAP7_75t_L g562 ( 
.A1(n_510),
.A2(n_473),
.B(n_499),
.Y(n_562)
);

AOI21xp5_ASAP7_75t_L g563 ( 
.A1(n_510),
.A2(n_522),
.B(n_518),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_567),
.B(n_585),
.Y(n_597)
);

XNOR2xp5_ASAP7_75t_L g598 ( 
.A(n_569),
.B(n_570),
.Y(n_598)
);

XOR2xp5_ASAP7_75t_L g570 ( 
.A(n_540),
.B(n_535),
.Y(n_570)
);

XNOR2xp5_ASAP7_75t_L g571 ( 
.A(n_551),
.B(n_554),
.Y(n_571)
);

XNOR2xp5_ASAP7_75t_L g599 ( 
.A(n_571),
.B(n_584),
.Y(n_599)
);

XOR2xp5_ASAP7_75t_L g591 ( 
.A(n_572),
.B(n_586),
.Y(n_591)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_541),
.Y(n_576)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_576),
.Y(n_588)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_541),
.Y(n_577)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_577),
.Y(n_589)
);

CKINVDCx20_ASAP7_75t_R g578 ( 
.A(n_544),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_SL g590 ( 
.A(n_578),
.B(n_580),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_579),
.B(n_581),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_552),
.B(n_537),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_545),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_549),
.B(n_520),
.Y(n_583)
);

CKINVDCx14_ASAP7_75t_R g602 ( 
.A(n_583),
.Y(n_602)
);

XNOR2xp5_ASAP7_75t_L g584 ( 
.A(n_547),
.B(n_559),
.Y(n_584)
);

MAJIxp5_ASAP7_75t_L g585 ( 
.A(n_547),
.B(n_537),
.C(n_499),
.Y(n_585)
);

XOR2xp5_ASAP7_75t_L g586 ( 
.A(n_540),
.B(n_442),
.Y(n_586)
);

AND2x2_ASAP7_75t_L g587 ( 
.A(n_574),
.B(n_563),
.Y(n_587)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_587),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_571),
.B(n_561),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_592),
.B(n_593),
.Y(n_617)
);

MAJIxp5_ASAP7_75t_L g593 ( 
.A(n_567),
.B(n_550),
.C(n_553),
.Y(n_593)
);

NOR2x1_ASAP7_75t_L g594 ( 
.A(n_575),
.B(n_543),
.Y(n_594)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_594),
.Y(n_612)
);

MAJIxp5_ASAP7_75t_L g595 ( 
.A(n_584),
.B(n_557),
.C(n_546),
.Y(n_595)
);

AOI21xp5_ASAP7_75t_L g611 ( 
.A1(n_595),
.A2(n_600),
.B(n_601),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_585),
.B(n_542),
.Y(n_596)
);

CKINVDCx14_ASAP7_75t_R g616 ( 
.A(n_596),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_573),
.B(n_548),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_569),
.B(n_565),
.Y(n_601)
);

MAJIxp5_ASAP7_75t_L g604 ( 
.A(n_582),
.B(n_555),
.C(n_562),
.Y(n_604)
);

MAJIxp5_ASAP7_75t_L g618 ( 
.A(n_604),
.B(n_566),
.C(n_574),
.Y(n_618)
);

XNOR2xp5_ASAP7_75t_L g605 ( 
.A(n_593),
.B(n_570),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_605),
.B(n_610),
.Y(n_623)
);

AOI22xp5_ASAP7_75t_L g607 ( 
.A1(n_602),
.A2(n_572),
.B1(n_564),
.B2(n_579),
.Y(n_607)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_607),
.Y(n_628)
);

XOR2xp5_ASAP7_75t_L g608 ( 
.A(n_598),
.B(n_568),
.Y(n_608)
);

XNOR2xp5_ASAP7_75t_L g627 ( 
.A(n_608),
.B(n_609),
.Y(n_627)
);

XOR2xp5_ASAP7_75t_L g609 ( 
.A(n_598),
.B(n_568),
.Y(n_609)
);

AOI22xp5_ASAP7_75t_L g610 ( 
.A1(n_588),
.A2(n_586),
.B1(n_549),
.B2(n_560),
.Y(n_610)
);

XNOR2xp5_ASAP7_75t_L g613 ( 
.A(n_604),
.B(n_599),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_613),
.B(n_618),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_590),
.B(n_583),
.Y(n_614)
);

OAI21x1_ASAP7_75t_L g620 ( 
.A1(n_614),
.A2(n_615),
.B(n_603),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_599),
.B(n_566),
.Y(n_615)
);

OAI21xp5_ASAP7_75t_L g619 ( 
.A1(n_611),
.A2(n_616),
.B(n_617),
.Y(n_619)
);

AOI21xp5_ASAP7_75t_L g630 ( 
.A1(n_619),
.A2(n_622),
.B(n_625),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_620),
.B(n_621),
.Y(n_635)
);

MAJIxp5_ASAP7_75t_L g621 ( 
.A(n_605),
.B(n_597),
.C(n_595),
.Y(n_621)
);

MAJIxp5_ASAP7_75t_L g622 ( 
.A(n_613),
.B(n_591),
.C(n_587),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_612),
.B(n_606),
.Y(n_625)
);

MAJIxp5_ASAP7_75t_L g626 ( 
.A(n_618),
.B(n_591),
.C(n_587),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_626),
.B(n_608),
.Y(n_633)
);

AOI21xp33_ASAP7_75t_SL g629 ( 
.A1(n_621),
.A2(n_594),
.B(n_610),
.Y(n_629)
);

AO21x1_ASAP7_75t_L g639 ( 
.A1(n_629),
.A2(n_631),
.B(n_634),
.Y(n_639)
);

OAI21xp5_ASAP7_75t_L g631 ( 
.A1(n_624),
.A2(n_603),
.B(n_589),
.Y(n_631)
);

OAI21xp5_ASAP7_75t_SL g632 ( 
.A1(n_626),
.A2(n_607),
.B(n_609),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_632),
.B(n_633),
.Y(n_636)
);

OAI21xp5_ASAP7_75t_L g634 ( 
.A1(n_623),
.A2(n_476),
.B(n_475),
.Y(n_634)
);

AOI21x1_ASAP7_75t_L g637 ( 
.A1(n_630),
.A2(n_622),
.B(n_628),
.Y(n_637)
);

OA21x2_ASAP7_75t_L g640 ( 
.A1(n_637),
.A2(n_437),
.B(n_439),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_635),
.B(n_627),
.Y(n_638)
);

AOI21xp5_ASAP7_75t_L g641 ( 
.A1(n_638),
.A2(n_450),
.B(n_455),
.Y(n_641)
);

NAND2x1_ASAP7_75t_SL g642 ( 
.A(n_640),
.B(n_641),
.Y(n_642)
);

AO21x1_ASAP7_75t_L g643 ( 
.A1(n_642),
.A2(n_636),
.B(n_639),
.Y(n_643)
);

MAJx2_ASAP7_75t_L g644 ( 
.A(n_643),
.B(n_457),
.C(n_558),
.Y(n_644)
);

XNOR2xp5_ASAP7_75t_L g645 ( 
.A(n_644),
.B(n_429),
.Y(n_645)
);


endmodule