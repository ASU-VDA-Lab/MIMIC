module fake_jpeg_16184_n_300 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_300);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_300;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_152;
wire n_73;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_288;
wire n_272;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_118;
wire n_82;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx6f_ASAP7_75t_SL g36 ( 
.A(n_7),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_4),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_15),
.B(n_39),
.Y(n_40)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_40),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

INVx2_ASAP7_75t_R g43 ( 
.A(n_36),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_43),
.B(n_27),
.Y(n_94)
);

INVx6_ASAP7_75t_SL g44 ( 
.A(n_35),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_44),
.B(n_48),
.Y(n_73)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_15),
.B(n_6),
.Y(n_46)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_46),
.Y(n_107)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

INVx11_ASAP7_75t_L g102 ( 
.A(n_47),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_25),
.B(n_39),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_25),
.B(n_6),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_50),
.B(n_52),
.Y(n_80)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_51),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_26),
.B(n_5),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

CKINVDCx6p67_ASAP7_75t_R g85 ( 
.A(n_54),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_26),
.B(n_5),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_55),
.B(n_56),
.Y(n_90)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

BUFx24_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_58),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_61),
.B(n_62),
.Y(n_93)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_64),
.B(n_34),
.Y(n_101)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_66),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_67),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_52),
.B(n_38),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_70),
.B(n_72),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_61),
.A2(n_23),
.B1(n_31),
.B2(n_30),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_71),
.A2(n_86),
.B1(n_88),
.B2(n_92),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_49),
.B(n_38),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_57),
.B(n_28),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_74),
.B(n_75),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_66),
.B(n_28),
.Y(n_75)
);

AOI21xp33_ASAP7_75t_L g81 ( 
.A1(n_43),
.A2(n_30),
.B(n_32),
.Y(n_81)
);

AOI21xp33_ASAP7_75t_L g145 ( 
.A1(n_81),
.A2(n_111),
.B(n_83),
.Y(n_145)
);

AND2x4_ASAP7_75t_L g83 ( 
.A(n_43),
.B(n_0),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_83),
.A2(n_104),
.B(n_86),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_62),
.A2(n_23),
.B1(n_31),
.B2(n_18),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_60),
.A2(n_22),
.B1(n_32),
.B2(n_18),
.Y(n_88)
);

NOR2x1_ASAP7_75t_L g89 ( 
.A(n_58),
.B(n_27),
.Y(n_89)
);

CKINVDCx14_ASAP7_75t_R g147 ( 
.A(n_89),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_63),
.A2(n_65),
.B1(n_47),
.B2(n_19),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_94),
.B(n_112),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_51),
.B(n_19),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_95),
.B(n_70),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_45),
.A2(n_22),
.B1(n_44),
.B2(n_29),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_96),
.A2(n_97),
.B1(n_110),
.B2(n_59),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_42),
.A2(n_34),
.B1(n_29),
.B2(n_17),
.Y(n_97)
);

BUFx12_ASAP7_75t_L g98 ( 
.A(n_56),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_98),
.B(n_3),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_101),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_64),
.B(n_34),
.Y(n_103)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_103),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_42),
.A2(n_29),
.B1(n_17),
.B2(n_8),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_67),
.B(n_17),
.Y(n_105)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_105),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_67),
.B(n_5),
.Y(n_108)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_108),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_42),
.A2(n_13),
.B1(n_14),
.B2(n_11),
.Y(n_110)
);

AOI21xp33_ASAP7_75t_SL g111 ( 
.A1(n_58),
.A2(n_0),
.B(n_1),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_41),
.B(n_0),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_72),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_114),
.B(n_115),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_99),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_100),
.Y(n_116)
);

BUFx2_ASAP7_75t_L g183 ( 
.A(n_116),
.Y(n_183)
);

BUFx12_ASAP7_75t_L g119 ( 
.A(n_98),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_119),
.B(n_122),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_120),
.A2(n_93),
.B(n_113),
.Y(n_158)
);

BUFx5_ASAP7_75t_L g121 ( 
.A(n_99),
.Y(n_121)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_121),
.Y(n_169)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_87),
.Y(n_122)
);

BUFx8_ASAP7_75t_L g123 ( 
.A(n_89),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_123),
.Y(n_188)
);

OAI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_83),
.A2(n_54),
.B1(n_53),
.B2(n_58),
.Y(n_124)
);

AO21x1_ASAP7_75t_L g160 ( 
.A1(n_124),
.A2(n_153),
.B(n_85),
.Y(n_160)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_100),
.Y(n_125)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_125),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_126),
.B(n_127),
.Y(n_165)
);

OAI22xp33_ASAP7_75t_L g132 ( 
.A1(n_84),
.A2(n_2),
.B1(n_4),
.B2(n_9),
.Y(n_132)
);

OAI22xp33_ASAP7_75t_L g164 ( 
.A1(n_132),
.A2(n_136),
.B1(n_140),
.B2(n_102),
.Y(n_164)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_68),
.Y(n_133)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_133),
.Y(n_175)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_68),
.Y(n_134)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_134),
.Y(n_181)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_69),
.Y(n_135)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_135),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_77),
.A2(n_91),
.B1(n_83),
.B2(n_69),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_80),
.B(n_4),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_137),
.B(n_141),
.Y(n_168)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_76),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_139),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_77),
.A2(n_9),
.B1(n_13),
.B2(n_14),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_74),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_107),
.B(n_2),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_143),
.B(n_147),
.Y(n_184)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_76),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_144),
.B(n_146),
.Y(n_172)
);

A2O1A1Ixp33_ASAP7_75t_L g174 ( 
.A1(n_145),
.A2(n_87),
.B(n_102),
.C(n_118),
.Y(n_174)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_75),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_84),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_148),
.B(n_149),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_106),
.B(n_2),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_79),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_150),
.B(n_151),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_104),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_152),
.A2(n_85),
.B(n_82),
.Y(n_173)
);

OA22x2_ASAP7_75t_L g153 ( 
.A1(n_91),
.A2(n_109),
.B1(n_94),
.B2(n_85),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_78),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_154),
.B(n_125),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_129),
.B(n_112),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_156),
.B(n_167),
.C(n_170),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_131),
.B(n_118),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_157),
.B(n_161),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_158),
.A2(n_173),
.B(n_185),
.Y(n_209)
);

OR2x2_ASAP7_75t_L g213 ( 
.A(n_160),
.B(n_176),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_131),
.B(n_90),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_131),
.B(n_78),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_163),
.B(n_176),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_164),
.B(n_171),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_152),
.B(n_73),
.C(n_79),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_118),
.B(n_98),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_130),
.B(n_82),
.C(n_85),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_171),
.B(n_177),
.C(n_121),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_174),
.B(n_117),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_153),
.B(n_123),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_142),
.B(n_151),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_180),
.B(n_122),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_184),
.B(n_186),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_153),
.B(n_132),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_138),
.B(n_128),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_153),
.B(n_123),
.Y(n_187)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_187),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_190),
.B(n_205),
.Y(n_224)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_166),
.Y(n_191)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_191),
.Y(n_227)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_166),
.Y(n_192)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_192),
.Y(n_235)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_175),
.Y(n_194)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_194),
.Y(n_237)
);

AOI322xp5_ASAP7_75t_SL g195 ( 
.A1(n_184),
.A2(n_117),
.A3(n_119),
.B1(n_133),
.B2(n_135),
.C1(n_134),
.C2(n_144),
.Y(n_195)
);

NOR3xp33_ASAP7_75t_L g230 ( 
.A(n_195),
.B(n_188),
.C(n_158),
.Y(n_230)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_175),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_197),
.B(n_198),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_183),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_181),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_199),
.B(n_201),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_183),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_181),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_202),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_203),
.B(n_204),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_155),
.B(n_115),
.Y(n_204)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_182),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_206),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_185),
.A2(n_119),
.B1(n_139),
.B2(n_177),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_208),
.A2(n_211),
.B1(n_185),
.B2(n_167),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_172),
.B(n_178),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_210),
.B(n_212),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_183),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_213),
.A2(n_216),
.B(n_157),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_182),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_214),
.B(n_215),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_169),
.B(n_159),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_163),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_209),
.A2(n_173),
.B(n_187),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_217),
.A2(n_213),
.B(n_193),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_218),
.A2(n_219),
.B(n_191),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_211),
.A2(n_189),
.B1(n_216),
.B2(n_207),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_220),
.A2(n_222),
.B1(n_232),
.B2(n_189),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_196),
.B(n_170),
.C(n_156),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_221),
.B(n_236),
.C(n_205),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_211),
.A2(n_160),
.B1(n_174),
.B2(n_164),
.Y(n_222)
);

OAI32xp33_ASAP7_75t_L g226 ( 
.A1(n_207),
.A2(n_161),
.A3(n_160),
.B1(n_179),
.B2(n_188),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_SL g240 ( 
.A(n_226),
.B(n_190),
.Y(n_240)
);

AOI221xp5_ASAP7_75t_L g245 ( 
.A1(n_230),
.A2(n_193),
.B1(n_214),
.B2(n_200),
.C(n_206),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_208),
.Y(n_231)
);

CKINVDCx14_ASAP7_75t_R g246 ( 
.A(n_231),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_209),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_196),
.B(n_165),
.C(n_168),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_239),
.A2(n_250),
.B1(n_256),
.B2(n_229),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_240),
.B(n_243),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_234),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_241),
.B(n_249),
.Y(n_268)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_238),
.Y(n_242)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_242),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_244),
.B(n_248),
.Y(n_262)
);

OA21x2_ASAP7_75t_SL g264 ( 
.A1(n_245),
.A2(n_249),
.B(n_241),
.Y(n_264)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_227),
.Y(n_247)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_247),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_224),
.B(n_197),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_233),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_231),
.A2(n_202),
.B1(n_199),
.B2(n_194),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_251),
.B(n_253),
.Y(n_266)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_227),
.Y(n_252)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_252),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_224),
.B(n_192),
.C(n_198),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_221),
.B(n_169),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_254),
.B(n_255),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_220),
.B(n_218),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_232),
.A2(n_201),
.B1(n_212),
.B2(n_162),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_260),
.A2(n_261),
.B1(n_243),
.B2(n_237),
.Y(n_275)
);

OAI321xp33_ASAP7_75t_L g261 ( 
.A1(n_240),
.A2(n_226),
.A3(n_217),
.B1(n_219),
.B2(n_222),
.C(n_223),
.Y(n_261)
);

FAx1_ASAP7_75t_L g263 ( 
.A(n_244),
.B(n_250),
.CI(n_255),
.CON(n_263),
.SN(n_263)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_263),
.A2(n_237),
.B(n_235),
.Y(n_278)
);

AOI31xp67_ASAP7_75t_L g270 ( 
.A1(n_264),
.A2(n_246),
.A3(n_236),
.B(n_225),
.Y(n_270)
);

INVx1_ASAP7_75t_SL g265 ( 
.A(n_256),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_265),
.B(n_228),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_270),
.B(n_275),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_268),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_271),
.B(n_276),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_266),
.B(n_253),
.C(n_254),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_272),
.B(n_273),
.C(n_279),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_266),
.B(n_248),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_274),
.A2(n_257),
.B1(n_265),
.B2(n_259),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_260),
.B(n_162),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_268),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_277),
.B(n_280),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_278),
.A2(n_263),
.B1(n_258),
.B2(n_262),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_267),
.B(n_235),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_259),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_278),
.B(n_262),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_281),
.A2(n_285),
.B(n_273),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_287),
.B(n_162),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_271),
.A2(n_263),
.B1(n_267),
.B2(n_269),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_288),
.B(n_279),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_289),
.B(n_290),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_284),
.B(n_272),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_291),
.B(n_292),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_281),
.A2(n_287),
.B1(n_288),
.B2(n_285),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_293),
.B(n_282),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_296),
.B(n_292),
.C(n_283),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_294),
.A2(n_286),
.B(n_283),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_297),
.B(n_298),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_295),
.Y(n_300)
);


endmodule