module fake_jpeg_15696_n_350 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_350);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_350;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_37),
.Y(n_76)
);

BUFx4f_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_20),
.B(n_8),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_48),
.B(n_16),
.Y(n_66)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_24),
.Y(n_49)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_44),
.A2(n_34),
.B1(n_30),
.B2(n_18),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_51),
.A2(n_57),
.B1(n_61),
.B2(n_62),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_17),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_52),
.B(n_53),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_17),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_50),
.B(n_33),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_55),
.B(n_33),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_44),
.A2(n_20),
.B1(n_31),
.B2(n_23),
.Y(n_57)
);

INVx4_ASAP7_75t_SL g59 ( 
.A(n_38),
.Y(n_59)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_59),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_40),
.A2(n_23),
.B1(n_22),
.B2(n_21),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_40),
.A2(n_28),
.B1(n_27),
.B2(n_22),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_42),
.A2(n_31),
.B1(n_28),
.B2(n_27),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_65),
.A2(n_73),
.B1(n_49),
.B2(n_12),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_66),
.B(n_25),
.Y(n_96)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_69),
.Y(n_104)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_49),
.A2(n_38),
.B1(n_13),
.B2(n_2),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_74),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_79),
.B(n_83),
.Y(n_134)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_81),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_55),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_84),
.B(n_96),
.Y(n_143)
);

CKINVDCx6p67_ASAP7_75t_R g85 ( 
.A(n_72),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g133 ( 
.A(n_85),
.Y(n_133)
);

HB1xp67_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

BUFx2_ASAP7_75t_L g136 ( 
.A(n_86),
.Y(n_136)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_87),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_88),
.Y(n_122)
);

OA22x2_ASAP7_75t_L g89 ( 
.A1(n_54),
.A2(n_38),
.B1(n_49),
.B2(n_36),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_89),
.A2(n_103),
.B1(n_112),
.B2(n_64),
.Y(n_124)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_90),
.B(n_94),
.Y(n_135)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_92),
.Y(n_119)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_68),
.Y(n_93)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_93),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_52),
.B(n_48),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_68),
.Y(n_95)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_95),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_53),
.B(n_25),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_100),
.Y(n_116)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_76),
.Y(n_98)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_98),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_SL g99 ( 
.A(n_65),
.B(n_25),
.C(n_33),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_SL g127 ( 
.A(n_99),
.B(n_110),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_60),
.B(n_75),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_57),
.B(n_25),
.Y(n_101)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_101),
.Y(n_137)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_58),
.Y(n_102)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_102),
.Y(n_125)
);

BUFx12_ASAP7_75t_L g105 ( 
.A(n_63),
.Y(n_105)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_105),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_59),
.A2(n_12),
.B1(n_15),
.B2(n_2),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_106),
.A2(n_11),
.B1(n_15),
.B2(n_3),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_74),
.B(n_47),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_107),
.A2(n_67),
.B(n_26),
.Y(n_141)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_59),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_108),
.Y(n_120)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_75),
.Y(n_109)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_109),
.Y(n_138)
);

AOI32xp33_ASAP7_75t_L g110 ( 
.A1(n_56),
.A2(n_47),
.A3(n_37),
.B1(n_39),
.B2(n_43),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_72),
.B(n_39),
.C(n_37),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_111),
.A2(n_77),
.B1(n_70),
.B2(n_64),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_69),
.A2(n_71),
.B1(n_77),
.B2(n_70),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_63),
.Y(n_113)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_113),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_67),
.B(n_16),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_114),
.Y(n_140)
);

INVx13_ASAP7_75t_L g115 ( 
.A(n_105),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_115),
.B(n_105),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_118),
.A2(n_142),
.B1(n_85),
.B2(n_9),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_124),
.A2(n_132),
.B1(n_102),
.B2(n_104),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_128),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_80),
.B(n_33),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_130),
.B(n_107),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_82),
.A2(n_43),
.B1(n_36),
.B2(n_67),
.Y(n_132)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_88),
.Y(n_139)
);

INVxp33_ASAP7_75t_L g164 ( 
.A(n_139),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_141),
.A2(n_145),
.B(n_10),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_80),
.A2(n_97),
.B1(n_84),
.B2(n_99),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_92),
.A2(n_9),
.B1(n_15),
.B2(n_3),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_126),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_146),
.B(n_160),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_124),
.A2(n_132),
.B1(n_116),
.B2(n_127),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_147),
.A2(n_173),
.B1(n_174),
.B2(n_125),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_148),
.B(n_151),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_116),
.B(n_100),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_149),
.B(n_151),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_150),
.A2(n_163),
.B1(n_172),
.B2(n_139),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_130),
.B(n_98),
.Y(n_151)
);

AOI21xp33_ASAP7_75t_L g152 ( 
.A1(n_142),
.A2(n_91),
.B(n_104),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_152),
.A2(n_154),
.B(n_157),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_143),
.B(n_79),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_153),
.B(n_156),
.Y(n_200)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_117),
.Y(n_155)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_155),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_143),
.B(n_109),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_137),
.A2(n_127),
.B(n_143),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_117),
.Y(n_158)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_158),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_141),
.B(n_111),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_159),
.B(n_168),
.C(n_136),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_126),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_129),
.Y(n_161)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_161),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_137),
.A2(n_91),
.B(n_78),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_162),
.A2(n_167),
.B(n_138),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_134),
.A2(n_87),
.B1(n_95),
.B2(n_93),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_R g210 ( 
.A(n_165),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_135),
.B(n_89),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_166),
.B(n_175),
.Y(n_204)
);

XOR2x2_ASAP7_75t_L g167 ( 
.A(n_118),
.B(n_89),
.Y(n_167)
);

MAJx2_ASAP7_75t_L g168 ( 
.A(n_140),
.B(n_89),
.C(n_81),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_122),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_169),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_129),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_170),
.B(n_136),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_119),
.A2(n_113),
.B1(n_85),
.B2(n_26),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_119),
.A2(n_85),
.B1(n_8),
.B2(n_3),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_140),
.B(n_0),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_131),
.Y(n_176)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_176),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_120),
.B(n_0),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_177),
.B(n_179),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_120),
.A2(n_125),
.B1(n_121),
.B2(n_123),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_178),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_121),
.B(n_10),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_182),
.B(n_162),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_184),
.A2(n_1),
.B1(n_206),
.B2(n_205),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_167),
.A2(n_131),
.B1(n_138),
.B2(n_123),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_186),
.A2(n_189),
.B1(n_201),
.B2(n_174),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_188),
.A2(n_209),
.B(n_213),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_190),
.B(n_173),
.Y(n_215)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_191),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_159),
.B(n_167),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_192),
.A2(n_7),
.B(n_4),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_L g193 ( 
.A1(n_150),
.A2(n_136),
.B1(n_133),
.B2(n_115),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_193),
.A2(n_174),
.B1(n_158),
.B2(n_160),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_159),
.B(n_157),
.C(n_156),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_195),
.B(n_199),
.C(n_205),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_155),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_197),
.B(n_164),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_149),
.B(n_0),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_198),
.B(n_211),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_153),
.B(n_147),
.C(n_148),
.Y(n_199)
);

OAI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_168),
.A2(n_133),
.B1(n_122),
.B2(n_144),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_161),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_203),
.B(n_208),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_152),
.B(n_122),
.C(n_133),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_173),
.A2(n_144),
.B1(n_1),
.B2(n_0),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_206),
.A2(n_6),
.B1(n_11),
.B2(n_13),
.Y(n_236)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_176),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_154),
.A2(n_26),
.B(n_16),
.Y(n_209)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_178),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_166),
.A2(n_7),
.B(n_13),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_177),
.B(n_0),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_214),
.B(n_1),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_215),
.B(n_222),
.C(n_226),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_210),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_216),
.B(n_232),
.Y(n_250)
);

O2A1O1Ixp33_ASAP7_75t_L g217 ( 
.A1(n_183),
.A2(n_171),
.B(n_168),
.C(n_170),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_217),
.A2(n_230),
.B(n_209),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_219),
.B(n_204),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_220),
.A2(n_229),
.B1(n_210),
.B2(n_200),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_195),
.B(n_162),
.C(n_178),
.Y(n_222)
);

INVxp67_ASAP7_75t_SL g248 ( 
.A(n_224),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_211),
.A2(n_175),
.B1(n_146),
.B2(n_179),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_225),
.A2(n_212),
.B1(n_193),
.B2(n_203),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_190),
.B(n_163),
.Y(n_226)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_227),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_189),
.A2(n_165),
.B1(n_172),
.B2(n_169),
.Y(n_229)
);

OAI21x1_ASAP7_75t_SL g230 ( 
.A1(n_188),
.A2(n_169),
.B(n_4),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_192),
.B(n_14),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_231),
.B(n_212),
.C(n_214),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_191),
.Y(n_232)
);

XNOR2x1_ASAP7_75t_L g233 ( 
.A(n_192),
.B(n_7),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_233),
.B(n_234),
.Y(n_246)
);

A2O1A1O1Ixp25_ASAP7_75t_L g235 ( 
.A1(n_192),
.A2(n_10),
.B(n_4),
.C(n_5),
.D(n_6),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_235),
.B(n_213),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_236),
.A2(n_237),
.B1(n_243),
.B2(n_198),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_184),
.A2(n_6),
.B1(n_11),
.B2(n_14),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_238),
.B(n_242),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_182),
.B(n_6),
.Y(n_239)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_239),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_197),
.B(n_11),
.Y(n_240)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_240),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_196),
.B(n_14),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_247),
.A2(n_252),
.B1(n_241),
.B2(n_233),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_228),
.Y(n_249)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_249),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_220),
.A2(n_199),
.B1(n_196),
.B2(n_200),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_251),
.A2(n_262),
.B1(n_243),
.B2(n_223),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_215),
.B(n_185),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_253),
.B(n_239),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_221),
.B(n_185),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_254),
.B(n_265),
.C(n_266),
.Y(n_271)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_255),
.Y(n_275)
);

AO21x1_ASAP7_75t_L g274 ( 
.A1(n_256),
.A2(n_257),
.B(n_219),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_218),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_260),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_229),
.A2(n_186),
.B1(n_204),
.B2(n_201),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_263),
.B(n_264),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_221),
.B(n_180),
.C(n_194),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_226),
.B(n_181),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_232),
.B(n_216),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_267),
.B(n_218),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_222),
.B(n_180),
.C(n_194),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_268),
.B(n_234),
.C(n_241),
.Y(n_281)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_270),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_274),
.B(n_285),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_266),
.B(n_231),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_276),
.B(n_283),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_277),
.B(n_279),
.Y(n_304)
);

AOI21xp33_ASAP7_75t_L g278 ( 
.A1(n_257),
.A2(n_230),
.B(n_223),
.Y(n_278)
);

CKINVDCx14_ASAP7_75t_R g291 ( 
.A(n_278),
.Y(n_291)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_244),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_280),
.A2(n_245),
.B1(n_253),
.B2(n_263),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_281),
.B(n_284),
.C(n_286),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_247),
.A2(n_217),
.B1(n_237),
.B2(n_224),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_282),
.A2(n_287),
.B1(n_289),
.B2(n_269),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_268),
.B(n_225),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_259),
.B(n_242),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_250),
.A2(n_181),
.B(n_235),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_285),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_250),
.A2(n_202),
.B(n_207),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_265),
.B(n_202),
.C(n_207),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_288),
.B(n_258),
.C(n_246),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_262),
.A2(n_208),
.B1(n_236),
.B2(n_187),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_SL g290 ( 
.A(n_283),
.B(n_254),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_290),
.B(n_295),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_284),
.B(n_259),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_292),
.B(n_300),
.C(n_302),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_SL g295 ( 
.A(n_281),
.B(n_251),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_275),
.A2(n_267),
.B1(n_248),
.B2(n_264),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_298),
.A2(n_287),
.B1(n_282),
.B2(n_277),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_299),
.B(n_286),
.Y(n_314)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_270),
.Y(n_301)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_301),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_273),
.B(n_246),
.Y(n_302)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_303),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_273),
.B(n_252),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_305),
.B(n_271),
.C(n_288),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g311 ( 
.A(n_306),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_304),
.B(n_272),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_309),
.B(n_316),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_310),
.B(n_320),
.Y(n_323)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_313),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_314),
.B(n_305),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_291),
.A2(n_271),
.B1(n_289),
.B2(n_274),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_315),
.A2(n_295),
.B1(n_290),
.B2(n_296),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g316 ( 
.A(n_294),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_300),
.B(n_276),
.C(n_258),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_317),
.B(n_292),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_298),
.B(n_261),
.Y(n_319)
);

OR2x2_ASAP7_75t_L g326 ( 
.A(n_319),
.B(n_293),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_302),
.B(n_238),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_321),
.B(n_328),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_322),
.B(n_307),
.C(n_317),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_315),
.A2(n_297),
.B(n_296),
.Y(n_324)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_324),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_313),
.B(n_187),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_325),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_326),
.B(n_327),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_312),
.B(n_293),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_332),
.B(n_323),
.C(n_310),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_326),
.B(n_319),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g342 ( 
.A1(n_333),
.A2(n_329),
.B(n_321),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_330),
.B(n_311),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_334),
.B(n_320),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_338),
.B(n_339),
.C(n_342),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_337),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_340),
.A2(n_341),
.B(n_336),
.Y(n_343)
);

OR2x2_ASAP7_75t_L g341 ( 
.A(n_331),
.B(n_308),
.Y(n_341)
);

OA21x2_ASAP7_75t_SL g345 ( 
.A1(n_343),
.A2(n_341),
.B(n_332),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_345),
.B(n_344),
.C(n_335),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_346),
.B(n_335),
.C(n_323),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_347),
.A2(n_307),
.B1(n_328),
.B2(n_314),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_SL g349 ( 
.A(n_348),
.B(n_318),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_349),
.B(n_318),
.Y(n_350)
);


endmodule