module real_jpeg_87_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_83;
wire n_78;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_93;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_92;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_85;
wire n_89;
wire n_16;

INVx2_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_1),
.B(n_31),
.Y(n_65)
);

AND2x2_ASAP7_75t_SL g91 ( 
.A(n_1),
.B(n_26),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_3),
.B(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_3),
.B(n_26),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_3),
.B(n_23),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_4),
.B(n_23),
.Y(n_22)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_4),
.B(n_19),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_4),
.B(n_56),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_5),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_6),
.B(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_6),
.B(n_31),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_6),
.B(n_23),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_6),
.B(n_19),
.Y(n_76)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_8),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_9),
.B(n_19),
.Y(n_18)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_9),
.B(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_9),
.B(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_10),
.B(n_31),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_68),
.Y(n_12)
);

OAI21xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_50),
.B(n_67),
.Y(n_13)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_38),
.B(n_49),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_33),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_16),
.B(n_33),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_24),
.Y(n_16)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_22),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_18),
.B(n_22),
.C(n_24),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_29),
.B1(n_30),
.B2(n_32),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_25),
.Y(n_32)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_29),
.B(n_32),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

INVx3_ASAP7_75t_SL g41 ( 
.A(n_31),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_36),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_34),
.B(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_34),
.A2(n_36),
.B1(n_37),
.B2(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_43),
.B(n_48),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_42),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_42),
.B(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_46),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_46),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_52),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_52),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_58),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_59),
.C(n_62),
.Y(n_71)
);

BUFx24_ASAP7_75t_SL g95 ( 
.A(n_53),
.Y(n_95)
);

FAx1_ASAP7_75t_SL g53 ( 
.A(n_54),
.B(n_55),
.CI(n_57),
.CON(n_53),
.SN(n_53)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_54),
.B(n_55),
.C(n_57),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_61),
.B2(n_62),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_63),
.A2(n_64),
.B1(n_65),
.B2(n_66),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_63),
.B(n_66),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_65),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_94),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_72),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_71),
.B(n_72),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_85),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_75),
.B1(n_83),
.B2(n_84),
.Y(n_73)
);

CKINVDCx14_ASAP7_75t_R g83 ( 
.A(n_74),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_75),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_77),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_79),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_SL g85 ( 
.A(n_86),
.B(n_87),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_89),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_91),
.B1(n_92),
.B2(n_93),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);


endmodule