module fake_netlist_5_89_n_2021 (n_137, n_168, n_164, n_191, n_91, n_82, n_122, n_194, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_188, n_190, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_196, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_2021);

input n_137;
input n_168;
input n_164;
input n_191;
input n_91;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_188;
input n_190;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_196;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_2021;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_1960;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_447;
wire n_247;
wire n_2001;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_2011;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_1949;
wire n_343;
wire n_1449;
wire n_308;
wire n_1946;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_1948;
wire n_1984;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1097;
wire n_1036;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_798;
wire n_350;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_1931;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_845;
wire n_663;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1986;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1971;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1891;
wire n_1662;
wire n_1481;
wire n_1942;
wire n_434;
wire n_1978;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_2009;
wire n_759;
wire n_1892;
wire n_806;
wire n_1997;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1963;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_526;
wire n_1916;
wire n_293;
wire n_677;
wire n_372;
wire n_244;
wire n_1333;
wire n_1121;
wire n_433;
wire n_314;
wire n_368;
wire n_604;
wire n_2007;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_1851;
wire n_758;
wire n_999;
wire n_1933;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_1874;
wire n_563;
wire n_1987;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_1989;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_2017;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1980;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_239;
wire n_630;
wire n_1902;
wire n_1941;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_2015;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1958;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_968;
wire n_315;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_1974;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1966;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1992;
wire n_1643;
wire n_883;
wire n_1983;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1400;
wire n_1342;
wire n_900;
wire n_856;
wire n_1793;
wire n_1976;
wire n_918;
wire n_942;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_2020;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1928;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_584;
wire n_681;
wire n_336;
wire n_1638;
wire n_1786;
wire n_430;
wire n_2002;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_1998;
wire n_304;
wire n_1338;
wire n_577;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1834;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_1968;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_421;
wire n_1988;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_2003;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_2008;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_2012;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_1999;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1985;
wire n_1898;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1944;
wire n_909;
wire n_1817;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_1981;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_2006;
wire n_1995;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_2014;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1962;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_685;
wire n_598;
wire n_608;
wire n_928;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_1975;
wire n_273;
wire n_1937;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_1936;
wire n_1956;
wire n_437;
wire n_1642;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1969;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_2013;
wire n_1990;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVx2_ASAP7_75t_L g199 ( 
.A(n_127),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_149),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_159),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_171),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_77),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_59),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_0),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_67),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_119),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_22),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_26),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_170),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_40),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_72),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_24),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_160),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_95),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_130),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_5),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_190),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_8),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_74),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_23),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_50),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_107),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_121),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_94),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_184),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_173),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_86),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_78),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_133),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_150),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_108),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_176),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_104),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_32),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_112),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_66),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_16),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_83),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_106),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_137),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_196),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_118),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_63),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_186),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_148),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_100),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_59),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_28),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_102),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_188),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_145),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_156),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_143),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_73),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_111),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_62),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_82),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_42),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_34),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_164),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_7),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_15),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_194),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_116),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_122),
.Y(n_266)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_44),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_61),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_54),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_75),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_198),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_17),
.Y(n_272)
);

CKINVDCx14_ASAP7_75t_R g273 ( 
.A(n_183),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_36),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_67),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_28),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_45),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_44),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_117),
.Y(n_279)
);

BUFx3_ASAP7_75t_L g280 ( 
.A(n_157),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_53),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_192),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_110),
.Y(n_283)
);

BUFx10_ASAP7_75t_L g284 ( 
.A(n_90),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_3),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_161),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_152),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_162),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_53),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_15),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_129),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_166),
.Y(n_292)
);

INVx2_ASAP7_75t_SL g293 ( 
.A(n_6),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_30),
.Y(n_294)
);

BUFx10_ASAP7_75t_L g295 ( 
.A(n_8),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_84),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_54),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_88),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_39),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_43),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_101),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_1),
.Y(n_302)
);

INVx1_ASAP7_75t_SL g303 ( 
.A(n_5),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_115),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_41),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_132),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_41),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_38),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_92),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_140),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_12),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_165),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_12),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_21),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_70),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_182),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_178),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_189),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_18),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_76),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_174),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_33),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_197),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_179),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_6),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_4),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_9),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_34),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_42),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_138),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_57),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_168),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_80),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_158),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_185),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_195),
.Y(n_336)
);

BUFx3_ASAP7_75t_L g337 ( 
.A(n_20),
.Y(n_337)
);

INVx1_ASAP7_75t_SL g338 ( 
.A(n_172),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_144),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_45),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_19),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_142),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_66),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_3),
.Y(n_344)
);

BUFx8_ASAP7_75t_SL g345 ( 
.A(n_11),
.Y(n_345)
);

INVx1_ASAP7_75t_SL g346 ( 
.A(n_98),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_81),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_191),
.Y(n_348)
);

BUFx3_ASAP7_75t_L g349 ( 
.A(n_131),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_99),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_69),
.Y(n_351)
);

HB1xp67_ASAP7_75t_L g352 ( 
.A(n_43),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_93),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_146),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_23),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_68),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_51),
.Y(n_357)
);

BUFx5_ASAP7_75t_L g358 ( 
.A(n_11),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_29),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_62),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_105),
.Y(n_361)
);

BUFx10_ASAP7_75t_L g362 ( 
.A(n_21),
.Y(n_362)
);

INVxp67_ASAP7_75t_SL g363 ( 
.A(n_135),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_60),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_40),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_39),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_153),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_17),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_147),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_36),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_50),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_123),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_167),
.Y(n_373)
);

BUFx3_ASAP7_75t_L g374 ( 
.A(n_1),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_32),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_154),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_57),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_103),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_58),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_134),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_33),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_48),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_51),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_65),
.Y(n_384)
);

BUFx10_ASAP7_75t_L g385 ( 
.A(n_0),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_85),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_14),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_125),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_18),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_46),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_61),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_2),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_10),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_120),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_65),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_109),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_212),
.Y(n_397)
);

INVxp67_ASAP7_75t_SL g398 ( 
.A(n_210),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_358),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_358),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_358),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_358),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_345),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_358),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_202),
.B(n_2),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_206),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_358),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_358),
.Y(n_408)
);

NOR2xp67_ASAP7_75t_L g409 ( 
.A(n_260),
.B(n_4),
.Y(n_409)
);

INVx1_ASAP7_75t_SL g410 ( 
.A(n_325),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_242),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_358),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_202),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_209),
.Y(n_414)
);

NOR2xp67_ASAP7_75t_L g415 ( 
.A(n_352),
.B(n_7),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_216),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_216),
.Y(n_417)
);

CKINVDCx16_ASAP7_75t_R g418 ( 
.A(n_312),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_218),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_213),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_258),
.Y(n_421)
);

HB1xp67_ASAP7_75t_L g422 ( 
.A(n_219),
.Y(n_422)
);

INVxp33_ASAP7_75t_L g423 ( 
.A(n_204),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_259),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_259),
.Y(n_425)
);

CKINVDCx14_ASAP7_75t_R g426 ( 
.A(n_273),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_237),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_286),
.Y(n_428)
);

CKINVDCx16_ASAP7_75t_R g429 ( 
.A(n_295),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_373),
.Y(n_430)
);

BUFx10_ASAP7_75t_L g431 ( 
.A(n_293),
.Y(n_431)
);

CKINVDCx16_ASAP7_75t_R g432 ( 
.A(n_295),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_244),
.Y(n_433)
);

INVx1_ASAP7_75t_SL g434 ( 
.A(n_327),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_248),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_249),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_200),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_257),
.Y(n_438)
);

BUFx6f_ASAP7_75t_SL g439 ( 
.A(n_284),
.Y(n_439)
);

OR2x2_ASAP7_75t_L g440 ( 
.A(n_204),
.B(n_9),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_201),
.Y(n_441)
);

INVxp67_ASAP7_75t_SL g442 ( 
.A(n_210),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_203),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_218),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_223),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_214),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_223),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_215),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_224),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_224),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_262),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_227),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_227),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_269),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_228),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_272),
.Y(n_456)
);

INVxp67_ASAP7_75t_SL g457 ( 
.A(n_241),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_276),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_220),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_228),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_229),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_229),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_232),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_277),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_232),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_233),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_225),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_281),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_285),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_233),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_289),
.Y(n_471)
);

HB1xp67_ASAP7_75t_L g472 ( 
.A(n_290),
.Y(n_472)
);

INVxp67_ASAP7_75t_SL g473 ( 
.A(n_241),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_199),
.B(n_10),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_294),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_234),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_234),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_300),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_243),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_226),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_243),
.B(n_13),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_302),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_308),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_231),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_355),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_311),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_245),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_245),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_313),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_239),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_250),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_319),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_199),
.B(n_13),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_328),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_331),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_250),
.B(n_14),
.Y(n_496)
);

CKINVDCx14_ASAP7_75t_R g497 ( 
.A(n_295),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_240),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_254),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_399),
.Y(n_500)
);

OR2x6_ASAP7_75t_L g501 ( 
.A(n_415),
.B(n_280),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g502 ( 
.A(n_398),
.B(n_280),
.Y(n_502)
);

OAI21x1_ASAP7_75t_L g503 ( 
.A1(n_400),
.A2(n_230),
.B(n_207),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_400),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_401),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_442),
.B(n_349),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_457),
.B(n_349),
.Y(n_507)
);

HB1xp67_ASAP7_75t_L g508 ( 
.A(n_422),
.Y(n_508)
);

AOI22x1_ASAP7_75t_SL g509 ( 
.A1(n_397),
.A2(n_329),
.B1(n_364),
.B2(n_222),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_402),
.Y(n_510)
);

BUFx2_ASAP7_75t_L g511 ( 
.A(n_406),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_404),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_407),
.Y(n_513)
);

AND2x4_ASAP7_75t_L g514 ( 
.A(n_408),
.B(n_207),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_412),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_473),
.B(n_396),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_424),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_424),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_425),
.Y(n_519)
);

OR2x6_ASAP7_75t_L g520 ( 
.A(n_474),
.B(n_293),
.Y(n_520)
);

AND2x4_ASAP7_75t_L g521 ( 
.A(n_413),
.B(n_416),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_425),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_406),
.B(n_338),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_485),
.Y(n_524)
);

INVx2_ASAP7_75t_SL g525 ( 
.A(n_431),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_417),
.B(n_267),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_485),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_419),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_444),
.Y(n_529)
);

INVx4_ASAP7_75t_L g530 ( 
.A(n_440),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_445),
.B(n_267),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_447),
.Y(n_532)
);

HB1xp67_ASAP7_75t_L g533 ( 
.A(n_414),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_449),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_450),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_414),
.B(n_346),
.Y(n_536)
);

NAND2xp33_ASAP7_75t_SL g537 ( 
.A(n_439),
.B(n_340),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_452),
.B(n_246),
.Y(n_538)
);

XNOR2xp5_ASAP7_75t_L g539 ( 
.A(n_410),
.B(n_217),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_453),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_455),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_460),
.Y(n_542)
);

HB1xp67_ASAP7_75t_L g543 ( 
.A(n_420),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_461),
.B(n_247),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_462),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_463),
.B(n_499),
.Y(n_546)
);

BUFx3_ASAP7_75t_L g547 ( 
.A(n_465),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_466),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_470),
.B(n_476),
.Y(n_549)
);

INVx2_ASAP7_75t_SL g550 ( 
.A(n_431),
.Y(n_550)
);

AND2x4_ASAP7_75t_L g551 ( 
.A(n_477),
.B(n_230),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_479),
.Y(n_552)
);

OA22x2_ASAP7_75t_SL g553 ( 
.A1(n_487),
.A2(n_208),
.B1(n_211),
.B2(n_205),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_488),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_491),
.Y(n_555)
);

AND2x6_ASAP7_75t_L g556 ( 
.A(n_405),
.B(n_347),
.Y(n_556)
);

BUFx6f_ASAP7_75t_L g557 ( 
.A(n_493),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_440),
.Y(n_558)
);

INVx4_ASAP7_75t_L g559 ( 
.A(n_439),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_481),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_496),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_431),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_420),
.B(n_254),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_409),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_423),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_426),
.B(n_251),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_472),
.Y(n_567)
);

BUFx6f_ASAP7_75t_L g568 ( 
.A(n_427),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_427),
.Y(n_569)
);

BUFx6f_ASAP7_75t_L g570 ( 
.A(n_433),
.Y(n_570)
);

BUFx6f_ASAP7_75t_L g571 ( 
.A(n_433),
.Y(n_571)
);

HB1xp67_ASAP7_75t_L g572 ( 
.A(n_435),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_497),
.B(n_274),
.Y(n_573)
);

AND2x4_ASAP7_75t_L g574 ( 
.A(n_435),
.B(n_236),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_436),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_436),
.B(n_274),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_438),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_438),
.B(n_252),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_451),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_557),
.B(n_451),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_502),
.B(n_454),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_512),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_546),
.Y(n_583)
);

AND2x6_ASAP7_75t_L g584 ( 
.A(n_557),
.B(n_236),
.Y(n_584)
);

NAND3xp33_ASAP7_75t_L g585 ( 
.A(n_560),
.B(n_456),
.C(n_454),
.Y(n_585)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_502),
.B(n_456),
.Y(n_586)
);

INVx4_ASAP7_75t_L g587 ( 
.A(n_504),
.Y(n_587)
);

INVx2_ASAP7_75t_SL g588 ( 
.A(n_565),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_512),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_546),
.Y(n_590)
);

INVx3_ASAP7_75t_L g591 ( 
.A(n_504),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_546),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_500),
.Y(n_593)
);

AO21x2_ASAP7_75t_L g594 ( 
.A1(n_503),
.A2(n_264),
.B(n_261),
.Y(n_594)
);

INVx4_ASAP7_75t_L g595 ( 
.A(n_504),
.Y(n_595)
);

INVx8_ASAP7_75t_L g596 ( 
.A(n_568),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_502),
.B(n_458),
.Y(n_597)
);

INVx3_ASAP7_75t_L g598 ( 
.A(n_504),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_512),
.Y(n_599)
);

BUFx2_ASAP7_75t_L g600 ( 
.A(n_565),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_517),
.Y(n_601)
);

INVx4_ASAP7_75t_L g602 ( 
.A(n_504),
.Y(n_602)
);

BUFx3_ASAP7_75t_L g603 ( 
.A(n_547),
.Y(n_603)
);

AND2x6_ASAP7_75t_L g604 ( 
.A(n_557),
.B(n_282),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_523),
.B(n_418),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_500),
.Y(n_606)
);

AOI22xp33_ASAP7_75t_L g607 ( 
.A1(n_560),
.A2(n_355),
.B1(n_374),
.B2(n_337),
.Y(n_607)
);

INVx4_ASAP7_75t_L g608 ( 
.A(n_504),
.Y(n_608)
);

BUFx10_ASAP7_75t_L g609 ( 
.A(n_536),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_505),
.Y(n_610)
);

INVx4_ASAP7_75t_L g611 ( 
.A(n_504),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_517),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_517),
.Y(n_613)
);

BUFx3_ASAP7_75t_L g614 ( 
.A(n_547),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_578),
.B(n_437),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_505),
.Y(n_616)
);

INVx4_ASAP7_75t_L g617 ( 
.A(n_557),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_525),
.B(n_429),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_510),
.Y(n_619)
);

INVx2_ASAP7_75t_SL g620 ( 
.A(n_576),
.Y(n_620)
);

INVx3_ASAP7_75t_L g621 ( 
.A(n_517),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_557),
.B(n_458),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_557),
.B(n_464),
.Y(n_623)
);

OAI22xp5_ASAP7_75t_L g624 ( 
.A1(n_561),
.A2(n_498),
.B1(n_441),
.B2(n_443),
.Y(n_624)
);

NOR2x1p5_ASAP7_75t_L g625 ( 
.A(n_559),
.B(n_403),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_557),
.B(n_464),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_549),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_549),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_516),
.B(n_468),
.Y(n_629)
);

INVx8_ASAP7_75t_L g630 ( 
.A(n_568),
.Y(n_630)
);

AND2x4_ASAP7_75t_L g631 ( 
.A(n_547),
.B(n_255),
.Y(n_631)
);

INVx3_ASAP7_75t_L g632 ( 
.A(n_517),
.Y(n_632)
);

HB1xp67_ASAP7_75t_L g633 ( 
.A(n_539),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_517),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_549),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_516),
.B(n_468),
.Y(n_636)
);

BUFx2_ASAP7_75t_L g637 ( 
.A(n_539),
.Y(n_637)
);

BUFx2_ASAP7_75t_L g638 ( 
.A(n_576),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_517),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_510),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_513),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_503),
.Y(n_642)
);

AND2x6_ASAP7_75t_L g643 ( 
.A(n_506),
.B(n_282),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_519),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_525),
.B(n_550),
.Y(n_645)
);

NAND2xp33_ASAP7_75t_L g646 ( 
.A(n_556),
.B(n_347),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_525),
.B(n_432),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_519),
.Y(n_648)
);

OR2x2_ASAP7_75t_L g649 ( 
.A(n_558),
.B(n_434),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_519),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_513),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_574),
.B(n_469),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_574),
.B(n_469),
.Y(n_653)
);

OR2x6_ASAP7_75t_L g654 ( 
.A(n_520),
.B(n_299),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_574),
.B(n_471),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_574),
.B(n_561),
.Y(n_656)
);

INVxp67_ASAP7_75t_L g657 ( 
.A(n_508),
.Y(n_657)
);

BUFx4f_ASAP7_75t_L g658 ( 
.A(n_568),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_522),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_522),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_515),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_515),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_522),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_524),
.Y(n_664)
);

CKINVDCx16_ASAP7_75t_R g665 ( 
.A(n_533),
.Y(n_665)
);

AND2x6_ASAP7_75t_L g666 ( 
.A(n_506),
.B(n_255),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_524),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_550),
.B(n_471),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_524),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_529),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_528),
.Y(n_671)
);

INVxp33_ASAP7_75t_L g672 ( 
.A(n_558),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_529),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_528),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_578),
.B(n_446),
.Y(n_675)
);

BUFx6f_ASAP7_75t_L g676 ( 
.A(n_503),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_529),
.Y(n_677)
);

BUFx6f_ASAP7_75t_L g678 ( 
.A(n_514),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_532),
.Y(n_679)
);

BUFx3_ASAP7_75t_L g680 ( 
.A(n_521),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_534),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_569),
.B(n_448),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_534),
.Y(n_683)
);

INVx4_ASAP7_75t_L g684 ( 
.A(n_514),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_SL g685 ( 
.A(n_559),
.B(n_403),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_532),
.Y(n_686)
);

INVx4_ASAP7_75t_L g687 ( 
.A(n_514),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_540),
.Y(n_688)
);

BUFx6f_ASAP7_75t_L g689 ( 
.A(n_514),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_574),
.B(n_475),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_540),
.Y(n_691)
);

OR2x2_ASAP7_75t_L g692 ( 
.A(n_558),
.B(n_475),
.Y(n_692)
);

INVxp67_ASAP7_75t_SL g693 ( 
.A(n_538),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_569),
.B(n_459),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_506),
.B(n_478),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_511),
.Y(n_696)
);

INVx2_ASAP7_75t_SL g697 ( 
.A(n_576),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_541),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_541),
.Y(n_699)
);

AOI22xp33_ASAP7_75t_L g700 ( 
.A1(n_530),
.A2(n_337),
.B1(n_299),
.B2(n_374),
.Y(n_700)
);

INVx3_ASAP7_75t_L g701 ( 
.A(n_514),
.Y(n_701)
);

INVx4_ASAP7_75t_L g702 ( 
.A(n_551),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_507),
.B(n_478),
.Y(n_703)
);

AND2x6_ASAP7_75t_L g704 ( 
.A(n_507),
.B(n_291),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_507),
.B(n_482),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_575),
.B(n_579),
.Y(n_706)
);

BUFx2_ASAP7_75t_L g707 ( 
.A(n_520),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_542),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_532),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_530),
.B(n_482),
.Y(n_710)
);

INVx1_ASAP7_75t_SL g711 ( 
.A(n_573),
.Y(n_711)
);

INVx6_ASAP7_75t_L g712 ( 
.A(n_521),
.Y(n_712)
);

OR2x6_ASAP7_75t_L g713 ( 
.A(n_520),
.B(n_205),
.Y(n_713)
);

AND2x6_ASAP7_75t_L g714 ( 
.A(n_573),
.B(n_291),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_550),
.B(n_483),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_575),
.B(n_579),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_542),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_545),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_545),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_552),
.Y(n_720)
);

AOI22xp5_ASAP7_75t_L g721 ( 
.A1(n_567),
.A2(n_480),
.B1(n_484),
.B2(n_467),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_552),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_535),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_554),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_563),
.B(n_483),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_530),
.B(n_490),
.Y(n_726)
);

OAI22xp33_ASAP7_75t_L g727 ( 
.A1(n_520),
.A2(n_303),
.B1(n_375),
.B2(n_389),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_535),
.Y(n_728)
);

INVx3_ASAP7_75t_L g729 ( 
.A(n_535),
.Y(n_729)
);

AND2x2_ASAP7_75t_L g730 ( 
.A(n_530),
.B(n_486),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_562),
.B(n_486),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_568),
.B(n_570),
.Y(n_732)
);

INVxp67_ASAP7_75t_L g733 ( 
.A(n_649),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_681),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_658),
.B(n_568),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_670),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_672),
.B(n_568),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_693),
.B(n_568),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_658),
.B(n_570),
.Y(n_739)
);

O2A1O1Ixp5_ASAP7_75t_L g740 ( 
.A1(n_701),
.A2(n_538),
.B(n_544),
.C(n_551),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_658),
.B(n_570),
.Y(n_741)
);

INVx2_ASAP7_75t_SL g742 ( 
.A(n_649),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_620),
.B(n_570),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_580),
.B(n_570),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_670),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_673),
.Y(n_746)
);

AOI21xp5_ASAP7_75t_L g747 ( 
.A1(n_622),
.A2(n_544),
.B(n_566),
.Y(n_747)
);

OAI221xp5_ASAP7_75t_L g748 ( 
.A1(n_656),
.A2(n_553),
.B1(n_520),
.B2(n_554),
.C(n_555),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_681),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_623),
.B(n_570),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_683),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_683),
.Y(n_752)
);

NOR2xp67_ASAP7_75t_L g753 ( 
.A(n_585),
.B(n_559),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_626),
.B(n_570),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_688),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_688),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_672),
.B(n_573),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_593),
.B(n_571),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_706),
.B(n_571),
.Y(n_759)
);

INVxp67_ASAP7_75t_L g760 ( 
.A(n_633),
.Y(n_760)
);

AND2x2_ASAP7_75t_L g761 ( 
.A(n_588),
.B(n_511),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_593),
.B(n_571),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_673),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_620),
.B(n_571),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_691),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_697),
.B(n_571),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_677),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_606),
.B(n_571),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_677),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_691),
.Y(n_770)
);

INVx2_ASAP7_75t_SL g771 ( 
.A(n_692),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_698),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_679),
.Y(n_773)
);

AOI22xp33_ASAP7_75t_L g774 ( 
.A1(n_666),
.A2(n_556),
.B1(n_520),
.B2(n_344),
.Y(n_774)
);

OAI22xp5_ASAP7_75t_L g775 ( 
.A1(n_695),
.A2(n_577),
.B1(n_571),
.B2(n_501),
.Y(n_775)
);

AOI22xp33_ASAP7_75t_L g776 ( 
.A1(n_666),
.A2(n_556),
.B1(n_322),
.B2(n_211),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_679),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_606),
.B(n_577),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_697),
.B(n_577),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_698),
.Y(n_780)
);

OR2x6_ASAP7_75t_L g781 ( 
.A(n_713),
.B(n_577),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_610),
.B(n_577),
.Y(n_782)
);

AND2x2_ASAP7_75t_L g783 ( 
.A(n_588),
.B(n_562),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_610),
.B(n_577),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_699),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_616),
.B(n_619),
.Y(n_786)
);

INVx5_ASAP7_75t_L g787 ( 
.A(n_642),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_716),
.B(n_703),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_616),
.B(n_577),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_619),
.B(n_556),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_699),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_705),
.B(n_567),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_686),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_686),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_702),
.B(n_347),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_708),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_640),
.B(n_556),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_708),
.Y(n_798)
);

BUFx3_ASAP7_75t_L g799 ( 
.A(n_603),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_640),
.B(n_556),
.Y(n_800)
);

BUFx6f_ASAP7_75t_L g801 ( 
.A(n_680),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_717),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_629),
.B(n_508),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_702),
.B(n_347),
.Y(n_804)
);

NAND2xp33_ASAP7_75t_L g805 ( 
.A(n_596),
.B(n_556),
.Y(n_805)
);

NAND2xp33_ASAP7_75t_L g806 ( 
.A(n_596),
.B(n_556),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_717),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_702),
.B(n_347),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_641),
.B(n_651),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_718),
.Y(n_810)
);

AND2x6_ASAP7_75t_SL g811 ( 
.A(n_682),
.B(n_208),
.Y(n_811)
);

NAND3xp33_ASAP7_75t_L g812 ( 
.A(n_692),
.B(n_492),
.C(n_489),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_718),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_609),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_709),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_701),
.Y(n_816)
);

INVx2_ASAP7_75t_SL g817 ( 
.A(n_600),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_600),
.B(n_543),
.Y(n_818)
);

OR2x6_ASAP7_75t_L g819 ( 
.A(n_713),
.B(n_572),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_617),
.B(n_521),
.Y(n_820)
);

AND2x4_ASAP7_75t_L g821 ( 
.A(n_603),
.B(n_526),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_641),
.B(n_556),
.Y(n_822)
);

BUFx2_ASAP7_75t_L g823 ( 
.A(n_638),
.Y(n_823)
);

AO22x2_ASAP7_75t_L g824 ( 
.A1(n_624),
.A2(n_509),
.B1(n_553),
.B2(n_380),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_661),
.B(n_501),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_662),
.B(n_501),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_636),
.B(n_489),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_701),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_581),
.B(n_564),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_617),
.B(n_501),
.Y(n_830)
);

NOR2xp33_ASAP7_75t_L g831 ( 
.A(n_725),
.B(n_492),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_617),
.B(n_501),
.Y(n_832)
);

AOI22xp33_ASAP7_75t_L g833 ( 
.A1(n_666),
.A2(n_238),
.B1(n_344),
.B2(n_221),
.Y(n_833)
);

INVx1_ASAP7_75t_SL g834 ( 
.A(n_696),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_678),
.B(n_521),
.Y(n_835)
);

BUFx3_ASAP7_75t_L g836 ( 
.A(n_614),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_678),
.B(n_521),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_709),
.Y(n_838)
);

INVx2_ASAP7_75t_SL g839 ( 
.A(n_581),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_671),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_711),
.B(n_494),
.Y(n_841)
);

OR2x6_ASAP7_75t_L g842 ( 
.A(n_713),
.B(n_501),
.Y(n_842)
);

INVxp67_ASAP7_75t_L g843 ( 
.A(n_731),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_666),
.B(n_704),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_674),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_723),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_666),
.B(n_564),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_666),
.B(n_566),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_719),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_723),
.Y(n_850)
);

BUFx3_ASAP7_75t_L g851 ( 
.A(n_614),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_704),
.B(n_551),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_720),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_704),
.B(n_551),
.Y(n_854)
);

AOI22xp33_ASAP7_75t_L g855 ( 
.A1(n_704),
.A2(n_221),
.B1(n_326),
.B2(n_322),
.Y(n_855)
);

INVx2_ASAP7_75t_SL g856 ( 
.A(n_586),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_728),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_728),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_678),
.B(n_559),
.Y(n_859)
);

OR2x6_ASAP7_75t_L g860 ( 
.A(n_713),
.B(n_526),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_704),
.B(n_722),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_678),
.B(n_551),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_704),
.B(n_724),
.Y(n_863)
);

O2A1O1Ixp33_ASAP7_75t_L g864 ( 
.A1(n_583),
.A2(n_592),
.B(n_627),
.C(n_590),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_680),
.B(n_494),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_643),
.B(n_495),
.Y(n_866)
);

INVx2_ASAP7_75t_SL g867 ( 
.A(n_586),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_643),
.B(n_495),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_644),
.Y(n_869)
);

NAND3xp33_ASAP7_75t_L g870 ( 
.A(n_597),
.B(n_537),
.C(n_531),
.Y(n_870)
);

AND2x6_ASAP7_75t_SL g871 ( 
.A(n_694),
.B(n_235),
.Y(n_871)
);

BUFx5_ASAP7_75t_L g872 ( 
.A(n_584),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_643),
.B(n_548),
.Y(n_873)
);

INVx1_ASAP7_75t_SL g874 ( 
.A(n_696),
.Y(n_874)
);

OR2x2_ASAP7_75t_L g875 ( 
.A(n_637),
.B(n_526),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_643),
.B(n_548),
.Y(n_876)
);

NAND3xp33_ASAP7_75t_L g877 ( 
.A(n_597),
.B(n_531),
.C(n_555),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_644),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_628),
.Y(n_879)
);

AOI22xp33_ASAP7_75t_L g880 ( 
.A1(n_643),
.A2(n_305),
.B1(n_238),
.B2(n_275),
.Y(n_880)
);

AOI22xp33_ASAP7_75t_L g881 ( 
.A1(n_643),
.A2(n_278),
.B1(n_314),
.B2(n_326),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_678),
.B(n_266),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_635),
.B(n_689),
.Y(n_883)
);

AND2x4_ASAP7_75t_L g884 ( 
.A(n_631),
.B(n_531),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_689),
.B(n_548),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_648),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_712),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_L g888 ( 
.A(n_638),
.B(n_439),
.Y(n_888)
);

BUFx4f_ASAP7_75t_L g889 ( 
.A(n_714),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_689),
.B(n_296),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_609),
.Y(n_891)
);

NOR2x1p5_ASAP7_75t_L g892 ( 
.A(n_652),
.B(n_341),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_689),
.B(n_296),
.Y(n_893)
);

BUFx6f_ASAP7_75t_L g894 ( 
.A(n_642),
.Y(n_894)
);

INVx2_ASAP7_75t_SL g895 ( 
.A(n_710),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_609),
.B(n_411),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_648),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_650),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_650),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_689),
.B(n_304),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_659),
.Y(n_901)
);

NOR2xp33_ASAP7_75t_L g902 ( 
.A(n_653),
.B(n_343),
.Y(n_902)
);

AOI221xp5_ASAP7_75t_L g903 ( 
.A1(n_727),
.A2(n_235),
.B1(n_368),
.B2(n_395),
.C(n_370),
.Y(n_903)
);

INVx8_ASAP7_75t_L g904 ( 
.A(n_714),
.Y(n_904)
);

INVxp67_ASAP7_75t_L g905 ( 
.A(n_637),
.Y(n_905)
);

NOR3xp33_ASAP7_75t_L g906 ( 
.A(n_831),
.B(n_665),
.C(n_615),
.Y(n_906)
);

AOI22xp33_ASAP7_75t_L g907 ( 
.A1(n_788),
.A2(n_712),
.B1(n_714),
.B2(n_684),
.Y(n_907)
);

AOI21xp33_ASAP7_75t_L g908 ( 
.A1(n_803),
.A2(n_605),
.B(n_675),
.Y(n_908)
);

O2A1O1Ixp33_ASAP7_75t_L g909 ( 
.A1(n_788),
.A2(n_690),
.B(n_655),
.C(n_732),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_744),
.A2(n_630),
.B(n_596),
.Y(n_910)
);

NOR2xp33_ASAP7_75t_L g911 ( 
.A(n_843),
.B(n_421),
.Y(n_911)
);

BUFx2_ASAP7_75t_L g912 ( 
.A(n_823),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_831),
.B(n_428),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_759),
.B(n_730),
.Y(n_914)
);

A2O1A1Ixp33_ASAP7_75t_L g915 ( 
.A1(n_759),
.A2(n_726),
.B(n_730),
.C(n_710),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_SL g916 ( 
.A(n_761),
.B(n_721),
.Y(n_916)
);

HB1xp67_ASAP7_75t_L g917 ( 
.A(n_817),
.Y(n_917)
);

OAI21x1_ASAP7_75t_L g918 ( 
.A1(n_790),
.A2(n_800),
.B(n_797),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_750),
.A2(n_630),
.B(n_596),
.Y(n_919)
);

NOR3xp33_ASAP7_75t_L g920 ( 
.A(n_803),
.B(n_760),
.C(n_905),
.Y(n_920)
);

BUFx6f_ASAP7_75t_L g921 ( 
.A(n_801),
.Y(n_921)
);

BUFx12f_ASAP7_75t_L g922 ( 
.A(n_742),
.Y(n_922)
);

OAI21xp5_ASAP7_75t_L g923 ( 
.A1(n_740),
.A2(n_687),
.B(n_684),
.Y(n_923)
);

NOR2xp33_ASAP7_75t_L g924 ( 
.A(n_827),
.B(n_430),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_754),
.A2(n_630),
.B(n_805),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_SL g926 ( 
.A(n_895),
.B(n_707),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_827),
.B(n_657),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_818),
.B(n_668),
.Y(n_928)
);

NAND2x1p5_ASAP7_75t_L g929 ( 
.A(n_787),
.B(n_684),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_737),
.B(n_738),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_737),
.B(n_630),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_806),
.A2(n_687),
.B(n_676),
.Y(n_932)
);

AND2x4_ASAP7_75t_L g933 ( 
.A(n_799),
.B(n_707),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_757),
.B(n_714),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_736),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_787),
.A2(n_687),
.B(n_676),
.Y(n_936)
);

AOI21x1_ASAP7_75t_L g937 ( 
.A1(n_848),
.A2(n_612),
.B(n_601),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_792),
.B(n_714),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_792),
.B(n_714),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_787),
.A2(n_676),
.B(n_642),
.Y(n_940)
);

O2A1O1Ixp33_ASAP7_75t_L g941 ( 
.A1(n_864),
.A2(n_645),
.B(n_715),
.C(n_631),
.Y(n_941)
);

A2O1A1Ixp33_ASAP7_75t_L g942 ( 
.A1(n_747),
.A2(n_631),
.B(n_618),
.C(n_647),
.Y(n_942)
);

OAI21xp33_ASAP7_75t_L g943 ( 
.A1(n_841),
.A2(n_829),
.B(n_733),
.Y(n_943)
);

OAI21xp33_ASAP7_75t_L g944 ( 
.A1(n_841),
.A2(n_607),
.B(n_700),
.Y(n_944)
);

OAI22xp5_ASAP7_75t_L g945 ( 
.A1(n_889),
.A2(n_712),
.B1(n_642),
.B2(n_676),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_816),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_783),
.B(n_734),
.Y(n_947)
);

AOI33xp33_ASAP7_75t_L g948 ( 
.A1(n_903),
.A2(n_278),
.A3(n_307),
.B1(n_395),
.B2(n_392),
.B3(n_391),
.Y(n_948)
);

NAND2x1_ASAP7_75t_L g949 ( 
.A(n_894),
.B(n_801),
.Y(n_949)
);

INVx3_ASAP7_75t_L g950 ( 
.A(n_801),
.Y(n_950)
);

A2O1A1Ixp33_ASAP7_75t_L g951 ( 
.A1(n_902),
.A2(n_334),
.B(n_335),
.C(n_304),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_787),
.A2(n_676),
.B(n_642),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_820),
.A2(n_646),
.B(n_595),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_749),
.B(n_712),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_828),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_751),
.B(n_729),
.Y(n_956)
);

INVx3_ASAP7_75t_L g957 ( 
.A(n_801),
.Y(n_957)
);

BUFx6f_ASAP7_75t_L g958 ( 
.A(n_894),
.Y(n_958)
);

A2O1A1Ixp33_ASAP7_75t_L g959 ( 
.A1(n_902),
.A2(n_335),
.B(n_342),
.C(n_354),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_736),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_820),
.A2(n_646),
.B(n_595),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_885),
.A2(n_595),
.B(n_587),
.Y(n_962)
);

NOR2xp33_ASAP7_75t_L g963 ( 
.A(n_771),
.B(n_685),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_752),
.B(n_729),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_839),
.B(n_654),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_856),
.B(n_654),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_755),
.B(n_729),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_883),
.A2(n_762),
.B(n_758),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_756),
.B(n_765),
.Y(n_969)
);

AOI22xp33_ASAP7_75t_L g970 ( 
.A1(n_833),
.A2(n_604),
.B1(n_584),
.B2(n_654),
.Y(n_970)
);

INVx2_ASAP7_75t_SL g971 ( 
.A(n_875),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_770),
.B(n_591),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_772),
.B(n_591),
.Y(n_973)
);

OR2x2_ASAP7_75t_L g974 ( 
.A(n_834),
.B(n_654),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_768),
.A2(n_602),
.B(n_587),
.Y(n_975)
);

AND2x2_ASAP7_75t_L g976 ( 
.A(n_867),
.B(n_625),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_780),
.B(n_591),
.Y(n_977)
);

AOI21x1_ASAP7_75t_L g978 ( 
.A1(n_795),
.A2(n_808),
.B(n_804),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_785),
.B(n_598),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_778),
.A2(n_602),
.B(n_587),
.Y(n_980)
);

NOR2xp33_ASAP7_75t_L g981 ( 
.A(n_812),
.B(n_509),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_782),
.A2(n_608),
.B(n_602),
.Y(n_982)
);

OAI21xp33_ASAP7_75t_L g983 ( 
.A1(n_879),
.A2(n_359),
.B(n_357),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_SL g984 ( 
.A(n_884),
.B(n_253),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_784),
.A2(n_789),
.B(n_739),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_745),
.Y(n_986)
);

AOI22xp5_ASAP7_75t_L g987 ( 
.A1(n_775),
.A2(n_604),
.B1(n_584),
.B2(n_363),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_791),
.B(n_598),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_796),
.B(n_598),
.Y(n_989)
);

AOI22xp5_ASAP7_75t_L g990 ( 
.A1(n_743),
.A2(n_604),
.B1(n_584),
.B2(n_594),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_798),
.B(n_582),
.Y(n_991)
);

NAND2xp33_ASAP7_75t_L g992 ( 
.A(n_894),
.B(n_584),
.Y(n_992)
);

O2A1O1Ixp33_ASAP7_75t_L g993 ( 
.A1(n_748),
.A2(n_669),
.B(n_667),
.C(n_664),
.Y(n_993)
);

A2O1A1Ixp33_ASAP7_75t_L g994 ( 
.A1(n_877),
.A2(n_380),
.B(n_386),
.C(n_356),
.Y(n_994)
);

OAI21xp5_ASAP7_75t_L g995 ( 
.A1(n_822),
.A2(n_589),
.B(n_582),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_735),
.A2(n_611),
.B(n_608),
.Y(n_996)
);

OAI21xp5_ASAP7_75t_L g997 ( 
.A1(n_847),
.A2(n_599),
.B(n_589),
.Y(n_997)
);

OAI321xp33_ASAP7_75t_L g998 ( 
.A1(n_870),
.A2(n_314),
.A3(n_275),
.B1(n_297),
.B2(n_305),
.C(n_392),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_L g999 ( 
.A(n_874),
.B(n_608),
.Y(n_999)
);

AOI22xp5_ASAP7_75t_L g1000 ( 
.A1(n_743),
.A2(n_604),
.B1(n_584),
.B2(n_594),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_852),
.A2(n_611),
.B(n_601),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_802),
.B(n_599),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_745),
.Y(n_1003)
);

AO21x1_ASAP7_75t_L g1004 ( 
.A1(n_735),
.A2(n_310),
.B(n_309),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_854),
.A2(n_611),
.B(n_612),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_807),
.B(n_604),
.Y(n_1006)
);

OAI21xp33_ASAP7_75t_L g1007 ( 
.A1(n_888),
.A2(n_845),
.B(n_840),
.Y(n_1007)
);

NOR2xp67_ASAP7_75t_L g1008 ( 
.A(n_814),
.B(n_659),
.Y(n_1008)
);

OR2x2_ASAP7_75t_L g1009 ( 
.A(n_896),
.B(n_594),
.Y(n_1009)
);

AOI21xp33_ASAP7_75t_L g1010 ( 
.A1(n_865),
.A2(n_309),
.B(n_361),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_810),
.B(n_604),
.Y(n_1011)
);

BUFx2_ASAP7_75t_L g1012 ( 
.A(n_860),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_739),
.A2(n_639),
.B(n_634),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_741),
.A2(n_639),
.B(n_634),
.Y(n_1014)
);

AND2x2_ASAP7_75t_L g1015 ( 
.A(n_821),
.B(n_362),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_830),
.A2(n_613),
.B(n_632),
.Y(n_1016)
);

O2A1O1Ixp33_ASAP7_75t_L g1017 ( 
.A1(n_764),
.A2(n_663),
.B(n_660),
.C(n_332),
.Y(n_1017)
);

AND2x4_ASAP7_75t_L g1018 ( 
.A(n_799),
.B(n_518),
.Y(n_1018)
);

NOR2xp33_ASAP7_75t_L g1019 ( 
.A(n_891),
.B(n_360),
.Y(n_1019)
);

O2A1O1Ixp33_ASAP7_75t_L g1020 ( 
.A1(n_766),
.A2(n_779),
.B(n_786),
.C(n_809),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_SL g1021 ( 
.A(n_884),
.B(n_256),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_813),
.B(n_660),
.Y(n_1022)
);

HB1xp67_ASAP7_75t_L g1023 ( 
.A(n_821),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_766),
.B(n_663),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_832),
.A2(n_613),
.B(n_632),
.Y(n_1025)
);

NOR2xp33_ASAP7_75t_SL g1026 ( 
.A(n_888),
.B(n_284),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_741),
.A2(n_632),
.B(n_621),
.Y(n_1027)
);

NOR2xp33_ASAP7_75t_L g1028 ( 
.A(n_836),
.B(n_366),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_862),
.A2(n_621),
.B(n_270),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_862),
.A2(n_621),
.B(n_271),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_894),
.A2(n_351),
.B(n_310),
.Y(n_1031)
);

BUFx2_ASAP7_75t_L g1032 ( 
.A(n_860),
.Y(n_1032)
);

AOI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_779),
.A2(n_333),
.B1(n_279),
.B2(n_283),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_835),
.A2(n_320),
.B(n_394),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_746),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_835),
.A2(n_320),
.B(n_394),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_SL g1037 ( 
.A(n_836),
.B(n_851),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_837),
.A2(n_354),
.B(n_356),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_849),
.B(n_853),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_746),
.Y(n_1040)
);

OAI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_861),
.A2(n_334),
.B(n_323),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_837),
.A2(n_323),
.B(n_332),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_763),
.Y(n_1043)
);

INVx3_ASAP7_75t_L g1044 ( 
.A(n_887),
.Y(n_1044)
);

BUFx6f_ASAP7_75t_L g1045 ( 
.A(n_851),
.Y(n_1045)
);

BUFx8_ASAP7_75t_SL g1046 ( 
.A(n_819),
.Y(n_1046)
);

AND2x2_ASAP7_75t_L g1047 ( 
.A(n_892),
.B(n_860),
.Y(n_1047)
);

OAI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_863),
.A2(n_342),
.B(n_386),
.Y(n_1048)
);

AOI22xp5_ASAP7_75t_L g1049 ( 
.A1(n_825),
.A2(n_378),
.B1(n_353),
.B2(n_265),
.Y(n_1049)
);

NOR3xp33_ASAP7_75t_L g1050 ( 
.A(n_866),
.B(n_361),
.C(n_379),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_763),
.Y(n_1051)
);

A2O1A1Ixp33_ASAP7_75t_L g1052 ( 
.A1(n_826),
.A2(n_263),
.B(n_268),
.C(n_527),
.Y(n_1052)
);

OAI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_873),
.A2(n_527),
.B(n_518),
.Y(n_1053)
);

AOI22xp5_ASAP7_75t_L g1054 ( 
.A1(n_868),
.A2(n_350),
.B1(n_287),
.B2(n_288),
.Y(n_1054)
);

OAI21xp33_ASAP7_75t_L g1055 ( 
.A1(n_833),
.A2(n_393),
.B(n_381),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_876),
.A2(n_348),
.B(n_292),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_767),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_880),
.B(n_298),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_767),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_769),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_880),
.B(n_301),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_844),
.A2(n_889),
.B(n_893),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_881),
.B(n_306),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_881),
.B(n_315),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_855),
.B(n_316),
.Y(n_1065)
);

BUFx6f_ASAP7_75t_L g1066 ( 
.A(n_781),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_890),
.A2(n_317),
.B(n_318),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_900),
.A2(n_369),
.B(n_321),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_769),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_SL g1070 ( 
.A(n_774),
.B(n_324),
.Y(n_1070)
);

A2O1A1Ixp33_ASAP7_75t_L g1071 ( 
.A1(n_855),
.A2(n_391),
.B(n_297),
.C(n_307),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_773),
.B(n_330),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_773),
.Y(n_1073)
);

NOR2xp67_ASAP7_75t_L g1074 ( 
.A(n_753),
.B(n_336),
.Y(n_1074)
);

AOI21xp33_ASAP7_75t_L g1075 ( 
.A1(n_842),
.A2(n_390),
.B(n_382),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_SL g1076 ( 
.A(n_774),
.B(n_339),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_795),
.A2(n_388),
.B(n_367),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_SL g1078 ( 
.A(n_776),
.B(n_872),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_777),
.Y(n_1079)
);

BUFx6f_ASAP7_75t_L g1080 ( 
.A(n_781),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_777),
.B(n_372),
.Y(n_1081)
);

BUFx6f_ASAP7_75t_L g1082 ( 
.A(n_781),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_793),
.Y(n_1083)
);

INVx3_ASAP7_75t_L g1084 ( 
.A(n_794),
.Y(n_1084)
);

AND2x6_ASAP7_75t_L g1085 ( 
.A(n_869),
.B(n_387),
.Y(n_1085)
);

NOR2xp33_ASAP7_75t_SL g1086 ( 
.A(n_819),
.B(n_284),
.Y(n_1086)
);

OAI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_804),
.A2(n_376),
.B(n_384),
.Y(n_1087)
);

NOR2xp33_ASAP7_75t_L g1088 ( 
.A(n_819),
.B(n_362),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_815),
.B(n_387),
.Y(n_1089)
);

INVx2_ASAP7_75t_SL g1090 ( 
.A(n_824),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_808),
.A2(n_365),
.B(n_384),
.Y(n_1091)
);

OAI321xp33_ASAP7_75t_L g1092 ( 
.A1(n_776),
.A2(n_370),
.A3(n_383),
.B1(n_377),
.B2(n_371),
.C(n_365),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_882),
.A2(n_368),
.B(n_383),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_815),
.Y(n_1094)
);

HB1xp67_ASAP7_75t_L g1095 ( 
.A(n_842),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_838),
.B(n_371),
.Y(n_1096)
);

BUFx6f_ASAP7_75t_L g1097 ( 
.A(n_842),
.Y(n_1097)
);

CKINVDCx14_ASAP7_75t_R g1098 ( 
.A(n_912),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_SL g1099 ( 
.A(n_908),
.B(n_872),
.Y(n_1099)
);

CKINVDCx16_ASAP7_75t_R g1100 ( 
.A(n_922),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_952),
.A2(n_904),
.B(n_859),
.Y(n_1101)
);

BUFx4f_ASAP7_75t_L g1102 ( 
.A(n_1066),
.Y(n_1102)
);

INVx1_ASAP7_75t_SL g1103 ( 
.A(n_928),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_914),
.B(n_838),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_930),
.B(n_846),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_1046),
.Y(n_1106)
);

AND2x2_ASAP7_75t_L g1107 ( 
.A(n_927),
.B(n_824),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_1057),
.Y(n_1108)
);

AOI22xp5_ASAP7_75t_L g1109 ( 
.A1(n_924),
.A2(n_824),
.B1(n_859),
.B2(n_882),
.Y(n_1109)
);

AND2x2_ASAP7_75t_L g1110 ( 
.A(n_971),
.B(n_362),
.Y(n_1110)
);

O2A1O1Ixp33_ASAP7_75t_L g1111 ( 
.A1(n_915),
.A2(n_377),
.B(n_858),
.C(n_857),
.Y(n_1111)
);

NOR2xp33_ASAP7_75t_L g1112 ( 
.A(n_913),
.B(n_811),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_1084),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_947),
.B(n_846),
.Y(n_1114)
);

NOR3xp33_ASAP7_75t_L g1115 ( 
.A(n_911),
.B(n_871),
.C(n_858),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_969),
.B(n_850),
.Y(n_1116)
);

INVx6_ASAP7_75t_L g1117 ( 
.A(n_1045),
.Y(n_1117)
);

AOI22xp5_ASAP7_75t_L g1118 ( 
.A1(n_906),
.A2(n_904),
.B1(n_850),
.B2(n_857),
.Y(n_1118)
);

NOR2xp33_ASAP7_75t_L g1119 ( 
.A(n_943),
.B(n_886),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_944),
.B(n_897),
.Y(n_1120)
);

NOR3xp33_ASAP7_75t_SL g1121 ( 
.A(n_981),
.B(n_385),
.C(n_19),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_1039),
.B(n_897),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_952),
.A2(n_904),
.B(n_901),
.Y(n_1123)
);

NAND2x1p5_ASAP7_75t_L g1124 ( 
.A(n_1066),
.B(n_901),
.Y(n_1124)
);

INVx3_ASAP7_75t_L g1125 ( 
.A(n_921),
.Y(n_1125)
);

AND2x2_ASAP7_75t_L g1126 ( 
.A(n_920),
.B(n_385),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_999),
.B(n_899),
.Y(n_1127)
);

NOR2xp33_ASAP7_75t_L g1128 ( 
.A(n_916),
.B(n_899),
.Y(n_1128)
);

NOR2xp33_ASAP7_75t_L g1129 ( 
.A(n_963),
.B(n_898),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1060),
.Y(n_1130)
);

OAI21x1_ASAP7_75t_SL g1131 ( 
.A1(n_941),
.A2(n_1004),
.B(n_1020),
.Y(n_1131)
);

BUFx6f_ASAP7_75t_L g1132 ( 
.A(n_1066),
.Y(n_1132)
);

BUFx2_ASAP7_75t_R g1133 ( 
.A(n_1012),
.Y(n_1133)
);

INVxp67_ASAP7_75t_L g1134 ( 
.A(n_917),
.Y(n_1134)
);

BUFx6f_ASAP7_75t_L g1135 ( 
.A(n_1080),
.Y(n_1135)
);

INVx5_ASAP7_75t_L g1136 ( 
.A(n_958),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_945),
.A2(n_898),
.B(n_886),
.Y(n_1137)
);

INVx3_ASAP7_75t_L g1138 ( 
.A(n_921),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_SL g1139 ( 
.A(n_1009),
.B(n_872),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_1084),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_940),
.A2(n_878),
.B(n_869),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1073),
.Y(n_1142)
);

NOR2xp33_ASAP7_75t_L g1143 ( 
.A(n_1019),
.B(n_1007),
.Y(n_1143)
);

AND2x4_ASAP7_75t_L g1144 ( 
.A(n_933),
.B(n_878),
.Y(n_1144)
);

A2O1A1Ixp33_ASAP7_75t_L g1145 ( 
.A1(n_909),
.A2(n_872),
.B(n_385),
.C(n_22),
.Y(n_1145)
);

AND2x2_ASAP7_75t_L g1146 ( 
.A(n_1015),
.B(n_16),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_938),
.B(n_20),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_968),
.B(n_939),
.Y(n_1148)
);

A2O1A1Ixp33_ASAP7_75t_L g1149 ( 
.A1(n_1010),
.A2(n_24),
.B(n_25),
.C(n_26),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_968),
.B(n_89),
.Y(n_1150)
);

A2O1A1Ixp33_ASAP7_75t_L g1151 ( 
.A1(n_942),
.A2(n_25),
.B(n_27),
.C(n_29),
.Y(n_1151)
);

BUFx2_ASAP7_75t_SL g1152 ( 
.A(n_1008),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_931),
.A2(n_91),
.B(n_187),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_936),
.A2(n_87),
.B(n_181),
.Y(n_1154)
);

OAI22xp5_ASAP7_75t_L g1155 ( 
.A1(n_907),
.A2(n_27),
.B1(n_30),
.B2(n_31),
.Y(n_1155)
);

A2O1A1Ixp33_ASAP7_75t_L g1156 ( 
.A1(n_1041),
.A2(n_31),
.B(n_35),
.C(n_37),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_925),
.A2(n_97),
.B(n_180),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_925),
.A2(n_1078),
.B(n_932),
.Y(n_1158)
);

OR2x2_ASAP7_75t_L g1159 ( 
.A(n_1023),
.B(n_974),
.Y(n_1159)
);

AND2x4_ASAP7_75t_L g1160 ( 
.A(n_933),
.B(n_1097),
.Y(n_1160)
);

OAI21xp33_ASAP7_75t_L g1161 ( 
.A1(n_1026),
.A2(n_35),
.B(n_37),
.Y(n_1161)
);

BUFx6f_ASAP7_75t_L g1162 ( 
.A(n_1080),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_929),
.A2(n_113),
.B(n_177),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1079),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1094),
.Y(n_1165)
);

INVxp67_ASAP7_75t_L g1166 ( 
.A(n_1028),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1018),
.B(n_38),
.Y(n_1167)
);

NOR2xp33_ASAP7_75t_L g1168 ( 
.A(n_1090),
.B(n_46),
.Y(n_1168)
);

O2A1O1Ixp33_ASAP7_75t_L g1169 ( 
.A1(n_951),
.A2(n_47),
.B(n_48),
.C(n_49),
.Y(n_1169)
);

INVx1_ASAP7_75t_SL g1170 ( 
.A(n_1018),
.Y(n_1170)
);

AOI21x1_ASAP7_75t_L g1171 ( 
.A1(n_937),
.A2(n_919),
.B(n_910),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1022),
.Y(n_1172)
);

NOR2xp33_ASAP7_75t_L g1173 ( 
.A(n_926),
.B(n_47),
.Y(n_1173)
);

NOR3xp33_ASAP7_75t_SL g1174 ( 
.A(n_1088),
.B(n_49),
.C(n_52),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_946),
.B(n_124),
.Y(n_1175)
);

AOI22xp33_ASAP7_75t_L g1176 ( 
.A1(n_1087),
.A2(n_52),
.B1(n_55),
.B2(n_56),
.Y(n_1176)
);

A2O1A1Ixp33_ASAP7_75t_SL g1177 ( 
.A1(n_1050),
.A2(n_126),
.B(n_175),
.C(n_169),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_SL g1178 ( 
.A(n_1080),
.B(n_114),
.Y(n_1178)
);

O2A1O1Ixp33_ASAP7_75t_L g1179 ( 
.A1(n_959),
.A2(n_55),
.B(n_56),
.C(n_58),
.Y(n_1179)
);

HB1xp67_ASAP7_75t_L g1180 ( 
.A(n_1095),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_SL g1181 ( 
.A(n_1082),
.B(n_136),
.Y(n_1181)
);

OAI21xp33_ASAP7_75t_L g1182 ( 
.A1(n_983),
.A2(n_60),
.B(n_63),
.Y(n_1182)
);

AOI21x1_ASAP7_75t_L g1183 ( 
.A1(n_910),
.A2(n_139),
.B(n_71),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_991),
.Y(n_1184)
);

AOI22xp33_ASAP7_75t_L g1185 ( 
.A1(n_1065),
.A2(n_64),
.B1(n_79),
.B2(n_96),
.Y(n_1185)
);

AO32x2_ASAP7_75t_L g1186 ( 
.A1(n_998),
.A2(n_64),
.A3(n_193),
.B1(n_141),
.B2(n_151),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1002),
.Y(n_1187)
);

OAI21x1_ASAP7_75t_L g1188 ( 
.A1(n_1013),
.A2(n_128),
.B(n_155),
.Y(n_1188)
);

NOR2xp67_ASAP7_75t_SL g1189 ( 
.A(n_1092),
.B(n_163),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_SL g1190 ( 
.A(n_1082),
.B(n_966),
.Y(n_1190)
);

INVxp67_ASAP7_75t_SL g1191 ( 
.A(n_958),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_935),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_955),
.B(n_934),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_929),
.A2(n_923),
.B(n_1062),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_960),
.B(n_986),
.Y(n_1195)
);

NOR2xp33_ASAP7_75t_L g1196 ( 
.A(n_1075),
.B(n_1086),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_1032),
.Y(n_1197)
);

HB1xp67_ASAP7_75t_L g1198 ( 
.A(n_965),
.Y(n_1198)
);

INVx2_ASAP7_75t_SL g1199 ( 
.A(n_976),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1062),
.A2(n_919),
.B(n_961),
.Y(n_1200)
);

AND2x4_ASAP7_75t_L g1201 ( 
.A(n_1097),
.B(n_1047),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1003),
.Y(n_1202)
);

OAI21xp33_ASAP7_75t_SL g1203 ( 
.A1(n_1048),
.A2(n_1053),
.B(n_1000),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_953),
.A2(n_961),
.B(n_985),
.Y(n_1204)
);

INVx3_ASAP7_75t_L g1205 ( 
.A(n_921),
.Y(n_1205)
);

AO21x1_ASAP7_75t_L g1206 ( 
.A1(n_985),
.A2(n_1036),
.B(n_1038),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_SL g1207 ( 
.A(n_1082),
.B(n_1049),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_950),
.B(n_957),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1035),
.Y(n_1209)
);

OR2x6_ASAP7_75t_SL g1210 ( 
.A(n_1058),
.B(n_1061),
.Y(n_1210)
);

A2O1A1Ixp33_ASAP7_75t_SL g1211 ( 
.A1(n_993),
.A2(n_1056),
.B(n_950),
.C(n_957),
.Y(n_1211)
);

AOI22xp5_ASAP7_75t_L g1212 ( 
.A1(n_1037),
.A2(n_1021),
.B1(n_984),
.B2(n_1054),
.Y(n_1212)
);

OAI22x1_ASAP7_75t_L g1213 ( 
.A1(n_990),
.A2(n_1070),
.B1(n_1076),
.B2(n_987),
.Y(n_1213)
);

OAI21xp33_ASAP7_75t_L g1214 ( 
.A1(n_1055),
.A2(n_948),
.B(n_1063),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_SL g1215 ( 
.A(n_958),
.B(n_1097),
.Y(n_1215)
);

O2A1O1Ixp33_ASAP7_75t_SL g1216 ( 
.A1(n_994),
.A2(n_1071),
.B(n_1052),
.C(n_1011),
.Y(n_1216)
);

INVx1_ASAP7_75t_SL g1217 ( 
.A(n_1072),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1040),
.Y(n_1218)
);

NOR2xp33_ASAP7_75t_L g1219 ( 
.A(n_954),
.B(n_1033),
.Y(n_1219)
);

INVxp67_ASAP7_75t_SL g1220 ( 
.A(n_949),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1043),
.B(n_1051),
.Y(n_1221)
);

OAI22xp5_ASAP7_75t_L g1222 ( 
.A1(n_970),
.A2(n_1064),
.B1(n_1089),
.B2(n_1096),
.Y(n_1222)
);

BUFx3_ASAP7_75t_L g1223 ( 
.A(n_1085),
.Y(n_1223)
);

BUFx12f_ASAP7_75t_L g1224 ( 
.A(n_1085),
.Y(n_1224)
);

INVx4_ASAP7_75t_L g1225 ( 
.A(n_1044),
.Y(n_1225)
);

OAI21x1_ASAP7_75t_L g1226 ( 
.A1(n_1013),
.A2(n_1014),
.B(n_1025),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_1059),
.Y(n_1227)
);

INVx2_ASAP7_75t_SL g1228 ( 
.A(n_1085),
.Y(n_1228)
);

INVx2_ASAP7_75t_L g1229 ( 
.A(n_1069),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1083),
.Y(n_1230)
);

OAI21x1_ASAP7_75t_SL g1231 ( 
.A1(n_1034),
.A2(n_1042),
.B(n_1031),
.Y(n_1231)
);

BUFx2_ASAP7_75t_L g1232 ( 
.A(n_1085),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_956),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1024),
.B(n_967),
.Y(n_1234)
);

INVxp67_ASAP7_75t_SL g1235 ( 
.A(n_992),
.Y(n_1235)
);

OAI22xp5_ASAP7_75t_L g1236 ( 
.A1(n_953),
.A2(n_964),
.B1(n_1006),
.B2(n_988),
.Y(n_1236)
);

OR2x2_ASAP7_75t_L g1237 ( 
.A(n_1081),
.B(n_972),
.Y(n_1237)
);

NOR2xp33_ASAP7_75t_R g1238 ( 
.A(n_978),
.B(n_989),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_973),
.Y(n_1239)
);

BUFx3_ASAP7_75t_L g1240 ( 
.A(n_1085),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_977),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_962),
.A2(n_975),
.B(n_980),
.Y(n_1242)
);

BUFx6f_ASAP7_75t_L g1243 ( 
.A(n_979),
.Y(n_1243)
);

AOI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_962),
.A2(n_975),
.B(n_980),
.Y(n_1244)
);

NAND3xp33_ASAP7_75t_SL g1245 ( 
.A(n_1093),
.B(n_1091),
.C(n_1068),
.Y(n_1245)
);

AOI22xp5_ASAP7_75t_L g1246 ( 
.A1(n_1074),
.A2(n_1067),
.B1(n_1068),
.B2(n_1056),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1091),
.B(n_997),
.Y(n_1247)
);

OAI22x1_ASAP7_75t_L g1248 ( 
.A1(n_1093),
.A2(n_1077),
.B1(n_1014),
.B2(n_1067),
.Y(n_1248)
);

OR2x2_ASAP7_75t_SL g1249 ( 
.A(n_1077),
.B(n_1030),
.Y(n_1249)
);

AOI21x1_ASAP7_75t_L g1250 ( 
.A1(n_1016),
.A2(n_996),
.B(n_982),
.Y(n_1250)
);

BUFx8_ASAP7_75t_L g1251 ( 
.A(n_1029),
.Y(n_1251)
);

NOR2xp33_ASAP7_75t_R g1252 ( 
.A(n_1017),
.B(n_1027),
.Y(n_1252)
);

BUFx8_ASAP7_75t_SL g1253 ( 
.A(n_1001),
.Y(n_1253)
);

AOI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_982),
.A2(n_996),
.B(n_1005),
.Y(n_1254)
);

O2A1O1Ixp33_ASAP7_75t_L g1255 ( 
.A1(n_995),
.A2(n_908),
.B(n_915),
.C(n_843),
.Y(n_1255)
);

AND2x4_ASAP7_75t_L g1256 ( 
.A(n_918),
.B(n_933),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_952),
.A2(n_787),
.B(n_658),
.Y(n_1257)
);

AND2x4_ASAP7_75t_L g1258 ( 
.A(n_933),
.B(n_1097),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1057),
.Y(n_1259)
);

OAI22xp5_ASAP7_75t_SL g1260 ( 
.A1(n_913),
.A2(n_924),
.B1(n_411),
.B2(n_421),
.Y(n_1260)
);

INVx2_ASAP7_75t_SL g1261 ( 
.A(n_1117),
.Y(n_1261)
);

OAI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1171),
.A2(n_1200),
.B(n_1242),
.Y(n_1262)
);

AOI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1148),
.A2(n_1203),
.B(n_1194),
.Y(n_1263)
);

NOR2xp67_ASAP7_75t_L g1264 ( 
.A(n_1212),
.B(n_1136),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_SL g1265 ( 
.A1(n_1235),
.A2(n_1255),
.B(n_1150),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1148),
.A2(n_1101),
.B(n_1204),
.Y(n_1266)
);

AND2x2_ASAP7_75t_L g1267 ( 
.A(n_1103),
.B(n_1107),
.Y(n_1267)
);

O2A1O1Ixp33_ASAP7_75t_L g1268 ( 
.A1(n_1143),
.A2(n_1112),
.B(n_1196),
.C(n_1161),
.Y(n_1268)
);

OAI21xp5_ASAP7_75t_SL g1269 ( 
.A1(n_1176),
.A2(n_1166),
.B(n_1109),
.Y(n_1269)
);

AO31x2_ASAP7_75t_L g1270 ( 
.A1(n_1206),
.A2(n_1244),
.A3(n_1248),
.B(n_1254),
.Y(n_1270)
);

NOR2xp33_ASAP7_75t_L g1271 ( 
.A(n_1103),
.B(n_1260),
.Y(n_1271)
);

A2O1A1Ixp33_ASAP7_75t_L g1272 ( 
.A1(n_1214),
.A2(n_1219),
.B(n_1128),
.C(n_1111),
.Y(n_1272)
);

AOI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1257),
.A2(n_1158),
.B(n_1247),
.Y(n_1273)
);

AO31x2_ASAP7_75t_L g1274 ( 
.A1(n_1145),
.A2(n_1213),
.A3(n_1236),
.B(n_1151),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1217),
.B(n_1172),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1217),
.B(n_1184),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1187),
.B(n_1129),
.Y(n_1277)
);

A2O1A1Ixp33_ASAP7_75t_L g1278 ( 
.A1(n_1182),
.A2(n_1173),
.B(n_1115),
.C(n_1119),
.Y(n_1278)
);

NOR2xp33_ASAP7_75t_L g1279 ( 
.A(n_1134),
.B(n_1170),
.Y(n_1279)
);

OR2x2_ASAP7_75t_L g1280 ( 
.A(n_1159),
.B(n_1170),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1233),
.B(n_1114),
.Y(n_1281)
);

NOR2xp67_ASAP7_75t_SL g1282 ( 
.A(n_1100),
.B(n_1136),
.Y(n_1282)
);

OAI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1147),
.A2(n_1222),
.B(n_1099),
.Y(n_1283)
);

BUFx6f_ASAP7_75t_L g1284 ( 
.A(n_1102),
.Y(n_1284)
);

OAI22xp33_ASAP7_75t_L g1285 ( 
.A1(n_1167),
.A2(n_1155),
.B1(n_1210),
.B2(n_1199),
.Y(n_1285)
);

OAI21x1_ASAP7_75t_L g1286 ( 
.A1(n_1250),
.A2(n_1226),
.B(n_1123),
.Y(n_1286)
);

AOI21xp5_ASAP7_75t_L g1287 ( 
.A1(n_1247),
.A2(n_1150),
.B(n_1222),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1108),
.Y(n_1288)
);

OAI21x1_ASAP7_75t_L g1289 ( 
.A1(n_1137),
.A2(n_1141),
.B(n_1188),
.Y(n_1289)
);

OAI22xp33_ASAP7_75t_L g1290 ( 
.A1(n_1155),
.A2(n_1197),
.B1(n_1198),
.B2(n_1237),
.Y(n_1290)
);

INVx2_ASAP7_75t_L g1291 ( 
.A(n_1192),
.Y(n_1291)
);

O2A1O1Ixp33_ASAP7_75t_L g1292 ( 
.A1(n_1156),
.A2(n_1149),
.B(n_1179),
.C(n_1169),
.Y(n_1292)
);

NAND3xp33_ASAP7_75t_L g1293 ( 
.A(n_1121),
.B(n_1174),
.C(n_1185),
.Y(n_1293)
);

A2O1A1Ixp33_ASAP7_75t_L g1294 ( 
.A1(n_1189),
.A2(n_1118),
.B(n_1193),
.C(n_1175),
.Y(n_1294)
);

NAND3xp33_ASAP7_75t_SL g1295 ( 
.A(n_1126),
.B(n_1146),
.C(n_1110),
.Y(n_1295)
);

INVx2_ASAP7_75t_L g1296 ( 
.A(n_1227),
.Y(n_1296)
);

NOR2xp33_ASAP7_75t_L g1297 ( 
.A(n_1180),
.B(n_1190),
.Y(n_1297)
);

INVxp67_ASAP7_75t_L g1298 ( 
.A(n_1133),
.Y(n_1298)
);

OAI21x1_ASAP7_75t_L g1299 ( 
.A1(n_1236),
.A2(n_1120),
.B(n_1131),
.Y(n_1299)
);

OAI21x1_ASAP7_75t_L g1300 ( 
.A1(n_1157),
.A2(n_1183),
.B(n_1231),
.Y(n_1300)
);

AOI221xp5_ASAP7_75t_SL g1301 ( 
.A1(n_1168),
.A2(n_1207),
.B1(n_1193),
.B2(n_1142),
.C(n_1259),
.Y(n_1301)
);

AND2x2_ASAP7_75t_L g1302 ( 
.A(n_1144),
.B(n_1160),
.Y(n_1302)
);

AOI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1105),
.A2(n_1104),
.B(n_1127),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1114),
.B(n_1122),
.Y(n_1304)
);

OAI21x1_ASAP7_75t_L g1305 ( 
.A1(n_1105),
.A2(n_1234),
.B(n_1139),
.Y(n_1305)
);

OAI21x1_ASAP7_75t_L g1306 ( 
.A1(n_1234),
.A2(n_1104),
.B(n_1175),
.Y(n_1306)
);

OAI22x1_ASAP7_75t_L g1307 ( 
.A1(n_1232),
.A2(n_1201),
.B1(n_1256),
.B2(n_1215),
.Y(n_1307)
);

NOR2xp33_ASAP7_75t_L g1308 ( 
.A(n_1144),
.B(n_1152),
.Y(n_1308)
);

AO21x2_ASAP7_75t_L g1309 ( 
.A1(n_1238),
.A2(n_1245),
.B(n_1246),
.Y(n_1309)
);

AOI22xp5_ASAP7_75t_L g1310 ( 
.A1(n_1239),
.A2(n_1241),
.B1(n_1201),
.B2(n_1178),
.Y(n_1310)
);

OAI21x1_ASAP7_75t_L g1311 ( 
.A1(n_1195),
.A2(n_1221),
.B(n_1154),
.Y(n_1311)
);

BUFx12f_ASAP7_75t_L g1312 ( 
.A(n_1106),
.Y(n_1312)
);

BUFx12f_ASAP7_75t_L g1313 ( 
.A(n_1117),
.Y(n_1313)
);

AOI21xp5_ASAP7_75t_L g1314 ( 
.A1(n_1211),
.A2(n_1116),
.B(n_1216),
.Y(n_1314)
);

NAND3xp33_ASAP7_75t_L g1315 ( 
.A(n_1251),
.B(n_1181),
.C(n_1153),
.Y(n_1315)
);

O2A1O1Ixp33_ASAP7_75t_L g1316 ( 
.A1(n_1177),
.A2(n_1130),
.B(n_1165),
.C(n_1164),
.Y(n_1316)
);

OAI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_1256),
.A2(n_1221),
.B(n_1209),
.Y(n_1317)
);

NAND3xp33_ASAP7_75t_L g1318 ( 
.A(n_1251),
.B(n_1243),
.C(n_1202),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1218),
.Y(n_1319)
);

OAI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1225),
.A2(n_1243),
.B1(n_1124),
.B2(n_1230),
.Y(n_1320)
);

NAND2x1_ASAP7_75t_L g1321 ( 
.A(n_1225),
.B(n_1205),
.Y(n_1321)
);

NOR2xp33_ASAP7_75t_SL g1322 ( 
.A(n_1160),
.B(n_1258),
.Y(n_1322)
);

NOR2xp33_ASAP7_75t_L g1323 ( 
.A(n_1258),
.B(n_1243),
.Y(n_1323)
);

O2A1O1Ixp5_ASAP7_75t_SL g1324 ( 
.A1(n_1125),
.A2(n_1205),
.B(n_1138),
.C(n_1208),
.Y(n_1324)
);

AOI21xp5_ASAP7_75t_L g1325 ( 
.A1(n_1220),
.A2(n_1136),
.B(n_1163),
.Y(n_1325)
);

AOI21xp33_ASAP7_75t_L g1326 ( 
.A1(n_1229),
.A2(n_1113),
.B(n_1140),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1191),
.Y(n_1327)
);

AO31x2_ASAP7_75t_L g1328 ( 
.A1(n_1249),
.A2(n_1186),
.A3(n_1252),
.B(n_1228),
.Y(n_1328)
);

AOI21xp5_ASAP7_75t_L g1329 ( 
.A1(n_1125),
.A2(n_1138),
.B(n_1253),
.Y(n_1329)
);

NOR2xp33_ASAP7_75t_L g1330 ( 
.A(n_1132),
.B(n_1135),
.Y(n_1330)
);

NOR2xp33_ASAP7_75t_L g1331 ( 
.A(n_1132),
.B(n_1135),
.Y(n_1331)
);

AOI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1223),
.A2(n_1240),
.B(n_1135),
.Y(n_1332)
);

O2A1O1Ixp33_ASAP7_75t_L g1333 ( 
.A1(n_1186),
.A2(n_1224),
.B(n_1132),
.C(n_1162),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1162),
.B(n_1186),
.Y(n_1334)
);

AOI211x1_ASAP7_75t_L g1335 ( 
.A1(n_1162),
.A2(n_1214),
.B(n_1155),
.C(n_1182),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1108),
.Y(n_1336)
);

CKINVDCx5p33_ASAP7_75t_R g1337 ( 
.A(n_1098),
.Y(n_1337)
);

OAI22xp33_ASAP7_75t_L g1338 ( 
.A1(n_1112),
.A2(n_908),
.B1(n_1026),
.B2(n_843),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1143),
.B(n_788),
.Y(n_1339)
);

O2A1O1Ixp33_ASAP7_75t_SL g1340 ( 
.A1(n_1151),
.A2(n_915),
.B(n_1156),
.C(n_959),
.Y(n_1340)
);

NOR2xp33_ASAP7_75t_L g1341 ( 
.A(n_1166),
.B(n_908),
.Y(n_1341)
);

AOI21xp5_ASAP7_75t_L g1342 ( 
.A1(n_1148),
.A2(n_658),
.B(n_630),
.Y(n_1342)
);

OAI22x1_ASAP7_75t_L g1343 ( 
.A1(n_1196),
.A2(n_1090),
.B1(n_1109),
.B2(n_1107),
.Y(n_1343)
);

NOR2xp33_ASAP7_75t_L g1344 ( 
.A(n_1166),
.B(n_908),
.Y(n_1344)
);

INVx1_ASAP7_75t_SL g1345 ( 
.A(n_1133),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1143),
.B(n_788),
.Y(n_1346)
);

NAND3xp33_ASAP7_75t_SL g1347 ( 
.A(n_1112),
.B(n_913),
.C(n_924),
.Y(n_1347)
);

BUFx2_ASAP7_75t_L g1348 ( 
.A(n_1098),
.Y(n_1348)
);

OAI21x1_ASAP7_75t_L g1349 ( 
.A1(n_1171),
.A2(n_1200),
.B(n_1242),
.Y(n_1349)
);

O2A1O1Ixp33_ASAP7_75t_L g1350 ( 
.A1(n_1143),
.A2(n_908),
.B(n_843),
.C(n_927),
.Y(n_1350)
);

OA21x2_ASAP7_75t_L g1351 ( 
.A1(n_1200),
.A2(n_1204),
.B(n_1226),
.Y(n_1351)
);

AND2x4_ASAP7_75t_L g1352 ( 
.A(n_1160),
.B(n_1258),
.Y(n_1352)
);

INVx2_ASAP7_75t_SL g1353 ( 
.A(n_1117),
.Y(n_1353)
);

AOI22x1_ASAP7_75t_SL g1354 ( 
.A1(n_1106),
.A2(n_814),
.B1(n_891),
.B2(n_696),
.Y(n_1354)
);

INVx1_ASAP7_75t_SL g1355 ( 
.A(n_1133),
.Y(n_1355)
);

INVx3_ASAP7_75t_L g1356 ( 
.A(n_1225),
.Y(n_1356)
);

AOI21xp5_ASAP7_75t_L g1357 ( 
.A1(n_1148),
.A2(n_658),
.B(n_630),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1143),
.B(n_788),
.Y(n_1358)
);

NOR2xp33_ASAP7_75t_L g1359 ( 
.A(n_1166),
.B(n_908),
.Y(n_1359)
);

BUFx2_ASAP7_75t_L g1360 ( 
.A(n_1098),
.Y(n_1360)
);

AOI21xp5_ASAP7_75t_L g1361 ( 
.A1(n_1148),
.A2(n_658),
.B(n_630),
.Y(n_1361)
);

AOI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1148),
.A2(n_658),
.B(n_630),
.Y(n_1362)
);

OAI21x1_ASAP7_75t_L g1363 ( 
.A1(n_1171),
.A2(n_1200),
.B(n_1242),
.Y(n_1363)
);

O2A1O1Ixp33_ASAP7_75t_L g1364 ( 
.A1(n_1143),
.A2(n_908),
.B(n_843),
.C(n_927),
.Y(n_1364)
);

AO31x2_ASAP7_75t_L g1365 ( 
.A1(n_1200),
.A2(n_1206),
.A3(n_1244),
.B(n_1242),
.Y(n_1365)
);

AOI211x1_ASAP7_75t_L g1366 ( 
.A1(n_1214),
.A2(n_1155),
.B(n_1182),
.C(n_1161),
.Y(n_1366)
);

OAI21x1_ASAP7_75t_L g1367 ( 
.A1(n_1171),
.A2(n_1200),
.B(n_1242),
.Y(n_1367)
);

A2O1A1Ixp33_ASAP7_75t_L g1368 ( 
.A1(n_1203),
.A2(n_908),
.B(n_1143),
.C(n_1196),
.Y(n_1368)
);

NOR2xp33_ASAP7_75t_L g1369 ( 
.A(n_1166),
.B(n_908),
.Y(n_1369)
);

OAI22xp5_ASAP7_75t_L g1370 ( 
.A1(n_1143),
.A2(n_759),
.B1(n_908),
.B2(n_843),
.Y(n_1370)
);

AOI21xp5_ASAP7_75t_L g1371 ( 
.A1(n_1148),
.A2(n_658),
.B(n_630),
.Y(n_1371)
);

O2A1O1Ixp33_ASAP7_75t_L g1372 ( 
.A1(n_1143),
.A2(n_908),
.B(n_843),
.C(n_927),
.Y(n_1372)
);

AND2x4_ASAP7_75t_L g1373 ( 
.A(n_1160),
.B(n_1258),
.Y(n_1373)
);

OAI21xp5_ASAP7_75t_L g1374 ( 
.A1(n_1203),
.A2(n_908),
.B(n_915),
.Y(n_1374)
);

A2O1A1Ixp33_ASAP7_75t_L g1375 ( 
.A1(n_1203),
.A2(n_908),
.B(n_1143),
.C(n_1196),
.Y(n_1375)
);

AO31x2_ASAP7_75t_L g1376 ( 
.A1(n_1200),
.A2(n_1206),
.A3(n_1244),
.B(n_1242),
.Y(n_1376)
);

OR2x2_ASAP7_75t_L g1377 ( 
.A(n_1103),
.B(n_875),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1103),
.B(n_761),
.Y(n_1378)
);

INVx1_ASAP7_75t_SL g1379 ( 
.A(n_1133),
.Y(n_1379)
);

NOR2xp67_ASAP7_75t_SL g1380 ( 
.A(n_1100),
.B(n_922),
.Y(n_1380)
);

A2O1A1Ixp33_ASAP7_75t_L g1381 ( 
.A1(n_1203),
.A2(n_908),
.B(n_1143),
.C(n_1196),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1108),
.Y(n_1382)
);

AOI21xp5_ASAP7_75t_L g1383 ( 
.A1(n_1148),
.A2(n_658),
.B(n_630),
.Y(n_1383)
);

AOI21xp5_ASAP7_75t_L g1384 ( 
.A1(n_1148),
.A2(n_658),
.B(n_630),
.Y(n_1384)
);

AOI21xp33_ASAP7_75t_L g1385 ( 
.A1(n_1143),
.A2(n_908),
.B(n_913),
.Y(n_1385)
);

AND2x4_ASAP7_75t_L g1386 ( 
.A(n_1160),
.B(n_1258),
.Y(n_1386)
);

AO31x2_ASAP7_75t_L g1387 ( 
.A1(n_1200),
.A2(n_1206),
.A3(n_1244),
.B(n_1242),
.Y(n_1387)
);

AOI22xp33_ASAP7_75t_L g1388 ( 
.A1(n_1196),
.A2(n_908),
.B1(n_913),
.B2(n_924),
.Y(n_1388)
);

OR2x2_ASAP7_75t_L g1389 ( 
.A(n_1103),
.B(n_875),
.Y(n_1389)
);

OAI21x1_ASAP7_75t_L g1390 ( 
.A1(n_1171),
.A2(n_1200),
.B(n_1242),
.Y(n_1390)
);

AO31x2_ASAP7_75t_L g1391 ( 
.A1(n_1200),
.A2(n_1206),
.A3(n_1244),
.B(n_1242),
.Y(n_1391)
);

AOI21xp5_ASAP7_75t_L g1392 ( 
.A1(n_1148),
.A2(n_658),
.B(n_630),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1108),
.Y(n_1393)
);

NAND2x1p5_ASAP7_75t_L g1394 ( 
.A(n_1102),
.B(n_1136),
.Y(n_1394)
);

OAI221xp5_ASAP7_75t_L g1395 ( 
.A1(n_1112),
.A2(n_908),
.B1(n_913),
.B2(n_924),
.C(n_605),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1108),
.Y(n_1396)
);

INVx5_ASAP7_75t_L g1397 ( 
.A(n_1136),
.Y(n_1397)
);

AOI21xp5_ASAP7_75t_L g1398 ( 
.A1(n_1148),
.A2(n_658),
.B(n_630),
.Y(n_1398)
);

NOR4xp25_ASAP7_75t_L g1399 ( 
.A(n_1161),
.B(n_908),
.C(n_1156),
.D(n_1155),
.Y(n_1399)
);

O2A1O1Ixp33_ASAP7_75t_L g1400 ( 
.A1(n_1143),
.A2(n_908),
.B(n_843),
.C(n_927),
.Y(n_1400)
);

OA21x2_ASAP7_75t_L g1401 ( 
.A1(n_1200),
.A2(n_1204),
.B(n_1226),
.Y(n_1401)
);

OR2x2_ASAP7_75t_L g1402 ( 
.A(n_1103),
.B(n_875),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1103),
.B(n_761),
.Y(n_1403)
);

A2O1A1Ixp33_ASAP7_75t_L g1404 ( 
.A1(n_1203),
.A2(n_908),
.B(n_1143),
.C(n_1196),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1103),
.B(n_761),
.Y(n_1405)
);

AOI21xp5_ASAP7_75t_L g1406 ( 
.A1(n_1148),
.A2(n_658),
.B(n_630),
.Y(n_1406)
);

O2A1O1Ixp33_ASAP7_75t_SL g1407 ( 
.A1(n_1151),
.A2(n_915),
.B(n_1156),
.C(n_959),
.Y(n_1407)
);

AO31x2_ASAP7_75t_L g1408 ( 
.A1(n_1200),
.A2(n_1206),
.A3(n_1244),
.B(n_1242),
.Y(n_1408)
);

AO31x2_ASAP7_75t_L g1409 ( 
.A1(n_1200),
.A2(n_1206),
.A3(n_1244),
.B(n_1242),
.Y(n_1409)
);

AOI21xp5_ASAP7_75t_L g1410 ( 
.A1(n_1148),
.A2(n_658),
.B(n_630),
.Y(n_1410)
);

OAI21x1_ASAP7_75t_SL g1411 ( 
.A1(n_1193),
.A2(n_1175),
.B(n_1131),
.Y(n_1411)
);

CKINVDCx5p33_ASAP7_75t_R g1412 ( 
.A(n_1098),
.Y(n_1412)
);

AOI21xp5_ASAP7_75t_L g1413 ( 
.A1(n_1148),
.A2(n_658),
.B(n_630),
.Y(n_1413)
);

CKINVDCx5p33_ASAP7_75t_R g1414 ( 
.A(n_1098),
.Y(n_1414)
);

NOR2xp33_ASAP7_75t_SL g1415 ( 
.A(n_1133),
.B(n_834),
.Y(n_1415)
);

CKINVDCx8_ASAP7_75t_R g1416 ( 
.A(n_1100),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1143),
.B(n_788),
.Y(n_1417)
);

OR2x2_ASAP7_75t_L g1418 ( 
.A(n_1103),
.B(n_875),
.Y(n_1418)
);

NAND3xp33_ASAP7_75t_L g1419 ( 
.A(n_1143),
.B(n_908),
.C(n_927),
.Y(n_1419)
);

OAI21xp33_ASAP7_75t_L g1420 ( 
.A1(n_1112),
.A2(n_908),
.B(n_927),
.Y(n_1420)
);

AOI21xp5_ASAP7_75t_L g1421 ( 
.A1(n_1148),
.A2(n_658),
.B(n_630),
.Y(n_1421)
);

BUFx2_ASAP7_75t_L g1422 ( 
.A(n_1098),
.Y(n_1422)
);

OAI21x1_ASAP7_75t_L g1423 ( 
.A1(n_1171),
.A2(n_1200),
.B(n_1242),
.Y(n_1423)
);

INVx1_ASAP7_75t_SL g1424 ( 
.A(n_1133),
.Y(n_1424)
);

AOI22xp5_ASAP7_75t_L g1425 ( 
.A1(n_1347),
.A2(n_1395),
.B1(n_1388),
.B2(n_1420),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1288),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1339),
.B(n_1346),
.Y(n_1427)
);

CKINVDCx11_ASAP7_75t_R g1428 ( 
.A(n_1416),
.Y(n_1428)
);

AOI22xp33_ASAP7_75t_L g1429 ( 
.A1(n_1385),
.A2(n_1420),
.B1(n_1293),
.B2(n_1419),
.Y(n_1429)
);

CKINVDCx20_ASAP7_75t_R g1430 ( 
.A(n_1337),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1336),
.Y(n_1431)
);

AOI22xp33_ASAP7_75t_L g1432 ( 
.A1(n_1293),
.A2(n_1419),
.B1(n_1338),
.B2(n_1369),
.Y(n_1432)
);

AOI22xp33_ASAP7_75t_L g1433 ( 
.A1(n_1341),
.A2(n_1359),
.B1(n_1344),
.B2(n_1370),
.Y(n_1433)
);

INVx6_ASAP7_75t_L g1434 ( 
.A(n_1284),
.Y(n_1434)
);

BUFx12f_ASAP7_75t_L g1435 ( 
.A(n_1412),
.Y(n_1435)
);

OAI22xp5_ASAP7_75t_L g1436 ( 
.A1(n_1358),
.A2(n_1417),
.B1(n_1277),
.B2(n_1333),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1296),
.Y(n_1437)
);

BUFx3_ASAP7_75t_L g1438 ( 
.A(n_1313),
.Y(n_1438)
);

CKINVDCx5p33_ASAP7_75t_R g1439 ( 
.A(n_1312),
.Y(n_1439)
);

CKINVDCx16_ASAP7_75t_R g1440 ( 
.A(n_1415),
.Y(n_1440)
);

AOI22xp33_ASAP7_75t_SL g1441 ( 
.A1(n_1271),
.A2(n_1374),
.B1(n_1275),
.B2(n_1276),
.Y(n_1441)
);

BUFx12f_ASAP7_75t_L g1442 ( 
.A(n_1414),
.Y(n_1442)
);

CKINVDCx11_ASAP7_75t_R g1443 ( 
.A(n_1345),
.Y(n_1443)
);

CKINVDCx11_ASAP7_75t_R g1444 ( 
.A(n_1355),
.Y(n_1444)
);

CKINVDCx5p33_ASAP7_75t_R g1445 ( 
.A(n_1354),
.Y(n_1445)
);

CKINVDCx5p33_ASAP7_75t_R g1446 ( 
.A(n_1348),
.Y(n_1446)
);

BUFx10_ASAP7_75t_L g1447 ( 
.A(n_1284),
.Y(n_1447)
);

BUFx12f_ASAP7_75t_L g1448 ( 
.A(n_1360),
.Y(n_1448)
);

OAI21xp5_ASAP7_75t_L g1449 ( 
.A1(n_1368),
.A2(n_1381),
.B(n_1375),
.Y(n_1449)
);

CKINVDCx6p67_ASAP7_75t_R g1450 ( 
.A(n_1397),
.Y(n_1450)
);

BUFx2_ASAP7_75t_L g1451 ( 
.A(n_1422),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1382),
.Y(n_1452)
);

INVx3_ASAP7_75t_L g1453 ( 
.A(n_1397),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1393),
.Y(n_1454)
);

AOI22xp5_ASAP7_75t_L g1455 ( 
.A1(n_1295),
.A2(n_1269),
.B1(n_1290),
.B2(n_1285),
.Y(n_1455)
);

AOI22xp33_ASAP7_75t_L g1456 ( 
.A1(n_1343),
.A2(n_1267),
.B1(n_1264),
.B2(n_1405),
.Y(n_1456)
);

CKINVDCx11_ASAP7_75t_R g1457 ( 
.A(n_1379),
.Y(n_1457)
);

AOI22xp33_ASAP7_75t_L g1458 ( 
.A1(n_1264),
.A2(n_1378),
.B1(n_1403),
.B2(n_1389),
.Y(n_1458)
);

AOI22xp5_ASAP7_75t_L g1459 ( 
.A1(n_1269),
.A2(n_1322),
.B1(n_1308),
.B2(n_1404),
.Y(n_1459)
);

AOI22xp33_ASAP7_75t_L g1460 ( 
.A1(n_1377),
.A2(n_1418),
.B1(n_1402),
.B2(n_1315),
.Y(n_1460)
);

AOI22xp33_ASAP7_75t_L g1461 ( 
.A1(n_1315),
.A2(n_1297),
.B1(n_1411),
.B2(n_1318),
.Y(n_1461)
);

OAI22xp33_ASAP7_75t_L g1462 ( 
.A1(n_1281),
.A2(n_1280),
.B1(n_1310),
.B2(n_1304),
.Y(n_1462)
);

CKINVDCx11_ASAP7_75t_R g1463 ( 
.A(n_1424),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1396),
.Y(n_1464)
);

CKINVDCx5p33_ASAP7_75t_R g1465 ( 
.A(n_1298),
.Y(n_1465)
);

BUFx12f_ASAP7_75t_L g1466 ( 
.A(n_1261),
.Y(n_1466)
);

OAI22xp5_ASAP7_75t_SL g1467 ( 
.A1(n_1366),
.A2(n_1399),
.B1(n_1335),
.B2(n_1318),
.Y(n_1467)
);

AOI22xp5_ASAP7_75t_L g1468 ( 
.A1(n_1278),
.A2(n_1323),
.B1(n_1302),
.B2(n_1380),
.Y(n_1468)
);

AOI22xp33_ASAP7_75t_SL g1469 ( 
.A1(n_1268),
.A2(n_1399),
.B1(n_1366),
.B2(n_1263),
.Y(n_1469)
);

BUFx2_ASAP7_75t_L g1470 ( 
.A(n_1352),
.Y(n_1470)
);

CKINVDCx6p67_ASAP7_75t_R g1471 ( 
.A(n_1352),
.Y(n_1471)
);

BUFx2_ASAP7_75t_L g1472 ( 
.A(n_1373),
.Y(n_1472)
);

OAI22xp33_ASAP7_75t_SL g1473 ( 
.A1(n_1310),
.A2(n_1319),
.B1(n_1400),
.B2(n_1350),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1327),
.Y(n_1474)
);

BUFx2_ASAP7_75t_L g1475 ( 
.A(n_1373),
.Y(n_1475)
);

BUFx3_ASAP7_75t_L g1476 ( 
.A(n_1353),
.Y(n_1476)
);

BUFx4f_ASAP7_75t_SL g1477 ( 
.A(n_1386),
.Y(n_1477)
);

BUFx4f_ASAP7_75t_L g1478 ( 
.A(n_1394),
.Y(n_1478)
);

BUFx12f_ASAP7_75t_L g1479 ( 
.A(n_1386),
.Y(n_1479)
);

CKINVDCx20_ASAP7_75t_R g1480 ( 
.A(n_1279),
.Y(n_1480)
);

AOI22xp33_ASAP7_75t_L g1481 ( 
.A1(n_1307),
.A2(n_1309),
.B1(n_1317),
.B2(n_1283),
.Y(n_1481)
);

AOI22xp33_ASAP7_75t_L g1482 ( 
.A1(n_1309),
.A2(n_1287),
.B1(n_1326),
.B2(n_1282),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1303),
.B(n_1335),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1305),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1272),
.B(n_1372),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1316),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1334),
.Y(n_1487)
);

OAI22x1_ASAP7_75t_L g1488 ( 
.A1(n_1330),
.A2(n_1331),
.B1(n_1364),
.B2(n_1301),
.Y(n_1488)
);

OAI22xp33_ASAP7_75t_R g1489 ( 
.A1(n_1292),
.A2(n_1407),
.B1(n_1340),
.B2(n_1265),
.Y(n_1489)
);

AOI22xp33_ASAP7_75t_L g1490 ( 
.A1(n_1320),
.A2(n_1329),
.B1(n_1314),
.B2(n_1299),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1332),
.B(n_1274),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1356),
.Y(n_1492)
);

INVx1_ASAP7_75t_SL g1493 ( 
.A(n_1321),
.Y(n_1493)
);

BUFx10_ASAP7_75t_L g1494 ( 
.A(n_1324),
.Y(n_1494)
);

OAI21xp5_ASAP7_75t_L g1495 ( 
.A1(n_1294),
.A2(n_1306),
.B(n_1266),
.Y(n_1495)
);

BUFx12f_ASAP7_75t_L g1496 ( 
.A(n_1325),
.Y(n_1496)
);

BUFx6f_ASAP7_75t_L g1497 ( 
.A(n_1311),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1328),
.Y(n_1498)
);

CKINVDCx20_ASAP7_75t_R g1499 ( 
.A(n_1351),
.Y(n_1499)
);

INVx2_ASAP7_75t_SL g1500 ( 
.A(n_1328),
.Y(n_1500)
);

AOI22xp33_ASAP7_75t_L g1501 ( 
.A1(n_1273),
.A2(n_1351),
.B1(n_1401),
.B2(n_1413),
.Y(n_1501)
);

INVx4_ASAP7_75t_L g1502 ( 
.A(n_1401),
.Y(n_1502)
);

AOI22xp33_ASAP7_75t_L g1503 ( 
.A1(n_1342),
.A2(n_1421),
.B1(n_1410),
.B2(n_1406),
.Y(n_1503)
);

BUFx4f_ASAP7_75t_SL g1504 ( 
.A(n_1274),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1274),
.B(n_1270),
.Y(n_1505)
);

OAI22xp33_ASAP7_75t_L g1506 ( 
.A1(n_1357),
.A2(n_1371),
.B1(n_1384),
.B2(n_1383),
.Y(n_1506)
);

AOI22xp5_ASAP7_75t_L g1507 ( 
.A1(n_1361),
.A2(n_1398),
.B1(n_1392),
.B2(n_1362),
.Y(n_1507)
);

AOI22xp33_ASAP7_75t_SL g1508 ( 
.A1(n_1300),
.A2(n_1289),
.B1(n_1367),
.B2(n_1423),
.Y(n_1508)
);

OAI22xp33_ASAP7_75t_L g1509 ( 
.A1(n_1270),
.A2(n_1376),
.B1(n_1408),
.B2(n_1391),
.Y(n_1509)
);

NAND2x1p5_ASAP7_75t_L g1510 ( 
.A(n_1286),
.B(n_1262),
.Y(n_1510)
);

AOI22xp33_ASAP7_75t_SL g1511 ( 
.A1(n_1349),
.A2(n_1363),
.B1(n_1390),
.B2(n_1376),
.Y(n_1511)
);

OAI22xp33_ASAP7_75t_L g1512 ( 
.A1(n_1365),
.A2(n_1376),
.B1(n_1387),
.B2(n_1391),
.Y(n_1512)
);

AOI22xp33_ASAP7_75t_L g1513 ( 
.A1(n_1387),
.A2(n_1391),
.B1(n_1408),
.B2(n_1409),
.Y(n_1513)
);

OAI22xp33_ASAP7_75t_L g1514 ( 
.A1(n_1387),
.A2(n_1346),
.B1(n_1358),
.B2(n_1339),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1408),
.Y(n_1515)
);

BUFx2_ASAP7_75t_R g1516 ( 
.A(n_1409),
.Y(n_1516)
);

AOI22xp33_ASAP7_75t_L g1517 ( 
.A1(n_1409),
.A2(n_1395),
.B1(n_1385),
.B2(n_908),
.Y(n_1517)
);

AND2x4_ASAP7_75t_L g1518 ( 
.A(n_1352),
.B(n_1373),
.Y(n_1518)
);

AOI22xp33_ASAP7_75t_L g1519 ( 
.A1(n_1395),
.A2(n_1385),
.B1(n_908),
.B2(n_1347),
.Y(n_1519)
);

AOI22xp33_ASAP7_75t_L g1520 ( 
.A1(n_1395),
.A2(n_1385),
.B1(n_908),
.B2(n_1347),
.Y(n_1520)
);

AOI22xp33_ASAP7_75t_SL g1521 ( 
.A1(n_1395),
.A2(n_1419),
.B1(n_913),
.B2(n_924),
.Y(n_1521)
);

OAI22xp5_ASAP7_75t_L g1522 ( 
.A1(n_1339),
.A2(n_1346),
.B1(n_1417),
.B2(n_1358),
.Y(n_1522)
);

OAI22xp5_ASAP7_75t_L g1523 ( 
.A1(n_1339),
.A2(n_1346),
.B1(n_1417),
.B2(n_1358),
.Y(n_1523)
);

INVx8_ASAP7_75t_L g1524 ( 
.A(n_1397),
.Y(n_1524)
);

INVx8_ASAP7_75t_L g1525 ( 
.A(n_1397),
.Y(n_1525)
);

INVx6_ASAP7_75t_L g1526 ( 
.A(n_1284),
.Y(n_1526)
);

BUFx12f_ASAP7_75t_L g1527 ( 
.A(n_1337),
.Y(n_1527)
);

INVx6_ASAP7_75t_L g1528 ( 
.A(n_1284),
.Y(n_1528)
);

BUFx12f_ASAP7_75t_L g1529 ( 
.A(n_1337),
.Y(n_1529)
);

AOI22xp33_ASAP7_75t_L g1530 ( 
.A1(n_1395),
.A2(n_1385),
.B1(n_908),
.B2(n_1347),
.Y(n_1530)
);

AOI22xp5_ASAP7_75t_L g1531 ( 
.A1(n_1347),
.A2(n_913),
.B1(n_924),
.B2(n_1112),
.Y(n_1531)
);

CKINVDCx11_ASAP7_75t_R g1532 ( 
.A(n_1416),
.Y(n_1532)
);

INVx6_ASAP7_75t_L g1533 ( 
.A(n_1284),
.Y(n_1533)
);

AOI22xp33_ASAP7_75t_L g1534 ( 
.A1(n_1395),
.A2(n_1385),
.B1(n_908),
.B2(n_1347),
.Y(n_1534)
);

CKINVDCx6p67_ASAP7_75t_R g1535 ( 
.A(n_1312),
.Y(n_1535)
);

INVx2_ASAP7_75t_SL g1536 ( 
.A(n_1313),
.Y(n_1536)
);

BUFx3_ASAP7_75t_L g1537 ( 
.A(n_1313),
.Y(n_1537)
);

AOI22xp33_ASAP7_75t_SL g1538 ( 
.A1(n_1395),
.A2(n_1419),
.B1(n_913),
.B2(n_924),
.Y(n_1538)
);

BUFx3_ASAP7_75t_L g1539 ( 
.A(n_1313),
.Y(n_1539)
);

INVx3_ASAP7_75t_L g1540 ( 
.A(n_1397),
.Y(n_1540)
);

OAI22xp5_ASAP7_75t_L g1541 ( 
.A1(n_1339),
.A2(n_1346),
.B1(n_1417),
.B2(n_1358),
.Y(n_1541)
);

OAI22xp5_ASAP7_75t_L g1542 ( 
.A1(n_1339),
.A2(n_1346),
.B1(n_1417),
.B2(n_1358),
.Y(n_1542)
);

INVx8_ASAP7_75t_L g1543 ( 
.A(n_1397),
.Y(n_1543)
);

BUFx8_ASAP7_75t_L g1544 ( 
.A(n_1312),
.Y(n_1544)
);

AOI22xp5_ASAP7_75t_L g1545 ( 
.A1(n_1347),
.A2(n_913),
.B1(n_924),
.B2(n_1112),
.Y(n_1545)
);

AOI22xp33_ASAP7_75t_L g1546 ( 
.A1(n_1395),
.A2(n_1385),
.B1(n_908),
.B2(n_1347),
.Y(n_1546)
);

OAI22xp33_ASAP7_75t_SL g1547 ( 
.A1(n_1395),
.A2(n_1026),
.B1(n_1346),
.B2(n_1339),
.Y(n_1547)
);

BUFx3_ASAP7_75t_L g1548 ( 
.A(n_1313),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1339),
.B(n_1346),
.Y(n_1549)
);

INVx1_ASAP7_75t_SL g1550 ( 
.A(n_1280),
.Y(n_1550)
);

CKINVDCx11_ASAP7_75t_R g1551 ( 
.A(n_1416),
.Y(n_1551)
);

CKINVDCx10_ASAP7_75t_R g1552 ( 
.A(n_1416),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1267),
.B(n_1378),
.Y(n_1553)
);

INVx6_ASAP7_75t_L g1554 ( 
.A(n_1284),
.Y(n_1554)
);

OAI22xp33_ASAP7_75t_L g1555 ( 
.A1(n_1339),
.A2(n_1358),
.B1(n_1346),
.B2(n_1417),
.Y(n_1555)
);

INVx1_ASAP7_75t_SL g1556 ( 
.A(n_1280),
.Y(n_1556)
);

OAI22xp33_ASAP7_75t_L g1557 ( 
.A1(n_1339),
.A2(n_1358),
.B1(n_1346),
.B2(n_1417),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1291),
.Y(n_1558)
);

OAI22xp5_ASAP7_75t_L g1559 ( 
.A1(n_1339),
.A2(n_1346),
.B1(n_1417),
.B2(n_1358),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1288),
.Y(n_1560)
);

OAI22xp33_ASAP7_75t_L g1561 ( 
.A1(n_1339),
.A2(n_1358),
.B1(n_1346),
.B2(n_1417),
.Y(n_1561)
);

AOI22xp33_ASAP7_75t_SL g1562 ( 
.A1(n_1547),
.A2(n_1449),
.B1(n_1467),
.B2(n_1485),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1498),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1487),
.B(n_1505),
.Y(n_1564)
);

INVx4_ASAP7_75t_L g1565 ( 
.A(n_1524),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1515),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1500),
.Y(n_1567)
);

BUFx2_ASAP7_75t_L g1568 ( 
.A(n_1491),
.Y(n_1568)
);

BUFx2_ASAP7_75t_L g1569 ( 
.A(n_1504),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1449),
.B(n_1553),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1483),
.Y(n_1571)
);

AO21x1_ASAP7_75t_L g1572 ( 
.A1(n_1485),
.A2(n_1486),
.B(n_1473),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1433),
.B(n_1517),
.Y(n_1573)
);

OR2x2_ASAP7_75t_L g1574 ( 
.A(n_1513),
.B(n_1550),
.Y(n_1574)
);

HB1xp67_ASAP7_75t_L g1575 ( 
.A(n_1550),
.Y(n_1575)
);

AO31x2_ASAP7_75t_L g1576 ( 
.A1(n_1502),
.A2(n_1483),
.A3(n_1484),
.B(n_1436),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1555),
.B(n_1557),
.Y(n_1577)
);

BUFx3_ASAP7_75t_L g1578 ( 
.A(n_1496),
.Y(n_1578)
);

BUFx3_ASAP7_75t_L g1579 ( 
.A(n_1524),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1504),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1516),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1497),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1516),
.Y(n_1583)
);

INVxp67_ASAP7_75t_L g1584 ( 
.A(n_1556),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_1497),
.Y(n_1585)
);

OAI21x1_ASAP7_75t_L g1586 ( 
.A1(n_1495),
.A2(n_1510),
.B(n_1501),
.Y(n_1586)
);

HB1xp67_ASAP7_75t_L g1587 ( 
.A(n_1556),
.Y(n_1587)
);

OAI21x1_ASAP7_75t_L g1588 ( 
.A1(n_1495),
.A2(n_1510),
.B(n_1503),
.Y(n_1588)
);

HB1xp67_ASAP7_75t_L g1589 ( 
.A(n_1452),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1499),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1426),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1431),
.Y(n_1592)
);

INVx3_ASAP7_75t_L g1593 ( 
.A(n_1494),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1429),
.B(n_1432),
.Y(n_1594)
);

AOI22xp5_ASAP7_75t_L g1595 ( 
.A1(n_1521),
.A2(n_1538),
.B1(n_1425),
.B2(n_1531),
.Y(n_1595)
);

OAI21x1_ASAP7_75t_L g1596 ( 
.A1(n_1507),
.A2(n_1490),
.B(n_1482),
.Y(n_1596)
);

O2A1O1Ixp33_ASAP7_75t_SL g1597 ( 
.A1(n_1545),
.A2(n_1561),
.B(n_1557),
.C(n_1555),
.Y(n_1597)
);

BUFx3_ASAP7_75t_L g1598 ( 
.A(n_1524),
.Y(n_1598)
);

HB1xp67_ASAP7_75t_L g1599 ( 
.A(n_1454),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1561),
.B(n_1514),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1560),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1509),
.Y(n_1602)
);

HB1xp67_ASAP7_75t_L g1603 ( 
.A(n_1464),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1509),
.Y(n_1604)
);

OAI21x1_ASAP7_75t_L g1605 ( 
.A1(n_1481),
.A2(n_1461),
.B(n_1456),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1494),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1474),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1514),
.B(n_1436),
.Y(n_1608)
);

BUFx3_ASAP7_75t_L g1609 ( 
.A(n_1525),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1512),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1469),
.B(n_1441),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1441),
.B(n_1522),
.Y(n_1612)
);

HB1xp67_ASAP7_75t_L g1613 ( 
.A(n_1488),
.Y(n_1613)
);

BUFx2_ASAP7_75t_L g1614 ( 
.A(n_1455),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1469),
.B(n_1437),
.Y(n_1615)
);

AND2x4_ASAP7_75t_L g1616 ( 
.A(n_1459),
.B(n_1492),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1512),
.Y(n_1617)
);

CKINVDCx5p33_ASAP7_75t_R g1618 ( 
.A(n_1552),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1489),
.Y(n_1619)
);

OA21x2_ASAP7_75t_L g1620 ( 
.A1(n_1519),
.A2(n_1520),
.B(n_1530),
.Y(n_1620)
);

OAI21x1_ASAP7_75t_L g1621 ( 
.A1(n_1508),
.A2(n_1458),
.B(n_1453),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1506),
.Y(n_1622)
);

INVxp67_ASAP7_75t_SL g1623 ( 
.A(n_1462),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1506),
.Y(n_1624)
);

HB1xp67_ASAP7_75t_L g1625 ( 
.A(n_1451),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1558),
.B(n_1427),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1511),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1511),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1462),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1508),
.Y(n_1630)
);

OAI21x1_ASAP7_75t_L g1631 ( 
.A1(n_1453),
.A2(n_1540),
.B(n_1546),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1522),
.Y(n_1632)
);

HB1xp67_ASAP7_75t_L g1633 ( 
.A(n_1470),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1523),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1523),
.Y(n_1635)
);

BUFx3_ASAP7_75t_L g1636 ( 
.A(n_1543),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1427),
.B(n_1549),
.Y(n_1637)
);

NOR2xp33_ASAP7_75t_L g1638 ( 
.A(n_1480),
.B(n_1549),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1559),
.Y(n_1639)
);

OAI21x1_ASAP7_75t_L g1640 ( 
.A1(n_1540),
.A2(n_1534),
.B(n_1460),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1493),
.Y(n_1641)
);

INVx2_ASAP7_75t_SL g1642 ( 
.A(n_1543),
.Y(n_1642)
);

AOI21xp33_ASAP7_75t_L g1643 ( 
.A1(n_1521),
.A2(n_1538),
.B(n_1542),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1541),
.B(n_1559),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1493),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1541),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1542),
.Y(n_1647)
);

BUFx3_ASAP7_75t_L g1648 ( 
.A(n_1450),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1472),
.B(n_1475),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1468),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1518),
.B(n_1471),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1518),
.B(n_1440),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1478),
.Y(n_1653)
);

INVx8_ASAP7_75t_L g1654 ( 
.A(n_1479),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1478),
.Y(n_1655)
);

OA21x2_ASAP7_75t_L g1656 ( 
.A1(n_1445),
.A2(n_1446),
.B(n_1536),
.Y(n_1656)
);

AO21x2_ASAP7_75t_L g1657 ( 
.A1(n_1477),
.A2(n_1447),
.B(n_1554),
.Y(n_1657)
);

INVx3_ASAP7_75t_L g1658 ( 
.A(n_1477),
.Y(n_1658)
);

INVx2_ASAP7_75t_SL g1659 ( 
.A(n_1447),
.Y(n_1659)
);

OAI21x1_ASAP7_75t_L g1660 ( 
.A1(n_1434),
.A2(n_1554),
.B(n_1528),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1434),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1434),
.Y(n_1662)
);

AOI22xp33_ASAP7_75t_L g1663 ( 
.A1(n_1448),
.A2(n_1463),
.B1(n_1457),
.B2(n_1444),
.Y(n_1663)
);

AO21x2_ASAP7_75t_L g1664 ( 
.A1(n_1608),
.A2(n_1554),
.B(n_1533),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1568),
.B(n_1476),
.Y(n_1665)
);

A2O1A1Ixp33_ASAP7_75t_L g1666 ( 
.A1(n_1595),
.A2(n_1548),
.B(n_1539),
.C(n_1438),
.Y(n_1666)
);

AO21x2_ASAP7_75t_L g1667 ( 
.A1(n_1608),
.A2(n_1533),
.B(n_1528),
.Y(n_1667)
);

O2A1O1Ixp33_ASAP7_75t_SL g1668 ( 
.A1(n_1643),
.A2(n_1430),
.B(n_1544),
.C(n_1551),
.Y(n_1668)
);

INVx1_ASAP7_75t_SL g1669 ( 
.A(n_1625),
.Y(n_1669)
);

AOI211xp5_ASAP7_75t_L g1670 ( 
.A1(n_1597),
.A2(n_1465),
.B(n_1537),
.C(n_1439),
.Y(n_1670)
);

AO32x1_ASAP7_75t_L g1671 ( 
.A1(n_1611),
.A2(n_1443),
.A3(n_1526),
.B1(n_1528),
.B2(n_1428),
.Y(n_1671)
);

AOI21xp5_ASAP7_75t_SL g1672 ( 
.A1(n_1595),
.A2(n_1532),
.B(n_1544),
.Y(n_1672)
);

A2O1A1Ixp33_ASAP7_75t_L g1673 ( 
.A1(n_1643),
.A2(n_1526),
.B(n_1535),
.C(n_1466),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1590),
.B(n_1435),
.Y(n_1674)
);

OAI211xp5_ASAP7_75t_L g1675 ( 
.A1(n_1562),
.A2(n_1442),
.B(n_1527),
.C(n_1529),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1564),
.B(n_1570),
.Y(n_1676)
);

OAI21xp5_ASAP7_75t_L g1677 ( 
.A1(n_1612),
.A2(n_1573),
.B(n_1577),
.Y(n_1677)
);

OAI21xp5_ASAP7_75t_L g1678 ( 
.A1(n_1612),
.A2(n_1573),
.B(n_1577),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1570),
.B(n_1591),
.Y(n_1679)
);

BUFx3_ASAP7_75t_L g1680 ( 
.A(n_1660),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1591),
.B(n_1592),
.Y(n_1681)
);

NOR2x1_ASAP7_75t_R g1682 ( 
.A(n_1618),
.B(n_1578),
.Y(n_1682)
);

OAI21xp33_ASAP7_75t_L g1683 ( 
.A1(n_1594),
.A2(n_1611),
.B(n_1644),
.Y(n_1683)
);

OAI22xp5_ASAP7_75t_L g1684 ( 
.A1(n_1614),
.A2(n_1594),
.B1(n_1650),
.B2(n_1644),
.Y(n_1684)
);

OR2x2_ASAP7_75t_L g1685 ( 
.A(n_1610),
.B(n_1617),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1591),
.B(n_1592),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1637),
.B(n_1575),
.Y(n_1687)
);

AOI221xp5_ASAP7_75t_L g1688 ( 
.A1(n_1614),
.A2(n_1600),
.B1(n_1650),
.B2(n_1572),
.C(n_1623),
.Y(n_1688)
);

BUFx2_ASAP7_75t_L g1689 ( 
.A(n_1582),
.Y(n_1689)
);

HB1xp67_ASAP7_75t_L g1690 ( 
.A(n_1587),
.Y(n_1690)
);

AOI21xp5_ASAP7_75t_L g1691 ( 
.A1(n_1600),
.A2(n_1596),
.B(n_1572),
.Y(n_1691)
);

OR2x2_ASAP7_75t_L g1692 ( 
.A(n_1610),
.B(n_1617),
.Y(n_1692)
);

OA21x2_ASAP7_75t_L g1693 ( 
.A1(n_1596),
.A2(n_1586),
.B(n_1588),
.Y(n_1693)
);

NOR2xp33_ASAP7_75t_R g1694 ( 
.A(n_1658),
.B(n_1653),
.Y(n_1694)
);

A2O1A1Ixp33_ASAP7_75t_L g1695 ( 
.A1(n_1605),
.A2(n_1640),
.B(n_1613),
.C(n_1619),
.Y(n_1695)
);

OR2x6_ASAP7_75t_L g1696 ( 
.A(n_1569),
.B(n_1621),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1601),
.Y(n_1697)
);

NOR2xp33_ASAP7_75t_L g1698 ( 
.A(n_1638),
.B(n_1652),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1627),
.B(n_1628),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1627),
.B(n_1628),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1607),
.Y(n_1701)
);

AOI22xp33_ASAP7_75t_L g1702 ( 
.A1(n_1620),
.A2(n_1616),
.B1(n_1578),
.B2(n_1629),
.Y(n_1702)
);

NOR2xp33_ASAP7_75t_L g1703 ( 
.A(n_1652),
.B(n_1637),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1584),
.B(n_1626),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1607),
.B(n_1632),
.Y(n_1705)
);

O2A1O1Ixp33_ASAP7_75t_SL g1706 ( 
.A1(n_1653),
.A2(n_1655),
.B(n_1583),
.C(n_1581),
.Y(n_1706)
);

AOI221xp5_ASAP7_75t_L g1707 ( 
.A1(n_1632),
.A2(n_1635),
.B1(n_1634),
.B2(n_1639),
.C(n_1646),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1626),
.B(n_1589),
.Y(n_1708)
);

BUFx3_ASAP7_75t_L g1709 ( 
.A(n_1660),
.Y(n_1709)
);

CKINVDCx5p33_ASAP7_75t_R g1710 ( 
.A(n_1663),
.Y(n_1710)
);

A2O1A1Ixp33_ASAP7_75t_L g1711 ( 
.A1(n_1605),
.A2(n_1640),
.B(n_1578),
.C(n_1646),
.Y(n_1711)
);

A2O1A1Ixp33_ASAP7_75t_L g1712 ( 
.A1(n_1639),
.A2(n_1647),
.B(n_1581),
.C(n_1583),
.Y(n_1712)
);

OAI21xp5_ASAP7_75t_L g1713 ( 
.A1(n_1620),
.A2(n_1631),
.B(n_1588),
.Y(n_1713)
);

OR2x2_ASAP7_75t_L g1714 ( 
.A(n_1574),
.B(n_1602),
.Y(n_1714)
);

CKINVDCx20_ASAP7_75t_R g1715 ( 
.A(n_1633),
.Y(n_1715)
);

BUFx3_ASAP7_75t_L g1716 ( 
.A(n_1660),
.Y(n_1716)
);

OA21x2_ASAP7_75t_L g1717 ( 
.A1(n_1586),
.A2(n_1630),
.B(n_1624),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1606),
.B(n_1615),
.Y(n_1718)
);

AOI221xp5_ASAP7_75t_SL g1719 ( 
.A1(n_1604),
.A2(n_1615),
.B1(n_1630),
.B2(n_1606),
.C(n_1580),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1599),
.B(n_1603),
.Y(n_1720)
);

AOI22xp5_ASAP7_75t_L g1721 ( 
.A1(n_1620),
.A2(n_1616),
.B1(n_1656),
.B2(n_1651),
.Y(n_1721)
);

NOR2x1_ASAP7_75t_SL g1722 ( 
.A(n_1657),
.B(n_1641),
.Y(n_1722)
);

OR2x2_ASAP7_75t_L g1723 ( 
.A(n_1622),
.B(n_1624),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1576),
.B(n_1571),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_SL g1725 ( 
.A(n_1688),
.B(n_1645),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1724),
.B(n_1566),
.Y(n_1726)
);

OR2x2_ASAP7_75t_L g1727 ( 
.A(n_1717),
.B(n_1576),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1717),
.B(n_1566),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1697),
.Y(n_1729)
);

INVx2_ASAP7_75t_L g1730 ( 
.A(n_1697),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1696),
.B(n_1576),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1696),
.B(n_1576),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1701),
.Y(n_1733)
);

BUFx2_ASAP7_75t_L g1734 ( 
.A(n_1680),
.Y(n_1734)
);

NOR2xp33_ASAP7_75t_L g1735 ( 
.A(n_1683),
.B(n_1656),
.Y(n_1735)
);

NOR2xp33_ASAP7_75t_L g1736 ( 
.A(n_1684),
.B(n_1656),
.Y(n_1736)
);

OR2x2_ASAP7_75t_L g1737 ( 
.A(n_1696),
.B(n_1576),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1693),
.B(n_1679),
.Y(n_1738)
);

AOI22xp33_ASAP7_75t_L g1739 ( 
.A1(n_1677),
.A2(n_1649),
.B1(n_1656),
.B2(n_1654),
.Y(n_1739)
);

OR2x2_ASAP7_75t_L g1740 ( 
.A(n_1714),
.B(n_1685),
.Y(n_1740)
);

INVx3_ASAP7_75t_L g1741 ( 
.A(n_1680),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1713),
.B(n_1563),
.Y(n_1742)
);

INVxp67_ASAP7_75t_L g1743 ( 
.A(n_1664),
.Y(n_1743)
);

BUFx2_ASAP7_75t_L g1744 ( 
.A(n_1709),
.Y(n_1744)
);

INVx2_ASAP7_75t_L g1745 ( 
.A(n_1681),
.Y(n_1745)
);

INVxp67_ASAP7_75t_L g1746 ( 
.A(n_1664),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1705),
.B(n_1593),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1686),
.Y(n_1748)
);

HB1xp67_ASAP7_75t_L g1749 ( 
.A(n_1664),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1676),
.B(n_1593),
.Y(n_1750)
);

AND2x4_ASAP7_75t_L g1751 ( 
.A(n_1716),
.B(n_1585),
.Y(n_1751)
);

OR2x2_ASAP7_75t_L g1752 ( 
.A(n_1714),
.B(n_1567),
.Y(n_1752)
);

NOR3xp33_ASAP7_75t_L g1753 ( 
.A(n_1725),
.B(n_1675),
.C(n_1666),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1729),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1729),
.Y(n_1755)
);

OAI221xp5_ASAP7_75t_L g1756 ( 
.A1(n_1739),
.A2(n_1670),
.B1(n_1678),
.B2(n_1672),
.C(n_1673),
.Y(n_1756)
);

AND2x4_ASAP7_75t_L g1757 ( 
.A(n_1741),
.B(n_1722),
.Y(n_1757)
);

INVx2_ASAP7_75t_L g1758 ( 
.A(n_1728),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1750),
.B(n_1718),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_SL g1760 ( 
.A(n_1735),
.B(n_1721),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1733),
.Y(n_1761)
);

BUFx3_ASAP7_75t_L g1762 ( 
.A(n_1734),
.Y(n_1762)
);

NAND3xp33_ASAP7_75t_SL g1763 ( 
.A(n_1739),
.B(n_1691),
.C(n_1695),
.Y(n_1763)
);

BUFx2_ASAP7_75t_L g1764 ( 
.A(n_1734),
.Y(n_1764)
);

BUFx2_ASAP7_75t_L g1765 ( 
.A(n_1734),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1733),
.Y(n_1766)
);

INVxp67_ASAP7_75t_L g1767 ( 
.A(n_1740),
.Y(n_1767)
);

OR2x2_ASAP7_75t_L g1768 ( 
.A(n_1740),
.B(n_1687),
.Y(n_1768)
);

OR2x2_ASAP7_75t_L g1769 ( 
.A(n_1740),
.B(n_1690),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1735),
.B(n_1669),
.Y(n_1770)
);

AND2x4_ASAP7_75t_L g1771 ( 
.A(n_1741),
.B(n_1722),
.Y(n_1771)
);

AND2x4_ASAP7_75t_L g1772 ( 
.A(n_1741),
.B(n_1667),
.Y(n_1772)
);

AND2x4_ASAP7_75t_L g1773 ( 
.A(n_1741),
.B(n_1667),
.Y(n_1773)
);

NOR2x1_ASAP7_75t_L g1774 ( 
.A(n_1725),
.B(n_1667),
.Y(n_1774)
);

OR2x2_ASAP7_75t_L g1775 ( 
.A(n_1740),
.B(n_1692),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1728),
.Y(n_1776)
);

INVx2_ASAP7_75t_L g1777 ( 
.A(n_1728),
.Y(n_1777)
);

NOR2x1_ASAP7_75t_L g1778 ( 
.A(n_1736),
.B(n_1711),
.Y(n_1778)
);

INVx2_ASAP7_75t_L g1779 ( 
.A(n_1728),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1750),
.B(n_1699),
.Y(n_1780)
);

AND2x2_ASAP7_75t_L g1781 ( 
.A(n_1745),
.B(n_1699),
.Y(n_1781)
);

OR2x2_ASAP7_75t_L g1782 ( 
.A(n_1747),
.B(n_1692),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1745),
.B(n_1700),
.Y(n_1783)
);

INVx3_ASAP7_75t_L g1784 ( 
.A(n_1741),
.Y(n_1784)
);

INVx4_ASAP7_75t_L g1785 ( 
.A(n_1751),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1745),
.B(n_1700),
.Y(n_1786)
);

AND2x2_ASAP7_75t_L g1787 ( 
.A(n_1745),
.B(n_1748),
.Y(n_1787)
);

NAND3xp33_ASAP7_75t_L g1788 ( 
.A(n_1736),
.B(n_1702),
.C(n_1719),
.Y(n_1788)
);

OAI322xp33_ASAP7_75t_L g1789 ( 
.A1(n_1752),
.A2(n_1704),
.A3(n_1672),
.B1(n_1708),
.B2(n_1720),
.C1(n_1723),
.C2(n_1703),
.Y(n_1789)
);

NAND3xp33_ASAP7_75t_L g1790 ( 
.A(n_1743),
.B(n_1712),
.C(n_1707),
.Y(n_1790)
);

OR2x2_ASAP7_75t_L g1791 ( 
.A(n_1747),
.B(n_1689),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_1730),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1748),
.B(n_1665),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1748),
.B(n_1665),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1758),
.Y(n_1795)
);

INVx1_ASAP7_75t_SL g1796 ( 
.A(n_1764),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1785),
.B(n_1738),
.Y(n_1797)
);

HB1xp67_ASAP7_75t_L g1798 ( 
.A(n_1754),
.Y(n_1798)
);

HB1xp67_ASAP7_75t_L g1799 ( 
.A(n_1754),
.Y(n_1799)
);

AND2x2_ASAP7_75t_L g1800 ( 
.A(n_1785),
.B(n_1738),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1785),
.B(n_1738),
.Y(n_1801)
);

INVx2_ASAP7_75t_L g1802 ( 
.A(n_1758),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1785),
.B(n_1738),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1767),
.B(n_1726),
.Y(n_1804)
);

OR2x2_ASAP7_75t_L g1805 ( 
.A(n_1758),
.B(n_1727),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1776),
.B(n_1731),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1776),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1755),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1755),
.Y(n_1809)
);

NAND2xp33_ASAP7_75t_R g1810 ( 
.A(n_1764),
.B(n_1694),
.Y(n_1810)
);

OR2x2_ASAP7_75t_L g1811 ( 
.A(n_1776),
.B(n_1727),
.Y(n_1811)
);

NOR2xp33_ASAP7_75t_L g1812 ( 
.A(n_1789),
.B(n_1710),
.Y(n_1812)
);

HB1xp67_ASAP7_75t_L g1813 ( 
.A(n_1761),
.Y(n_1813)
);

OR2x2_ASAP7_75t_L g1814 ( 
.A(n_1777),
.B(n_1727),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1774),
.B(n_1726),
.Y(n_1815)
);

INVx2_ASAP7_75t_L g1816 ( 
.A(n_1777),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1777),
.B(n_1731),
.Y(n_1817)
);

AND2x2_ASAP7_75t_L g1818 ( 
.A(n_1779),
.B(n_1731),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1774),
.B(n_1726),
.Y(n_1819)
);

HB1xp67_ASAP7_75t_L g1820 ( 
.A(n_1766),
.Y(n_1820)
);

OR2x2_ASAP7_75t_L g1821 ( 
.A(n_1779),
.B(n_1727),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1790),
.B(n_1726),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1787),
.B(n_1731),
.Y(n_1823)
);

INVx2_ASAP7_75t_L g1824 ( 
.A(n_1792),
.Y(n_1824)
);

OR2x2_ASAP7_75t_L g1825 ( 
.A(n_1775),
.B(n_1749),
.Y(n_1825)
);

BUFx6f_ASAP7_75t_L g1826 ( 
.A(n_1762),
.Y(n_1826)
);

AOI22xp33_ASAP7_75t_L g1827 ( 
.A1(n_1753),
.A2(n_1710),
.B1(n_1698),
.B2(n_1715),
.Y(n_1827)
);

OR2x2_ASAP7_75t_L g1828 ( 
.A(n_1775),
.B(n_1749),
.Y(n_1828)
);

BUFx2_ASAP7_75t_L g1829 ( 
.A(n_1762),
.Y(n_1829)
);

INVx2_ASAP7_75t_L g1830 ( 
.A(n_1792),
.Y(n_1830)
);

NOR2xp33_ASAP7_75t_SL g1831 ( 
.A(n_1812),
.B(n_1756),
.Y(n_1831)
);

OR2x2_ASAP7_75t_L g1832 ( 
.A(n_1822),
.B(n_1770),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1812),
.B(n_1788),
.Y(n_1833)
);

OR2x2_ASAP7_75t_L g1834 ( 
.A(n_1822),
.B(n_1760),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1798),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1827),
.B(n_1778),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1827),
.B(n_1778),
.Y(n_1837)
);

OR2x2_ASAP7_75t_L g1838 ( 
.A(n_1815),
.B(n_1769),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_L g1839 ( 
.A(n_1815),
.B(n_1793),
.Y(n_1839)
);

OR2x2_ASAP7_75t_L g1840 ( 
.A(n_1819),
.B(n_1769),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1798),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1799),
.Y(n_1842)
);

AND2x2_ASAP7_75t_L g1843 ( 
.A(n_1829),
.B(n_1759),
.Y(n_1843)
);

INVx1_ASAP7_75t_SL g1844 ( 
.A(n_1829),
.Y(n_1844)
);

NOR3x1_ASAP7_75t_L g1845 ( 
.A(n_1819),
.B(n_1763),
.C(n_1765),
.Y(n_1845)
);

OR2x2_ASAP7_75t_L g1846 ( 
.A(n_1804),
.B(n_1768),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1799),
.Y(n_1847)
);

INVx2_ASAP7_75t_L g1848 ( 
.A(n_1824),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1804),
.B(n_1793),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1813),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_L g1851 ( 
.A(n_1796),
.B(n_1794),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_1796),
.B(n_1794),
.Y(n_1852)
);

INVx2_ASAP7_75t_L g1853 ( 
.A(n_1824),
.Y(n_1853)
);

NOR2x1p5_ASAP7_75t_L g1854 ( 
.A(n_1826),
.B(n_1648),
.Y(n_1854)
);

INVx2_ASAP7_75t_SL g1855 ( 
.A(n_1826),
.Y(n_1855)
);

AND2x2_ASAP7_75t_L g1856 ( 
.A(n_1823),
.B(n_1759),
.Y(n_1856)
);

AND2x4_ASAP7_75t_L g1857 ( 
.A(n_1826),
.B(n_1757),
.Y(n_1857)
);

OR2x2_ASAP7_75t_L g1858 ( 
.A(n_1825),
.B(n_1782),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_L g1859 ( 
.A(n_1826),
.B(n_1780),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1813),
.Y(n_1860)
);

NAND2x1p5_ASAP7_75t_L g1861 ( 
.A(n_1826),
.B(n_1765),
.Y(n_1861)
);

NOR2xp67_ASAP7_75t_L g1862 ( 
.A(n_1826),
.B(n_1784),
.Y(n_1862)
);

INVx2_ASAP7_75t_L g1863 ( 
.A(n_1824),
.Y(n_1863)
);

NOR2x1p5_ASAP7_75t_L g1864 ( 
.A(n_1826),
.B(n_1648),
.Y(n_1864)
);

BUFx3_ASAP7_75t_L g1865 ( 
.A(n_1808),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1823),
.B(n_1780),
.Y(n_1866)
);

OR2x2_ASAP7_75t_L g1867 ( 
.A(n_1825),
.B(n_1782),
.Y(n_1867)
);

INVx2_ASAP7_75t_L g1868 ( 
.A(n_1830),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1820),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1820),
.Y(n_1870)
);

INVx2_ASAP7_75t_L g1871 ( 
.A(n_1830),
.Y(n_1871)
);

AND2x2_ASAP7_75t_L g1872 ( 
.A(n_1823),
.B(n_1781),
.Y(n_1872)
);

INVx2_ASAP7_75t_SL g1873 ( 
.A(n_1808),
.Y(n_1873)
);

OAI22xp5_ASAP7_75t_L g1874 ( 
.A1(n_1825),
.A2(n_1768),
.B1(n_1715),
.B2(n_1737),
.Y(n_1874)
);

OR2x2_ASAP7_75t_L g1875 ( 
.A(n_1828),
.B(n_1791),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1809),
.Y(n_1876)
);

AND2x2_ASAP7_75t_L g1877 ( 
.A(n_1843),
.B(n_1797),
.Y(n_1877)
);

AND3x2_ASAP7_75t_L g1878 ( 
.A(n_1831),
.B(n_1674),
.C(n_1744),
.Y(n_1878)
);

AND2x2_ASAP7_75t_L g1879 ( 
.A(n_1843),
.B(n_1797),
.Y(n_1879)
);

INVx2_ASAP7_75t_L g1880 ( 
.A(n_1861),
.Y(n_1880)
);

HB1xp67_ASAP7_75t_L g1881 ( 
.A(n_1844),
.Y(n_1881)
);

AND2x2_ASAP7_75t_SL g1882 ( 
.A(n_1845),
.B(n_1674),
.Y(n_1882)
);

NOR2xp33_ASAP7_75t_L g1883 ( 
.A(n_1833),
.B(n_1682),
.Y(n_1883)
);

NOR2x1_ASAP7_75t_L g1884 ( 
.A(n_1854),
.B(n_1762),
.Y(n_1884)
);

OR2x2_ASAP7_75t_L g1885 ( 
.A(n_1834),
.B(n_1828),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_L g1886 ( 
.A(n_1836),
.B(n_1781),
.Y(n_1886)
);

NOR2xp33_ASAP7_75t_L g1887 ( 
.A(n_1837),
.B(n_1668),
.Y(n_1887)
);

OR2x2_ASAP7_75t_L g1888 ( 
.A(n_1834),
.B(n_1838),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1864),
.B(n_1797),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_L g1890 ( 
.A(n_1832),
.B(n_1783),
.Y(n_1890)
);

AND2x2_ASAP7_75t_SL g1891 ( 
.A(n_1857),
.B(n_1737),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1876),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1859),
.B(n_1783),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1873),
.Y(n_1894)
);

AND2x2_ASAP7_75t_L g1895 ( 
.A(n_1857),
.B(n_1800),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1873),
.Y(n_1896)
);

OR2x2_ASAP7_75t_L g1897 ( 
.A(n_1838),
.B(n_1828),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1865),
.Y(n_1898)
);

AND3x2_ASAP7_75t_L g1899 ( 
.A(n_1857),
.B(n_1841),
.C(n_1835),
.Y(n_1899)
);

INVx2_ASAP7_75t_L g1900 ( 
.A(n_1861),
.Y(n_1900)
);

INVxp67_ASAP7_75t_SL g1901 ( 
.A(n_1862),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1865),
.Y(n_1902)
);

INVx3_ASAP7_75t_L g1903 ( 
.A(n_1855),
.Y(n_1903)
);

AOI22xp33_ASAP7_75t_L g1904 ( 
.A1(n_1874),
.A2(n_1732),
.B1(n_1757),
.B2(n_1771),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1855),
.B(n_1786),
.Y(n_1905)
);

OR2x2_ASAP7_75t_L g1906 ( 
.A(n_1840),
.B(n_1795),
.Y(n_1906)
);

AND2x2_ASAP7_75t_L g1907 ( 
.A(n_1856),
.B(n_1800),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1851),
.B(n_1852),
.Y(n_1908)
);

CKINVDCx16_ASAP7_75t_R g1909 ( 
.A(n_1856),
.Y(n_1909)
);

BUFx2_ASAP7_75t_SL g1910 ( 
.A(n_1842),
.Y(n_1910)
);

AND2x2_ASAP7_75t_L g1911 ( 
.A(n_1872),
.B(n_1800),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1847),
.Y(n_1912)
);

AND2x4_ASAP7_75t_L g1913 ( 
.A(n_1872),
.B(n_1801),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1850),
.Y(n_1914)
);

O2A1O1Ixp33_ASAP7_75t_L g1915 ( 
.A1(n_1881),
.A2(n_1887),
.B(n_1902),
.C(n_1898),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1892),
.Y(n_1916)
);

AOI22xp5_ASAP7_75t_L g1917 ( 
.A1(n_1882),
.A2(n_1810),
.B1(n_1732),
.B2(n_1771),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1892),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1912),
.Y(n_1919)
);

HB1xp67_ASAP7_75t_L g1920 ( 
.A(n_1903),
.Y(n_1920)
);

AOI21xp33_ASAP7_75t_L g1921 ( 
.A1(n_1882),
.A2(n_1869),
.B(n_1860),
.Y(n_1921)
);

OAI21xp33_ASAP7_75t_L g1922 ( 
.A1(n_1882),
.A2(n_1840),
.B(n_1870),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1912),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_L g1924 ( 
.A(n_1898),
.B(n_1866),
.Y(n_1924)
);

AOI21xp33_ASAP7_75t_L g1925 ( 
.A1(n_1901),
.A2(n_1853),
.B(n_1848),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1914),
.Y(n_1926)
);

OAI22xp33_ASAP7_75t_L g1927 ( 
.A1(n_1909),
.A2(n_1737),
.B1(n_1671),
.B2(n_1875),
.Y(n_1927)
);

OR2x2_ASAP7_75t_L g1928 ( 
.A(n_1888),
.B(n_1886),
.Y(n_1928)
);

INVx2_ASAP7_75t_L g1929 ( 
.A(n_1909),
.Y(n_1929)
);

OAI221xp5_ASAP7_75t_L g1930 ( 
.A1(n_1884),
.A2(n_1875),
.B1(n_1867),
.B2(n_1858),
.C(n_1846),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_L g1931 ( 
.A(n_1902),
.B(n_1839),
.Y(n_1931)
);

XNOR2x2_ASAP7_75t_L g1932 ( 
.A(n_1899),
.B(n_1858),
.Y(n_1932)
);

AOI22xp33_ASAP7_75t_L g1933 ( 
.A1(n_1910),
.A2(n_1732),
.B1(n_1737),
.B2(n_1742),
.Y(n_1933)
);

AOI21xp33_ASAP7_75t_L g1934 ( 
.A1(n_1880),
.A2(n_1853),
.B(n_1848),
.Y(n_1934)
);

OA22x2_ASAP7_75t_L g1935 ( 
.A1(n_1878),
.A2(n_1772),
.B1(n_1773),
.B2(n_1771),
.Y(n_1935)
);

AOI21xp33_ASAP7_75t_SL g1936 ( 
.A1(n_1883),
.A2(n_1867),
.B(n_1654),
.Y(n_1936)
);

INVx2_ASAP7_75t_L g1937 ( 
.A(n_1891),
.Y(n_1937)
);

AND2x2_ASAP7_75t_L g1938 ( 
.A(n_1889),
.B(n_1849),
.Y(n_1938)
);

AOI211xp5_ASAP7_75t_L g1939 ( 
.A1(n_1914),
.A2(n_1888),
.B(n_1900),
.C(n_1880),
.Y(n_1939)
);

AOI21xp5_ASAP7_75t_SL g1940 ( 
.A1(n_1900),
.A2(n_1648),
.B(n_1598),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1910),
.Y(n_1941)
);

XNOR2xp5_ASAP7_75t_L g1942 ( 
.A(n_1932),
.B(n_1891),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1920),
.Y(n_1943)
);

AOI322xp5_ASAP7_75t_L g1944 ( 
.A1(n_1922),
.A2(n_1921),
.A3(n_1933),
.B1(n_1927),
.B2(n_1929),
.C1(n_1941),
.C2(n_1917),
.Y(n_1944)
);

OAI21xp33_ASAP7_75t_L g1945 ( 
.A1(n_1929),
.A2(n_1891),
.B(n_1889),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1920),
.Y(n_1946)
);

AND2x2_ASAP7_75t_L g1947 ( 
.A(n_1937),
.B(n_1895),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1916),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_L g1949 ( 
.A(n_1939),
.B(n_1877),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1918),
.Y(n_1950)
);

OAI21xp5_ASAP7_75t_L g1951 ( 
.A1(n_1915),
.A2(n_1908),
.B(n_1904),
.Y(n_1951)
);

OAI21xp5_ASAP7_75t_L g1952 ( 
.A1(n_1930),
.A2(n_1896),
.B(n_1894),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1919),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1923),
.Y(n_1954)
);

AOI221xp5_ASAP7_75t_L g1955 ( 
.A1(n_1927),
.A2(n_1896),
.B1(n_1894),
.B2(n_1903),
.C(n_1885),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1926),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_SL g1957 ( 
.A(n_1937),
.B(n_1903),
.Y(n_1957)
);

OAI21xp33_ASAP7_75t_L g1958 ( 
.A1(n_1924),
.A2(n_1895),
.B(n_1885),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1928),
.Y(n_1959)
);

AOI211xp5_ASAP7_75t_L g1960 ( 
.A1(n_1936),
.A2(n_1897),
.B(n_1879),
.C(n_1877),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1931),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1938),
.Y(n_1962)
);

INVx2_ASAP7_75t_L g1963 ( 
.A(n_1935),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_SL g1964 ( 
.A(n_1942),
.B(n_1935),
.Y(n_1964)
);

A2O1A1Ixp33_ASAP7_75t_L g1965 ( 
.A1(n_1944),
.A2(n_1933),
.B(n_1925),
.C(n_1934),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1946),
.Y(n_1966)
);

AND2x2_ASAP7_75t_L g1967 ( 
.A(n_1947),
.B(n_1879),
.Y(n_1967)
);

NOR2xp33_ASAP7_75t_L g1968 ( 
.A(n_1942),
.B(n_1940),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_L g1969 ( 
.A(n_1962),
.B(n_1907),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1946),
.Y(n_1970)
);

OAI21xp5_ASAP7_75t_SL g1971 ( 
.A1(n_1951),
.A2(n_1913),
.B(n_1911),
.Y(n_1971)
);

AOI21xp33_ASAP7_75t_L g1972 ( 
.A1(n_1945),
.A2(n_1897),
.B(n_1906),
.Y(n_1972)
);

AOI22xp5_ASAP7_75t_L g1973 ( 
.A1(n_1949),
.A2(n_1905),
.B1(n_1913),
.B2(n_1911),
.Y(n_1973)
);

INVx1_ASAP7_75t_SL g1974 ( 
.A(n_1947),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1943),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1966),
.Y(n_1976)
);

AOI221xp5_ASAP7_75t_L g1977 ( 
.A1(n_1964),
.A2(n_1952),
.B1(n_1955),
.B2(n_1963),
.C(n_1957),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1970),
.Y(n_1978)
);

OAI211xp5_ASAP7_75t_L g1979 ( 
.A1(n_1965),
.A2(n_1957),
.B(n_1960),
.C(n_1963),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1974),
.Y(n_1980)
);

XOR2xp5_ASAP7_75t_L g1981 ( 
.A(n_1973),
.B(n_1959),
.Y(n_1981)
);

NAND2xp33_ASAP7_75t_L g1982 ( 
.A(n_1967),
.B(n_1958),
.Y(n_1982)
);

NOR4xp25_ASAP7_75t_L g1983 ( 
.A(n_1975),
.B(n_1950),
.C(n_1956),
.D(n_1954),
.Y(n_1983)
);

AOI221xp5_ASAP7_75t_L g1984 ( 
.A1(n_1968),
.A2(n_1961),
.B1(n_1953),
.B2(n_1948),
.C(n_1913),
.Y(n_1984)
);

AOI322xp5_ASAP7_75t_L g1985 ( 
.A1(n_1968),
.A2(n_1913),
.A3(n_1907),
.B1(n_1890),
.B2(n_1893),
.C1(n_1818),
.C2(n_1806),
.Y(n_1985)
);

A2O1A1Ixp33_ASAP7_75t_L g1986 ( 
.A1(n_1977),
.A2(n_1971),
.B(n_1972),
.C(n_1969),
.Y(n_1986)
);

AOI22xp5_ASAP7_75t_L g1987 ( 
.A1(n_1979),
.A2(n_1871),
.B1(n_1868),
.B2(n_1863),
.Y(n_1987)
);

AOI221xp5_ASAP7_75t_L g1988 ( 
.A1(n_1983),
.A2(n_1906),
.B1(n_1871),
.B2(n_1868),
.C(n_1863),
.Y(n_1988)
);

NAND3xp33_ASAP7_75t_SL g1989 ( 
.A(n_1984),
.B(n_1803),
.C(n_1801),
.Y(n_1989)
);

NAND3xp33_ASAP7_75t_L g1990 ( 
.A(n_1980),
.B(n_1706),
.C(n_1659),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_L g1991 ( 
.A(n_1981),
.B(n_1801),
.Y(n_1991)
);

OAI221xp5_ASAP7_75t_L g1992 ( 
.A1(n_1986),
.A2(n_1982),
.B1(n_1978),
.B2(n_1976),
.C(n_1985),
.Y(n_1992)
);

AND2x2_ASAP7_75t_L g1993 ( 
.A(n_1991),
.B(n_1803),
.Y(n_1993)
);

AOI211xp5_ASAP7_75t_L g1994 ( 
.A1(n_1989),
.A2(n_1659),
.B(n_1771),
.C(n_1757),
.Y(n_1994)
);

OAI211xp5_ASAP7_75t_L g1995 ( 
.A1(n_1987),
.A2(n_1654),
.B(n_1565),
.C(n_1658),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1990),
.Y(n_1996)
);

AND4x1_ASAP7_75t_L g1997 ( 
.A(n_1988),
.B(n_1803),
.C(n_1661),
.D(n_1662),
.Y(n_1997)
);

NAND3x1_ASAP7_75t_L g1998 ( 
.A(n_1991),
.B(n_1817),
.C(n_1806),
.Y(n_1998)
);

AND2x4_ASAP7_75t_L g1999 ( 
.A(n_1996),
.B(n_1830),
.Y(n_1999)
);

NAND4xp75_ASAP7_75t_L g2000 ( 
.A(n_1993),
.B(n_1642),
.C(n_1806),
.D(n_1818),
.Y(n_2000)
);

INVx1_ASAP7_75t_SL g2001 ( 
.A(n_1998),
.Y(n_2001)
);

INVx3_ASAP7_75t_L g2002 ( 
.A(n_1997),
.Y(n_2002)
);

AND2x4_ASAP7_75t_L g2003 ( 
.A(n_1992),
.B(n_1995),
.Y(n_2003)
);

AND2x2_ASAP7_75t_L g2004 ( 
.A(n_1994),
.B(n_1817),
.Y(n_2004)
);

NAND3xp33_ASAP7_75t_L g2005 ( 
.A(n_2003),
.B(n_1746),
.C(n_1743),
.Y(n_2005)
);

HB1xp67_ASAP7_75t_L g2006 ( 
.A(n_2001),
.Y(n_2006)
);

O2A1O1Ixp33_ASAP7_75t_L g2007 ( 
.A1(n_2001),
.A2(n_1802),
.B(n_1816),
.C(n_1795),
.Y(n_2007)
);

AND2x4_ASAP7_75t_L g2008 ( 
.A(n_2002),
.B(n_1795),
.Y(n_2008)
);

OAI22xp33_ASAP7_75t_L g2009 ( 
.A1(n_2006),
.A2(n_2002),
.B1(n_2003),
.B2(n_2004),
.Y(n_2009)
);

AO22x2_ASAP7_75t_L g2010 ( 
.A1(n_2009),
.A2(n_2008),
.B1(n_1999),
.B2(n_2005),
.Y(n_2010)
);

OA22x2_ASAP7_75t_L g2011 ( 
.A1(n_2010),
.A2(n_1999),
.B1(n_2007),
.B2(n_2000),
.Y(n_2011)
);

NAND5xp2_ASAP7_75t_L g2012 ( 
.A(n_2010),
.B(n_1999),
.C(n_1654),
.D(n_1651),
.E(n_1661),
.Y(n_2012)
);

HB1xp67_ASAP7_75t_L g2013 ( 
.A(n_2011),
.Y(n_2013)
);

OAI22xp5_ASAP7_75t_SL g2014 ( 
.A1(n_2012),
.A2(n_1598),
.B1(n_1636),
.B2(n_1579),
.Y(n_2014)
);

AO22x2_ASAP7_75t_L g2015 ( 
.A1(n_2013),
.A2(n_1802),
.B1(n_1807),
.B2(n_1816),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_2014),
.Y(n_2016)
);

AOI21xp5_ASAP7_75t_L g2017 ( 
.A1(n_2016),
.A2(n_1654),
.B(n_1802),
.Y(n_2017)
);

NAND2xp33_ASAP7_75t_SL g2018 ( 
.A(n_2017),
.B(n_2015),
.Y(n_2018)
);

OAI21xp5_ASAP7_75t_L g2019 ( 
.A1(n_2018),
.A2(n_1816),
.B(n_1807),
.Y(n_2019)
);

OAI221xp5_ASAP7_75t_R g2020 ( 
.A1(n_2019),
.A2(n_1805),
.B1(n_1821),
.B2(n_1811),
.C(n_1814),
.Y(n_2020)
);

AOI211xp5_ASAP7_75t_L g2021 ( 
.A1(n_2020),
.A2(n_1636),
.B(n_1609),
.C(n_1598),
.Y(n_2021)
);


endmodule