module fake_jpeg_13689_n_443 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_443);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_443;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx24_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_9),
.B(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx6f_ASAP7_75t_SL g39 ( 
.A(n_4),
.Y(n_39)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

CKINVDCx14_ASAP7_75t_R g41 ( 
.A(n_10),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_9),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_15),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_29),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_47),
.B(n_59),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_48),
.Y(n_127)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_49),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_50),
.Y(n_133)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx3_ASAP7_75t_SL g126 ( 
.A(n_52),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_29),
.B(n_15),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_53),
.B(n_14),
.Y(n_119)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_54),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g122 ( 
.A(n_55),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_56),
.Y(n_124)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_57),
.Y(n_94)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_58),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_34),
.Y(n_59)
);

INVx11_ASAP7_75t_SL g60 ( 
.A(n_19),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_60),
.Y(n_95)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_61),
.B(n_64),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_62),
.Y(n_103)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_27),
.Y(n_63)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_63),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_19),
.Y(n_64)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_65),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_28),
.Y(n_66)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_66),
.Y(n_125)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_16),
.Y(n_67)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_67),
.Y(n_96)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_68),
.B(n_70),
.Y(n_113)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_27),
.Y(n_69)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_69),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_45),
.B(n_15),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_28),
.Y(n_71)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_71),
.Y(n_132)
);

BUFx8_ASAP7_75t_L g72 ( 
.A(n_25),
.Y(n_72)
);

NAND2x1_ASAP7_75t_SL g120 ( 
.A(n_72),
.B(n_73),
.Y(n_120)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_31),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_74),
.Y(n_118)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g111 ( 
.A(n_75),
.B(n_84),
.Y(n_111)
);

BUFx12_ASAP7_75t_L g76 ( 
.A(n_39),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_76),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_77),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_34),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_78),
.B(n_80),
.Y(n_108)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_27),
.Y(n_79)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_79),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_34),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_34),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_81),
.B(n_83),
.Y(n_110)
);

BUFx10_ASAP7_75t_L g82 ( 
.A(n_28),
.Y(n_82)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_82),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_32),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_18),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_85),
.B(n_86),
.Y(n_112)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_32),
.Y(n_86)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_22),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_87),
.B(n_89),
.Y(n_116)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_41),
.Y(n_88)
);

AOI21xp33_ASAP7_75t_L g142 ( 
.A1(n_88),
.A2(n_3),
.B(n_4),
.Y(n_142)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_22),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_26),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_90),
.B(n_36),
.Y(n_117)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_91),
.B(n_20),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_92),
.B(n_142),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_88),
.A2(n_20),
.B1(n_17),
.B2(n_32),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_97),
.A2(n_98),
.B1(n_105),
.B2(n_135),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_54),
.A2(n_20),
.B1(n_17),
.B2(n_21),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_67),
.B(n_46),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_101),
.B(n_106),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_48),
.A2(n_17),
.B1(n_45),
.B2(n_42),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_102),
.A2(n_107),
.B1(n_129),
.B2(n_131),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_58),
.A2(n_46),
.B1(n_43),
.B2(n_26),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_91),
.B(n_43),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_50),
.A2(n_42),
.B1(n_33),
.B2(n_37),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_52),
.A2(n_33),
.B1(n_37),
.B2(n_23),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_115),
.A2(n_123),
.B1(n_60),
.B2(n_62),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_117),
.B(n_71),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_119),
.B(n_121),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_87),
.B(n_30),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_86),
.A2(n_30),
.B1(n_24),
.B2(n_23),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_73),
.B(n_24),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_128),
.B(n_68),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_63),
.A2(n_36),
.B1(n_35),
.B2(n_41),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_83),
.A2(n_35),
.B1(n_1),
.B2(n_2),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_65),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_49),
.B(n_1),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_136),
.B(n_5),
.Y(n_170)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_95),
.Y(n_144)
);

BUFx2_ASAP7_75t_L g204 ( 
.A(n_144),
.Y(n_204)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_127),
.Y(n_145)
);

INVx3_ASAP7_75t_SL g196 ( 
.A(n_145),
.Y(n_196)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_96),
.Y(n_146)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_146),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_116),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_148),
.B(n_149),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_108),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_123),
.A2(n_79),
.B1(n_69),
.B2(n_57),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_150),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_112),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_151),
.B(n_152),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_110),
.Y(n_152)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_127),
.Y(n_153)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_153),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_92),
.A2(n_56),
.B1(n_77),
.B2(n_74),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_154),
.A2(n_102),
.B1(n_126),
.B2(n_133),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_156),
.B(n_165),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_158),
.A2(n_100),
.B1(n_140),
.B2(n_125),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_115),
.A2(n_82),
.B1(n_55),
.B2(n_66),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_160),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_101),
.B(n_71),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_161),
.A2(n_190),
.B(n_120),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_104),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_162),
.B(n_169),
.Y(n_202)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_95),
.Y(n_163)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_163),
.Y(n_213)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_96),
.Y(n_164)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_164),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_99),
.B(n_66),
.Y(n_165)
);

INVx8_ASAP7_75t_L g166 ( 
.A(n_127),
.Y(n_166)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_166),
.Y(n_228)
);

BUFx4f_ASAP7_75t_SL g167 ( 
.A(n_120),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g229 ( 
.A(n_167),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_134),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_168),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_119),
.B(n_82),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_170),
.B(n_174),
.Y(n_203)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_134),
.Y(n_171)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_171),
.Y(n_198)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_124),
.Y(n_172)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_172),
.Y(n_219)
);

OR2x2_ASAP7_75t_L g173 ( 
.A(n_106),
.B(n_75),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_173),
.B(n_179),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_136),
.B(n_5),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_126),
.A2(n_76),
.B1(n_72),
.B2(n_7),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_175),
.A2(n_189),
.B1(n_126),
.B2(n_141),
.Y(n_195)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_93),
.Y(n_176)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_176),
.Y(n_199)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_93),
.Y(n_177)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_177),
.Y(n_221)
);

BUFx12f_ASAP7_75t_L g178 ( 
.A(n_103),
.Y(n_178)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_178),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_113),
.B(n_76),
.C(n_72),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_138),
.Y(n_180)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_180),
.Y(n_211)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_122),
.Y(n_181)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_181),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_120),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_182),
.B(n_184),
.Y(n_231)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_138),
.Y(n_183)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_183),
.Y(n_215)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_118),
.Y(n_185)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_185),
.Y(n_220)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_122),
.Y(n_186)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_186),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_113),
.B(n_5),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_187),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_113),
.B(n_6),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_188),
.B(n_8),
.Y(n_222)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_118),
.Y(n_189)
);

OR2x2_ASAP7_75t_L g190 ( 
.A(n_107),
.B(n_6),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_193),
.A2(n_164),
.B1(n_177),
.B2(n_133),
.Y(n_245)
);

OAI32xp33_ASAP7_75t_L g194 ( 
.A1(n_157),
.A2(n_111),
.A3(n_131),
.B1(n_130),
.B2(n_137),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_194),
.B(n_222),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_195),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_157),
.A2(n_111),
.B1(n_137),
.B2(n_133),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_201),
.A2(n_224),
.B1(n_161),
.B2(n_151),
.Y(n_236)
);

O2A1O1Ixp33_ASAP7_75t_L g205 ( 
.A1(n_155),
.A2(n_167),
.B(n_161),
.C(n_158),
.Y(n_205)
);

O2A1O1Ixp33_ASAP7_75t_L g259 ( 
.A1(n_205),
.A2(n_122),
.B(n_124),
.C(n_178),
.Y(n_259)
);

AOI211xp5_ASAP7_75t_L g206 ( 
.A1(n_155),
.A2(n_167),
.B(n_152),
.C(n_173),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_206),
.A2(n_159),
.B(n_148),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_207),
.B(n_179),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_143),
.A2(n_141),
.B1(n_100),
.B2(n_132),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_217),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_155),
.A2(n_125),
.B(n_132),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_223),
.A2(n_180),
.B(n_183),
.Y(n_247)
);

OAI22xp33_ASAP7_75t_L g224 ( 
.A1(n_147),
.A2(n_190),
.B1(n_143),
.B2(n_154),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_225),
.A2(n_172),
.B1(n_103),
.B2(n_176),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_170),
.B(n_94),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_226),
.B(n_174),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_233),
.Y(n_288)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_198),
.Y(n_234)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_234),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_209),
.Y(n_235)
);

INVx3_ASAP7_75t_SL g300 ( 
.A(n_235),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_236),
.A2(n_244),
.B1(n_252),
.B2(n_266),
.Y(n_296)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_198),
.Y(n_237)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_237),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_239),
.B(n_243),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_192),
.B(n_162),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_240),
.B(n_242),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_241),
.B(n_204),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_200),
.B(n_149),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_197),
.B(n_171),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_245),
.A2(n_259),
.B1(n_214),
.B2(n_218),
.Y(n_271)
);

INVx3_ASAP7_75t_SL g246 ( 
.A(n_196),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_246),
.A2(n_250),
.B1(n_269),
.B2(n_270),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_247),
.B(n_257),
.Y(n_303)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_191),
.Y(n_248)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_248),
.Y(n_290)
);

AO21x1_ASAP7_75t_SL g250 ( 
.A1(n_205),
.A2(n_114),
.B(n_140),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_203),
.B(n_216),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_251),
.B(n_253),
.C(n_258),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_224),
.A2(n_146),
.B1(n_185),
.B2(n_189),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_203),
.B(n_144),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_202),
.B(n_163),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_254),
.B(n_255),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_230),
.B(n_130),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_208),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_256),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_229),
.B(n_94),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_231),
.B(n_114),
.Y(n_258)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_191),
.Y(n_260)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_260),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_218),
.A2(n_186),
.B(n_181),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_261),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_226),
.B(n_166),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_262),
.B(n_265),
.Y(n_274)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_199),
.Y(n_263)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_263),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_194),
.B(n_153),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_201),
.A2(n_145),
.B1(n_109),
.B2(n_139),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_210),
.Y(n_267)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_267),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_206),
.A2(n_139),
.B1(n_109),
.B2(n_122),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_268),
.A2(n_178),
.B1(n_232),
.B2(n_11),
.Y(n_304)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_229),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_199),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_271),
.B(n_304),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_265),
.A2(n_214),
.B1(n_193),
.B2(n_230),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_277),
.A2(n_282),
.B1(n_286),
.B2(n_287),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_251),
.B(n_223),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_279),
.B(n_281),
.C(n_283),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_233),
.B(n_207),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_249),
.A2(n_208),
.B1(n_209),
.B2(n_219),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_233),
.B(n_211),
.C(n_215),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_236),
.A2(n_219),
.B1(n_196),
.B2(n_228),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_258),
.A2(n_196),
.B1(n_228),
.B2(n_211),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_262),
.A2(n_215),
.B1(n_222),
.B2(n_220),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_289),
.A2(n_293),
.B1(n_301),
.B2(n_246),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_253),
.B(n_227),
.C(n_212),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_291),
.B(n_295),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_245),
.A2(n_220),
.B1(n_213),
.B2(n_204),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_239),
.B(n_227),
.C(n_212),
.Y(n_295)
);

INVx1_ASAP7_75t_SL g320 ( 
.A(n_297),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_264),
.A2(n_213),
.B1(n_210),
.B2(n_221),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_241),
.B(n_221),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_302),
.B(n_247),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_280),
.B(n_238),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_305),
.B(n_309),
.Y(n_336)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_272),
.Y(n_306)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_306),
.Y(n_344)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_308),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_273),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_275),
.Y(n_310)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_310),
.Y(n_358)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_290),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_311),
.B(n_312),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_299),
.B(n_268),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_278),
.A2(n_264),
.B(n_261),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_313),
.A2(n_315),
.B(n_330),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_285),
.B(n_237),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_314),
.B(n_317),
.Y(n_335)
);

XNOR2x1_ASAP7_75t_L g345 ( 
.A(n_315),
.B(n_276),
.Y(n_345)
);

AO21x2_ASAP7_75t_L g316 ( 
.A1(n_284),
.A2(n_250),
.B(n_259),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_316),
.A2(n_271),
.B1(n_288),
.B2(n_282),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_295),
.B(n_234),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_274),
.B(n_270),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_318),
.B(n_322),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_276),
.B(n_252),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_319),
.B(n_279),
.C(n_257),
.Y(n_355)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_292),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_277),
.A2(n_244),
.B1(n_266),
.B2(n_263),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_323),
.A2(n_248),
.B1(n_246),
.B2(n_289),
.Y(n_352)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_294),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g339 ( 
.A(n_324),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_303),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_325),
.B(n_327),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_274),
.B(n_260),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_326),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_303),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_298),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_328),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_302),
.B(n_269),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_329),
.B(n_332),
.Y(n_351)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_293),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_286),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_333),
.B(n_301),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_334),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_320),
.A2(n_303),
.B(n_288),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g361 ( 
.A1(n_337),
.A2(n_341),
.B(n_318),
.Y(n_361)
);

AO21x1_ASAP7_75t_L g338 ( 
.A1(n_330),
.A2(n_297),
.B(n_287),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_338),
.A2(n_342),
.B(n_313),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_320),
.A2(n_296),
.B(n_283),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_321),
.B(n_331),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_343),
.B(n_347),
.C(n_355),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_345),
.B(n_307),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_321),
.B(n_281),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_330),
.A2(n_291),
.B1(n_257),
.B2(n_300),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_348),
.A2(n_352),
.B1(n_306),
.B2(n_300),
.Y(n_379)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_354),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_331),
.B(n_232),
.C(n_267),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_357),
.B(n_308),
.C(n_324),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_360),
.B(n_361),
.Y(n_394)
);

NOR2x1_ASAP7_75t_L g363 ( 
.A(n_335),
.B(n_314),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_363),
.B(n_365),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_346),
.A2(n_316),
.B1(n_332),
.B2(n_333),
.Y(n_364)
);

AOI322xp5_ASAP7_75t_L g380 ( 
.A1(n_364),
.A2(n_367),
.A3(n_378),
.B1(n_334),
.B2(n_338),
.C1(n_351),
.C2(n_352),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_336),
.B(n_317),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_340),
.Y(n_366)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_366),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_346),
.A2(n_316),
.B1(n_326),
.B2(n_307),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_349),
.B(n_319),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_369),
.B(n_372),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_353),
.B(n_328),
.Y(n_370)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_370),
.Y(n_386)
);

BUFx2_ASAP7_75t_L g371 ( 
.A(n_356),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_371),
.B(n_376),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_339),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_340),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_373),
.B(n_379),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_374),
.B(n_357),
.C(n_343),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_375),
.B(n_347),
.C(n_341),
.Y(n_395)
);

INVxp67_ASAP7_75t_SL g376 ( 
.A(n_350),
.Y(n_376)
);

OAI21xp33_ASAP7_75t_L g377 ( 
.A1(n_335),
.A2(n_316),
.B(n_322),
.Y(n_377)
);

HB1xp67_ASAP7_75t_L g387 ( 
.A(n_377),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_338),
.A2(n_316),
.B1(n_323),
.B2(n_310),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_380),
.A2(n_362),
.B1(n_359),
.B2(n_348),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_381),
.B(n_395),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_368),
.B(n_355),
.C(n_345),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_384),
.B(n_389),
.Y(n_400)
);

BUFx2_ASAP7_75t_L g385 ( 
.A(n_362),
.Y(n_385)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_385),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_374),
.B(n_353),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_366),
.B(n_358),
.Y(n_391)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_391),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_373),
.B(n_358),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_392),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_381),
.B(n_368),
.C(n_375),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_398),
.B(n_399),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_395),
.B(n_361),
.C(n_359),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_402),
.B(n_403),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_384),
.B(n_360),
.C(n_367),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_393),
.B(n_363),
.Y(n_404)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_404),
.Y(n_418)
);

BUFx24_ASAP7_75t_SL g406 ( 
.A(n_390),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_406),
.B(n_400),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_394),
.B(n_342),
.C(n_364),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_407),
.B(n_402),
.C(n_403),
.Y(n_409)
);

FAx1_ASAP7_75t_SL g408 ( 
.A(n_387),
.B(n_337),
.CI(n_370),
.CON(n_408),
.SN(n_408)
);

O2A1O1Ixp33_ASAP7_75t_SL g413 ( 
.A1(n_408),
.A2(n_378),
.B(n_388),
.C(n_391),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_409),
.B(n_410),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_401),
.B(n_398),
.C(n_407),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_411),
.B(n_412),
.C(n_417),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_401),
.B(n_394),
.C(n_388),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_413),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_396),
.B(n_385),
.Y(n_415)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_415),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_405),
.B(n_383),
.C(n_382),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_397),
.B(n_386),
.C(n_392),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_419),
.B(n_408),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_SL g430 ( 
.A(n_421),
.B(n_426),
.Y(n_430)
);

NAND3xp33_ASAP7_75t_SL g423 ( 
.A(n_416),
.B(n_408),
.C(n_344),
.Y(n_423)
);

AOI22xp33_ASAP7_75t_L g434 ( 
.A1(n_423),
.A2(n_428),
.B1(n_8),
.B2(n_10),
.Y(n_434)
);

OAI21xp5_ASAP7_75t_L g425 ( 
.A1(n_414),
.A2(n_371),
.B(n_344),
.Y(n_425)
);

CKINVDCx16_ASAP7_75t_R g429 ( 
.A(n_425),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_418),
.B(n_235),
.Y(n_426)
);

A2O1A1Ixp33_ASAP7_75t_SL g428 ( 
.A1(n_413),
.A2(n_356),
.B(n_178),
.C(n_11),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_422),
.B(n_415),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_431),
.B(n_433),
.Y(n_435)
);

OR2x2_ASAP7_75t_L g432 ( 
.A(n_424),
.B(n_356),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_SL g436 ( 
.A1(n_432),
.A2(n_434),
.B(n_428),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_SL g433 ( 
.A(n_420),
.B(n_13),
.Y(n_433)
);

AOI31xp33_ASAP7_75t_L g438 ( 
.A1(n_436),
.A2(n_437),
.A3(n_427),
.B(n_435),
.Y(n_438)
);

BUFx24_ASAP7_75t_SL g437 ( 
.A(n_430),
.Y(n_437)
);

MAJx2_ASAP7_75t_L g440 ( 
.A(n_438),
.B(n_439),
.C(n_434),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_L g439 ( 
.A1(n_435),
.A2(n_429),
.B(n_428),
.Y(n_439)
);

O2A1O1Ixp33_ASAP7_75t_SL g441 ( 
.A1(n_440),
.A2(n_8),
.B(n_10),
.C(n_11),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_L g442 ( 
.A1(n_441),
.A2(n_10),
.B(n_12),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_442),
.B(n_12),
.Y(n_443)
);


endmodule