module fake_jpeg_2963_n_43 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_43);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_43;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_15;

INVx1_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

BUFx3_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx2_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_12),
.B(n_16),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_17),
.B(n_13),
.Y(n_21)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_19),
.B(n_14),
.Y(n_23)
);

OR2x2_ASAP7_75t_L g20 ( 
.A(n_19),
.B(n_15),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_20),
.B(n_21),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_23),
.B(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_20),
.Y(n_25)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_22),
.A2(n_18),
.B1(n_14),
.B2(n_2),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_26),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_L g30 ( 
.A(n_27),
.B(n_7),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_30),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_L g29 ( 
.A1(n_24),
.A2(n_3),
.B(n_4),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_L g34 ( 
.A1(n_29),
.A2(n_26),
.B(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_31),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_32),
.B(n_34),
.Y(n_36)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

XOR2xp5_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_8),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_38),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_SL g40 ( 
.A1(n_36),
.A2(n_4),
.B(n_9),
.Y(n_40)
);

XOR2xp5_ASAP7_75t_L g41 ( 
.A(n_40),
.B(n_37),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_41),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_42),
.B(n_39),
.C(n_10),
.Y(n_43)
);


endmodule