module fake_netlist_5_1426_n_26 (n_8, n_4, n_5, n_7, n_0, n_9, n_2, n_3, n_6, n_1, n_26);

input n_8;
input n_4;
input n_5;
input n_7;
input n_0;
input n_9;
input n_2;
input n_3;
input n_6;
input n_1;

output n_26;

wire n_16;
wire n_12;
wire n_25;
wire n_18;
wire n_22;
wire n_10;
wire n_24;
wire n_21;
wire n_11;
wire n_17;
wire n_19;
wire n_15;
wire n_14;
wire n_23;
wire n_13;
wire n_20;

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_7),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

BUFx3_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

INVx4_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

AOI22xp5_ASAP7_75t_L g15 ( 
.A1(n_14),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_15)
);

AO31x2_ASAP7_75t_L g16 ( 
.A1(n_14),
.A2(n_0),
.A3(n_2),
.B(n_3),
.Y(n_16)
);

NAND3xp33_ASAP7_75t_L g17 ( 
.A(n_14),
.B(n_4),
.C(n_6),
.Y(n_17)
);

AND2x2_ASAP7_75t_L g18 ( 
.A(n_15),
.B(n_13),
.Y(n_18)
);

AO21x2_ASAP7_75t_L g19 ( 
.A1(n_17),
.A2(n_11),
.B(n_12),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_19),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_19),
.Y(n_21)
);

AOI221xp5_ASAP7_75t_L g22 ( 
.A1(n_20),
.A2(n_18),
.B1(n_12),
.B2(n_11),
.C(n_13),
.Y(n_22)
);

AOI311xp33_ASAP7_75t_L g23 ( 
.A1(n_21),
.A2(n_18),
.A3(n_16),
.B(n_14),
.C(n_4),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_22),
.A2(n_10),
.B1(n_8),
.B2(n_9),
.Y(n_24)
);

OAI321xp33_ASAP7_75t_L g25 ( 
.A1(n_24),
.A2(n_10),
.A3(n_23),
.B1(n_15),
.B2(n_22),
.C(n_17),
.Y(n_25)
);

OR2x2_ASAP7_75t_L g26 ( 
.A(n_25),
.B(n_10),
.Y(n_26)
);


endmodule