module fake_jpeg_5414_n_137 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_137);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_137;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_9),
.Y(n_12)
);

BUFx5_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_6),
.B(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx4_ASAP7_75t_SL g27 ( 
.A(n_23),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_29),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_33),
.Y(n_34)
);

OAI22xp33_ASAP7_75t_L g35 ( 
.A1(n_30),
.A2(n_22),
.B1(n_21),
.B2(n_19),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_35),
.A2(n_31),
.B1(n_33),
.B2(n_22),
.Y(n_46)
);

BUFx4f_ASAP7_75t_SL g39 ( 
.A(n_27),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_39),
.Y(n_49)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_29),
.B(n_25),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_15),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_47),
.Y(n_62)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_40),
.A2(n_27),
.B1(n_26),
.B2(n_19),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_41),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_50),
.B(n_54),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_35),
.A2(n_31),
.B1(n_33),
.B2(n_44),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_51),
.A2(n_55),
.B1(n_59),
.B2(n_34),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_42),
.A2(n_26),
.B1(n_21),
.B2(n_15),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_52),
.A2(n_14),
.B1(n_12),
.B2(n_16),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_53),
.B(n_20),
.Y(n_69)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

OA22x2_ASAP7_75t_L g55 ( 
.A1(n_39),
.A2(n_32),
.B1(n_30),
.B2(n_31),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_45),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_56),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_42),
.B(n_25),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_58),
.A2(n_16),
.B(n_39),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_44),
.A2(n_33),
.B1(n_12),
.B2(n_14),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_61),
.B(n_68),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_65),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

NAND2x1p5_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_41),
.Y(n_66)
);

OAI21xp33_ASAP7_75t_L g79 ( 
.A1(n_66),
.A2(n_72),
.B(n_47),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_53),
.B(n_38),
.Y(n_67)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_69),
.B(n_70),
.Y(n_77)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_56),
.A2(n_55),
.B(n_50),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_46),
.A2(n_34),
.B1(n_32),
.B2(n_30),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_49),
.C(n_41),
.Y(n_86)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_74),
.B(n_57),
.Y(n_85)
);

OA21x2_ASAP7_75t_L g95 ( 
.A1(n_79),
.A2(n_82),
.B(n_63),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_75),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_80),
.B(n_89),
.Y(n_99)
);

AND2x4_ASAP7_75t_L g82 ( 
.A(n_66),
.B(n_41),
.Y(n_82)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_84),
.B(n_85),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_86),
.A2(n_71),
.B1(n_73),
.B2(n_68),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_60),
.B(n_49),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_87),
.B(n_65),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_29),
.C(n_36),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_88),
.B(n_28),
.C(n_29),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_74),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_83),
.A2(n_71),
.B1(n_66),
.B2(n_70),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_93),
.Y(n_109)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_87),
.Y(n_93)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_94),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_95),
.A2(n_97),
.B1(n_24),
.B2(n_29),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_96),
.B(n_98),
.C(n_100),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_76),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_88),
.B(n_61),
.C(n_29),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_81),
.B(n_77),
.Y(n_101)
);

OA21x2_ASAP7_75t_SL g110 ( 
.A1(n_101),
.A2(n_11),
.B(n_8),
.Y(n_110)
);

AOI322xp5_ASAP7_75t_L g103 ( 
.A1(n_95),
.A2(n_79),
.A3(n_82),
.B1(n_78),
.B2(n_86),
.C1(n_28),
.C2(n_54),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_103),
.B(n_108),
.C(n_111),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_96),
.A2(n_78),
.B1(n_82),
.B2(n_36),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_104),
.B(n_0),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_107),
.A2(n_32),
.B1(n_24),
.B2(n_37),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_98),
.B(n_28),
.C(n_37),
.Y(n_108)
);

AOI321xp33_ASAP7_75t_L g112 ( 
.A1(n_110),
.A2(n_99),
.A3(n_91),
.B1(n_8),
.B2(n_95),
.C(n_92),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_100),
.B(n_24),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_112),
.A2(n_114),
.B(n_117),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_106),
.B(n_90),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_113),
.B(n_105),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_106),
.B(n_24),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_115),
.A2(n_118),
.B1(n_109),
.B2(n_105),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_SL g117 ( 
.A(n_104),
.B(n_0),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_118),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_119),
.B(n_123),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_120),
.B(n_122),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_116),
.B(n_108),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_118),
.A2(n_102),
.B(n_111),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_124),
.B(n_0),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_119),
.A2(n_102),
.B1(n_1),
.B2(n_2),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_125),
.A2(n_127),
.B(n_129),
.Y(n_130)
);

OAI21x1_ASAP7_75t_SL g129 ( 
.A1(n_121),
.A2(n_5),
.B(n_2),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_128),
.B(n_4),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_131),
.B(n_132),
.C(n_125),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_126),
.B(n_1),
.Y(n_132)
);

NAND3xp33_ASAP7_75t_L g135 ( 
.A(n_133),
.B(n_134),
.C(n_130),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_132),
.B(n_3),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_4),
.Y(n_136)
);

BUFx24_ASAP7_75t_SL g137 ( 
.A(n_136),
.Y(n_137)
);


endmodule