module fake_jpeg_16990_n_294 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_294);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_294;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_273;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_288;
wire n_272;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_7),
.B(n_1),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_15),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_19),
.B(n_0),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_44),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_43),
.B(n_20),
.Y(n_45)
);

BUFx12f_ASAP7_75t_SL g44 ( 
.A(n_27),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_45),
.Y(n_102)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_44),
.A2(n_27),
.B1(n_35),
.B2(n_30),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_48),
.A2(n_27),
.B1(n_24),
.B2(n_32),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_22),
.Y(n_51)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_41),
.A2(n_35),
.B1(n_31),
.B2(n_29),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_53),
.A2(n_62),
.B1(n_23),
.B2(n_29),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_22),
.Y(n_54)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_58),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_34),
.Y(n_59)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_60),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_61),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_36),
.A2(n_35),
.B1(n_31),
.B2(n_23),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_36),
.B(n_34),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_63),
.B(n_65),
.Y(n_69)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_67),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_68),
.B(n_73),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_55),
.A2(n_31),
.B1(n_23),
.B2(n_29),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_70),
.A2(n_81),
.B1(n_85),
.B2(n_89),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_19),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_71),
.B(n_87),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_72),
.A2(n_74),
.B1(n_84),
.B2(n_5),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_28),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_57),
.A2(n_24),
.B1(n_32),
.B2(n_28),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_75),
.Y(n_110)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_76),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_57),
.A2(n_25),
.B1(n_33),
.B2(n_24),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_82),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_53),
.A2(n_26),
.B1(n_37),
.B2(n_21),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_L g85 ( 
.A1(n_52),
.A2(n_37),
.B1(n_26),
.B2(n_33),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_47),
.B(n_18),
.Y(n_87)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_88),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_62),
.A2(n_26),
.B1(n_25),
.B2(n_21),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_47),
.B(n_18),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_90),
.B(n_91),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_49),
.B(n_18),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_64),
.A2(n_26),
.B1(n_2),
.B2(n_3),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_92),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_113)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_93),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_49),
.B(n_18),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_94),
.B(n_95),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_50),
.B(n_0),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_64),
.A2(n_11),
.B1(n_3),
.B2(n_4),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_96),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_103)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_97),
.B(n_98),
.Y(n_127)
);

INVx1_ASAP7_75t_SL g98 ( 
.A(n_61),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_61),
.B(n_0),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_99),
.B(n_20),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_58),
.B(n_4),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_100),
.B(n_21),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_103),
.A2(n_126),
.B1(n_12),
.B2(n_13),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_69),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_104),
.B(n_114),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_107),
.B(n_128),
.Y(n_155)
);

O2A1O1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_67),
.A2(n_65),
.B(n_58),
.C(n_56),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_108),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_109),
.B(n_115),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_113),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_85),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_71),
.B(n_20),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g117 ( 
.A(n_81),
.B(n_56),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_117),
.B(n_99),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_95),
.B(n_91),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_120),
.A2(n_99),
.B1(n_68),
.B2(n_102),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_75),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_121),
.B(n_123),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_122),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_66),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_78),
.A2(n_7),
.B1(n_10),
.B2(n_11),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_77),
.B(n_11),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_83),
.B(n_12),
.Y(n_129)
);

NOR3xp33_ASAP7_75t_L g152 ( 
.A(n_129),
.B(n_96),
.C(n_14),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_131),
.B(n_109),
.C(n_115),
.Y(n_168)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_110),
.Y(n_132)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_132),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_133),
.A2(n_153),
.B(n_157),
.Y(n_169)
);

OAI21xp33_ASAP7_75t_SL g180 ( 
.A1(n_134),
.A2(n_103),
.B(n_126),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_110),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_135),
.B(n_149),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_130),
.B(n_90),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_139),
.B(n_147),
.Y(n_170)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_127),
.Y(n_141)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_141),
.Y(n_176)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_127),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_142),
.Y(n_162)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_124),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_144),
.Y(n_184)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_124),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_145),
.Y(n_161)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_116),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_146),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_130),
.B(n_120),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_106),
.B(n_76),
.Y(n_148)
);

CKINVDCx14_ASAP7_75t_R g163 ( 
.A(n_148),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_106),
.B(n_80),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_120),
.B(n_87),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_151),
.B(n_158),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_152),
.B(n_156),
.Y(n_171)
);

OAI21xp33_ASAP7_75t_L g153 ( 
.A1(n_111),
.A2(n_94),
.B(n_14),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_116),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_154),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_117),
.Y(n_156)
);

A2O1A1O1Ixp25_ASAP7_75t_L g157 ( 
.A1(n_117),
.A2(n_70),
.B(n_82),
.C(n_101),
.D(n_16),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_120),
.B(n_119),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_112),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_159),
.Y(n_173)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_112),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_160),
.Y(n_186)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_159),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_166),
.B(n_167),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_133),
.A2(n_105),
.B(n_111),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_168),
.B(n_179),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_143),
.B(n_119),
.C(n_105),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_175),
.B(n_155),
.C(n_140),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_138),
.A2(n_114),
.B1(n_122),
.B2(n_125),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_178),
.A2(n_180),
.B1(n_183),
.B2(n_185),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_156),
.A2(n_108),
.B(n_107),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_139),
.B(n_123),
.Y(n_181)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_181),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_147),
.B(n_125),
.Y(n_182)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_182),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_138),
.A2(n_108),
.B1(n_118),
.B2(n_97),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_137),
.A2(n_136),
.B1(n_151),
.B2(n_158),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_131),
.B(n_128),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_187),
.B(n_190),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_137),
.A2(n_118),
.B1(n_88),
.B2(n_98),
.Y(n_188)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_188),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_141),
.A2(n_101),
.B1(n_86),
.B2(n_93),
.Y(n_189)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_189),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_142),
.A2(n_86),
.B1(n_79),
.B2(n_129),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_175),
.B(n_143),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_192),
.B(n_193),
.C(n_202),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_174),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_194),
.B(n_198),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_174),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_181),
.B(n_135),
.Y(n_199)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_199),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_170),
.B(n_155),
.Y(n_200)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_200),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_168),
.B(n_160),
.C(n_154),
.Y(n_202)
);

XNOR2x1_ASAP7_75t_SL g203 ( 
.A(n_167),
.B(n_157),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_203),
.B(n_190),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_170),
.B(n_132),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_205),
.B(n_207),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_177),
.B(n_145),
.Y(n_207)
);

BUFx24_ASAP7_75t_SL g208 ( 
.A(n_162),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_208),
.B(n_165),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_166),
.B(n_146),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_209),
.B(n_212),
.Y(n_232)
);

AOI322xp5_ASAP7_75t_L g210 ( 
.A1(n_169),
.A2(n_150),
.A3(n_134),
.B1(n_144),
.B2(n_79),
.C1(n_16),
.C2(n_15),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_210),
.B(n_169),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_177),
.B(n_150),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_185),
.B(n_13),
.C(n_14),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_213),
.B(n_187),
.C(n_171),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_176),
.B(n_13),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_214),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_199),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_215),
.B(n_221),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_216),
.B(n_218),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_192),
.B(n_179),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_217),
.B(n_191),
.Y(n_234)
);

INVxp33_ASAP7_75t_L g218 ( 
.A(n_214),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_212),
.B(n_176),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_222),
.A2(n_225),
.B(n_201),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_206),
.A2(n_182),
.B(n_186),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_226),
.B(n_229),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_228),
.B(n_230),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_191),
.B(n_178),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_195),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_211),
.A2(n_183),
.B1(n_163),
.B2(n_188),
.Y(n_231)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_231),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_234),
.B(n_243),
.C(n_244),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_230),
.A2(n_197),
.B1(n_211),
.B2(n_201),
.Y(n_235)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_235),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_225),
.A2(n_197),
.B(n_204),
.Y(n_238)
);

INVx1_ASAP7_75t_SL g260 ( 
.A(n_238),
.Y(n_260)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_222),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_240),
.B(n_248),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_223),
.B(n_200),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_242),
.B(n_233),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_217),
.B(n_202),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_229),
.B(n_193),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_224),
.B(n_205),
.C(n_207),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_245),
.B(n_220),
.C(n_219),
.Y(n_262)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_227),
.Y(n_246)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_246),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_218),
.B(n_173),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_249),
.B(n_226),
.Y(n_253)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_253),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_245),
.B(n_224),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_254),
.B(n_255),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_236),
.B(n_216),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_237),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_256),
.B(n_259),
.Y(n_268)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_258),
.Y(n_270)
);

OR2x2_ASAP7_75t_L g259 ( 
.A(n_238),
.B(n_232),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_235),
.B(n_189),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_261),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_262),
.B(n_243),
.C(n_249),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_264),
.A2(n_250),
.B(n_222),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_260),
.A2(n_240),
.B(n_241),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_265),
.B(n_253),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_262),
.B(n_250),
.C(n_234),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_267),
.B(n_271),
.Y(n_276)
);

AO21x1_ASAP7_75t_L g271 ( 
.A1(n_260),
.A2(n_203),
.B(n_219),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_257),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_272),
.B(n_164),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_268),
.A2(n_252),
.B1(n_247),
.B2(n_259),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_273),
.B(n_275),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_274),
.B(n_277),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_266),
.B(n_186),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_264),
.B(n_251),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_278),
.B(n_279),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_270),
.A2(n_228),
.B1(n_196),
.B2(n_164),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_280),
.A2(n_276),
.B(n_265),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_282),
.A2(n_285),
.B(n_213),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_278),
.A2(n_263),
.B(n_269),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_274),
.B(n_196),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_286),
.B(n_172),
.C(n_161),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_283),
.A2(n_267),
.B1(n_172),
.B2(n_271),
.Y(n_287)
);

OAI321xp33_ASAP7_75t_L g292 ( 
.A1(n_287),
.A2(n_288),
.A3(n_290),
.B1(n_239),
.B2(n_161),
.C(n_184),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_284),
.B(n_244),
.Y(n_289)
);

A2O1A1Ixp33_ASAP7_75t_L g291 ( 
.A1(n_289),
.A2(n_281),
.B(n_239),
.C(n_173),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_291),
.B(n_292),
.C(n_289),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_293),
.B(n_15),
.Y(n_294)
);


endmodule