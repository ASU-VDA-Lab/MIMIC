module fake_jpeg_1378_n_150 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_150);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_150;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_0),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_24),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

HB1xp67_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_16),
.Y(n_44)
);

BUFx16f_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_21),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_35),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_36),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_11),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_27),
.Y(n_54)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

HB1xp67_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_61),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

BUFx10_ASAP7_75t_L g64 ( 
.A(n_60),
.Y(n_64)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_45),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_57),
.A2(n_42),
.B1(n_48),
.B2(n_41),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_60),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_53),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_71),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_60),
.B(n_39),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_56),
.A2(n_48),
.B1(n_43),
.B2(n_54),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_72),
.A2(n_47),
.B1(n_49),
.B2(n_46),
.Y(n_86)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_74),
.Y(n_97)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_76),
.Y(n_88)
);

OR2x2_ASAP7_75t_SL g76 ( 
.A(n_70),
.B(n_53),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_77),
.B(n_83),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_78),
.A2(n_86),
.B1(n_44),
.B2(n_47),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_66),
.B(n_40),
.C(n_50),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_82),
.Y(n_91)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_63),
.A2(n_54),
.B1(n_43),
.B2(n_62),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_84),
.A2(n_72),
.B1(n_64),
.B2(n_2),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_51),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_85),
.B(n_87),
.Y(n_94)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_64),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_89),
.B(n_101),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_90),
.A2(n_22),
.B1(n_30),
.B2(n_29),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_0),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_93),
.B(n_95),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_1),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_1),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_98),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_2),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_78),
.A2(n_64),
.B1(n_4),
.B2(n_5),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_99),
.A2(n_100),
.B1(n_7),
.B2(n_9),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_74),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_100)
);

OA22x2_ASAP7_75t_L g101 ( 
.A1(n_86),
.A2(n_20),
.B1(n_33),
.B2(n_32),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_75),
.B(n_3),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_102),
.B(n_103),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_6),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_92),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_104),
.B(n_106),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_88),
.A2(n_7),
.B(n_8),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_105),
.A2(n_12),
.B(n_13),
.Y(n_123)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_97),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_94),
.Y(n_107)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_107),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_SL g108 ( 
.A(n_91),
.B(n_99),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_108),
.B(n_113),
.Y(n_127)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_109),
.Y(n_125)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_100),
.Y(n_112)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_112),
.Y(n_131)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_101),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_114),
.B(n_118),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_101),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_92),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_119),
.B(n_15),
.Y(n_130)
);

CKINVDCx11_ASAP7_75t_R g120 ( 
.A(n_92),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_120),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_108),
.B(n_18),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_123),
.B(n_117),
.C(n_115),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_105),
.A2(n_13),
.B(n_34),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_129),
.B(n_116),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_130),
.A2(n_132),
.B1(n_110),
.B2(n_113),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_116),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_133),
.B(n_134),
.Y(n_139)
);

BUFx24_ASAP7_75t_SL g138 ( 
.A(n_135),
.Y(n_138)
);

AO221x1_ASAP7_75t_L g136 ( 
.A1(n_128),
.A2(n_28),
.B1(n_106),
.B2(n_111),
.C(n_124),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_136),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_121),
.B(n_122),
.C(n_127),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_SL g141 ( 
.A(n_137),
.B(n_126),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_141),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_140),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_143),
.A2(n_125),
.B(n_131),
.Y(n_144)
);

AO21x1_ASAP7_75t_L g145 ( 
.A1(n_144),
.A2(n_123),
.B(n_129),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_133),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_142),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_147),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_148),
.A2(n_139),
.B(n_138),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_132),
.Y(n_150)
);


endmodule