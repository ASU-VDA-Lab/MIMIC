module fake_jpeg_7314_n_341 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_341);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_341;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_15),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx11_ASAP7_75t_SL g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx6_ASAP7_75t_SL g34 ( 
.A(n_14),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_8),
.B(n_15),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_39),
.Y(n_68)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_40),
.B(n_41),
.Y(n_76)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx4_ASAP7_75t_SL g42 ( 
.A(n_34),
.Y(n_42)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_45),
.A2(n_25),
.B1(n_26),
.B2(n_47),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g46 ( 
.A(n_18),
.Y(n_46)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_6),
.Y(n_51)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_52),
.B(n_55),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_53),
.Y(n_104)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_47),
.A2(n_26),
.B1(n_25),
.B2(n_32),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_56),
.A2(n_67),
.B1(n_71),
.B2(n_17),
.Y(n_101)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_58),
.B(n_70),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_17),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_62),
.B(n_22),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_66),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_38),
.A2(n_26),
.B1(n_16),
.B2(n_20),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_40),
.B(n_25),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_69),
.B(n_57),
.Y(n_97)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_38),
.A2(n_26),
.B1(n_25),
.B2(n_32),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_41),
.A2(n_20),
.B1(n_21),
.B2(n_16),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_73),
.A2(n_19),
.B1(n_28),
.B2(n_22),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_74),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_73),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_77),
.B(n_81),
.Y(n_121)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_74),
.Y(n_79)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_79),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_76),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_82),
.B(n_83),
.Y(n_145)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_84),
.A2(n_108),
.B1(n_109),
.B2(n_115),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_59),
.A2(n_49),
.B1(n_48),
.B2(n_45),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_85),
.A2(n_46),
.B1(n_75),
.B2(n_36),
.Y(n_128)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_86),
.B(n_88),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_66),
.Y(n_87)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_87),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_65),
.B(n_28),
.Y(n_88)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g132 ( 
.A(n_89),
.Y(n_132)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_69),
.Y(n_90)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_90),
.Y(n_124)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_52),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_91),
.Y(n_123)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_55),
.Y(n_92)
);

INVx4_ASAP7_75t_SL g134 ( 
.A(n_92),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_65),
.B(n_21),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_93),
.B(n_99),
.Y(n_143)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_58),
.Y(n_94)
);

HB1xp67_ASAP7_75t_L g120 ( 
.A(n_94),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_70),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_95),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_74),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_96),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_97),
.A2(n_100),
.B(n_18),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_61),
.B(n_17),
.Y(n_99)
);

NAND2xp33_ASAP7_75t_SL g100 ( 
.A(n_60),
.B(n_45),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_101),
.A2(n_24),
.B1(n_37),
.B2(n_31),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_72),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_102),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_103),
.A2(n_105),
.B1(n_36),
.B2(n_35),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_64),
.A2(n_19),
.B1(n_32),
.B2(n_28),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_72),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g153 ( 
.A(n_106),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_57),
.B(n_22),
.Y(n_107)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_107),
.Y(n_126)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_72),
.Y(n_108)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_64),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_61),
.Y(n_110)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_110),
.Y(n_133)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_63),
.Y(n_111)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_111),
.Y(n_146)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_63),
.Y(n_113)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_113),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_60),
.B(n_43),
.C(n_44),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_114),
.B(n_40),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_68),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_68),
.Y(n_116)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_116),
.Y(n_148)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_117),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_118),
.A2(n_129),
.B1(n_152),
.B2(n_30),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_127),
.A2(n_97),
.B(n_114),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_128),
.A2(n_108),
.B1(n_80),
.B2(n_84),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_104),
.A2(n_75),
.B1(n_36),
.B2(n_46),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_104),
.A2(n_23),
.B(n_29),
.Y(n_130)
);

A2O1A1Ixp33_ASAP7_75t_L g181 ( 
.A1(n_130),
.A2(n_141),
.B(n_147),
.C(n_13),
.Y(n_181)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_79),
.Y(n_131)
);

INVxp67_ASAP7_75t_SL g159 ( 
.A(n_131),
.Y(n_159)
);

NAND2xp33_ASAP7_75t_SL g156 ( 
.A(n_135),
.B(n_97),
.Y(n_156)
);

AND2x2_ASAP7_75t_SL g137 ( 
.A(n_99),
.B(n_29),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_137),
.B(n_82),
.Y(n_157)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_92),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_139),
.Y(n_160)
);

FAx1_ASAP7_75t_L g141 ( 
.A(n_117),
.B(n_42),
.CI(n_18),
.CON(n_141),
.SN(n_141)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_103),
.A2(n_37),
.B1(n_31),
.B2(n_29),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_144),
.A2(n_85),
.B1(n_109),
.B2(n_80),
.Y(n_155)
);

AOI32xp33_ASAP7_75t_L g147 ( 
.A1(n_100),
.A2(n_50),
.A3(n_42),
.B1(n_24),
.B2(n_31),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_78),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_151),
.B(n_93),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_154),
.B(n_156),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_155),
.A2(n_167),
.B1(n_186),
.B2(n_131),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_157),
.B(n_158),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_150),
.B(n_113),
.Y(n_158)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_161),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_145),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_162),
.B(n_169),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_163),
.A2(n_181),
.B1(n_187),
.B2(n_182),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_128),
.A2(n_89),
.B1(n_94),
.B2(n_112),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_164),
.A2(n_172),
.B1(n_182),
.B2(n_140),
.Y(n_198)
);

AO22x1_ASAP7_75t_L g165 ( 
.A1(n_141),
.A2(n_98),
.B1(n_37),
.B2(n_24),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_165),
.B(n_166),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_150),
.B(n_37),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_152),
.A2(n_98),
.B1(n_102),
.B2(n_106),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_137),
.B(n_0),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_168),
.B(n_176),
.Y(n_206)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_137),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_143),
.B(n_126),
.Y(n_170)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_170),
.Y(n_196)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_121),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_171),
.B(n_173),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_141),
.A2(n_96),
.B1(n_50),
.B2(n_87),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_143),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_144),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_174),
.B(n_175),
.Y(n_204)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_149),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_119),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_127),
.B(n_0),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_177),
.B(n_179),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g211 ( 
.A1(n_178),
.A2(n_133),
.B1(n_132),
.B2(n_142),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_126),
.B(n_0),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_122),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_180),
.B(n_183),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_135),
.A2(n_6),
.B1(n_12),
.B2(n_11),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_122),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_127),
.B(n_1),
.Y(n_184)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_184),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_124),
.B(n_1),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_185),
.B(n_146),
.Y(n_202)
);

OA22x2_ASAP7_75t_L g186 ( 
.A1(n_140),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_130),
.A2(n_13),
.B1(n_11),
.B2(n_10),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_154),
.B(n_118),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_189),
.B(n_190),
.C(n_205),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_184),
.B(n_157),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_191),
.B(n_203),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_172),
.A2(n_125),
.B1(n_146),
.B2(n_133),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_193),
.A2(n_199),
.B1(n_211),
.B2(n_220),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_198),
.B(n_207),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_202),
.B(n_208),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_158),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_173),
.B(n_148),
.C(n_123),
.Y(n_205)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_166),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_159),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_169),
.B(n_148),
.C(n_132),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_209),
.B(n_213),
.C(n_216),
.Y(n_244)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_179),
.Y(n_210)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_210),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_181),
.A2(n_134),
.B1(n_136),
.B2(n_142),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_212),
.A2(n_218),
.B1(n_186),
.B2(n_175),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_168),
.B(n_120),
.C(n_134),
.Y(n_213)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_163),
.Y(n_215)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_215),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_164),
.B(n_139),
.C(n_153),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_174),
.A2(n_153),
.B1(n_138),
.B2(n_3),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_180),
.Y(n_219)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_219),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_176),
.A2(n_11),
.B1(n_10),
.B2(n_9),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_219),
.Y(n_221)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_221),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_217),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_223),
.B(n_242),
.Y(n_250)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_217),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_225),
.B(n_226),
.Y(n_256)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_194),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_201),
.A2(n_165),
.B(n_171),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_229),
.A2(n_237),
.B1(n_206),
.B2(n_214),
.Y(n_259)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_194),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_230),
.B(n_233),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_200),
.B(n_189),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_231),
.B(n_236),
.C(n_213),
.Y(n_260)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_204),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_195),
.B(n_214),
.Y(n_234)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_234),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_235),
.A2(n_246),
.B1(n_198),
.B2(n_212),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_200),
.B(n_177),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_201),
.A2(n_165),
.B(n_177),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_218),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_238),
.B(n_240),
.Y(n_258)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_188),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_216),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_206),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_243),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_199),
.A2(n_167),
.B1(n_155),
.B2(n_186),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_205),
.Y(n_247)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_247),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_248),
.A2(n_255),
.B1(n_263),
.B2(n_268),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_221),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_251),
.B(n_267),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_231),
.B(n_190),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_253),
.B(n_260),
.C(n_262),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_224),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_254),
.B(n_269),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_246),
.A2(n_196),
.B1(n_197),
.B2(n_208),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_259),
.B(n_229),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_239),
.A2(n_209),
.B1(n_192),
.B2(n_186),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_261),
.A2(n_222),
.B1(n_233),
.B2(n_228),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_232),
.B(n_202),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_242),
.A2(n_160),
.B1(n_183),
.B2(n_185),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_225),
.B(n_185),
.Y(n_265)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_265),
.Y(n_276)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_234),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_235),
.A2(n_238),
.B1(n_241),
.B2(n_230),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_245),
.Y(n_269)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_258),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_271),
.B(n_275),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_SL g295 ( 
.A(n_273),
.B(n_248),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_258),
.B(n_226),
.Y(n_274)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_274),
.Y(n_290)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_257),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_268),
.A2(n_237),
.B(n_227),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_277),
.A2(n_287),
.B(n_265),
.Y(n_301)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_257),
.Y(n_278)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_278),
.Y(n_292)
);

INVx1_ASAP7_75t_SL g280 ( 
.A(n_256),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_280),
.B(n_285),
.Y(n_289)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_281),
.Y(n_296)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_256),
.Y(n_282)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_282),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_260),
.B(n_232),
.C(n_244),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_283),
.B(n_284),
.C(n_262),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_253),
.B(n_244),
.C(n_227),
.Y(n_284)
);

INVxp33_ASAP7_75t_L g285 ( 
.A(n_250),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_252),
.B(n_240),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_286),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_249),
.B(n_236),
.Y(n_287)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_291),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_284),
.B(n_266),
.C(n_263),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_293),
.B(n_273),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_279),
.A2(n_266),
.B1(n_267),
.B2(n_249),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_294),
.A2(n_298),
.B1(n_272),
.B2(n_138),
.Y(n_309)
);

MAJx2_ASAP7_75t_L g310 ( 
.A(n_295),
.B(n_299),
.C(n_302),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_279),
.A2(n_280),
.B1(n_276),
.B2(n_261),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_272),
.B(n_255),
.Y(n_299)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_301),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_276),
.A2(n_264),
.B(n_251),
.Y(n_302)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_304),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_295),
.A2(n_270),
.B1(n_285),
.B2(n_281),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_306),
.A2(n_307),
.B1(n_308),
.B2(n_298),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_296),
.A2(n_270),
.B1(n_274),
.B2(n_277),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_290),
.A2(n_288),
.B1(n_287),
.B2(n_283),
.Y(n_308)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_309),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_297),
.B(n_5),
.Y(n_311)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_311),
.Y(n_321)
);

BUFx2_ASAP7_75t_L g312 ( 
.A(n_289),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_SL g322 ( 
.A1(n_312),
.A2(n_301),
.B1(n_293),
.B2(n_299),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_294),
.B(n_5),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_314),
.B(n_289),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_315),
.B(n_323),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_313),
.A2(n_302),
.B(n_300),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_317),
.A2(n_319),
.B(n_310),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_305),
.A2(n_303),
.B(n_292),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_320),
.B(n_307),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_322),
.Y(n_324)
);

BUFx24_ASAP7_75t_SL g323 ( 
.A(n_308),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_316),
.B(n_291),
.C(n_306),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_325),
.B(n_328),
.Y(n_332)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_327),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_321),
.B(n_312),
.Y(n_328)
);

INVxp33_ASAP7_75t_L g330 ( 
.A(n_329),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_324),
.A2(n_318),
.B(n_322),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_333),
.A2(n_310),
.B(n_326),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_334),
.A2(n_335),
.B(n_331),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_332),
.B(n_1),
.Y(n_335)
);

NOR3xp33_ASAP7_75t_SL g337 ( 
.A(n_336),
.B(n_330),
.C(n_3),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_2),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_2),
.C(n_4),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_339),
.A2(n_5),
.B(n_2),
.Y(n_340)
);

AOI21x1_ASAP7_75t_SL g341 ( 
.A1(n_340),
.A2(n_4),
.B(n_337),
.Y(n_341)
);


endmodule