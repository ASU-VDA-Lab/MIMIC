module fake_jpeg_13606_n_645 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_645);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_645;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_352;
wire n_350;
wire n_150;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_18),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_8),
.B(n_1),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_17),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_18),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_9),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_14),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_14),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_18),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_8),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_10),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_6),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_2),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_7),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_0),
.Y(n_61)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

INVx13_ASAP7_75t_L g150 ( 
.A(n_62),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_32),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_63),
.B(n_70),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_61),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_64),
.Y(n_153)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_26),
.Y(n_65)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_65),
.Y(n_167)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_66),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g132 ( 
.A(n_67),
.Y(n_132)
);

BUFx12_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

BUFx24_ASAP7_75t_L g208 ( 
.A(n_68),
.Y(n_208)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_69),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_32),
.B(n_9),
.Y(n_70)
);

BUFx12_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g177 ( 
.A(n_71),
.Y(n_177)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_28),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g161 ( 
.A(n_72),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_47),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_73),
.B(n_78),
.Y(n_147)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_35),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_74),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

INVx6_ASAP7_75t_L g184 ( 
.A(n_75),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_42),
.B(n_10),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_76),
.B(n_104),
.Y(n_137)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_77),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_47),
.Y(n_78)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_28),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_79),
.Y(n_135)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_24),
.Y(n_80)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_80),
.Y(n_191)
);

AND2x2_ASAP7_75t_SL g81 ( 
.A(n_23),
.B(n_0),
.Y(n_81)
);

AND2x2_ASAP7_75t_SL g164 ( 
.A(n_81),
.B(n_124),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_52),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_82),
.B(n_89),
.Y(n_154)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_21),
.Y(n_83)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_83),
.Y(n_141)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_26),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g179 ( 
.A(n_84),
.Y(n_179)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_31),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_85),
.Y(n_148)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_21),
.Y(n_86)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_86),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_87),
.Y(n_186)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g133 ( 
.A(n_88),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_58),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_37),
.Y(n_90)
);

INVx8_ASAP7_75t_L g159 ( 
.A(n_90),
.Y(n_159)
);

BUFx12_ASAP7_75t_L g91 ( 
.A(n_20),
.Y(n_91)
);

INVx6_ASAP7_75t_SL g188 ( 
.A(n_91),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_33),
.B(n_10),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_92),
.B(n_93),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_33),
.B(n_8),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_58),
.Y(n_94)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_94),
.Y(n_174)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_20),
.Y(n_95)
);

INVx11_ASAP7_75t_L g131 ( 
.A(n_95),
.Y(n_131)
);

BUFx2_ASAP7_75t_L g96 ( 
.A(n_31),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_96),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_40),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_97),
.B(n_100),
.Y(n_155)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_60),
.Y(n_98)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_98),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_37),
.Y(n_99)
);

INVx8_ASAP7_75t_L g176 ( 
.A(n_99),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_34),
.B(n_8),
.Y(n_100)
);

BUFx4f_ASAP7_75t_SL g101 ( 
.A(n_39),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g171 ( 
.A(n_101),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_23),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_102),
.Y(n_189)
);

BUFx5_ASAP7_75t_L g103 ( 
.A(n_39),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_103),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_40),
.B(n_11),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_41),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_105),
.B(n_108),
.Y(n_160)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_27),
.Y(n_106)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_106),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_51),
.A2(n_11),
.B1(n_2),
.B2(n_3),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_107),
.A2(n_59),
.B1(n_49),
.B2(n_48),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_34),
.B(n_43),
.Y(n_108)
);

BUFx12_ASAP7_75t_L g109 ( 
.A(n_55),
.Y(n_109)
);

BUFx12_ASAP7_75t_L g190 ( 
.A(n_109),
.Y(n_190)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_23),
.Y(n_110)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_110),
.Y(n_212)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_37),
.Y(n_111)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_111),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_45),
.Y(n_112)
);

INVx8_ASAP7_75t_L g205 ( 
.A(n_112),
.Y(n_205)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_41),
.Y(n_113)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_113),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_45),
.Y(n_114)
);

BUFx2_ASAP7_75t_L g145 ( 
.A(n_114),
.Y(n_145)
);

INVx3_ASAP7_75t_SL g115 ( 
.A(n_22),
.Y(n_115)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_115),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_46),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_116),
.B(n_125),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_29),
.Y(n_117)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_117),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_45),
.Y(n_118)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_118),
.Y(n_200)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_27),
.Y(n_119)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_119),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_56),
.Y(n_120)
);

INVx5_ASAP7_75t_L g213 ( 
.A(n_120),
.Y(n_213)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_60),
.Y(n_121)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_121),
.Y(n_210)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_30),
.Y(n_122)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_122),
.Y(n_216)
);

BUFx12f_ASAP7_75t_L g123 ( 
.A(n_53),
.Y(n_123)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_123),
.Y(n_138)
);

INVx2_ASAP7_75t_SL g124 ( 
.A(n_29),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_43),
.B(n_11),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_56),
.Y(n_126)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_126),
.Y(n_195)
);

INVx11_ASAP7_75t_L g127 ( 
.A(n_55),
.Y(n_127)
);

INVx11_ASAP7_75t_L g165 ( 
.A(n_127),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_56),
.Y(n_128)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_128),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_48),
.B(n_59),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_129),
.B(n_36),
.Y(n_175)
);

BUFx4f_ASAP7_75t_L g130 ( 
.A(n_29),
.Y(n_130)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_130),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_139),
.A2(n_44),
.B1(n_36),
.B2(n_179),
.Y(n_255)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_110),
.Y(n_143)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_143),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_65),
.B(n_49),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_144),
.B(n_158),
.Y(n_229)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_130),
.Y(n_149)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_149),
.Y(n_242)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_130),
.Y(n_156)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_156),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_71),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_157),
.B(n_170),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_84),
.B(n_38),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_106),
.B(n_38),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_162),
.B(n_183),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_66),
.A2(n_51),
.B1(n_46),
.B2(n_57),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_163),
.A2(n_178),
.B1(n_214),
.B2(n_25),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_96),
.A2(n_22),
.B1(n_25),
.B2(n_53),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_168),
.A2(n_115),
.B1(n_102),
.B2(n_117),
.Y(n_250)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_88),
.Y(n_169)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_169),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_71),
.Y(n_170)
);

INVx11_ASAP7_75t_L g172 ( 
.A(n_95),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_172),
.Y(n_272)
);

INVx11_ASAP7_75t_L g173 ( 
.A(n_127),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_173),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_175),
.B(n_193),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_104),
.A2(n_51),
.B1(n_57),
.B2(n_24),
.Y(n_178)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_67),
.Y(n_182)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_182),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_119),
.B(n_50),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_91),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_91),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_198),
.B(n_215),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_122),
.B(n_30),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_199),
.B(n_202),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_81),
.B(n_50),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_201),
.B(n_124),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_81),
.B(n_54),
.Y(n_202)
);

INVx11_ASAP7_75t_L g203 ( 
.A(n_62),
.Y(n_203)
);

CKINVDCx14_ASAP7_75t_R g262 ( 
.A(n_203),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_123),
.B(n_54),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_207),
.B(n_72),
.Y(n_254)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_123),
.Y(n_209)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_209),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_L g214 ( 
.A1(n_69),
.A2(n_57),
.B1(n_25),
.B2(n_22),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_109),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_164),
.B(n_83),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_217),
.B(n_239),
.C(n_274),
.Y(n_294)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_147),
.Y(n_218)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_218),
.Y(n_305)
);

INVx5_ASAP7_75t_L g219 ( 
.A(n_177),
.Y(n_219)
);

INVxp67_ASAP7_75t_SL g311 ( 
.A(n_219),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_L g220 ( 
.A1(n_214),
.A2(n_111),
.B1(n_121),
.B2(n_98),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_220),
.A2(n_244),
.B1(n_250),
.B2(n_251),
.Y(n_293)
);

INVx6_ASAP7_75t_L g221 ( 
.A(n_153),
.Y(n_221)
);

INVx6_ASAP7_75t_L g345 ( 
.A(n_221),
.Y(n_345)
);

INVx13_ASAP7_75t_L g222 ( 
.A(n_188),
.Y(n_222)
);

INVx13_ASAP7_75t_L g346 ( 
.A(n_222),
.Y(n_346)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_167),
.Y(n_224)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_224),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_153),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_225),
.Y(n_304)
);

INVx5_ASAP7_75t_L g226 ( 
.A(n_177),
.Y(n_226)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_226),
.Y(n_329)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_187),
.Y(n_228)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_228),
.Y(n_314)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_134),
.Y(n_230)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_230),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_160),
.B(n_77),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_234),
.B(n_240),
.Y(n_333)
);

INVx5_ASAP7_75t_L g235 ( 
.A(n_177),
.Y(n_235)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_235),
.Y(n_340)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_136),
.Y(n_236)
);

INVx4_ASAP7_75t_L g344 ( 
.A(n_236),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_137),
.A2(n_113),
.B1(n_74),
.B2(n_128),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_237),
.A2(n_245),
.B1(n_259),
.B2(n_268),
.Y(n_300)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_196),
.Y(n_238)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_238),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_164),
.B(n_86),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_154),
.Y(n_240)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_216),
.Y(n_243)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_243),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_L g244 ( 
.A1(n_163),
.A2(n_75),
.B1(n_87),
.B2(n_64),
.Y(n_244)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_136),
.Y(n_246)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_246),
.Y(n_325)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_149),
.Y(n_247)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_247),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_248),
.B(n_256),
.Y(n_298)
);

INVx4_ASAP7_75t_L g249 ( 
.A(n_156),
.Y(n_249)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_249),
.Y(n_307)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_135),
.A2(n_24),
.B1(n_80),
.B2(n_29),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_254),
.B(n_273),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_255),
.A2(n_279),
.B1(n_289),
.B2(n_292),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_155),
.B(n_94),
.Y(n_256)
);

BUFx3_ASAP7_75t_L g257 ( 
.A(n_132),
.Y(n_257)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_257),
.Y(n_318)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_141),
.Y(n_258)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_258),
.Y(n_342)
);

OAI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_168),
.A2(n_126),
.B1(n_120),
.B2(n_118),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_184),
.Y(n_260)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_260),
.Y(n_319)
);

INVx5_ASAP7_75t_L g261 ( 
.A(n_132),
.Y(n_261)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_261),
.Y(n_320)
);

OR2x2_ASAP7_75t_SL g263 ( 
.A(n_151),
.B(n_140),
.Y(n_263)
);

NAND2x1_ASAP7_75t_SL g316 ( 
.A(n_263),
.B(n_281),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_166),
.B(n_179),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_264),
.B(n_283),
.Y(n_303)
);

BUFx12f_ASAP7_75t_L g265 ( 
.A(n_189),
.Y(n_265)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_265),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_142),
.A2(n_44),
.B1(n_114),
.B2(n_112),
.Y(n_266)
);

OAI21xp33_ASAP7_75t_L g335 ( 
.A1(n_266),
.A2(n_280),
.B(n_208),
.Y(n_335)
);

INVx4_ASAP7_75t_L g267 ( 
.A(n_203),
.Y(n_267)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_267),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_184),
.A2(n_90),
.B1(n_99),
.B2(n_109),
.Y(n_268)
);

INVx8_ASAP7_75t_L g271 ( 
.A(n_186),
.Y(n_271)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_271),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_190),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_174),
.B(n_103),
.Y(n_274)
);

INVx5_ASAP7_75t_L g276 ( 
.A(n_132),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_276),
.B(n_277),
.Y(n_324)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_180),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_186),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_278),
.B(n_282),
.Y(n_343)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_135),
.A2(n_101),
.B1(n_85),
.B2(n_79),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_148),
.A2(n_101),
.B1(n_68),
.B2(n_4),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_171),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_190),
.Y(n_282)
);

INVx6_ASAP7_75t_L g283 ( 
.A(n_159),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_192),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_284),
.B(n_286),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g285 ( 
.A(n_194),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_285),
.Y(n_302)
);

INVx8_ASAP7_75t_L g286 ( 
.A(n_181),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_210),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_287),
.B(n_288),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_212),
.B(n_12),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_L g289 ( 
.A1(n_145),
.A2(n_204),
.B1(n_195),
.B2(n_205),
.Y(n_289)
);

INVx4_ASAP7_75t_SL g290 ( 
.A(n_208),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_290),
.B(n_291),
.Y(n_317)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_143),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_L g292 ( 
.A1(n_145),
.A2(n_12),
.B1(n_2),
.B2(n_4),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_255),
.A2(n_181),
.B1(n_211),
.B2(n_206),
.Y(n_295)
);

OA21x2_ASAP7_75t_L g361 ( 
.A1(n_295),
.A2(n_332),
.B(n_334),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_217),
.B(n_191),
.C(n_182),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_297),
.B(n_327),
.C(n_347),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_233),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_299),
.B(n_309),
.Y(n_366)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_250),
.A2(n_173),
.B(n_172),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g368 ( 
.A1(n_301),
.A2(n_226),
.B(n_219),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_231),
.B(n_204),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_306),
.B(n_310),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_281),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_229),
.B(n_195),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_237),
.A2(n_211),
.B1(n_206),
.B2(n_176),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_322),
.A2(n_300),
.B1(n_310),
.B2(n_306),
.Y(n_377)
);

AO22x1_ASAP7_75t_SL g326 ( 
.A1(n_217),
.A2(n_131),
.B1(n_165),
.B2(n_208),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_326),
.B(n_328),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_239),
.B(n_131),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_239),
.B(n_252),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_230),
.B(n_263),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_330),
.B(n_339),
.Y(n_388)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_274),
.B(n_290),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_331),
.B(n_335),
.Y(n_389)
);

OA22x2_ASAP7_75t_L g332 ( 
.A1(n_266),
.A2(n_165),
.B1(n_176),
.B2(n_205),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_251),
.A2(n_159),
.B1(n_200),
.B2(n_213),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_227),
.B(n_213),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_274),
.B(n_169),
.C(n_133),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_280),
.B(n_190),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_348),
.B(n_241),
.C(n_269),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_222),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_349),
.B(n_235),
.Y(n_371)
);

OAI22xp33_ASAP7_75t_SL g350 ( 
.A1(n_279),
.A2(n_197),
.B1(n_148),
.B2(n_133),
.Y(n_350)
);

OAI22xp33_ASAP7_75t_SL g355 ( 
.A1(n_350),
.A2(n_185),
.B1(n_272),
.B2(n_267),
.Y(n_355)
);

AOI32xp33_ASAP7_75t_L g352 ( 
.A1(n_272),
.A2(n_265),
.A3(n_253),
.B1(n_223),
.B2(n_197),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_SL g364 ( 
.A1(n_352),
.A2(n_331),
.B(n_301),
.Y(n_364)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_296),
.Y(n_353)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_353),
.Y(n_402)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_296),
.Y(n_354)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_354),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_355),
.A2(n_377),
.B1(n_392),
.B2(n_293),
.Y(n_400)
);

INVx13_ASAP7_75t_L g356 ( 
.A(n_346),
.Y(n_356)
);

INVx1_ASAP7_75t_SL g423 ( 
.A(n_356),
.Y(n_423)
);

INVx13_ASAP7_75t_L g357 ( 
.A(n_346),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_357),
.Y(n_407)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_342),
.Y(n_358)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_358),
.Y(n_413)
);

NAND3xp33_ASAP7_75t_L g359 ( 
.A(n_298),
.B(n_262),
.C(n_275),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_SL g429 ( 
.A(n_359),
.B(n_380),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_343),
.Y(n_360)
);

OAI21xp33_ASAP7_75t_L g415 ( 
.A1(n_360),
.A2(n_362),
.B(n_370),
.Y(n_415)
);

CKINVDCx14_ASAP7_75t_R g362 ( 
.A(n_331),
.Y(n_362)
);

INVx8_ASAP7_75t_L g363 ( 
.A(n_304),
.Y(n_363)
);

INVx4_ASAP7_75t_L g425 ( 
.A(n_363),
.Y(n_425)
);

INVxp67_ASAP7_75t_L g438 ( 
.A(n_364),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_330),
.B(n_241),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_365),
.B(n_371),
.Y(n_409)
);

AND2x6_ASAP7_75t_L g367 ( 
.A(n_316),
.B(n_150),
.Y(n_367)
);

AOI32xp33_ASAP7_75t_L g435 ( 
.A1(n_367),
.A2(n_373),
.A3(n_378),
.B1(n_394),
.B2(n_265),
.Y(n_435)
);

AOI21xp5_ASAP7_75t_L g434 ( 
.A1(n_368),
.A2(n_276),
.B(n_320),
.Y(n_434)
);

NOR2x1_ASAP7_75t_R g370 ( 
.A(n_294),
.B(n_275),
.Y(n_370)
);

AOI22xp33_ASAP7_75t_SL g372 ( 
.A1(n_334),
.A2(n_283),
.B1(n_185),
.B2(n_270),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_L g428 ( 
.A1(n_372),
.A2(n_317),
.B(n_347),
.Y(n_428)
);

AND2x6_ASAP7_75t_L g373 ( 
.A(n_316),
.B(n_150),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_317),
.Y(n_374)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_374),
.Y(n_427)
);

INVx13_ASAP7_75t_L g375 ( 
.A(n_311),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_375),
.Y(n_417)
);

INVx13_ASAP7_75t_L g376 ( 
.A(n_329),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_376),
.Y(n_419)
);

AND2x6_ASAP7_75t_L g378 ( 
.A(n_326),
.B(n_161),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_314),
.Y(n_379)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_379),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_305),
.B(n_232),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_333),
.B(n_232),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_382),
.B(n_383),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_303),
.B(n_270),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_315),
.Y(n_384)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_384),
.Y(n_410)
);

BUFx3_ASAP7_75t_L g385 ( 
.A(n_329),
.Y(n_385)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_385),
.Y(n_421)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_321),
.Y(n_386)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_386),
.Y(n_416)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_325),
.Y(n_390)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_390),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_391),
.B(n_393),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_300),
.A2(n_200),
.B1(n_278),
.B2(n_260),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_348),
.B(n_242),
.Y(n_393)
);

AND2x6_ASAP7_75t_L g394 ( 
.A(n_326),
.B(n_261),
.Y(n_394)
);

INVx13_ASAP7_75t_L g395 ( 
.A(n_340),
.Y(n_395)
);

AO21x2_ASAP7_75t_L g408 ( 
.A1(n_395),
.A2(n_351),
.B(n_340),
.Y(n_408)
);

NAND3xp33_ASAP7_75t_L g396 ( 
.A(n_313),
.B(n_242),
.C(n_269),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_396),
.B(n_398),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_312),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_397),
.B(n_341),
.Y(n_411)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_319),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_336),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_399),
.B(n_366),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_400),
.A2(n_403),
.B1(n_405),
.B2(n_420),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_377),
.A2(n_337),
.B1(n_295),
.B2(n_335),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_369),
.B(n_294),
.C(n_388),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_404),
.B(n_414),
.C(n_433),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_361),
.A2(n_392),
.B1(n_387),
.B2(n_381),
.Y(n_405)
);

A2O1A1Ixp33_ASAP7_75t_SL g462 ( 
.A1(n_408),
.A2(n_434),
.B(n_356),
.C(n_375),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_SL g463 ( 
.A(n_411),
.B(n_399),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_369),
.B(n_328),
.Y(n_414)
);

AOI22xp33_ASAP7_75t_L g420 ( 
.A1(n_397),
.A2(n_332),
.B1(n_308),
.B2(n_317),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_387),
.A2(n_322),
.B1(n_297),
.B2(n_332),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_422),
.B(n_426),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_381),
.B(n_327),
.Y(n_426)
);

INVxp67_ASAP7_75t_L g454 ( 
.A(n_428),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_360),
.B(n_339),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_430),
.B(n_436),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_361),
.A2(n_332),
.B1(n_345),
.B2(n_319),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_431),
.A2(n_400),
.B1(n_403),
.B2(n_405),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_388),
.B(n_324),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_SL g457 ( 
.A1(n_435),
.A2(n_357),
.B(n_356),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_361),
.A2(n_271),
.B1(n_286),
.B2(n_221),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_437),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_439),
.A2(n_447),
.B1(n_453),
.B2(n_464),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_R g440 ( 
.A(n_415),
.B(n_373),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_440),
.B(n_457),
.Y(n_491)
);

AOI21xp5_ASAP7_75t_L g442 ( 
.A1(n_438),
.A2(n_368),
.B(n_364),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_L g480 ( 
.A1(n_442),
.A2(n_444),
.B(n_462),
.Y(n_480)
);

O2A1O1Ixp33_ASAP7_75t_L g444 ( 
.A1(n_438),
.A2(n_394),
.B(n_389),
.C(n_378),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_401),
.Y(n_445)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_445),
.Y(n_484)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_401),
.Y(n_446)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_446),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_431),
.A2(n_361),
.B1(n_365),
.B2(n_391),
.Y(n_447)
);

OAI21xp5_ASAP7_75t_L g448 ( 
.A1(n_434),
.A2(n_389),
.B(n_374),
.Y(n_448)
);

AO21x1_ASAP7_75t_L g485 ( 
.A1(n_448),
.A2(n_451),
.B(n_452),
.Y(n_485)
);

OAI32xp33_ASAP7_75t_L g449 ( 
.A1(n_426),
.A2(n_370),
.A3(n_367),
.B1(n_358),
.B2(n_379),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_449),
.B(n_456),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_428),
.B(n_389),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_427),
.B(n_393),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_404),
.A2(n_393),
.B1(n_386),
.B2(n_384),
.Y(n_453)
);

AND2x6_ASAP7_75t_L g456 ( 
.A(n_414),
.B(n_357),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_433),
.B(n_390),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_459),
.B(n_472),
.C(n_307),
.Y(n_498)
);

CKINVDCx16_ASAP7_75t_R g460 ( 
.A(n_430),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_460),
.B(n_423),
.Y(n_483)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_410),
.Y(n_461)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_461),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_SL g478 ( 
.A(n_463),
.B(n_471),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_L g464 ( 
.A1(n_436),
.A2(n_363),
.B1(n_345),
.B2(n_304),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_410),
.Y(n_465)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_465),
.Y(n_488)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_416),
.Y(n_466)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_466),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_422),
.A2(n_363),
.B1(n_398),
.B2(n_354),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_467),
.A2(n_419),
.B1(n_416),
.B2(n_418),
.Y(n_477)
);

AOI21xp5_ASAP7_75t_SL g468 ( 
.A1(n_432),
.A2(n_409),
.B(n_429),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_L g494 ( 
.A1(n_468),
.A2(n_408),
.B(n_320),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_424),
.B(n_417),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_469),
.Y(n_490)
);

INVx13_ASAP7_75t_L g470 ( 
.A(n_423),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_470),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_411),
.B(n_302),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_406),
.B(n_353),
.C(n_323),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_413),
.B(n_385),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_SL g508 ( 
.A(n_473),
.B(n_236),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_402),
.B(n_344),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_474),
.B(n_338),
.Y(n_503)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_455),
.B(n_406),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g520 ( 
.A(n_476),
.B(n_479),
.Y(n_520)
);

OAI22xp5_ASAP7_75t_L g513 ( 
.A1(n_477),
.A2(n_450),
.B1(n_466),
.B2(n_465),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_SL g479 ( 
.A(n_455),
.B(n_418),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_439),
.A2(n_425),
.B1(n_412),
.B2(n_421),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_SL g511 ( 
.A1(n_482),
.A2(n_487),
.B1(n_495),
.B2(n_507),
.Y(n_511)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_483),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_441),
.A2(n_425),
.B1(n_421),
.B2(n_408),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_443),
.A2(n_408),
.B1(n_407),
.B2(n_225),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_489),
.A2(n_499),
.B1(n_464),
.B2(n_484),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_459),
.B(n_307),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g533 ( 
.A(n_492),
.B(n_493),
.Y(n_533)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_453),
.B(n_407),
.Y(n_493)
);

AOI21xp33_ASAP7_75t_L g528 ( 
.A1(n_494),
.A2(n_462),
.B(n_452),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_447),
.A2(n_408),
.B1(n_323),
.B2(n_318),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_469),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_497),
.B(n_508),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_498),
.B(n_500),
.C(n_506),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_443),
.A2(n_318),
.B1(n_338),
.B2(n_344),
.Y(n_499)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_449),
.B(n_395),
.Y(n_500)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_503),
.Y(n_512)
);

MAJx2_ASAP7_75t_L g504 ( 
.A(n_451),
.B(n_375),
.C(n_395),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_504),
.B(n_448),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_469),
.B(n_0),
.Y(n_505)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_505),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_472),
.B(n_376),
.C(n_249),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_467),
.A2(n_376),
.B1(n_146),
.B2(n_257),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_SL g545 ( 
.A(n_510),
.B(n_492),
.Y(n_545)
);

AOI22xp5_ASAP7_75t_L g563 ( 
.A1(n_513),
.A2(n_138),
.B1(n_0),
.B2(n_6),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_490),
.B(n_450),
.Y(n_514)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_514),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_480),
.B(n_444),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_515),
.B(n_526),
.Y(n_559)
);

HB1xp67_ASAP7_75t_L g516 ( 
.A(n_494),
.Y(n_516)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_516),
.Y(n_542)
);

OAI22xp5_ASAP7_75t_L g517 ( 
.A1(n_475),
.A2(n_458),
.B1(n_463),
.B2(n_440),
.Y(n_517)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_517),
.Y(n_551)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_503),
.Y(n_518)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_518),
.Y(n_558)
);

OAI22xp5_ASAP7_75t_L g553 ( 
.A1(n_522),
.A2(n_534),
.B1(n_487),
.B2(n_507),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_476),
.B(n_452),
.C(n_454),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_523),
.B(n_479),
.C(n_506),
.Y(n_539)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_481),
.Y(n_524)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_524),
.Y(n_561)
);

OAI22xp5_ASAP7_75t_SL g525 ( 
.A1(n_475),
.A2(n_454),
.B1(n_442),
.B2(n_456),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_L g541 ( 
.A1(n_525),
.A2(n_532),
.B1(n_536),
.B2(n_489),
.Y(n_541)
);

AOI21xp5_ASAP7_75t_SL g526 ( 
.A1(n_480),
.A2(n_457),
.B(n_451),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_481),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_527),
.B(n_529),
.Y(n_556)
);

HB1xp67_ASAP7_75t_L g543 ( 
.A(n_528),
.Y(n_543)
);

OAI21xp5_ASAP7_75t_L g529 ( 
.A1(n_502),
.A2(n_491),
.B(n_485),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_478),
.B(n_458),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_531),
.B(n_538),
.Y(n_562)
);

OAI22xp5_ASAP7_75t_SL g532 ( 
.A1(n_495),
.A2(n_468),
.B1(n_461),
.B2(n_446),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g534 ( 
.A1(n_500),
.A2(n_445),
.B1(n_462),
.B2(n_474),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_477),
.B(n_462),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g555 ( 
.A(n_535),
.Y(n_555)
);

OAI22xp5_ASAP7_75t_SL g536 ( 
.A1(n_502),
.A2(n_462),
.B1(n_470),
.B2(n_146),
.Y(n_536)
);

OAI21xp5_ASAP7_75t_SL g537 ( 
.A1(n_485),
.A2(n_152),
.B(n_189),
.Y(n_537)
);

INVxp33_ASAP7_75t_L g554 ( 
.A(n_537),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_498),
.B(n_152),
.Y(n_538)
);

XNOR2xp5_ASAP7_75t_L g574 ( 
.A(n_539),
.B(n_544),
.Y(n_574)
);

INVxp67_ASAP7_75t_L g580 ( 
.A(n_541),
.Y(n_580)
);

XNOR2xp5_ASAP7_75t_L g544 ( 
.A(n_519),
.B(n_493),
.Y(n_544)
);

XNOR2xp5_ASAP7_75t_SL g579 ( 
.A(n_545),
.B(n_547),
.Y(n_579)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_519),
.B(n_504),
.C(n_499),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_546),
.B(n_550),
.Y(n_571)
);

XOR2xp5_ASAP7_75t_L g547 ( 
.A(n_523),
.B(n_482),
.Y(n_547)
);

BUFx6f_ASAP7_75t_L g548 ( 
.A(n_509),
.Y(n_548)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_548),
.Y(n_564)
);

AOI22xp33_ASAP7_75t_SL g549 ( 
.A1(n_511),
.A2(n_496),
.B1(n_486),
.B2(n_501),
.Y(n_549)
);

CKINVDCx16_ASAP7_75t_R g582 ( 
.A(n_549),
.Y(n_582)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_520),
.B(n_501),
.C(n_488),
.Y(n_550)
);

XOR2xp5_ASAP7_75t_L g552 ( 
.A(n_520),
.B(n_533),
.Y(n_552)
);

XOR2xp5_ASAP7_75t_L g566 ( 
.A(n_552),
.B(n_533),
.Y(n_566)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_553),
.Y(n_572)
);

AOI22xp5_ASAP7_75t_L g557 ( 
.A1(n_511),
.A2(n_488),
.B1(n_486),
.B2(n_505),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_557),
.B(n_560),
.Y(n_570)
);

OAI22xp5_ASAP7_75t_L g560 ( 
.A1(n_522),
.A2(n_209),
.B1(n_138),
.B2(n_6),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_563),
.B(n_532),
.Y(n_573)
);

INVx13_ASAP7_75t_L g565 ( 
.A(n_540),
.Y(n_565)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_565),
.Y(n_592)
);

XNOR2xp5_ASAP7_75t_SL g590 ( 
.A(n_566),
.B(n_561),
.Y(n_590)
);

AOI321xp33_ASAP7_75t_L g567 ( 
.A1(n_556),
.A2(n_529),
.A3(n_530),
.B1(n_526),
.B2(n_515),
.C(n_514),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_567),
.B(n_568),
.Y(n_602)
);

MAJIxp5_ASAP7_75t_L g568 ( 
.A(n_550),
.B(n_525),
.C(n_515),
.Y(n_568)
);

OAI21xp5_ASAP7_75t_SL g569 ( 
.A1(n_559),
.A2(n_535),
.B(n_534),
.Y(n_569)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_569),
.Y(n_596)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_573),
.Y(n_600)
);

XNOR2xp5_ASAP7_75t_L g575 ( 
.A(n_547),
.B(n_546),
.Y(n_575)
);

XNOR2xp5_ASAP7_75t_L g586 ( 
.A(n_575),
.B(n_577),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_SL g576 ( 
.A(n_562),
.B(n_521),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_SL g598 ( 
.A(n_576),
.B(n_578),
.Y(n_598)
);

XOR2xp5_ASAP7_75t_L g577 ( 
.A(n_544),
.B(n_510),
.Y(n_577)
);

CKINVDCx20_ASAP7_75t_R g578 ( 
.A(n_556),
.Y(n_578)
);

MAJIxp5_ASAP7_75t_L g581 ( 
.A(n_539),
.B(n_552),
.C(n_543),
.Y(n_581)
);

MAJIxp5_ASAP7_75t_L g588 ( 
.A(n_581),
.B(n_558),
.C(n_541),
.Y(n_588)
);

OAI21xp5_ASAP7_75t_L g583 ( 
.A1(n_559),
.A2(n_536),
.B(n_518),
.Y(n_583)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_583),
.Y(n_601)
);

XOR2xp5_ASAP7_75t_L g584 ( 
.A(n_545),
.B(n_559),
.Y(n_584)
);

XOR2xp5_ASAP7_75t_L g597 ( 
.A(n_584),
.B(n_563),
.Y(n_597)
);

AOI22xp5_ASAP7_75t_SL g585 ( 
.A1(n_580),
.A2(n_554),
.B1(n_551),
.B2(n_555),
.Y(n_585)
);

OAI22xp5_ASAP7_75t_SL g606 ( 
.A1(n_585),
.A2(n_583),
.B1(n_580),
.B2(n_568),
.Y(n_606)
);

OAI21xp5_ASAP7_75t_SL g587 ( 
.A1(n_571),
.A2(n_554),
.B(n_542),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_587),
.B(n_588),
.Y(n_611)
);

MAJIxp5_ASAP7_75t_L g589 ( 
.A(n_575),
.B(n_557),
.C(n_512),
.Y(n_589)
);

MAJIxp5_ASAP7_75t_L g612 ( 
.A(n_589),
.B(n_594),
.C(n_579),
.Y(n_612)
);

XNOR2xp5_ASAP7_75t_SL g605 ( 
.A(n_590),
.B(n_597),
.Y(n_605)
);

BUFx3_ASAP7_75t_L g591 ( 
.A(n_572),
.Y(n_591)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_591),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_564),
.B(n_548),
.Y(n_593)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_593),
.Y(n_607)
);

MAJIxp5_ASAP7_75t_L g594 ( 
.A(n_574),
.B(n_537),
.C(n_527),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_582),
.B(n_574),
.Y(n_595)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_595),
.Y(n_616)
);

XNOR2xp5_ASAP7_75t_SL g599 ( 
.A(n_579),
.B(n_524),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_599),
.B(n_584),
.Y(n_603)
);

OAI21x1_ASAP7_75t_L g619 ( 
.A1(n_603),
.A2(n_586),
.B(n_599),
.Y(n_619)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_606),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_592),
.B(n_573),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_608),
.B(n_609),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_600),
.B(n_588),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_598),
.B(n_581),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_610),
.B(n_613),
.Y(n_620)
);

OR2x2_ASAP7_75t_L g621 ( 
.A(n_612),
.B(n_614),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_602),
.B(n_570),
.Y(n_613)
);

OAI22xp5_ASAP7_75t_SL g614 ( 
.A1(n_585),
.A2(n_570),
.B1(n_567),
.B2(n_569),
.Y(n_614)
);

NOR5xp2_ASAP7_75t_L g615 ( 
.A(n_590),
.B(n_565),
.C(n_577),
.D(n_566),
.E(n_14),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_615),
.Y(n_623)
);

MAJx2_ASAP7_75t_L g617 ( 
.A(n_611),
.B(n_586),
.C(n_594),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_SL g628 ( 
.A(n_617),
.B(n_622),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_619),
.B(n_624),
.Y(n_630)
);

O2A1O1Ixp33_ASAP7_75t_SL g622 ( 
.A1(n_614),
.A2(n_601),
.B(n_596),
.C(n_591),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_607),
.B(n_589),
.Y(n_624)
);

AOI21xp5_ASAP7_75t_SL g625 ( 
.A1(n_616),
.A2(n_597),
.B(n_7),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_625),
.B(n_604),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_609),
.B(n_2),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_626),
.B(n_7),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_629),
.B(n_631),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_620),
.B(n_608),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_632),
.B(n_634),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_618),
.B(n_606),
.Y(n_633)
);

AOI21xp5_ASAP7_75t_L g638 ( 
.A1(n_633),
.A2(n_621),
.B(n_618),
.Y(n_638)
);

AOI322xp5_ASAP7_75t_L g634 ( 
.A1(n_627),
.A2(n_612),
.A3(n_605),
.B1(n_68),
.B2(n_15),
.C1(n_7),
.C2(n_17),
.Y(n_634)
);

INVxp33_ASAP7_75t_L g636 ( 
.A(n_630),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_636),
.B(n_638),
.Y(n_640)
);

OAI22x1_ASAP7_75t_L g639 ( 
.A1(n_637),
.A2(n_623),
.B1(n_628),
.B2(n_633),
.Y(n_639)
);

OAI21xp5_ASAP7_75t_SL g641 ( 
.A1(n_639),
.A2(n_635),
.B(n_605),
.Y(n_641)
);

OAI21xp5_ASAP7_75t_SL g642 ( 
.A1(n_641),
.A2(n_640),
.B(n_14),
.Y(n_642)
);

MAJIxp5_ASAP7_75t_L g643 ( 
.A(n_642),
.B(n_11),
.C(n_15),
.Y(n_643)
);

BUFx24_ASAP7_75t_SL g644 ( 
.A(n_643),
.Y(n_644)
);

O2A1O1Ixp5_ASAP7_75t_L g645 ( 
.A1(n_644),
.A2(n_16),
.B(n_17),
.C(n_638),
.Y(n_645)
);


endmodule