module real_jpeg_10966_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_43;
wire n_37;
wire n_21;
wire n_35;
wire n_33;
wire n_38;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_44;
wire n_46;
wire n_23;
wire n_11;
wire n_14;
wire n_47;
wire n_45;
wire n_25;
wire n_42;
wire n_7;
wire n_22;
wire n_18;
wire n_39;
wire n_40;
wire n_36;
wire n_41;
wire n_27;
wire n_32;
wire n_20;
wire n_19;
wire n_26;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

OR2x2_ASAP7_75t_SL g30 ( 
.A(n_1),
.B(n_31),
.Y(n_30)
);

OR2x2_ASAP7_75t_SL g38 ( 
.A(n_1),
.B(n_3),
.Y(n_38)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_2),
.B(n_4),
.Y(n_14)
);

OR2x2_ASAP7_75t_L g19 ( 
.A(n_3),
.B(n_20),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

OA21x2_ASAP7_75t_L g23 ( 
.A1(n_5),
.A2(n_10),
.B(n_14),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g6 ( 
.A(n_7),
.Y(n_6)
);

OAI211xp5_ASAP7_75t_L g7 ( 
.A1(n_8),
.A2(n_15),
.B(n_21),
.C(n_41),
.Y(n_7)
);

AOI221xp5_ASAP7_75t_L g21 ( 
.A1(n_8),
.A2(n_22),
.B1(n_24),
.B2(n_27),
.C(n_32),
.Y(n_21)
);

OA21x2_ASAP7_75t_L g8 ( 
.A1(n_9),
.A2(n_10),
.B(n_14),
.Y(n_8)
);

AO21x1_ASAP7_75t_L g34 ( 
.A1(n_9),
.A2(n_17),
.B(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_9),
.B(n_17),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_9),
.B(n_18),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g10 ( 
.A(n_11),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_13),
.Y(n_11)
);

AOI221xp5_ASAP7_75t_L g41 ( 
.A1(n_12),
.A2(n_23),
.B1(n_42),
.B2(n_43),
.C(n_45),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_12),
.B(n_18),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g15 ( 
.A(n_16),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_19),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_17),
.B(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_17),
.B(n_29),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_SL g36 ( 
.A1(n_17),
.A2(n_37),
.B(n_39),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_17),
.B(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_17),
.B(n_30),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_18),
.Y(n_17)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

OR2x2_ASAP7_75t_SL g40 ( 
.A(n_20),
.B(n_31),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_36),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_46),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_44),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);


endmodule