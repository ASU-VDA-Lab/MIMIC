module fake_jpeg_8314_n_319 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_319);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_319;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_292;
wire n_213;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx8_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx6f_ASAP7_75t_SL g32 ( 
.A(n_9),
.Y(n_32)
);

INVx11_ASAP7_75t_SL g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_32),
.Y(n_34)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_42),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_28),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_38),
.B(n_43),
.Y(n_51)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_17),
.B(n_0),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_43),
.A2(n_20),
.B1(n_29),
.B2(n_19),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_44),
.A2(n_46),
.B1(n_58),
.B2(n_20),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_43),
.A2(n_29),
.B1(n_20),
.B2(n_19),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_22),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_52),
.B(n_64),
.Y(n_84)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

AOI21xp33_ASAP7_75t_L g57 ( 
.A1(n_38),
.A2(n_21),
.B(n_22),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_57),
.A2(n_16),
.B(n_18),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_35),
.A2(n_20),
.B1(n_29),
.B2(n_19),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_38),
.B(n_21),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_43),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_66),
.A2(n_37),
.B(n_18),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_67),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_48),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_69),
.B(n_71),
.Y(n_116)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_49),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_73),
.B(n_82),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_76),
.A2(n_78),
.B1(n_86),
.B2(n_36),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_47),
.A2(n_36),
.B1(n_31),
.B2(n_24),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_80),
.B(n_30),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_81),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_49),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_44),
.B(n_41),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_91),
.Y(n_94)
);

NOR3xp33_ASAP7_75t_L g85 ( 
.A(n_49),
.B(n_23),
.C(n_27),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_85),
.B(n_90),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_47),
.A2(n_36),
.B1(n_31),
.B2(n_24),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

AOI21xp33_ASAP7_75t_L g89 ( 
.A1(n_54),
.A2(n_23),
.B(n_27),
.Y(n_89)
);

NAND3xp33_ASAP7_75t_L g112 ( 
.A(n_89),
.B(n_8),
.C(n_15),
.Y(n_112)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_53),
.B(n_41),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_55),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_92),
.A2(n_42),
.B1(n_39),
.B2(n_34),
.Y(n_107)
);

OA22x2_ASAP7_75t_L g93 ( 
.A1(n_55),
.A2(n_39),
.B1(n_34),
.B2(n_36),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_93),
.A2(n_65),
.B1(n_62),
.B2(n_60),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_84),
.B(n_23),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_95),
.B(n_112),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_83),
.B(n_37),
.C(n_39),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_96),
.B(n_40),
.C(n_41),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_98),
.A2(n_118),
.B1(n_68),
.B2(n_88),
.Y(n_141)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_91),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_99),
.B(n_101),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_80),
.B(n_45),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_100),
.B(n_111),
.Y(n_143)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_87),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_93),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_102),
.B(n_103),
.Y(n_136)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_93),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_87),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_104),
.B(n_110),
.Y(n_142)
);

XNOR2x1_ASAP7_75t_SL g147 ( 
.A(n_105),
.B(n_113),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_107),
.A2(n_109),
.B1(n_114),
.B2(n_74),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_81),
.A2(n_39),
.B1(n_42),
.B2(n_34),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_93),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_66),
.B(n_41),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_66),
.A2(n_42),
.B1(n_61),
.B2(n_18),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_115),
.A2(n_72),
.B1(n_42),
.B2(n_79),
.Y(n_126)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_90),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_87),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_119),
.B(n_88),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_116),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_121),
.B(n_123),
.Y(n_155)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_114),
.Y(n_123)
);

BUFx2_ASAP7_75t_L g124 ( 
.A(n_108),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_124),
.Y(n_170)
);

OAI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_102),
.A2(n_53),
.B1(n_75),
.B2(n_77),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_125),
.A2(n_126),
.B1(n_127),
.B2(n_128),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_103),
.A2(n_72),
.B1(n_61),
.B2(n_71),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_110),
.A2(n_75),
.B1(n_77),
.B2(n_74),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_130),
.B(n_133),
.C(n_144),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_105),
.A2(n_24),
.B(n_16),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_131),
.A2(n_140),
.B(n_30),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_132),
.B(n_137),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_97),
.A2(n_70),
.B1(n_41),
.B2(n_40),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_133),
.A2(n_134),
.B1(n_135),
.B2(n_144),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_97),
.A2(n_70),
.B1(n_40),
.B2(n_16),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_94),
.A2(n_40),
.B1(n_31),
.B2(n_67),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_95),
.Y(n_137)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_138),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_120),
.Y(n_139)
);

INVx13_ASAP7_75t_L g181 ( 
.A(n_139),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_94),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_141),
.A2(n_150),
.B1(n_118),
.B2(n_106),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_111),
.A2(n_68),
.B1(n_26),
.B2(n_17),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_100),
.B(n_28),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_145),
.B(n_146),
.Y(n_153)
);

OR2x2_ASAP7_75t_L g146 ( 
.A(n_117),
.B(n_0),
.Y(n_146)
);

OR2x2_ASAP7_75t_L g148 ( 
.A(n_100),
.B(n_0),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_148),
.B(n_149),
.Y(n_157)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_115),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_109),
.A2(n_26),
.B1(n_17),
.B2(n_28),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_138),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_151),
.B(n_160),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_147),
.B(n_113),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_154),
.B(n_158),
.C(n_161),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_123),
.B(n_96),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_156),
.A2(n_172),
.B(n_173),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_140),
.B(n_99),
.Y(n_159)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_159),
.Y(n_198)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_122),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_143),
.B(n_106),
.C(n_119),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_122),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_163),
.B(n_171),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_164),
.A2(n_124),
.B1(n_8),
.B2(n_10),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_148),
.B(n_120),
.Y(n_165)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_165),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_149),
.A2(n_107),
.B1(n_104),
.B2(n_101),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_167),
.A2(n_169),
.B1(n_175),
.B2(n_180),
.Y(n_185)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_142),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_168),
.B(n_178),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_132),
.A2(n_26),
.B1(n_25),
.B2(n_30),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_143),
.A2(n_30),
.B(n_25),
.Y(n_172)
);

OAI21xp33_ASAP7_75t_L g173 ( 
.A1(n_145),
.A2(n_147),
.B(n_148),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_131),
.A2(n_30),
.B(n_25),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_174),
.A2(n_176),
.B(n_121),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_136),
.A2(n_142),
.B1(n_130),
.B2(n_150),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_131),
.A2(n_33),
.B(n_26),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_136),
.B(n_108),
.C(n_33),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_177),
.B(n_108),
.Y(n_199)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_128),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_124),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_179),
.B(n_127),
.Y(n_191)
);

AO22x1_ASAP7_75t_SL g180 ( 
.A1(n_126),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_180)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_159),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_184),
.B(n_201),
.Y(n_220)
);

AND2x4_ASAP7_75t_L g187 ( 
.A(n_151),
.B(n_135),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_187),
.A2(n_193),
.B(n_203),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_153),
.B(n_137),
.Y(n_188)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_188),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_189),
.B(n_190),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_167),
.Y(n_190)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_191),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_157),
.A2(n_129),
.B(n_146),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_182),
.A2(n_134),
.B1(n_146),
.B2(n_129),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_194),
.A2(n_169),
.B1(n_171),
.B2(n_164),
.Y(n_227)
);

OAI32xp33_ASAP7_75t_L g197 ( 
.A1(n_157),
.A2(n_9),
.A3(n_15),
.B1(n_14),
.B2(n_12),
.Y(n_197)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_197),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_199),
.B(n_210),
.C(n_174),
.Y(n_219)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_200),
.Y(n_214)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_155),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_154),
.B(n_7),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_202),
.B(n_176),
.Y(n_225)
);

OA21x2_ASAP7_75t_L g203 ( 
.A1(n_180),
.A2(n_1),
.B(n_2),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_180),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_204),
.B(n_206),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_153),
.B(n_1),
.Y(n_205)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_205),
.Y(n_224)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_177),
.Y(n_206)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_152),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_208),
.B(n_156),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_170),
.B(n_5),
.Y(n_209)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_209),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_161),
.B(n_5),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_190),
.A2(n_152),
.B1(n_162),
.B2(n_158),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_216),
.A2(n_218),
.B1(n_226),
.B2(n_231),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_186),
.A2(n_162),
.B1(n_181),
.B2(n_166),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_219),
.B(n_221),
.C(n_229),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_196),
.B(n_175),
.C(n_172),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_192),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_222),
.B(n_232),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_225),
.B(n_189),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_186),
.A2(n_181),
.B1(n_163),
.B2(n_160),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_227),
.A2(n_187),
.B1(n_193),
.B2(n_197),
.Y(n_249)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_228),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_196),
.B(n_195),
.C(n_202),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_195),
.B(n_199),
.C(n_198),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_230),
.B(n_235),
.C(n_187),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_198),
.A2(n_165),
.B1(n_156),
.B2(n_3),
.Y(n_231)
);

NAND3xp33_ASAP7_75t_L g232 ( 
.A(n_188),
.B(n_10),
.C(n_12),
.Y(n_232)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_183),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_234),
.B(n_207),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_207),
.B(n_210),
.C(n_185),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_236),
.B(n_237),
.C(n_250),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_230),
.B(n_185),
.Y(n_237)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_238),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_215),
.B(n_204),
.Y(n_239)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_239),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_218),
.B(n_194),
.Y(n_242)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_242),
.Y(n_264)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_220),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_244),
.B(n_245),
.Y(n_268)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_226),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_224),
.B(n_205),
.Y(n_246)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_246),
.Y(n_271)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_231),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_247),
.B(n_248),
.Y(n_258)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_223),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_249),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_224),
.B(n_211),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_251),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_221),
.B(n_187),
.C(n_203),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_252),
.B(n_219),
.C(n_229),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_212),
.B(n_203),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_253),
.B(n_255),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_216),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_240),
.A2(n_228),
.B1(n_217),
.B2(n_211),
.Y(n_261)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_261),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_241),
.A2(n_217),
.B(n_233),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_263),
.A2(n_245),
.B(n_233),
.Y(n_274)
);

HB1xp67_ASAP7_75t_L g265 ( 
.A(n_240),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_265),
.B(n_266),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_251),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_267),
.B(n_243),
.C(n_250),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_243),
.B(n_235),
.C(n_225),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_269),
.B(n_246),
.C(n_249),
.Y(n_285)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_268),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_273),
.A2(n_279),
.B(n_283),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_274),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_259),
.B(n_244),
.Y(n_275)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_275),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_276),
.B(n_277),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_269),
.B(n_237),
.C(n_252),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_264),
.B(n_247),
.Y(n_278)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_278),
.Y(n_296)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_268),
.Y(n_279)
);

INVxp67_ASAP7_75t_SL g280 ( 
.A(n_270),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_280),
.B(n_281),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_260),
.B(n_254),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_257),
.B(n_236),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_282),
.B(n_285),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_256),
.B(n_214),
.Y(n_283)
);

FAx1_ASAP7_75t_SL g289 ( 
.A(n_285),
.B(n_227),
.CI(n_271),
.CON(n_289),
.SN(n_289)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_289),
.B(n_11),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_R g291 ( 
.A(n_280),
.B(n_256),
.Y(n_291)
);

NOR2xp67_ASAP7_75t_L g305 ( 
.A(n_291),
.B(n_295),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_272),
.A2(n_258),
.B(n_262),
.Y(n_292)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_292),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_274),
.A2(n_263),
.B1(n_261),
.B2(n_213),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_295),
.A2(n_4),
.B(n_1),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_288),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_297),
.B(n_303),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_293),
.B(n_257),
.C(n_282),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_298),
.B(n_304),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_296),
.A2(n_284),
.B1(n_267),
.B2(n_11),
.Y(n_299)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_299),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_300),
.A2(n_305),
.B(n_286),
.Y(n_308)
);

AOI221xp5_ASAP7_75t_L g302 ( 
.A1(n_287),
.A2(n_14),
.B1(n_2),
.B2(n_3),
.C(n_4),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_302),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_289),
.B(n_14),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_308),
.A2(n_310),
.B(n_298),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_301),
.B(n_290),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_312),
.A2(n_313),
.B(n_314),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_306),
.B(n_293),
.C(n_294),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_309),
.A2(n_302),
.B(n_3),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_315),
.A2(n_307),
.B(n_309),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_316),
.B(n_311),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_3),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_4),
.Y(n_319)
);


endmodule