module fake_jpeg_20784_n_169 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_169);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_169;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_7),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx11_ASAP7_75t_SL g52 ( 
.A(n_8),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_9),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

BUFx10_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_3),
.Y(n_58)
);

BUFx4f_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_20),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_14),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_16),
.Y(n_65)
);

INVx11_ASAP7_75t_SL g66 ( 
.A(n_45),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_0),
.B(n_29),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_6),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_17),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_2),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_10),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_22),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_11),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_2),
.Y(n_75)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_4),
.Y(n_76)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_73),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_73),
.Y(n_78)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_78),
.Y(n_95)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_79),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_80),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_82),
.Y(n_87)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_83),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_0),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_84),
.B(n_71),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_84),
.B(n_49),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_90),
.B(n_91),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_69),
.Y(n_91)
);

INVx13_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_92),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_75),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_93),
.B(n_97),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_94),
.B(n_57),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_79),
.B(n_60),
.Y(n_97)
);

INVx13_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_100),
.A2(n_105),
.B1(n_110),
.B2(n_95),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_101),
.B(n_57),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_89),
.A2(n_62),
.B1(n_63),
.B2(n_64),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_102),
.A2(n_106),
.B1(n_70),
.B2(n_59),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_95),
.A2(n_66),
.B1(n_52),
.B2(n_51),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_86),
.A2(n_67),
.B1(n_50),
.B2(n_54),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_97),
.B(n_72),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_107),
.B(n_71),
.Y(n_124)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_88),
.Y(n_108)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_108),
.Y(n_122)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_109),
.Y(n_113)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_96),
.Y(n_111)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_111),
.Y(n_123)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_85),
.Y(n_112)
);

CKINVDCx14_ASAP7_75t_R g120 ( 
.A(n_112),
.Y(n_120)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_109),
.Y(n_114)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_114),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_115),
.B(n_118),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_98),
.Y(n_117)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_117),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_104),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_105),
.Y(n_119)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_119),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_121),
.A2(n_99),
.B1(n_60),
.B2(n_76),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_124),
.B(n_58),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_100),
.A2(n_52),
.B1(n_85),
.B2(n_61),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_125),
.A2(n_126),
.B1(n_110),
.B2(n_103),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_127),
.A2(n_130),
.B1(n_137),
.B2(n_139),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_128),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_101),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_129),
.B(n_136),
.C(n_18),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_121),
.A2(n_125),
.B1(n_122),
.B2(n_123),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_116),
.A2(n_53),
.B(n_55),
.Y(n_134)
);

XOR2x2_ASAP7_75t_L g141 ( 
.A(n_134),
.B(n_117),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_135),
.B(n_9),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_113),
.B(n_58),
.C(n_74),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_120),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_113),
.A2(n_1),
.B1(n_5),
.B2(n_6),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_141),
.A2(n_143),
.B1(n_145),
.B2(n_147),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_138),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_133),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_144),
.Y(n_151)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_132),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_146),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_135),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_147)
);

OAI21xp33_ASAP7_75t_SL g148 ( 
.A1(n_134),
.A2(n_13),
.B(n_15),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_148),
.A2(n_131),
.B1(n_136),
.B2(n_25),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_149),
.B(n_129),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_153),
.B(n_154),
.C(n_148),
.Y(n_155)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_155),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_151),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_156),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_158),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_157),
.C(n_150),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_160),
.A2(n_140),
.B1(n_152),
.B2(n_141),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_142),
.Y(n_162)
);

OAI21x1_ASAP7_75t_L g163 ( 
.A1(n_162),
.A2(n_152),
.B(n_24),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_19),
.C(n_26),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_164),
.A2(n_27),
.B(n_28),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_165),
.A2(n_30),
.B(n_32),
.Y(n_166)
);

O2A1O1Ixp33_ASAP7_75t_SL g167 ( 
.A1(n_166),
.A2(n_33),
.B(n_34),
.C(n_39),
.Y(n_167)
);

OAI21x1_ASAP7_75t_L g168 ( 
.A1(n_167),
.A2(n_40),
.B(n_41),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_168),
.A2(n_43),
.B(n_46),
.Y(n_169)
);


endmodule