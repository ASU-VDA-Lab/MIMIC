module fake_jpeg_27861_n_272 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_272);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_272;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_175;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_96;

INVx4_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

INVx6_ASAP7_75t_SL g32 ( 
.A(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_23),
.B(n_1),
.Y(n_37)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_46),
.Y(n_50)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_32),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_34),
.Y(n_62)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx3_ASAP7_75t_SL g77 ( 
.A(n_42),
.Y(n_77)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_43),
.B(n_27),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

CKINVDCx6p67_ASAP7_75t_R g72 ( 
.A(n_45),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_17),
.B(n_1),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

NAND2xp33_ASAP7_75t_SL g49 ( 
.A(n_37),
.B(n_34),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_49),
.B(n_68),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_41),
.A2(n_20),
.B1(n_16),
.B2(n_29),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_51),
.A2(n_56),
.B1(n_21),
.B2(n_30),
.Y(n_97)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_53),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_54),
.Y(n_94)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_55),
.B(n_62),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_41),
.A2(n_16),
.B1(n_29),
.B2(n_27),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_40),
.A2(n_16),
.B1(n_29),
.B2(n_31),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_58),
.A2(n_64),
.B1(n_66),
.B2(n_67),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_59),
.B(n_1),
.Y(n_108)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_63),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_38),
.A2(n_31),
.B1(n_26),
.B2(n_24),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_73),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_37),
.A2(n_26),
.B1(n_22),
.B2(n_24),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_37),
.A2(n_22),
.B1(n_19),
.B2(n_33),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_43),
.A2(n_33),
.B1(n_19),
.B2(n_35),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_69),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_46),
.A2(n_35),
.B1(n_18),
.B2(n_25),
.Y(n_70)
);

OA22x2_ASAP7_75t_L g81 ( 
.A1(n_70),
.A2(n_32),
.B1(n_18),
.B2(n_28),
.Y(n_81)
);

INVx5_ASAP7_75t_SL g73 ( 
.A(n_44),
.Y(n_73)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_75),
.Y(n_85)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_76),
.B(n_34),
.Y(n_87)
);

AND2x2_ASAP7_75t_SL g78 ( 
.A(n_49),
.B(n_45),
.Y(n_78)
);

OR2x2_ASAP7_75t_SL g122 ( 
.A(n_78),
.B(n_82),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_81),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_142)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_50),
.B(n_71),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_86),
.B(n_92),
.Y(n_128)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_87),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_50),
.B(n_34),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_89),
.B(n_90),
.Y(n_113)
);

NAND3xp33_ASAP7_75t_SL g90 ( 
.A(n_73),
.B(n_30),
.C(n_28),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_71),
.B(n_28),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_52),
.B(n_25),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_93),
.B(n_96),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_52),
.B(n_25),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_101),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_55),
.B(n_21),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_98),
.B(n_109),
.Y(n_119)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_63),
.Y(n_100)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_100),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_54),
.B(n_30),
.Y(n_101)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_60),
.Y(n_103)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_103),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_61),
.B(n_30),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_104),
.B(n_108),
.Y(n_126)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_60),
.Y(n_105)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_105),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_57),
.A2(n_47),
.B1(n_75),
.B2(n_65),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_106),
.A2(n_72),
.B1(n_77),
.B2(n_5),
.Y(n_129)
);

BUFx2_ASAP7_75t_L g107 ( 
.A(n_69),
.Y(n_107)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_107),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_48),
.B(n_2),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_47),
.Y(n_110)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_110),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_48),
.B(n_2),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_111),
.B(n_112),
.Y(n_125)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_57),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_79),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_114),
.B(n_115),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_107),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_82),
.A2(n_77),
.B1(n_53),
.B2(n_74),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_117),
.A2(n_112),
.B1(n_100),
.B2(n_110),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_86),
.B(n_61),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_118),
.B(n_78),
.C(n_80),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_85),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_121),
.B(n_123),
.Y(n_164)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_95),
.Y(n_123)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_95),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_127),
.B(n_134),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_129),
.A2(n_142),
.B1(n_99),
.B2(n_102),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_91),
.A2(n_72),
.B1(n_4),
.B2(n_5),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_130),
.A2(n_141),
.B1(n_144),
.B2(n_81),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_107),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_108),
.B(n_72),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_137),
.Y(n_162)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_93),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_138),
.B(n_139),
.Y(n_173)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_96),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_84),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_140),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_91),
.A2(n_72),
.B1(n_5),
.B2(n_6),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_92),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_143),
.B(n_105),
.Y(n_157)
);

AO22x1_ASAP7_75t_SL g144 ( 
.A1(n_80),
.A2(n_3),
.B1(n_8),
.B2(n_9),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_83),
.B(n_9),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_145),
.B(n_10),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_114),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_146),
.B(n_153),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_130),
.A2(n_78),
.B(n_80),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_148),
.A2(n_154),
.B(n_170),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_118),
.B(n_128),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_149),
.B(n_151),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_150),
.A2(n_123),
.B1(n_127),
.B2(n_14),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_152),
.A2(n_159),
.B1(n_169),
.B2(n_124),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_115),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_141),
.A2(n_101),
.B(n_94),
.Y(n_154)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_117),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_156),
.B(n_157),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_122),
.A2(n_101),
.B(n_81),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_158),
.A2(n_163),
.B(n_165),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_136),
.B(n_143),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_160),
.B(n_161),
.Y(n_192)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_125),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_122),
.A2(n_81),
.B(n_103),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_113),
.A2(n_116),
.B(n_140),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_138),
.B(n_88),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_167),
.B(n_168),
.Y(n_197)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_135),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_139),
.A2(n_99),
.B1(n_102),
.B2(n_88),
.Y(n_169)
);

O2A1O1Ixp33_ASAP7_75t_L g170 ( 
.A1(n_121),
.A2(n_94),
.B(n_95),
.C(n_11),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_116),
.A2(n_9),
.B(n_10),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_171),
.A2(n_11),
.B(n_13),
.Y(n_194)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_135),
.Y(n_172)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_172),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_174),
.B(n_126),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_176),
.A2(n_184),
.B1(n_190),
.B2(n_150),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_177),
.B(n_194),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_173),
.B(n_126),
.Y(n_178)
);

OR2x2_ASAP7_75t_L g215 ( 
.A(n_178),
.B(n_174),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_156),
.A2(n_129),
.B1(n_124),
.B2(n_120),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_179),
.A2(n_191),
.B1(n_195),
.B2(n_196),
.Y(n_198)
);

OA21x2_ASAP7_75t_L g180 ( 
.A1(n_154),
.A2(n_132),
.B(n_131),
.Y(n_180)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_180),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_149),
.B(n_151),
.C(n_173),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_181),
.B(n_147),
.C(n_164),
.Y(n_216)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_153),
.Y(n_182)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_182),
.Y(n_206)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_166),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_183),
.B(n_146),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_159),
.A2(n_120),
.B1(n_132),
.B2(n_131),
.Y(n_184)
);

AO22x1_ASAP7_75t_SL g188 ( 
.A1(n_163),
.A2(n_144),
.B1(n_134),
.B2(n_133),
.Y(n_188)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_188),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_152),
.A2(n_119),
.B1(n_144),
.B2(n_133),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_148),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_158),
.A2(n_15),
.B1(n_167),
.B2(n_157),
.Y(n_196)
);

INVxp67_ASAP7_75t_SL g199 ( 
.A(n_182),
.Y(n_199)
);

CKINVDCx14_ASAP7_75t_R g220 ( 
.A(n_199),
.Y(n_220)
);

OAI322xp33_ASAP7_75t_L g200 ( 
.A1(n_192),
.A2(n_160),
.A3(n_161),
.B1(n_162),
.B2(n_165),
.C1(n_171),
.C2(n_147),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_200),
.B(n_185),
.Y(n_218)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_201),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_193),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_202),
.B(n_203),
.Y(n_219)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_197),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_179),
.A2(n_196),
.B1(n_176),
.B2(n_195),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_204),
.A2(n_215),
.B1(n_190),
.B2(n_184),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_192),
.B(n_155),
.Y(n_208)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_208),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_210),
.A2(n_180),
.B1(n_183),
.B2(n_188),
.Y(n_226)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_197),
.Y(n_211)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_211),
.Y(n_227)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_187),
.Y(n_212)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_212),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_191),
.Y(n_213)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_213),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_186),
.B(n_155),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_214),
.B(n_185),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_216),
.B(n_186),
.C(n_181),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_217),
.B(n_230),
.C(n_201),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_218),
.B(n_221),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_205),
.A2(n_189),
.B(n_180),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_222),
.A2(n_198),
.B(n_206),
.Y(n_240)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_224),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_226),
.A2(n_209),
.B1(n_205),
.B2(n_204),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_214),
.B(n_189),
.C(n_187),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_216),
.B(n_164),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g244 ( 
.A(n_231),
.B(n_194),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_232),
.A2(n_237),
.B1(n_225),
.B2(n_228),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_233),
.B(n_244),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_224),
.A2(n_210),
.B1(n_202),
.B2(n_209),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_234),
.B(n_222),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_223),
.B(n_208),
.Y(n_236)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_236),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_229),
.A2(n_198),
.B1(n_207),
.B2(n_178),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_231),
.B(n_206),
.C(n_188),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_238),
.B(n_230),
.C(n_226),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_220),
.B(n_215),
.Y(n_239)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_239),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_240),
.B(n_242),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_219),
.B(n_175),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_241),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_219),
.B(n_175),
.Y(n_242)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_245),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_246),
.B(n_243),
.C(n_244),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_247),
.B(n_253),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_233),
.B(n_217),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_253),
.B(n_238),
.C(n_240),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_255),
.B(n_257),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_256),
.A2(n_246),
.B(n_249),
.Y(n_261)
);

NAND4xp25_ASAP7_75t_L g257 ( 
.A(n_252),
.B(n_218),
.C(n_234),
.D(n_177),
.Y(n_257)
);

AOI31xp67_ASAP7_75t_SL g259 ( 
.A1(n_250),
.A2(n_227),
.A3(n_170),
.B(n_168),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_259),
.B(n_170),
.Y(n_263)
);

XNOR2x1_ASAP7_75t_L g260 ( 
.A(n_255),
.B(n_235),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_260),
.B(n_261),
.C(n_264),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_263),
.A2(n_232),
.B1(n_172),
.B2(n_247),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_254),
.B(n_248),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_265),
.B(n_266),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_262),
.A2(n_258),
.B(n_251),
.Y(n_266)
);

A2O1A1Ixp33_ASAP7_75t_L g268 ( 
.A1(n_267),
.A2(n_251),
.B(n_235),
.C(n_221),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_268),
.B(n_169),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_270),
.B(n_269),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_271),
.B(n_166),
.Y(n_272)
);


endmodule