module fake_jpeg_24159_n_250 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_250);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_250;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_96;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

INVx11_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_34),
.Y(n_38)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_31),
.B(n_16),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_18),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_17),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_32),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_39),
.B(n_47),
.Y(n_61)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_40),
.B(n_49),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_0),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_52),
.Y(n_68)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_31),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_32),
.Y(n_47)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_36),
.A2(n_21),
.B1(n_17),
.B2(n_16),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_50),
.A2(n_30),
.B1(n_36),
.B2(n_34),
.Y(n_73)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_51),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_31),
.B(n_20),
.Y(n_52)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_53),
.A2(n_17),
.B1(n_16),
.B2(n_21),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_57),
.A2(n_63),
.B(n_66),
.Y(n_87)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_42),
.Y(n_58)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_44),
.A2(n_17),
.B1(n_23),
.B2(n_20),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_64),
.Y(n_90)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_44),
.A2(n_23),
.B1(n_20),
.B2(n_30),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_70),
.Y(n_89)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_71),
.B(n_38),
.Y(n_77)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_72),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_73),
.A2(n_48),
.B1(n_41),
.B2(n_37),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_71),
.A2(n_50),
.B1(n_51),
.B2(n_54),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_74),
.A2(n_75),
.B1(n_93),
.B2(n_58),
.Y(n_101)
);

AOI22x1_ASAP7_75t_L g75 ( 
.A1(n_68),
.A2(n_44),
.B1(n_29),
.B2(n_37),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_SL g76 ( 
.A(n_68),
.B(n_38),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_76),
.B(n_61),
.C(n_69),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_77),
.B(n_83),
.Y(n_103)
);

OAI32xp33_ASAP7_75t_L g80 ( 
.A1(n_73),
.A2(n_40),
.A3(n_49),
.B1(n_23),
.B2(n_28),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_80),
.B(n_81),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_55),
.B(n_47),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_55),
.B(n_39),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_60),
.B(n_41),
.Y(n_86)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_86),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_91),
.A2(n_65),
.B1(n_45),
.B2(n_64),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_60),
.A2(n_45),
.B1(n_41),
.B2(n_48),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_76),
.Y(n_115)
);

O2A1O1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_93),
.A2(n_61),
.B(n_37),
.C(n_35),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_95),
.A2(n_97),
.B(n_99),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_86),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_96),
.B(n_106),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_75),
.A2(n_62),
.B1(n_59),
.B2(n_67),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_98),
.A2(n_99),
.B1(n_101),
.B2(n_105),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_87),
.A2(n_35),
.B1(n_29),
.B2(n_43),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_72),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_102),
.B(n_111),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g104 ( 
.A(n_82),
.Y(n_104)
);

INVx13_ASAP7_75t_L g118 ( 
.A(n_104),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_75),
.A2(n_58),
.B1(n_35),
.B2(n_29),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_81),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_87),
.A2(n_43),
.B1(n_26),
.B2(n_25),
.Y(n_107)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_107),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_77),
.A2(n_24),
.B1(n_27),
.B2(n_15),
.Y(n_108)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_108),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_80),
.A2(n_24),
.B1(n_27),
.B2(n_15),
.Y(n_110)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_110),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_85),
.B(n_22),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_83),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_112),
.B(n_78),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_85),
.B(n_22),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_113),
.B(n_78),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_122),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_103),
.B(n_112),
.Y(n_116)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_116),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_119),
.A2(n_125),
.B(n_127),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_120),
.B(n_129),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_109),
.B(n_74),
.Y(n_122)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_123),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_96),
.A2(n_109),
.B(n_100),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_103),
.A2(n_22),
.B(n_25),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_104),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_108),
.B(n_100),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_130),
.B(n_133),
.Y(n_137)
);

AOI22x1_ASAP7_75t_L g131 ( 
.A1(n_97),
.A2(n_88),
.B1(n_92),
.B2(n_79),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_131),
.A2(n_88),
.B1(n_95),
.B2(n_90),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_94),
.B(n_92),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_132),
.B(n_106),
.C(n_101),
.Y(n_135)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_104),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_135),
.B(n_140),
.C(n_146),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_116),
.B(n_107),
.Y(n_138)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_138),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_117),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_139),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_132),
.B(n_105),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_114),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_142),
.B(n_144),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_127),
.B(n_104),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_125),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_145),
.B(n_149),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_115),
.B(n_110),
.C(n_98),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_148),
.A2(n_151),
.B1(n_152),
.B2(n_154),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_118),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_118),
.B(n_79),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_150),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_124),
.A2(n_128),
.B1(n_131),
.B2(n_126),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_124),
.A2(n_84),
.B1(n_90),
.B2(n_89),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_122),
.B(n_84),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_153),
.B(n_119),
.C(n_121),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_128),
.A2(n_89),
.B1(n_25),
.B2(n_26),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_137),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_156),
.B(n_160),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_141),
.B(n_126),
.Y(n_158)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_158),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_142),
.B(n_133),
.Y(n_159)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_159),
.Y(n_180)
);

OR2x2_ASAP7_75t_L g160 ( 
.A(n_145),
.B(n_131),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_141),
.B(n_129),
.Y(n_163)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_163),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_164),
.B(n_172),
.C(n_146),
.Y(n_177)
);

HB1xp67_ASAP7_75t_L g165 ( 
.A(n_152),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_165),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_139),
.B(n_121),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_167),
.A2(n_173),
.B(n_135),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_138),
.A2(n_26),
.B1(n_70),
.B2(n_18),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_168),
.A2(n_171),
.B1(n_14),
.B2(n_1),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_151),
.A2(n_70),
.B1(n_18),
.B2(n_24),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_134),
.B(n_18),
.C(n_24),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_143),
.B(n_27),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_136),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_174),
.B(n_154),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_173),
.A2(n_143),
.B1(n_147),
.B2(n_140),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_175),
.A2(n_191),
.B1(n_168),
.B2(n_158),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_177),
.B(n_179),
.Y(n_193)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_178),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_161),
.B(n_134),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_179),
.B(n_183),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_161),
.B(n_153),
.C(n_147),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_181),
.B(n_186),
.C(n_166),
.Y(n_196)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_182),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_164),
.B(n_15),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_172),
.B(n_15),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_184),
.B(n_171),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_163),
.B(n_24),
.C(n_15),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_187),
.B(n_156),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_157),
.B(n_14),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_189),
.B(n_14),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_167),
.A2(n_14),
.B1(n_1),
.B2(n_2),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_193),
.B(n_200),
.Y(n_208)
);

OAI211xp5_ASAP7_75t_SL g194 ( 
.A1(n_175),
.A2(n_160),
.B(n_169),
.C(n_162),
.Y(n_194)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_194),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_195),
.A2(n_176),
.B1(n_190),
.B2(n_186),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_196),
.B(n_201),
.C(n_205),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_197),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_180),
.B(n_166),
.Y(n_199)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_199),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_177),
.B(n_170),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_188),
.A2(n_155),
.B(n_162),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_203),
.A2(n_181),
.B(n_183),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_185),
.A2(n_160),
.B1(n_169),
.B2(n_3),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_204),
.B(n_206),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_189),
.B(n_8),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_207),
.A2(n_218),
.B1(n_211),
.B2(n_215),
.Y(n_228)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_209),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_204),
.Y(n_214)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_214),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_196),
.B(n_0),
.C(n_2),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_215),
.B(n_198),
.C(n_205),
.Y(n_220)
);

NOR3xp33_ASAP7_75t_L g217 ( 
.A(n_192),
.B(n_8),
.C(n_12),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_217),
.B(n_10),
.Y(n_219)
);

A2O1A1Ixp33_ASAP7_75t_L g218 ( 
.A1(n_201),
.A2(n_8),
.B(n_12),
.C(n_4),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_219),
.B(n_221),
.Y(n_231)
);

FAx1_ASAP7_75t_SL g235 ( 
.A(n_220),
.B(n_224),
.CI(n_5),
.CON(n_235),
.SN(n_235)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_217),
.B(n_202),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_214),
.A2(n_198),
.B(n_193),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_222),
.A2(n_4),
.B(n_5),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_210),
.B(n_6),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_216),
.B(n_6),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_225),
.B(n_227),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_213),
.B(n_7),
.Y(n_227)
);

A2O1A1Ixp33_ASAP7_75t_SL g230 ( 
.A1(n_228),
.A2(n_208),
.B(n_9),
.C(n_4),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_226),
.A2(n_212),
.B(n_218),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_229),
.B(n_233),
.C(n_231),
.Y(n_237)
);

AOI31xp67_ASAP7_75t_L g240 ( 
.A1(n_230),
.A2(n_235),
.A3(n_224),
.B(n_11),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_223),
.B(n_5),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_234),
.B(n_236),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_220),
.B(n_9),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_237),
.A2(n_239),
.B(n_242),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_230),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_240),
.B(n_241),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_229),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_232),
.B(n_222),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_238),
.A2(n_11),
.B(n_13),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_244),
.B(n_13),
.C(n_0),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_243),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_246),
.B(n_247),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_248),
.B(n_245),
.C(n_2),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_249),
.B(n_2),
.Y(n_250)
);


endmodule