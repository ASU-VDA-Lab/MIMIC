module fake_jpeg_9926_n_93 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_93);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_93;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_82;

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_31),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_18),
.Y(n_39)
);

INVx11_ASAP7_75t_SL g40 ( 
.A(n_14),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

BUFx16f_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_17),
.B(n_25),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_0),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_46),
.B(n_52),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_0),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_50),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_42),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_53),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_35),
.A2(n_20),
.B1(n_33),
.B2(n_32),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_49),
.A2(n_35),
.B1(n_43),
.B2(n_37),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_1),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_51),
.A2(n_43),
.B1(n_37),
.B2(n_41),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_34),
.B(n_2),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_45),
.B(n_2),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_54),
.B(n_3),
.Y(n_64)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_55),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_55),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_58),
.B(n_64),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_60),
.B(n_67),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_47),
.A2(n_44),
.B1(n_39),
.B2(n_21),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_3),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_69),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_51),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_70),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_6),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_47),
.A2(n_23),
.B1(n_8),
.B2(n_9),
.Y(n_73)
);

AOI32xp33_ASAP7_75t_L g82 ( 
.A1(n_81),
.A2(n_77),
.A3(n_63),
.B1(n_75),
.B2(n_59),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_82),
.B(n_83),
.C(n_74),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_77),
.A2(n_69),
.B1(n_66),
.B2(n_71),
.Y(n_83)
);

AOI221xp5_ASAP7_75t_L g85 ( 
.A1(n_84),
.A2(n_73),
.B1(n_75),
.B2(n_78),
.C(n_61),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_85),
.B(n_65),
.Y(n_86)
);

AO21x1_ASAP7_75t_L g87 ( 
.A1(n_86),
.A2(n_72),
.B(n_76),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_87),
.A2(n_80),
.B1(n_57),
.B2(n_79),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_88),
.B(n_80),
.Y(n_89)
);

AOI322xp5_ASAP7_75t_L g90 ( 
.A1(n_89),
.A2(n_62),
.A3(n_79),
.B1(n_11),
.B2(n_12),
.C1(n_13),
.C2(n_16),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_90),
.B(n_28),
.C(n_10),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_L g92 ( 
.A1(n_91),
.A2(n_29),
.B1(n_22),
.B2(n_24),
.Y(n_92)
);

NAND2x1_ASAP7_75t_L g93 ( 
.A(n_92),
.B(n_26),
.Y(n_93)
);


endmodule