module fake_jpeg_15177_n_353 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_353);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_353;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx24_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx2_ASAP7_75t_SL g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx24_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_8),
.Y(n_39)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx4_ASAP7_75t_SL g40 ( 
.A(n_22),
.Y(n_40)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

AND2x2_ASAP7_75t_SL g41 ( 
.A(n_19),
.B(n_24),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_47),
.Y(n_57)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_38),
.Y(n_56)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_24),
.B(n_0),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_28),
.B(n_9),
.Y(n_48)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_28),
.A2(n_9),
.B1(n_15),
.B2(n_14),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_49),
.A2(n_30),
.B1(n_27),
.B2(n_25),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_52),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_52),
.Y(n_55)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_40),
.A2(n_28),
.B1(n_36),
.B2(n_25),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_58),
.A2(n_49),
.B1(n_40),
.B2(n_27),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_47),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_61),
.B(n_68),
.Y(n_98)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_63),
.A2(n_26),
.B1(n_35),
.B2(n_17),
.Y(n_89)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_67),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_41),
.B(n_36),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_41),
.B(n_30),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_72),
.B(n_41),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_71),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_73),
.B(n_78),
.Y(n_118)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_74),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_61),
.A2(n_46),
.B1(n_51),
.B2(n_45),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_75),
.A2(n_103),
.B1(n_43),
.B2(n_29),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_76),
.B(n_82),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_77),
.A2(n_97),
.B1(n_102),
.B2(n_114),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_79),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_57),
.B(n_41),
.Y(n_82)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_84),
.Y(n_128)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_85),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_59),
.A2(n_40),
.B1(n_45),
.B2(n_33),
.Y(n_86)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_86),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_R g87 ( 
.A(n_63),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_87),
.B(n_99),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_89),
.A2(n_21),
.B1(n_32),
.B2(n_22),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_90),
.Y(n_135)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_91),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_57),
.B(n_51),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_92),
.B(n_94),
.Y(n_141)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_93),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_72),
.B(n_46),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_59),
.A2(n_35),
.B1(n_33),
.B2(n_17),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_95),
.A2(n_112),
.B1(n_113),
.B2(n_22),
.Y(n_124)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_62),
.Y(n_96)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_96),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_69),
.A2(n_48),
.B1(n_39),
.B2(n_26),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_69),
.B(n_32),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_65),
.B(n_43),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_100),
.B(n_104),
.Y(n_144)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_53),
.Y(n_101)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_101),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_65),
.A2(n_42),
.B1(n_18),
.B2(n_38),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_64),
.A2(n_42),
.B1(n_18),
.B2(n_38),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_60),
.B(n_1),
.Y(n_104)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_66),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_105),
.B(n_107),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_53),
.Y(n_106)
);

INVxp67_ASAP7_75t_SL g133 ( 
.A(n_106),
.Y(n_133)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_64),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_60),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_108),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_68),
.A2(n_37),
.B(n_50),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_109),
.B(n_44),
.C(n_22),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_71),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_110),
.B(n_111),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_71),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_57),
.A2(n_44),
.B1(n_18),
.B2(n_38),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_59),
.A2(n_18),
.B1(n_11),
.B2(n_12),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_61),
.A2(n_21),
.B1(n_44),
.B2(n_32),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_71),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_115),
.B(n_50),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_57),
.B(n_1),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_116),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_117),
.B(n_104),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_123),
.B(n_82),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_124),
.A2(n_132),
.B1(n_142),
.B2(n_104),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_126),
.B(n_138),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g149 ( 
.A(n_130),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_112),
.A2(n_43),
.B1(n_21),
.B2(n_32),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_92),
.A2(n_43),
.B1(n_32),
.B2(n_37),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_134),
.A2(n_107),
.B1(n_84),
.B2(n_105),
.Y(n_158)
);

NAND3xp33_ASAP7_75t_L g139 ( 
.A(n_94),
.B(n_13),
.C(n_16),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_139),
.Y(n_152)
);

OAI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_101),
.A2(n_32),
.B1(n_31),
.B2(n_23),
.Y(n_142)
);

NAND2x1_ASAP7_75t_L g147 ( 
.A(n_109),
.B(n_29),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_147),
.A2(n_125),
.B(n_144),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_148),
.A2(n_154),
.B1(n_167),
.B2(n_174),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_150),
.B(n_126),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_120),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_151),
.B(n_161),
.Y(n_180)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_131),
.Y(n_153)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_153),
.Y(n_181)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_131),
.Y(n_155)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_155),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_143),
.A2(n_76),
.B(n_108),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_156),
.A2(n_157),
.B(n_159),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_147),
.B(n_100),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_158),
.A2(n_132),
.B1(n_137),
.B2(n_128),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_141),
.B(n_116),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_135),
.Y(n_160)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_160),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_119),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_120),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_162),
.B(n_170),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_141),
.B(n_76),
.Y(n_163)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_163),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_127),
.B(n_98),
.C(n_81),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_SL g178 ( 
.A(n_164),
.B(n_169),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_141),
.B(n_116),
.Y(n_165)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_165),
.Y(n_194)
);

AO21x1_ASAP7_75t_L g176 ( 
.A1(n_166),
.A2(n_171),
.B(n_172),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_147),
.A2(n_124),
.B1(n_125),
.B2(n_123),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g168 ( 
.A(n_135),
.Y(n_168)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_168),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_127),
.B(n_144),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_121),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_121),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_145),
.Y(n_173)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_173),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_128),
.A2(n_81),
.B1(n_96),
.B2(n_85),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_144),
.A2(n_80),
.B1(n_83),
.B2(n_93),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_175),
.A2(n_136),
.B1(n_138),
.B2(n_146),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_177),
.B(n_182),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_153),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_150),
.B(n_169),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_183),
.B(n_165),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_166),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_184),
.B(n_186),
.Y(n_217)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_155),
.Y(n_185)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_185),
.Y(n_227)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_157),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_157),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_188),
.B(n_191),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_189),
.A2(n_193),
.B(n_200),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_175),
.Y(n_191)
);

OA21x2_ASAP7_75t_L g193 ( 
.A1(n_149),
.A2(n_122),
.B(n_118),
.Y(n_193)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_173),
.Y(n_198)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_198),
.Y(n_212)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_160),
.Y(n_199)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_199),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_149),
.A2(n_136),
.B1(n_146),
.B2(n_130),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_200),
.A2(n_203),
.B1(n_137),
.B2(n_80),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_151),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_202),
.B(n_205),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_157),
.A2(n_137),
.B1(n_134),
.B2(n_88),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_204),
.B(n_111),
.C(n_129),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_162),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_160),
.Y(n_206)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_206),
.Y(n_218)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_168),
.Y(n_207)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_207),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_184),
.B(n_163),
.Y(n_209)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_209),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_210),
.B(n_90),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_192),
.A2(n_167),
.B1(n_158),
.B2(n_148),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_211),
.A2(n_213),
.B1(n_207),
.B2(n_91),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_191),
.A2(n_159),
.B1(n_156),
.B2(n_154),
.Y(n_213)
);

A2O1A1Ixp33_ASAP7_75t_L g214 ( 
.A1(n_190),
.A2(n_171),
.B(n_152),
.C(n_164),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_214),
.B(n_216),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_197),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_186),
.A2(n_172),
.B(n_170),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_219),
.A2(n_233),
.B(n_236),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_183),
.B(n_78),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_221),
.B(n_222),
.C(n_226),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_176),
.B(n_145),
.Y(n_223)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_223),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_181),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_224),
.B(n_228),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_178),
.B(n_129),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_181),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_229),
.B(n_232),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_178),
.B(n_204),
.C(n_201),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_231),
.B(n_234),
.C(n_210),
.Y(n_242)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_176),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_201),
.B(n_79),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_190),
.B(n_83),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_235),
.B(n_106),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_194),
.A2(n_88),
.B(n_37),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_185),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_237),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_223),
.A2(n_188),
.B1(n_189),
.B2(n_203),
.Y(n_239)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_239),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_221),
.B(n_177),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_240),
.B(n_241),
.C(n_242),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_231),
.B(n_234),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_232),
.A2(n_194),
.B1(n_193),
.B2(n_196),
.Y(n_244)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_244),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_211),
.A2(n_193),
.B1(n_180),
.B2(n_187),
.Y(n_247)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_247),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_226),
.B(n_187),
.C(n_195),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_249),
.B(n_250),
.C(n_253),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_208),
.A2(n_220),
.B1(n_217),
.B2(n_233),
.Y(n_251)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_251),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_222),
.B(n_179),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_254),
.B(n_218),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_219),
.A2(n_31),
.B(n_23),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_255),
.B(n_236),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_209),
.B(n_213),
.C(n_235),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_256),
.B(n_258),
.C(n_259),
.Y(n_283)
);

NOR3xp33_ASAP7_75t_SL g257 ( 
.A(n_214),
.B(n_15),
.C(n_16),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_257),
.B(n_15),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_229),
.B(n_74),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_237),
.B(n_168),
.C(n_140),
.Y(n_259)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_262),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_212),
.A2(n_140),
.B1(n_133),
.B2(n_3),
.Y(n_263)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_263),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_245),
.B(n_212),
.Y(n_265)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_265),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_269),
.B(n_252),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_252),
.A2(n_251),
.B(n_246),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_272),
.A2(n_243),
.B1(n_249),
.B2(n_247),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_261),
.B(n_225),
.Y(n_273)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_273),
.Y(n_293)
);

AND2x2_ASAP7_75t_SL g275 ( 
.A(n_248),
.B(n_227),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_275),
.B(n_282),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_260),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_277),
.B(n_215),
.Y(n_292)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_258),
.Y(n_278)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_278),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_279),
.B(n_257),
.Y(n_287)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_239),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_280),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_281),
.A2(n_20),
.B1(n_31),
.B2(n_23),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_244),
.B(n_218),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_256),
.B(n_215),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_284),
.B(n_250),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_285),
.B(n_295),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_287),
.B(n_299),
.Y(n_317)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_288),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_267),
.B(n_241),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_289),
.B(n_297),
.C(n_300),
.Y(n_305)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_292),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_270),
.A2(n_259),
.B1(n_238),
.B2(n_242),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_294),
.A2(n_295),
.B1(n_303),
.B2(n_275),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_270),
.A2(n_238),
.B1(n_253),
.B2(n_240),
.Y(n_295)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_296),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_271),
.B(n_230),
.C(n_140),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_273),
.B(n_230),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_271),
.B(n_283),
.C(n_284),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_283),
.B(n_263),
.C(n_37),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_301),
.B(n_302),
.C(n_269),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_267),
.B(n_278),
.C(n_265),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_293),
.B(n_274),
.Y(n_304)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_304),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_307),
.B(n_308),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_286),
.B(n_274),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_309),
.A2(n_314),
.B(n_316),
.Y(n_328)
);

OAI221xp5_ASAP7_75t_L g310 ( 
.A1(n_298),
.A2(n_272),
.B1(n_282),
.B2(n_275),
.C(n_266),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_310),
.B(n_302),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_290),
.A2(n_268),
.B1(n_280),
.B2(n_264),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_311),
.A2(n_290),
.B1(n_296),
.B2(n_301),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_297),
.B(n_264),
.C(n_268),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_312),
.B(n_313),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_300),
.B(n_266),
.C(n_276),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_294),
.B(n_276),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_317),
.B(n_291),
.Y(n_322)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_322),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_323),
.B(n_326),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_306),
.A2(n_285),
.B(n_288),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_324),
.B(n_1),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_325),
.B(n_329),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_313),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_312),
.A2(n_289),
.B(n_11),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_327),
.B(n_305),
.C(n_29),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_315),
.B(n_9),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_320),
.B(n_318),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_332),
.B(n_338),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_326),
.A2(n_314),
.B1(n_307),
.B2(n_305),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_333),
.B(n_1),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_334),
.B(n_337),
.C(n_29),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_336),
.A2(n_2),
.B(n_3),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_321),
.A2(n_12),
.B1(n_16),
.B2(n_14),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_319),
.B(n_327),
.Y(n_338)
);

AOI21x1_ASAP7_75t_L g339 ( 
.A1(n_336),
.A2(n_324),
.B(n_328),
.Y(n_339)
);

OAI21x1_ASAP7_75t_L g346 ( 
.A1(n_339),
.A2(n_342),
.B(n_334),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_340),
.A2(n_343),
.B(n_330),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_341),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_335),
.A2(n_7),
.B(n_13),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g348 ( 
.A1(n_346),
.A2(n_347),
.B(n_344),
.Y(n_348)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_348),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_349),
.A2(n_331),
.B1(n_345),
.B2(n_333),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_350),
.B(n_7),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g352 ( 
.A1(n_351),
.A2(n_2),
.B(n_4),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_352),
.A2(n_5),
.B(n_6),
.Y(n_353)
);


endmodule