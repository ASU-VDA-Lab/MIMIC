module fake_jpeg_21538_n_105 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_105);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_105;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

INVx8_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

BUFx16f_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_26),
.Y(n_36)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_20),
.B(n_5),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_27),
.B(n_30),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_28),
.B(n_29),
.Y(n_32)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_14),
.B(n_0),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_L g31 ( 
.A(n_30),
.B(n_11),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_31),
.B(n_37),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_26),
.A2(n_21),
.B1(n_13),
.B2(n_20),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_33),
.A2(n_34),
.B1(n_40),
.B2(n_11),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_26),
.A2(n_13),
.B1(n_22),
.B2(n_18),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_24),
.B(n_22),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_29),
.A2(n_13),
.B1(n_1),
.B2(n_2),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_27),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_41),
.B(n_42),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_38),
.B(n_16),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_43),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_37),
.A2(n_29),
.B1(n_28),
.B2(n_24),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_28),
.Y(n_47)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_48),
.A2(n_50),
.B(n_34),
.Y(n_61)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_40),
.A2(n_17),
.B1(n_16),
.B2(n_12),
.Y(n_50)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_51),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_17),
.Y(n_52)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_60),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_61),
.A2(n_48),
.B1(n_45),
.B2(n_46),
.Y(n_68)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_62),
.B(n_51),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_63),
.B(n_46),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_65),
.B(n_66),
.Y(n_74)
);

CKINVDCx14_ASAP7_75t_R g67 ( 
.A(n_61),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_67),
.B(n_73),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_42),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_72),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_56),
.A2(n_47),
.B(n_41),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_59),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_36),
.C(n_35),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_71),
.B(n_55),
.C(n_54),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_33),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_59),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_75),
.B(n_79),
.C(n_19),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_68),
.B(n_25),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_76),
.A2(n_25),
.B(n_23),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_64),
.B(n_53),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_81),
.B(n_82),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_53),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_77),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_83),
.B(n_86),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_76),
.A2(n_70),
.B(n_0),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_85),
.B(n_89),
.Y(n_94)
);

FAx1_ASAP7_75t_SL g90 ( 
.A(n_87),
.B(n_80),
.CI(n_74),
.CON(n_90),
.SN(n_90)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_80),
.A2(n_19),
.B1(n_12),
.B2(n_8),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_88),
.B(n_4),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_12),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_90),
.B(n_91),
.C(n_89),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_23),
.C(n_19),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_92),
.B(n_6),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_96),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_93),
.B(n_4),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_94),
.Y(n_97)
);

OAI21x1_ASAP7_75t_L g101 ( 
.A1(n_97),
.A2(n_90),
.B(n_91),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_98),
.B(n_9),
.Y(n_100)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_100),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_101),
.A2(n_97),
.B(n_9),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_102),
.A2(n_10),
.B1(n_99),
.B2(n_103),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_10),
.Y(n_105)
);


endmodule