module real_jpeg_20967_n_10 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9, n_10);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_9;

output n_10;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_11;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_13;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_139;
wire n_33;
wire n_65;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

INVx13_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_1),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_1),
.A2(n_21),
.B1(n_22),
.B2(n_29),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_1),
.A2(n_29),
.B1(n_44),
.B2(n_45),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_1),
.A2(n_2),
.B1(n_29),
.B2(n_81),
.Y(n_80)
);

A2O1A1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_2),
.A2(n_23),
.B(n_35),
.C(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_2),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_2),
.A2(n_6),
.B1(n_35),
.B2(n_81),
.Y(n_83)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_3),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_6),
.B(n_19),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_6),
.A2(n_27),
.B1(n_28),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_6),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_6),
.A2(n_21),
.B1(n_22),
.B2(n_35),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_6),
.A2(n_35),
.B1(n_44),
.B2(n_45),
.Y(n_55)
);

AOI21xp33_ASAP7_75t_SL g60 ( 
.A1(n_6),
.A2(n_40),
.B(n_45),
.Y(n_60)
);

AOI21xp33_ASAP7_75t_SL g71 ( 
.A1(n_6),
.A2(n_7),
.B(n_22),
.Y(n_71)
);

AOI21xp33_ASAP7_75t_L g107 ( 
.A1(n_6),
.A2(n_8),
.B(n_28),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_7),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_20)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

OAI22xp33_ASAP7_75t_L g51 ( 
.A1(n_8),
.A2(n_44),
.B1(n_45),
.B2(n_52),
.Y(n_51)
);

INVx6_ASAP7_75t_SL g52 ( 
.A(n_8),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_8),
.A2(n_27),
.B1(n_28),
.B2(n_52),
.Y(n_53)
);

BUFx3_ASAP7_75t_SL g45 ( 
.A(n_9),
.Y(n_45)
);

XOR2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_99),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_SL g11 ( 
.A(n_12),
.B(n_97),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_66),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_13),
.B(n_66),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_49),
.C(n_56),
.Y(n_13)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_14),
.B(n_139),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g14 ( 
.A1(n_15),
.A2(n_16),
.B1(n_37),
.B2(n_38),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_16),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_24),
.B2(n_36),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_17),
.B(n_36),
.C(n_38),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_18),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_19),
.A2(n_80),
.B(n_82),
.Y(n_79)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

A2O1A1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_20),
.A2(n_81),
.B(n_85),
.C(n_86),
.Y(n_84)
);

A2O1A1Ixp33_ASAP7_75t_L g39 ( 
.A1(n_21),
.A2(n_40),
.B(n_42),
.C(n_43),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_21),
.B(n_40),
.Y(n_42)
);

INVx4_ASAP7_75t_SL g21 ( 
.A(n_22),
.Y(n_21)
);

A2O1A1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_22),
.A2(n_35),
.B(n_41),
.C(n_60),
.Y(n_59)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_23),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_24),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_24),
.B(n_104),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_24),
.B(n_104),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_30),
.B(n_32),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_26),
.A2(n_31),
.B1(n_33),
.B2(n_34),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_27),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_27),
.B(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_28),
.B(n_31),
.Y(n_33)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_31),
.B(n_35),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_34),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_33),
.B(n_65),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

A2O1A1Ixp33_ASAP7_75t_L g106 ( 
.A1(n_35),
.A2(n_45),
.B(n_52),
.C(n_107),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_35),
.B(n_53),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_35),
.B(n_43),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_36),
.B(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_43),
.B1(n_46),
.B2(n_48),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_39),
.B(n_48),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_40),
.A2(n_41),
.B1(n_44),
.B2(n_45),
.Y(n_43)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_43),
.Y(n_93)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_47),
.A2(n_93),
.B(n_94),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_49),
.A2(n_125),
.B1(n_126),
.B2(n_127),
.Y(n_124)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_49),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_49),
.B(n_72),
.C(n_126),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_49),
.A2(n_56),
.B1(n_57),
.B2(n_127),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_50),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_50),
.B(n_53),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_50),
.B(n_55),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_53),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_53),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_54),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_58),
.B(n_61),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_58),
.A2(n_59),
.B1(n_61),
.B2(n_62),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_64),
.Y(n_62)
);

XOR2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_77),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_69),
.B1(n_75),
.B2(n_76),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_72),
.B1(n_73),
.B2(n_74),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_70),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_72),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_72),
.B(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_72),
.B(n_118),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_72),
.A2(n_74),
.B1(n_124),
.B2(n_128),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_79),
.B1(n_87),
.B2(n_96),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_81),
.B(n_85),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_84),
.Y(n_82)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_87),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_89),
.B1(n_92),
.B2(n_95),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_91),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_92),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_92),
.A2(n_95),
.B1(n_108),
.B2(n_112),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_92),
.B(n_108),
.C(n_133),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_100),
.A2(n_136),
.B(n_140),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_130),
.B(n_135),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_102),
.A2(n_121),
.B(n_129),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_113),
.B(n_120),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_106),
.B1(n_108),
.B2(n_112),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_106),
.B(n_108),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_108),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_110),
.B(n_111),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_117),
.B(n_119),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_123),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_122),
.B(n_123),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_124),
.Y(n_128)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_132),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_131),
.B(n_132),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_134),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_138),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_137),
.B(n_138),
.Y(n_140)
);


endmodule