module fake_jpeg_4873_n_327 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_327);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_327;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_15),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx5p33_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_37),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx3_ASAP7_75t_SL g36 ( 
.A(n_29),
.Y(n_36)
);

INVx3_ASAP7_75t_SL g58 ( 
.A(n_36),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_39),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_42),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_27),
.B(n_0),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_44),
.Y(n_51)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_47),
.B(n_52),
.Y(n_77)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_27),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_54),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_27),
.Y(n_55)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_56),
.B(n_57),
.Y(n_78)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_63),
.Y(n_80)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_64),
.B(n_66),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_18),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_67),
.B(n_68),
.Y(n_90)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_51),
.A2(n_32),
.B1(n_23),
.B2(n_28),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_69),
.A2(n_26),
.B1(n_17),
.B2(n_31),
.Y(n_108)
);

CKINVDCx12_ASAP7_75t_R g70 ( 
.A(n_58),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_70),
.B(n_88),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_43),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_71),
.B(n_86),
.Y(n_105)
);

INVx3_ASAP7_75t_SL g72 ( 
.A(n_58),
.Y(n_72)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_72),
.Y(n_95)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_73),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_45),
.B(n_43),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_79),
.B(n_83),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_45),
.B(n_22),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_19),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_47),
.B(n_19),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_50),
.B(n_19),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_53),
.B(n_32),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_87),
.A2(n_93),
.B1(n_32),
.B2(n_23),
.Y(n_100)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_60),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_89),
.B(n_92),
.Y(n_115)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_60),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_62),
.A2(n_32),
.B1(n_23),
.B2(n_28),
.Y(n_93)
);

HB1xp67_ASAP7_75t_L g94 ( 
.A(n_46),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_94),
.B(n_66),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_78),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_96),
.B(n_97),
.Y(n_129)
);

CKINVDCx5p33_ASAP7_75t_R g97 ( 
.A(n_73),
.Y(n_97)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_72),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_98),
.B(n_103),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_100),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_102),
.B(n_114),
.Y(n_146)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_83),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_79),
.A2(n_57),
.B(n_64),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_104),
.A2(n_24),
.B(n_59),
.Y(n_148)
);

INVx2_ASAP7_75t_SL g106 ( 
.A(n_72),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_106),
.B(n_107),
.Y(n_145)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_84),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_108),
.A2(n_18),
.B1(n_21),
.B2(n_17),
.Y(n_141)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_88),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_110),
.A2(n_118),
.B1(n_120),
.B2(n_92),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_71),
.B(n_63),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_111),
.B(n_87),
.Y(n_127)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_90),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_112),
.B(n_116),
.Y(n_144)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_85),
.Y(n_113)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_113),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_82),
.B(n_86),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_77),
.Y(n_116)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_89),
.Y(n_118)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_119),
.Y(n_124)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_85),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_75),
.A2(n_28),
.B1(n_68),
.B2(n_56),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_121),
.A2(n_122),
.B1(n_91),
.B2(n_100),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_71),
.A2(n_34),
.B1(n_53),
.B2(n_41),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_115),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_123),
.B(n_126),
.Y(n_160)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_99),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_127),
.B(n_105),
.C(n_112),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_103),
.B(n_81),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_128),
.B(n_131),
.Y(n_154)
);

OAI32xp33_ASAP7_75t_L g131 ( 
.A1(n_99),
.A2(n_75),
.A3(n_81),
.B1(n_69),
.B2(n_82),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_108),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_132),
.B(n_133),
.Y(n_163)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_110),
.Y(n_133)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_118),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_135),
.A2(n_140),
.B1(n_101),
.B2(n_52),
.Y(n_172)
);

INVx13_ASAP7_75t_L g136 ( 
.A(n_95),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_136),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_137),
.A2(n_139),
.B1(n_95),
.B2(n_105),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_111),
.B(n_87),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_138),
.A2(n_148),
.B(n_24),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_122),
.A2(n_91),
.B1(n_80),
.B2(n_34),
.Y(n_139)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_97),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_141),
.Y(n_175)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_104),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_142),
.B(n_143),
.Y(n_156)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_114),
.Y(n_143)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_147),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_149),
.B(n_151),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_150),
.B(n_169),
.C(n_176),
.Y(n_188)
);

BUFx24_ASAP7_75t_SL g151 ( 
.A(n_128),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_134),
.A2(n_96),
.B1(n_107),
.B2(n_98),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_152),
.A2(n_156),
.B(n_166),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_143),
.B(n_102),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_153),
.B(n_157),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_126),
.B(n_116),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_155),
.B(n_159),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_132),
.B(n_109),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_142),
.B(n_106),
.Y(n_159)
);

BUFx5_ASAP7_75t_L g161 ( 
.A(n_135),
.Y(n_161)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_161),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_134),
.A2(n_106),
.B1(n_117),
.B2(n_113),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_162),
.A2(n_168),
.B1(n_125),
.B2(n_123),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_146),
.B(n_44),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_164),
.B(n_165),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_131),
.B(n_39),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_166),
.A2(n_173),
.B(n_18),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_127),
.B(n_39),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_167),
.B(n_124),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_137),
.A2(n_120),
.B1(n_101),
.B2(n_41),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_138),
.B(n_44),
.Y(n_169)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_130),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_171),
.B(n_174),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_172),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_148),
.A2(n_22),
.B(n_30),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_145),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_138),
.B(n_39),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_160),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_177),
.B(n_180),
.Y(n_204)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_178),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_176),
.B(n_129),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_179),
.B(n_203),
.Y(n_207)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_155),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_163),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_183),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_165),
.A2(n_139),
.B1(n_146),
.B2(n_140),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_186),
.A2(n_194),
.B1(n_170),
.B2(n_149),
.Y(n_205)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_162),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_187),
.B(n_197),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_189),
.A2(n_184),
.B1(n_187),
.B2(n_199),
.Y(n_225)
);

NOR4xp25_ASAP7_75t_L g215 ( 
.A(n_190),
.B(n_175),
.C(n_173),
.D(n_152),
.Y(n_215)
);

OR2x2_ASAP7_75t_L g191 ( 
.A(n_157),
.B(n_156),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_191),
.B(n_150),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_193),
.B(n_164),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_170),
.A2(n_125),
.B1(n_133),
.B2(n_124),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_154),
.B(n_144),
.Y(n_195)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_195),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_174),
.B(n_141),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_159),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_198),
.B(n_200),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_154),
.B(n_136),
.Y(n_199)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_199),
.Y(n_211)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_168),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_153),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_201),
.B(n_26),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_169),
.B(n_136),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_205),
.A2(n_189),
.B1(n_185),
.B2(n_184),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_202),
.B(n_171),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_210),
.B(n_218),
.Y(n_238)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_182),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_212),
.B(n_214),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_213),
.Y(n_235)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_182),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_215),
.A2(n_219),
.B(n_221),
.Y(n_244)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_217),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_183),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_193),
.Y(n_219)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_178),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_203),
.B(n_167),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_222),
.B(n_207),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_180),
.B(n_175),
.Y(n_223)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_223),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_198),
.B(n_158),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_224),
.B(n_225),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_200),
.A2(n_21),
.B1(n_161),
.B2(n_17),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_226),
.A2(n_216),
.B1(n_26),
.B2(n_31),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_181),
.B(n_21),
.Y(n_227)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_227),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_228),
.A2(n_201),
.B1(n_191),
.B2(n_177),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_207),
.B(n_188),
.C(n_179),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_229),
.B(n_242),
.C(n_247),
.Y(n_255)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_230),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_231),
.B(n_233),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_232),
.A2(n_236),
.B1(n_246),
.B2(n_238),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_222),
.B(n_188),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_206),
.A2(n_195),
.B1(n_185),
.B2(n_186),
.Y(n_236)
);

INVx11_ASAP7_75t_L g240 ( 
.A(n_224),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_240),
.B(n_243),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_225),
.B(n_190),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_241),
.B(n_16),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_212),
.B(n_196),
.C(n_65),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_206),
.A2(n_192),
.B1(n_22),
.B2(n_30),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_214),
.B(n_65),
.C(n_192),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_211),
.A2(n_24),
.B1(n_30),
.B2(n_31),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_248),
.A2(n_204),
.B(n_209),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_211),
.B(n_65),
.C(n_39),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_250),
.B(n_221),
.C(n_226),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_248),
.B(n_213),
.Y(n_251)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_251),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_239),
.B(n_223),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_252),
.A2(n_257),
.B(n_261),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_245),
.B(n_237),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_253),
.B(n_262),
.C(n_241),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_245),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_254),
.B(n_263),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_233),
.B(n_220),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_256),
.B(n_268),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_229),
.B(n_208),
.C(n_217),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_259),
.B(n_267),
.C(n_76),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_235),
.B(n_208),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_234),
.B(n_217),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_264),
.A2(n_244),
.B(n_258),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_240),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_266),
.B(n_243),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_231),
.B(n_247),
.C(n_242),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_269),
.A2(n_280),
.B(n_38),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_260),
.A2(n_236),
.B1(n_232),
.B2(n_262),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_274),
.A2(n_268),
.B1(n_33),
.B2(n_20),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_275),
.A2(n_276),
.B(n_277),
.Y(n_292)
);

A2O1A1O1Ixp25_ASAP7_75t_L g277 ( 
.A1(n_253),
.A2(n_250),
.B(n_249),
.C(n_16),
.D(n_76),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_278),
.B(n_281),
.C(n_282),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_267),
.A2(n_76),
.B(n_25),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_279),
.A2(n_283),
.B(n_16),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_266),
.B(n_76),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_265),
.B(n_25),
.C(n_74),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_265),
.B(n_74),
.C(n_38),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_255),
.B(n_74),
.C(n_38),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_273),
.B(n_255),
.Y(n_284)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_284),
.Y(n_300)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_285),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_270),
.B(n_272),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_286),
.B(n_296),
.C(n_35),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_287),
.A2(n_289),
.B(n_290),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_271),
.Y(n_289)
);

A2O1A1Ixp33_ASAP7_75t_L g290 ( 
.A1(n_277),
.A2(n_11),
.B(n_15),
.C(n_14),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_L g291 ( 
.A1(n_283),
.A2(n_11),
.B1(n_15),
.B2(n_14),
.Y(n_291)
);

OAI22x1_ASAP7_75t_L g298 ( 
.A1(n_291),
.A2(n_294),
.B1(n_290),
.B2(n_285),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_282),
.B(n_48),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_293),
.B(n_295),
.Y(n_299)
);

INVxp67_ASAP7_75t_SL g294 ( 
.A(n_278),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_270),
.B(n_48),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_292),
.B(n_41),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_297),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_L g309 ( 
.A1(n_298),
.A2(n_303),
.B1(n_306),
.B2(n_300),
.Y(n_309)
);

OAI21x1_ASAP7_75t_L g301 ( 
.A1(n_286),
.A2(n_288),
.B(n_289),
.Y(n_301)
);

OAI21x1_ASAP7_75t_L g307 ( 
.A1(n_301),
.A2(n_61),
.B(n_35),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_288),
.A2(n_9),
.B1(n_13),
.B2(n_10),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_302),
.A2(n_8),
.B1(n_14),
.B2(n_4),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_304),
.B(n_33),
.C(n_2),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_289),
.B(n_0),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_305),
.A2(n_1),
.B(n_2),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_307),
.A2(n_309),
.B(n_312),
.Y(n_319)
);

AOI322xp5_ASAP7_75t_L g315 ( 
.A1(n_308),
.A2(n_311),
.A3(n_298),
.B1(n_7),
.B2(n_4),
.C1(n_5),
.C2(n_6),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_299),
.B(n_20),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_297),
.B(n_35),
.Y(n_313)
);

OR2x2_ASAP7_75t_L g318 ( 
.A(n_313),
.B(n_7),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_314),
.A2(n_6),
.B(n_10),
.Y(n_317)
);

NOR2x1_ASAP7_75t_L g321 ( 
.A(n_315),
.B(n_317),
.Y(n_321)
);

HB1xp67_ASAP7_75t_L g316 ( 
.A(n_309),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_316),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_320),
.B(n_310),
.Y(n_322)
);

OAI311xp33_ASAP7_75t_L g323 ( 
.A1(n_322),
.A2(n_321),
.A3(n_318),
.B1(n_319),
.C1(n_314),
.Y(n_323)
);

AOI322xp5_ASAP7_75t_L g324 ( 
.A1(n_323),
.A2(n_33),
.A3(n_7),
.B1(n_4),
.B2(n_5),
.C1(n_8),
.C2(n_10),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_324),
.B(n_5),
.C(n_8),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_1),
.C(n_2),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_2),
.Y(n_327)
);


endmodule