module fake_jpeg_25244_n_168 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_168);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_168;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx4_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_36),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_40),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_16),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

BUFx16f_ASAP7_75t_L g52 ( 
.A(n_10),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

HB1xp67_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_38),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_7),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_12),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_14),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_11),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_5),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_67),
.B(n_0),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_71),
.B(n_66),
.Y(n_76)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g81 ( 
.A(n_73),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_46),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_50),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_72),
.A2(n_44),
.B1(n_62),
.B2(n_57),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_75),
.B(n_82),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_76),
.B(n_84),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_79),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_73),
.B(n_47),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_70),
.B(n_58),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_85),
.B(n_86),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_71),
.A2(n_49),
.B1(n_51),
.B2(n_62),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_71),
.B(n_65),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_87),
.B(n_66),
.Y(n_96)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_83),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_95),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_91),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_63),
.C(n_45),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_92),
.B(n_96),
.Y(n_108)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

INVx6_ASAP7_75t_SL g94 ( 
.A(n_79),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_94),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_78),
.Y(n_95)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_98),
.Y(n_114)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_75),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_99),
.B(n_102),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_77),
.B(n_56),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_101),
.B(n_64),
.Y(n_106)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_78),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g103 ( 
.A(n_81),
.Y(n_103)
);

NOR2x1_ASAP7_75t_L g105 ( 
.A(n_103),
.B(n_104),
.Y(n_105)
);

BUFx2_ASAP7_75t_SL g104 ( 
.A(n_81),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_106),
.B(n_48),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_67),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_112),
.B(n_115),
.C(n_97),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_90),
.A2(n_59),
.B(n_55),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_108),
.B(n_92),
.Y(n_116)
);

OAI21xp33_ASAP7_75t_L g135 ( 
.A1(n_116),
.A2(n_60),
.B(n_111),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_119),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_118),
.B(n_121),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_112),
.B(n_91),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_108),
.B(n_0),
.Y(n_120)
);

INVx1_ASAP7_75t_SL g137 ( 
.A(n_120),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_110),
.B(n_1),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_110),
.B(n_1),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_122),
.B(n_54),
.Y(n_131)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_107),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_123),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_107),
.B(n_53),
.C(n_100),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_124),
.B(n_114),
.C(n_93),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_105),
.A2(n_98),
.B1(n_102),
.B2(n_53),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_125),
.A2(n_89),
.B1(n_60),
.B2(n_52),
.Y(n_139)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_113),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_126),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_116),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_128),
.B(n_133),
.Y(n_149)
);

NAND2xp33_ASAP7_75t_SL g129 ( 
.A(n_118),
.B(n_103),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_129),
.B(n_4),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_131),
.B(n_132),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_116),
.B(n_54),
.Y(n_132)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_135),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_123),
.A2(n_109),
.B(n_52),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_138),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_139),
.A2(n_140),
.B1(n_141),
.B2(n_2),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_116),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_140)
);

O2A1O1Ixp33_ASAP7_75t_L g141 ( 
.A1(n_123),
.A2(n_20),
.B(n_39),
.C(n_34),
.Y(n_141)
);

CKINVDCx14_ASAP7_75t_R g155 ( 
.A(n_142),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_127),
.B(n_3),
.Y(n_143)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_143),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_145),
.B(n_147),
.C(n_148),
.Y(n_153)
);

FAx1_ASAP7_75t_SL g147 ( 
.A(n_128),
.B(n_5),
.CI(n_6),
.CON(n_147),
.SN(n_147)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_141),
.A2(n_23),
.B1(n_32),
.B2(n_31),
.Y(n_148)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_136),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_150),
.B(n_134),
.C(n_130),
.Y(n_154)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_154),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_155),
.B(n_146),
.C(n_149),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_157),
.A2(n_151),
.B1(n_153),
.B2(n_152),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_147),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_145),
.C(n_156),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_160),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_138),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_162),
.B(n_143),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_163),
.A2(n_137),
.B(n_144),
.Y(n_164)
);

OAI321xp33_ASAP7_75t_L g165 ( 
.A1(n_164),
.A2(n_135),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.C(n_10),
.Y(n_165)
);

OAI321xp33_ASAP7_75t_L g166 ( 
.A1(n_165),
.A2(n_6),
.A3(n_8),
.B1(n_9),
.B2(n_11),
.C(n_12),
.Y(n_166)
);

AOI221xp5_ASAP7_75t_L g167 ( 
.A1(n_166),
.A2(n_15),
.B1(n_18),
.B2(n_19),
.C(n_22),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_167),
.A2(n_24),
.B(n_26),
.Y(n_168)
);


endmodule