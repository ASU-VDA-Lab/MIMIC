module real_jpeg_32695_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_215;
wire n_176;
wire n_166;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_373;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_14;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

BUFx12f_ASAP7_75t_L g106 ( 
.A(n_0),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_0),
.Y(n_124)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_0),
.Y(n_222)
);

AOI22x1_ASAP7_75t_L g161 ( 
.A1(n_1),
.A2(n_112),
.B1(n_162),
.B2(n_163),
.Y(n_161)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_1),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_2),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_3),
.Y(n_66)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_4),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_4),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_4),
.Y(n_119)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_4),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_5),
.A2(n_42),
.B1(n_44),
.B2(n_45),
.Y(n_41)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

OA22x2_ASAP7_75t_L g93 ( 
.A1(n_5),
.A2(n_44),
.B1(n_94),
.B2(n_97),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_5),
.A2(n_44),
.B1(n_112),
.B2(n_116),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_5),
.A2(n_44),
.B1(n_200),
.B2(n_203),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_6),
.Y(n_69)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_6),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_6),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g304 ( 
.A(n_6),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_8),
.A2(n_212),
.B1(n_213),
.B2(n_215),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_8),
.Y(n_212)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_9),
.Y(n_183)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_9),
.Y(n_190)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_10),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_10),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_11),
.A2(n_32),
.B1(n_33),
.B2(n_37),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_11),
.Y(n_32)
);

OAI22x1_ASAP7_75t_SL g76 ( 
.A1(n_11),
.A2(n_32),
.B1(n_77),
.B2(n_81),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_11),
.A2(n_32),
.B1(n_126),
.B2(n_128),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_11),
.B(n_133),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_11),
.A2(n_32),
.B1(n_172),
.B2(n_176),
.Y(n_171)
);

NAND2xp33_ASAP7_75t_SL g258 ( 
.A(n_11),
.B(n_19),
.Y(n_258)
);

INVx2_ASAP7_75t_R g300 ( 
.A(n_11),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_11),
.B(n_61),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_11),
.B(n_198),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_241),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_239),
.Y(n_13)
);

OR2x2_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_223),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_15),
.B(n_223),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_153),
.Y(n_15)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_59),
.C(n_98),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_17),
.A2(n_59),
.B1(n_227),
.B2(n_228),
.Y(n_226)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_17),
.Y(n_228)
);

OA22x2_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_30),
.B1(n_41),
.B2(n_48),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_18),
.A2(n_41),
.B(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2x1_ASAP7_75t_L g49 ( 
.A(n_19),
.B(n_50),
.Y(n_49)
);

AO22x2_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_22),
.B1(n_25),
.B2(n_27),
.Y(n_19)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_21),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_21),
.Y(n_151)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_24),
.Y(n_83)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_25),
.Y(n_152)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_31),
.B(n_49),
.Y(n_157)
);

OAI211xp5_ASAP7_75t_SL g280 ( 
.A1(n_32),
.A2(n_281),
.B(n_284),
.C(n_287),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_32),
.B(n_318),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_32),
.B(n_323),
.Y(n_322)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_40),
.Y(n_146)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_46),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_53),
.B1(n_55),
.B2(n_56),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g134 ( 
.A(n_57),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_59),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_59),
.A2(n_227),
.B1(n_360),
.B2(n_361),
.Y(n_359)
);

OA22x2_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_75),
.B1(n_84),
.B2(n_93),
.Y(n_59)
);

AOI21x1_ASAP7_75t_L g158 ( 
.A1(n_60),
.A2(n_75),
.B(n_84),
.Y(n_158)
);

OA22x2_ASAP7_75t_L g234 ( 
.A1(n_60),
.A2(n_75),
.B1(n_84),
.B2(n_93),
.Y(n_234)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NAND2x1p5_ASAP7_75t_L g84 ( 
.A(n_62),
.B(n_85),
.Y(n_84)
);

AOI22x1_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_67),
.B1(n_70),
.B2(n_72),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_66),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_69),
.Y(n_178)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_74),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_74),
.Y(n_192)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_79),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_80),
.Y(n_139)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_83),
.Y(n_87)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_88),
.B1(n_89),
.B2(n_92),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_91),
.Y(n_286)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx2_ASAP7_75t_SL g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_99),
.B(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

OAI21xp33_ASAP7_75t_L g254 ( 
.A1(n_100),
.A2(n_101),
.B(n_131),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_131),
.Y(n_100)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_101),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_110),
.B(n_120),
.Y(n_101)
);

OA22x2_ASAP7_75t_L g347 ( 
.A1(n_102),
.A2(n_110),
.B1(n_276),
.B2(n_348),
.Y(n_347)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_103),
.A2(n_161),
.B1(n_210),
.B2(n_218),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_103),
.B(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_104),
.B(n_125),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_107),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g334 ( 
.A(n_105),
.B(n_300),
.Y(n_334)
);

INVx4_ASAP7_75t_SL g105 ( 
.A(n_106),
.Y(n_105)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_109),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_109),
.Y(n_130)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_109),
.Y(n_217)
);

INVx3_ASAP7_75t_L g321 ( 
.A(n_109),
.Y(n_321)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_111),
.B(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_115),
.Y(n_214)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx6_ASAP7_75t_L g165 ( 
.A(n_119),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_119),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_125),
.Y(n_120)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_124),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_124),
.Y(n_263)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_125),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

AO22x1_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_135),
.B1(n_143),
.B2(n_147),
.Y(n_131)
);

INVx1_ASAP7_75t_SL g133 ( 
.A(n_134),
.Y(n_133)
);

NAND2xp33_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_140),
.Y(n_135)
);

BUFx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_138),
.Y(n_289)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx11_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

BUFx12f_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_152),
.Y(n_147)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_206),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_159),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_158),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_156),
.Y(n_235)
);

AND2x4_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_170),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_160),
.A2(n_170),
.B1(n_230),
.B2(n_231),
.Y(n_229)
);

INVxp67_ASAP7_75t_SL g231 ( 
.A(n_160),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_166),
.B(n_169),
.Y(n_160)
);

BUFx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

BUFx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

OA22x2_ASAP7_75t_L g194 ( 
.A1(n_165),
.A2(n_195),
.B1(n_196),
.B2(n_197),
.Y(n_194)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_165),
.Y(n_197)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_169),
.B(n_261),
.Y(n_260)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_170),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_170),
.A2(n_230),
.B1(n_234),
.B2(n_251),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_170),
.A2(n_230),
.B1(n_315),
.B2(n_316),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g356 ( 
.A(n_170),
.Y(n_356)
);

AO22x2_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_179),
.B1(n_198),
.B2(n_199),
.Y(n_170)
);

AO22x2_ASAP7_75t_L g208 ( 
.A1(n_171),
.A2(n_179),
.B1(n_198),
.B2(n_199),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_171),
.B(n_237),
.Y(n_236)
);

INVx3_ASAP7_75t_L g325 ( 
.A(n_172),
.Y(n_325)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_178),
.Y(n_283)
);

AOI21x1_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_186),
.B(n_193),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_180),
.A2(n_317),
.B1(n_322),
.B2(n_326),
.Y(n_316)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

OAI21xp33_ASAP7_75t_SL g238 ( 
.A1(n_181),
.A2(n_187),
.B(n_194),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_184),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_183),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_183),
.Y(n_196)
);

INVx5_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_191),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_192),
.Y(n_202)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_192),
.Y(n_205)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_194),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_194),
.B(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

XOR2x2_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_209),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_207),
.B(n_308),
.C(n_310),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_207),
.A2(n_208),
.B1(n_363),
.B2(n_364),
.Y(n_362)
);

INVx2_ASAP7_75t_SL g207 ( 
.A(n_208),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_208),
.B(n_346),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_208),
.B(n_364),
.C(n_368),
.Y(n_367)
);

INVxp33_ASAP7_75t_SL g210 ( 
.A(n_211),
.Y(n_210)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx2_ASAP7_75t_SL g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_221),
.Y(n_279)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_229),
.C(n_232),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_225),
.B(n_246),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_227),
.B(n_257),
.C(n_259),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_229),
.B(n_233),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_230),
.B(n_315),
.Y(n_344)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.C(n_236),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_234),
.A2(n_236),
.B1(n_251),
.B2(n_252),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_234),
.Y(n_251)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_234),
.Y(n_355)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_235),
.Y(n_249)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_236),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_264),
.B(n_372),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_247),
.Y(n_244)
);

NOR2x1_ASAP7_75t_L g373 ( 
.A(n_245),
.B(n_247),
.Y(n_373)
);

MAJx2_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_253),
.C(n_255),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_SL g369 ( 
.A(n_248),
.B(n_370),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_254),
.B(n_256),
.Y(n_370)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_257),
.A2(n_258),
.B1(n_259),
.B2(n_260),
.Y(n_361)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_259),
.B(n_314),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_259),
.B(n_314),
.Y(n_342)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_260),
.B(n_333),
.Y(n_332)
);

BUFx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

BUFx2_ASAP7_75t_R g349 ( 
.A(n_263),
.Y(n_349)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

BUFx2_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

AO21x2_ASAP7_75t_L g266 ( 
.A1(n_267),
.A2(n_366),
.B(n_371),
.Y(n_266)
);

AO21x1_ASAP7_75t_L g267 ( 
.A1(n_268),
.A2(n_352),
.B(n_365),
.Y(n_267)
);

OAI21x1_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_311),
.B(n_351),
.Y(n_268)
);

NOR2xp67_ASAP7_75t_SL g269 ( 
.A(n_270),
.B(n_307),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_270),
.B(n_307),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_272),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_305),
.Y(n_272)
);

NAND3xp33_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_280),
.C(n_290),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

OAI21xp33_ASAP7_75t_L g305 ( 
.A1(n_275),
.A2(n_291),
.B(n_306),
.Y(n_305)
);

OAI21xp33_ASAP7_75t_SL g363 ( 
.A1(n_275),
.A2(n_291),
.B(n_306),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_280),
.Y(n_306)
);

INVx4_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_299),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx8_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_301),
.Y(n_299)
);

INVx4_ASAP7_75t_SL g301 ( 
.A(n_302),
.Y(n_301)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_309),
.B(n_331),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_309),
.B(n_331),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_310),
.B(n_347),
.Y(n_346)
);

AOI21x1_ASAP7_75t_L g311 ( 
.A1(n_312),
.A2(n_343),
.B(n_350),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_313),
.A2(n_329),
.B(n_342),
.Y(n_312)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx2_ASAP7_75t_SL g318 ( 
.A(n_319),
.Y(n_318)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx4_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_330),
.A2(n_332),
.B(n_341),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_334),
.B(n_335),
.Y(n_333)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

OR2x2_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_345),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_344),
.B(n_345),
.Y(n_350)
);

INVx1_ASAP7_75t_SL g348 ( 
.A(n_349),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_358),
.Y(n_352)
);

NOR2xp67_ASAP7_75t_L g365 ( 
.A(n_353),
.B(n_358),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_356),
.C(n_357),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_362),
.Y(n_358)
);

HB1xp67_ASAP7_75t_L g368 ( 
.A(n_359),
.Y(n_368)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_363),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_369),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_367),
.B(n_369),
.Y(n_371)
);

INVxp67_ASAP7_75t_SL g372 ( 
.A(n_373),
.Y(n_372)
);


endmodule