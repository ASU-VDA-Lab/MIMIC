module real_aes_9744_n_281 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_281);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_281;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_1199;
wire n_951;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_1537;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1589;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1346;
wire n_1383;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_1600;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1583;
wire n_360;
wire n_1284;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1628;
wire n_1587;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1615;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1510;
wire n_1495;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_1488;
wire n_337;
wire n_1572;
wire n_1514;
wire n_480;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1616;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1542;
wire n_1392;
wire n_665;
wire n_991;
wire n_667;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_1260;
wire n_328;
wire n_1606;
wire n_355;
wire n_1129;
wire n_1285;
wire n_1014;
wire n_742;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1594;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_1269;
wire n_677;
wire n_378;
wire n_591;
wire n_1518;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_1361;
wire n_510;
wire n_1358;
wire n_1577;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1612;
wire n_1479;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_1614;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_733;
wire n_402;
wire n_602;
wire n_1404;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_286;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1620;
wire n_985;
wire n_777;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_334;
wire n_1179;
wire n_1171;
wire n_569;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1580;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_1023;
wire n_419;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_282;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_300;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1133;
wire n_1593;
wire n_313;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_285;
wire n_1377;
wire n_800;
wire n_778;
wire n_1175;
wire n_1170;
wire n_522;
wire n_1475;
wire n_943;
wire n_977;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1268;
wire n_1113;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_936;
wire n_581;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_502;
wire n_769;
wire n_434;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1603;
wire n_1450;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_288;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1605;
wire n_1592;
wire n_1056;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_295;
wire n_845;
wire n_1619;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1617;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1466;
wire n_921;
wire n_1396;
wire n_640;
wire n_1176;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_1211;
wire n_650;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1480;
wire n_1101;
wire n_1251;
wire n_1076;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1596;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_364;
wire n_319;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_317;
wire n_1595;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1541;
wire n_1272;
wire n_408;
wire n_892;
wire n_372;
wire n_578;
wire n_938;
wire n_327;
wire n_774;
wire n_559;
wire n_1584;
wire n_466;
wire n_1277;
wire n_1049;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_1527;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_1100;
wire n_398;
wire n_1519;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_302;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1573;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_1300;
wire n_575;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_1630;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_1097;
wire n_703;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
AOI21xp33_ASAP7_75t_L g1083 ( .A1(n_0), .A2(n_566), .B(n_771), .Y(n_1083) );
INVx1_ASAP7_75t_L g1103 ( .A(n_0), .Y(n_1103) );
INVx1_ASAP7_75t_L g892 ( .A(n_1), .Y(n_892) );
OAI221xp5_ASAP7_75t_L g921 ( .A1(n_1), .A2(n_28), .B1(n_922), .B2(n_923), .C(n_924), .Y(n_921) );
AOI22xp33_ASAP7_75t_L g1314 ( .A1(n_2), .A2(n_69), .B1(n_1278), .B2(n_1305), .Y(n_1314) );
AOI222xp33_ASAP7_75t_L g1517 ( .A1(n_2), .A2(n_1518), .B1(n_1564), .B2(n_1568), .C1(n_1623), .C2(n_1627), .Y(n_1517) );
XNOR2xp5_ASAP7_75t_L g1522 ( .A(n_2), .B(n_1523), .Y(n_1522) );
HB1xp67_ASAP7_75t_L g295 ( .A(n_3), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_3), .B(n_215), .Y(n_318) );
AND2x2_ASAP7_75t_L g339 ( .A(n_3), .B(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g385 ( .A(n_3), .Y(n_385) );
CKINVDCx5p33_ASAP7_75t_R g537 ( .A(n_4), .Y(n_537) );
OAI221xp5_ASAP7_75t_L g1125 ( .A1(n_5), .A2(n_494), .B1(n_515), .B2(n_1126), .C(n_1132), .Y(n_1125) );
INVx1_ASAP7_75t_L g1147 ( .A(n_5), .Y(n_1147) );
XNOR2x2_ASAP7_75t_L g829 ( .A(n_6), .B(n_830), .Y(n_829) );
OAI22xp33_ASAP7_75t_L g1545 ( .A1(n_7), .A2(n_94), .B1(n_751), .B2(n_754), .Y(n_1545) );
INVx1_ASAP7_75t_L g1557 ( .A(n_7), .Y(n_1557) );
AOI221xp5_ASAP7_75t_L g1123 ( .A1(n_8), .A2(n_57), .B1(n_343), .B2(n_364), .C(n_530), .Y(n_1123) );
INVx1_ASAP7_75t_L g1152 ( .A(n_8), .Y(n_1152) );
INVx1_ASAP7_75t_L g1118 ( .A(n_9), .Y(n_1118) );
AOI22xp33_ASAP7_75t_L g1149 ( .A1(n_9), .A2(n_58), .B1(n_408), .B2(n_433), .Y(n_1149) );
INVx1_ASAP7_75t_L g978 ( .A(n_10), .Y(n_978) );
AO22x2_ASAP7_75t_L g1156 ( .A1(n_11), .A2(n_1157), .B1(n_1213), .B2(n_1214), .Y(n_1156) );
CKINVDCx14_ASAP7_75t_R g1213 ( .A(n_11), .Y(n_1213) );
AOI22xp33_ASAP7_75t_L g710 ( .A1(n_12), .A2(n_91), .B1(n_711), .B2(n_712), .Y(n_710) );
OAI22xp5_ASAP7_75t_L g747 ( .A1(n_12), .A2(n_31), .B1(n_490), .B2(n_517), .Y(n_747) );
AOI22xp33_ASAP7_75t_SL g895 ( .A1(n_13), .A2(n_246), .B1(n_748), .B2(n_896), .Y(n_895) );
AOI221xp5_ASAP7_75t_L g931 ( .A1(n_13), .A2(n_75), .B1(n_450), .B2(n_770), .C(n_932), .Y(n_931) );
CKINVDCx5p33_ASAP7_75t_R g539 ( .A(n_14), .Y(n_539) );
AOI22xp33_ASAP7_75t_L g897 ( .A1(n_15), .A2(n_75), .B1(n_898), .B2(n_900), .Y(n_897) );
AOI22xp33_ASAP7_75t_L g933 ( .A1(n_15), .A2(n_246), .B1(n_774), .B2(n_788), .Y(n_933) );
AOI22xp5_ASAP7_75t_L g1308 ( .A1(n_16), .A2(n_81), .B1(n_1304), .B2(n_1305), .Y(n_1308) );
INVx1_ASAP7_75t_L g1533 ( .A(n_17), .Y(n_1533) );
AOI221xp5_ASAP7_75t_L g768 ( .A1(n_18), .A2(n_241), .B1(n_769), .B2(n_770), .C(n_771), .Y(n_768) );
INVx1_ASAP7_75t_L g801 ( .A(n_18), .Y(n_801) );
OAI221xp5_ASAP7_75t_L g1065 ( .A1(n_19), .A2(n_1014), .B1(n_1066), .B2(n_1070), .C(n_1074), .Y(n_1065) );
AOI22xp33_ASAP7_75t_L g1097 ( .A1(n_19), .A2(n_193), .B1(n_741), .B2(n_1098), .Y(n_1097) );
CKINVDCx5p33_ASAP7_75t_R g1133 ( .A(n_20), .Y(n_1133) );
INVx1_ASAP7_75t_L g502 ( .A(n_21), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_21), .A2(n_243), .B1(n_587), .B2(n_588), .Y(n_586) );
INVx2_ASAP7_75t_L g399 ( .A(n_22), .Y(n_399) );
OR2x2_ASAP7_75t_L g412 ( .A(n_22), .B(n_397), .Y(n_412) );
AOI221xp5_ASAP7_75t_L g739 ( .A1(n_23), .A2(n_166), .B1(n_530), .B2(n_740), .C(n_741), .Y(n_739) );
OAI22xp5_ASAP7_75t_L g757 ( .A1(n_23), .A2(n_240), .B1(n_562), .B2(n_758), .Y(n_757) );
AO22x1_ASAP7_75t_L g1113 ( .A1(n_24), .A2(n_1114), .B1(n_1154), .B2(n_1155), .Y(n_1113) );
INVx1_ASAP7_75t_L g1155 ( .A(n_24), .Y(n_1155) );
AOI22xp33_ASAP7_75t_L g706 ( .A1(n_25), .A2(n_66), .B1(n_641), .B2(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g734 ( .A(n_25), .Y(n_734) );
OAI22xp5_ASAP7_75t_L g1025 ( .A1(n_26), .A2(n_253), .B1(n_923), .B2(n_1026), .Y(n_1025) );
OAI221xp5_ASAP7_75t_L g1040 ( .A1(n_26), .A2(n_253), .B1(n_805), .B2(n_1041), .C(n_1042), .Y(n_1040) );
AOI22xp5_ASAP7_75t_L g1307 ( .A1(n_27), .A2(n_140), .B1(n_1294), .B2(n_1300), .Y(n_1307) );
INVx1_ASAP7_75t_L g891 ( .A(n_28), .Y(n_891) );
AOI221xp5_ASAP7_75t_L g621 ( .A1(n_29), .A2(n_110), .B1(n_597), .B2(n_622), .C(n_624), .Y(n_621) );
INVx1_ASAP7_75t_L g655 ( .A(n_29), .Y(n_655) );
OR2x2_ASAP7_75t_L g317 ( .A(n_30), .B(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g338 ( .A(n_30), .Y(n_338) );
BUFx2_ASAP7_75t_L g360 ( .A(n_30), .Y(n_360) );
BUFx2_ASAP7_75t_L g393 ( .A(n_30), .Y(n_393) );
OAI222xp33_ASAP7_75t_L g750 ( .A1(n_31), .A2(n_166), .B1(n_170), .B2(n_391), .C1(n_751), .C2(n_754), .Y(n_750) );
INVx1_ASAP7_75t_L g1340 ( .A(n_32), .Y(n_1340) );
OAI22xp33_ASAP7_75t_L g1244 ( .A1(n_33), .A2(n_182), .B1(n_881), .B2(n_882), .Y(n_1244) );
INVx1_ASAP7_75t_L g1269 ( .A(n_33), .Y(n_1269) );
INVx1_ASAP7_75t_L g1160 ( .A(n_34), .Y(n_1160) );
AOI21xp33_ASAP7_75t_L g1204 ( .A1(n_34), .A2(n_408), .B(n_1205), .Y(n_1204) );
AOI221xp5_ASAP7_75t_L g635 ( .A1(n_35), .A2(n_172), .B1(n_591), .B2(n_636), .C(n_638), .Y(n_635) );
INVx1_ASAP7_75t_L g678 ( .A(n_35), .Y(n_678) );
CKINVDCx5p33_ASAP7_75t_R g1172 ( .A(n_36), .Y(n_1172) );
CKINVDCx5p33_ASAP7_75t_R g528 ( .A(n_37), .Y(n_528) );
OAI22xp5_ASAP7_75t_L g777 ( .A1(n_38), .A2(n_74), .B1(n_415), .B2(n_778), .Y(n_777) );
OAI221xp5_ASAP7_75t_L g803 ( .A1(n_38), .A2(n_74), .B1(n_670), .B2(n_804), .C(n_805), .Y(n_803) );
AOI22xp33_ASAP7_75t_L g1082 ( .A1(n_39), .A2(n_151), .B1(n_408), .B2(n_433), .Y(n_1082) );
INVx1_ASAP7_75t_L g1104 ( .A(n_39), .Y(n_1104) );
INVx1_ASAP7_75t_L g980 ( .A(n_40), .Y(n_980) );
INVx1_ASAP7_75t_L g1364 ( .A(n_41), .Y(n_1364) );
AOI22xp33_ASAP7_75t_L g1017 ( .A1(n_42), .A2(n_221), .B1(n_711), .B2(n_1018), .Y(n_1017) );
INVx1_ASAP7_75t_L g1047 ( .A(n_42), .Y(n_1047) );
OAI221xp5_ASAP7_75t_L g1206 ( .A1(n_43), .A2(n_236), .B1(n_420), .B2(n_1207), .C(n_1208), .Y(n_1206) );
INVx1_ASAP7_75t_L g1211 ( .A(n_43), .Y(n_1211) );
AOI22xp33_ASAP7_75t_SL g1592 ( .A1(n_44), .A2(n_111), .B1(n_1593), .B2(n_1594), .Y(n_1592) );
AOI221xp5_ASAP7_75t_L g1614 ( .A1(n_44), .A2(n_72), .B1(n_455), .B2(n_1615), .C(n_1617), .Y(n_1614) );
AOI22xp33_ASAP7_75t_L g903 ( .A1(n_45), .A2(n_54), .B1(n_904), .B2(n_906), .Y(n_903) );
INVx1_ASAP7_75t_L g935 ( .A(n_45), .Y(n_935) );
INVx1_ASAP7_75t_L g1131 ( .A(n_46), .Y(n_1131) );
AOI22xp33_ASAP7_75t_L g1142 ( .A1(n_46), .A2(n_156), .B1(n_432), .B2(n_433), .Y(n_1142) );
OAI22xp5_ASAP7_75t_L g1124 ( .A1(n_47), .A2(n_173), .B1(n_546), .B2(n_744), .Y(n_1124) );
OAI22xp5_ASAP7_75t_SL g1139 ( .A1(n_47), .A2(n_173), .B1(n_575), .B2(n_580), .Y(n_1139) );
AOI22xp33_ASAP7_75t_L g834 ( .A1(n_48), .A2(n_52), .B1(n_835), .B2(n_837), .Y(n_834) );
OAI22xp5_ASAP7_75t_L g886 ( .A1(n_48), .A2(n_71), .B1(n_562), .B2(n_758), .Y(n_886) );
CKINVDCx5p33_ASAP7_75t_R g630 ( .A(n_49), .Y(n_630) );
INVx1_ASAP7_75t_L g720 ( .A(n_50), .Y(n_720) );
OAI221xp5_ASAP7_75t_L g743 ( .A1(n_50), .A2(n_92), .B1(n_546), .B2(n_744), .C(n_746), .Y(n_743) );
AOI22xp33_ASAP7_75t_L g1241 ( .A1(n_51), .A2(n_84), .B1(n_461), .B2(n_1242), .Y(n_1241) );
OAI22xp5_ASAP7_75t_L g1246 ( .A1(n_51), .A2(n_84), .B1(n_485), .B2(n_487), .Y(n_1246) );
INVxp67_ASAP7_75t_SL g884 ( .A(n_52), .Y(n_884) );
AOI22xp33_ASAP7_75t_L g1293 ( .A1(n_53), .A2(n_105), .B1(n_1294), .B2(n_1300), .Y(n_1293) );
INVx1_ASAP7_75t_L g930 ( .A(n_54), .Y(n_930) );
OAI22xp33_ASAP7_75t_L g1084 ( .A1(n_55), .A2(n_193), .B1(n_470), .B2(n_474), .Y(n_1084) );
AOI22xp33_ASAP7_75t_L g1095 ( .A1(n_55), .A2(n_275), .B1(n_1092), .B2(n_1096), .Y(n_1095) );
INVx1_ASAP7_75t_L g856 ( .A(n_56), .Y(n_856) );
OAI22xp5_ASAP7_75t_L g1153 ( .A1(n_57), .A2(n_115), .B1(n_559), .B2(n_562), .Y(n_1153) );
INVx1_ASAP7_75t_L g1119 ( .A(n_58), .Y(n_1119) );
XNOR2xp5_ASAP7_75t_L g1569 ( .A(n_59), .B(n_1570), .Y(n_1569) );
AOI22xp33_ASAP7_75t_SL g362 ( .A1(n_60), .A2(n_116), .B1(n_363), .B2(n_366), .Y(n_362) );
AOI221xp5_ASAP7_75t_L g447 ( .A1(n_60), .A2(n_145), .B1(n_448), .B2(n_451), .C(n_455), .Y(n_447) );
AOI221xp5_ASAP7_75t_L g1016 ( .A1(n_61), .A2(n_80), .B1(n_450), .B2(n_638), .C(n_770), .Y(n_1016) );
INVxp67_ASAP7_75t_SL g1050 ( .A(n_61), .Y(n_1050) );
AO22x2_ASAP7_75t_L g480 ( .A1(n_62), .A2(n_481), .B1(n_482), .B2(n_609), .Y(n_480) );
INVx1_ASAP7_75t_L g609 ( .A(n_62), .Y(n_609) );
INVx1_ASAP7_75t_L g956 ( .A(n_63), .Y(n_956) );
AOI22xp33_ASAP7_75t_L g1230 ( .A1(n_64), .A2(n_152), .B1(n_1231), .B2(n_1232), .Y(n_1230) );
INVxp67_ASAP7_75t_SL g1254 ( .A(n_64), .Y(n_1254) );
CKINVDCx5p33_ASAP7_75t_R g541 ( .A(n_65), .Y(n_541) );
INVx1_ASAP7_75t_L g732 ( .A(n_66), .Y(n_732) );
OAI221xp5_ASAP7_75t_L g959 ( .A1(n_67), .A2(n_232), .B1(n_661), .B2(n_666), .C(n_669), .Y(n_959) );
OAI22xp5_ASAP7_75t_L g987 ( .A1(n_67), .A2(n_232), .B1(n_420), .B2(n_988), .Y(n_987) );
INVxp67_ASAP7_75t_L g970 ( .A(n_68), .Y(n_970) );
AOI22xp33_ASAP7_75t_L g1000 ( .A1(n_68), .A2(n_128), .B1(n_458), .B2(n_1001), .Y(n_1000) );
AOI22xp33_ASAP7_75t_L g625 ( .A1(n_70), .A2(n_197), .B1(n_626), .B2(n_627), .Y(n_625) );
INVx1_ASAP7_75t_L g653 ( .A(n_70), .Y(n_653) );
AOI221xp5_ASAP7_75t_L g840 ( .A1(n_71), .A2(n_203), .B1(n_530), .B2(n_841), .C(n_843), .Y(n_840) );
AOI22xp33_ASAP7_75t_L g1589 ( .A1(n_72), .A2(n_139), .B1(n_1590), .B2(n_1591), .Y(n_1589) );
AOI22xp5_ASAP7_75t_L g1316 ( .A1(n_73), .A2(n_120), .B1(n_1294), .B2(n_1300), .Y(n_1316) );
INVxp33_ASAP7_75t_SL g331 ( .A(n_76), .Y(n_331) );
AOI22xp33_ASAP7_75t_SL g431 ( .A1(n_76), .A2(n_217), .B1(n_432), .B2(n_433), .Y(n_431) );
OAI22xp5_ASAP7_75t_L g484 ( .A1(n_77), .A2(n_205), .B1(n_485), .B2(n_487), .Y(n_484) );
AOI22xp33_ASAP7_75t_SL g598 ( .A1(n_77), .A2(n_205), .B1(n_599), .B2(n_600), .Y(n_598) );
AOI22xp33_ASAP7_75t_L g787 ( .A1(n_78), .A2(n_268), .B1(n_788), .B2(n_789), .Y(n_787) );
INVx1_ASAP7_75t_L g811 ( .A(n_78), .Y(n_811) );
CKINVDCx5p33_ASAP7_75t_R g525 ( .A(n_79), .Y(n_525) );
INVxp67_ASAP7_75t_SL g1054 ( .A(n_80), .Y(n_1054) );
INVxp67_ASAP7_75t_SL g324 ( .A(n_82), .Y(n_324) );
OAI221xp5_ASAP7_75t_L g414 ( .A1(n_82), .A2(n_225), .B1(n_415), .B2(n_420), .C(n_424), .Y(n_414) );
AOI22xp33_ASAP7_75t_SL g1597 ( .A1(n_83), .A2(n_95), .B1(n_377), .B2(n_1598), .Y(n_1597) );
INVx1_ASAP7_75t_L g1613 ( .A(n_83), .Y(n_1613) );
INVx1_ASAP7_75t_L g1584 ( .A(n_85), .Y(n_1584) );
AOI221xp5_ASAP7_75t_L g1608 ( .A1(n_85), .A2(n_108), .B1(n_1609), .B2(n_1610), .C(n_1611), .Y(n_1608) );
CKINVDCx5p33_ASAP7_75t_R g544 ( .A(n_86), .Y(n_544) );
CKINVDCx5p33_ASAP7_75t_R g642 ( .A(n_87), .Y(n_642) );
AOI22xp33_ASAP7_75t_L g1596 ( .A1(n_88), .A2(n_231), .B1(n_686), .B2(n_1594), .Y(n_1596) );
INVx1_ASAP7_75t_L g1622 ( .A(n_88), .Y(n_1622) );
INVx1_ASAP7_75t_L g397 ( .A(n_89), .Y(n_397) );
INVx1_ASAP7_75t_L g440 ( .A(n_89), .Y(n_440) );
INVx1_ASAP7_75t_L g1011 ( .A(n_90), .Y(n_1011) );
INVx1_ASAP7_75t_L g742 ( .A(n_91), .Y(n_742) );
INVx1_ASAP7_75t_L g719 ( .A(n_92), .Y(n_719) );
INVx1_ASAP7_75t_L g1237 ( .A(n_93), .Y(n_1237) );
OAI221xp5_ASAP7_75t_L g1247 ( .A1(n_93), .A2(n_494), .B1(n_861), .B2(n_1248), .C(n_1251), .Y(n_1247) );
AOI221xp5_ASAP7_75t_L g1559 ( .A1(n_94), .A2(n_227), .B1(n_343), .B2(n_347), .C(n_1560), .Y(n_1559) );
INVx1_ASAP7_75t_L g1621 ( .A(n_95), .Y(n_1621) );
INVx1_ASAP7_75t_L g1071 ( .A(n_96), .Y(n_1071) );
AOI22xp33_ASAP7_75t_L g1089 ( .A1(n_96), .A2(n_171), .B1(n_741), .B2(n_1090), .Y(n_1089) );
INVx1_ASAP7_75t_L g1262 ( .A(n_97), .Y(n_1262) );
OAI22xp5_ASAP7_75t_L g1271 ( .A1(n_97), .A2(n_125), .B1(n_559), .B2(n_562), .Y(n_1271) );
OAI221xp5_ASAP7_75t_L g519 ( .A1(n_98), .A2(n_520), .B1(n_523), .B2(n_532), .C(n_540), .Y(n_519) );
AOI22xp33_ASAP7_75t_SL g593 ( .A1(n_98), .A2(n_134), .B1(n_594), .B2(n_597), .Y(n_593) );
AOI22xp5_ASAP7_75t_L g1313 ( .A1(n_99), .A2(n_126), .B1(n_1294), .B2(n_1300), .Y(n_1313) );
INVx1_ASAP7_75t_L g859 ( .A(n_100), .Y(n_859) );
AOI221xp5_ASAP7_75t_L g865 ( .A1(n_100), .A2(n_272), .B1(n_590), .B2(n_866), .C(n_868), .Y(n_865) );
AOI22xp33_ASAP7_75t_L g1330 ( .A1(n_101), .A2(n_226), .B1(n_1294), .B2(n_1300), .Y(n_1330) );
INVxp67_ASAP7_75t_L g965 ( .A(n_102), .Y(n_965) );
AOI221xp5_ASAP7_75t_L g995 ( .A1(n_102), .A2(n_124), .B1(n_455), .B2(n_996), .C(n_998), .Y(n_995) );
INVxp33_ASAP7_75t_SL g345 ( .A(n_103), .Y(n_345) );
AOI21xp33_ASAP7_75t_L g435 ( .A1(n_103), .A2(n_436), .B(n_438), .Y(n_435) );
AOI22xp5_ASAP7_75t_L g1303 ( .A1(n_104), .A2(n_144), .B1(n_1304), .B2(n_1305), .Y(n_1303) );
OAI22xp5_ASAP7_75t_L g1061 ( .A1(n_105), .A2(n_1062), .B1(n_1108), .B2(n_1109), .Y(n_1061) );
INVxp67_ASAP7_75t_SL g1108 ( .A(n_105), .Y(n_1108) );
INVx1_ASAP7_75t_L g1535 ( .A(n_106), .Y(n_1535) );
OAI221xp5_ASAP7_75t_L g1550 ( .A1(n_106), .A2(n_494), .B1(n_861), .B2(n_1551), .C(n_1553), .Y(n_1550) );
INVx1_ASAP7_75t_L g1322 ( .A(n_107), .Y(n_1322) );
INVx1_ASAP7_75t_L g1579 ( .A(n_108), .Y(n_1579) );
AOI22xp33_ASAP7_75t_SL g708 ( .A1(n_109), .A2(n_176), .B1(n_607), .B2(n_709), .Y(n_708) );
AOI21xp33_ASAP7_75t_L g730 ( .A1(n_109), .A2(n_554), .B(n_673), .Y(n_730) );
INVx1_ASAP7_75t_L g657 ( .A(n_110), .Y(n_657) );
AOI22xp33_ASAP7_75t_L g1618 ( .A1(n_111), .A2(n_139), .B1(n_594), .B2(n_1619), .Y(n_1618) );
AOI221xp5_ASAP7_75t_L g1263 ( .A1(n_112), .A2(n_125), .B1(n_375), .B2(n_377), .C(n_1264), .Y(n_1263) );
OAI22xp5_ASAP7_75t_L g1272 ( .A1(n_112), .A2(n_209), .B1(n_751), .B2(n_754), .Y(n_1272) );
AOI22xp33_ASAP7_75t_L g1022 ( .A1(n_113), .A2(n_247), .B1(n_1023), .B2(n_1024), .Y(n_1022) );
INVx1_ASAP7_75t_L g1038 ( .A(n_113), .Y(n_1038) );
AOI22xp33_ASAP7_75t_L g374 ( .A1(n_114), .A2(n_175), .B1(n_375), .B2(n_377), .Y(n_374) );
INVxp33_ASAP7_75t_SL g468 ( .A(n_114), .Y(n_468) );
AOI22xp33_ASAP7_75t_L g1121 ( .A1(n_115), .A2(n_135), .B1(n_738), .B2(n_1122), .Y(n_1121) );
AOI22xp33_ASAP7_75t_L g457 ( .A1(n_116), .A2(n_119), .B1(n_458), .B2(n_460), .Y(n_457) );
INVxp33_ASAP7_75t_L g952 ( .A(n_117), .Y(n_952) );
AOI221xp5_ASAP7_75t_L g989 ( .A1(n_117), .A2(n_155), .B1(n_588), .B2(n_990), .C(n_991), .Y(n_989) );
AOI221xp5_ASAP7_75t_L g1021 ( .A1(n_118), .A2(n_230), .B1(n_566), .B2(n_770), .C(n_771), .Y(n_1021) );
INVx1_ASAP7_75t_L g1037 ( .A(n_118), .Y(n_1037) );
AOI22xp33_ASAP7_75t_L g368 ( .A1(n_119), .A2(n_145), .B1(n_369), .B2(n_370), .Y(n_368) );
INVx1_ASAP7_75t_L g513 ( .A(n_121), .Y(n_513) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_121), .A2(n_143), .B1(n_590), .B2(n_591), .Y(n_589) );
INVx1_ASAP7_75t_L g287 ( .A(n_122), .Y(n_287) );
INVx1_ASAP7_75t_L g479 ( .A(n_123), .Y(n_479) );
AO22x1_ASAP7_75t_SL g1319 ( .A1(n_123), .A2(n_233), .B1(n_1294), .B2(n_1300), .Y(n_1319) );
INVxp67_ASAP7_75t_L g967 ( .A(n_124), .Y(n_967) );
CKINVDCx5p33_ASAP7_75t_R g792 ( .A(n_127), .Y(n_792) );
INVx1_ASAP7_75t_L g962 ( .A(n_128), .Y(n_962) );
AOI22xp33_ASAP7_75t_L g373 ( .A1(n_129), .A2(n_192), .B1(n_369), .B2(n_370), .Y(n_373) );
INVxp67_ASAP7_75t_SL g413 ( .A(n_129), .Y(n_413) );
INVx1_ASAP7_75t_L g826 ( .A(n_130), .Y(n_826) );
AOI22xp33_ASAP7_75t_L g901 ( .A1(n_131), .A2(n_204), .B1(n_835), .B2(n_902), .Y(n_901) );
INVx1_ASAP7_75t_L g936 ( .A(n_131), .Y(n_936) );
CKINVDCx5p33_ASAP7_75t_R g1169 ( .A(n_132), .Y(n_1169) );
AOI22xp33_ASAP7_75t_L g772 ( .A1(n_133), .A2(n_206), .B1(n_773), .B2(n_774), .Y(n_772) );
INVx1_ASAP7_75t_L g798 ( .A(n_133), .Y(n_798) );
OAI221xp5_ASAP7_75t_L g493 ( .A1(n_134), .A2(n_494), .B1(n_496), .B2(n_505), .C(n_515), .Y(n_493) );
INVx1_ASAP7_75t_L g1151 ( .A(n_135), .Y(n_1151) );
INVx1_ASAP7_75t_L g954 ( .A(n_136), .Y(n_954) );
AO221x2_ASAP7_75t_L g1334 ( .A1(n_137), .A2(n_270), .B1(n_1278), .B2(n_1335), .C(n_1336), .Y(n_1334) );
INVx1_ASAP7_75t_L g1536 ( .A(n_138), .Y(n_1536) );
OAI211xp5_ASAP7_75t_SL g1554 ( .A1(n_138), .A2(n_520), .B(n_1555), .C(n_1561), .Y(n_1554) );
INVx1_ASAP7_75t_L g341 ( .A(n_141), .Y(n_341) );
INVx1_ASAP7_75t_L g863 ( .A(n_142), .Y(n_863) );
INVx1_ASAP7_75t_L g510 ( .A(n_143), .Y(n_510) );
CKINVDCx5p33_ASAP7_75t_R g910 ( .A(n_146), .Y(n_910) );
CKINVDCx5p33_ASAP7_75t_R g1175 ( .A(n_147), .Y(n_1175) );
INVx1_ASAP7_75t_L g938 ( .A(n_148), .Y(n_938) );
XNOR2xp5_ASAP7_75t_L g699 ( .A(n_149), .B(n_700), .Y(n_699) );
CKINVDCx5p33_ASAP7_75t_R g1078 ( .A(n_150), .Y(n_1078) );
OAI22xp5_ASAP7_75t_L g1105 ( .A1(n_151), .A2(n_261), .B1(n_1106), .B2(n_1107), .Y(n_1105) );
INVxp67_ASAP7_75t_SL g1258 ( .A(n_152), .Y(n_1258) );
INVx1_ASAP7_75t_L g1600 ( .A(n_153), .Y(n_1600) );
CKINVDCx5p33_ASAP7_75t_R g791 ( .A(n_154), .Y(n_791) );
INVxp33_ASAP7_75t_L g957 ( .A(n_155), .Y(n_957) );
INVx1_ASAP7_75t_L g1129 ( .A(n_156), .Y(n_1129) );
INVx1_ASAP7_75t_L g908 ( .A(n_157), .Y(n_908) );
AOI22xp33_ASAP7_75t_L g926 ( .A1(n_157), .A2(n_242), .B1(n_409), .B2(n_629), .Y(n_926) );
INVx1_ASAP7_75t_L g1240 ( .A(n_158), .Y(n_1240) );
OAI211xp5_ASAP7_75t_SL g1259 ( .A1(n_158), .A2(n_520), .B(n_1260), .C(n_1265), .Y(n_1259) );
INVx1_ASAP7_75t_L g1161 ( .A(n_159), .Y(n_1161) );
AOI22xp33_ASAP7_75t_SL g1202 ( .A1(n_159), .A2(n_207), .B1(n_433), .B2(n_1203), .Y(n_1202) );
AOI22xp5_ASAP7_75t_L g1331 ( .A1(n_160), .A2(n_263), .B1(n_1304), .B2(n_1305), .Y(n_1331) );
CKINVDCx5p33_ASAP7_75t_R g1532 ( .A(n_161), .Y(n_1532) );
CKINVDCx5p33_ASAP7_75t_R g1583 ( .A(n_162), .Y(n_1583) );
OAI22xp33_ASAP7_75t_L g1541 ( .A1(n_163), .A2(n_238), .B1(n_882), .B2(n_1542), .Y(n_1541) );
INVx1_ASAP7_75t_L g1563 ( .A(n_163), .Y(n_1563) );
OAI22xp5_ASAP7_75t_L g846 ( .A1(n_164), .A2(n_188), .B1(n_546), .B2(n_744), .Y(n_846) );
OAI221xp5_ASAP7_75t_L g880 ( .A1(n_164), .A2(n_188), .B1(n_606), .B2(n_881), .C(n_882), .Y(n_880) );
CKINVDCx5p33_ASAP7_75t_R g782 ( .A(n_165), .Y(n_782) );
INVx1_ASAP7_75t_L g1538 ( .A(n_167), .Y(n_1538) );
OAI22xp5_ASAP7_75t_L g1549 ( .A1(n_167), .A2(n_267), .B1(n_485), .B2(n_487), .Y(n_1549) );
INVx1_ASAP7_75t_L g1015 ( .A(n_168), .Y(n_1015) );
CKINVDCx5p33_ASAP7_75t_R g549 ( .A(n_169), .Y(n_549) );
AOI22xp33_ASAP7_75t_L g736 ( .A1(n_170), .A2(n_240), .B1(n_737), .B2(n_738), .Y(n_736) );
INVx1_ASAP7_75t_L g1068 ( .A(n_171), .Y(n_1068) );
INVx1_ASAP7_75t_L g683 ( .A(n_172), .Y(n_683) );
AOI22xp33_ASAP7_75t_SL g714 ( .A1(n_174), .A2(n_183), .B1(n_461), .B2(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g724 ( .A(n_174), .Y(n_724) );
INVxp67_ASAP7_75t_SL g446 ( .A(n_175), .Y(n_446) );
INVx1_ASAP7_75t_L g729 ( .A(n_176), .Y(n_729) );
OAI22xp5_ASAP7_75t_L g1184 ( .A1(n_177), .A2(n_235), .B1(n_390), .B2(n_1106), .Y(n_1184) );
AOI22xp33_ASAP7_75t_SL g1197 ( .A1(n_177), .A2(n_202), .B1(n_408), .B2(n_433), .Y(n_1197) );
AOI221xp5_ASAP7_75t_L g783 ( .A1(n_178), .A2(n_244), .B1(n_638), .B2(n_784), .C(n_786), .Y(n_783) );
INVx1_ASAP7_75t_L g817 ( .A(n_178), .Y(n_817) );
AOI21xp33_ASAP7_75t_L g1073 ( .A1(n_179), .A2(n_432), .B(n_455), .Y(n_1073) );
AOI22xp33_ASAP7_75t_L g1091 ( .A1(n_179), .A2(n_260), .B1(n_1092), .B2(n_1093), .Y(n_1091) );
OAI22xp5_ASAP7_75t_L g1181 ( .A1(n_180), .A2(n_202), .B1(n_1182), .B2(n_1183), .Y(n_1181) );
INVx1_ASAP7_75t_L g1193 ( .A(n_180), .Y(n_1193) );
CKINVDCx5p33_ASAP7_75t_R g1219 ( .A(n_181), .Y(n_1219) );
INVx1_ASAP7_75t_L g1268 ( .A(n_182), .Y(n_1268) );
INVx1_ASAP7_75t_L g725 ( .A(n_183), .Y(n_725) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_184), .Y(n_289) );
AND3x2_ASAP7_75t_L g1282 ( .A(n_184), .B(n_287), .C(n_1283), .Y(n_1282) );
NAND2xp5_ASAP7_75t_L g1299 ( .A(n_184), .B(n_287), .Y(n_1299) );
CKINVDCx5p33_ASAP7_75t_R g1170 ( .A(n_185), .Y(n_1170) );
OA332x1_ASAP7_75t_L g1158 ( .A1(n_186), .A2(n_672), .A3(n_1159), .B1(n_1164), .B2(n_1168), .B3(n_1171), .C1(n_1177), .C2(n_1178), .Y(n_1158) );
AOI21xp5_ASAP7_75t_L g1198 ( .A1(n_186), .A2(n_771), .B(n_1199), .Y(n_1198) );
AOI22xp33_ASAP7_75t_L g1317 ( .A1(n_187), .A2(n_252), .B1(n_1278), .B2(n_1305), .Y(n_1317) );
INVx2_ASAP7_75t_L g300 ( .A(n_189), .Y(n_300) );
INVx1_ASAP7_75t_L g1027 ( .A(n_190), .Y(n_1027) );
INVx1_ASAP7_75t_L g975 ( .A(n_191), .Y(n_975) );
INVxp33_ASAP7_75t_SL g472 ( .A(n_192), .Y(n_472) );
OAI22xp33_ASAP7_75t_L g1544 ( .A1(n_194), .A2(n_227), .B1(n_559), .B2(n_562), .Y(n_1544) );
INVx1_ASAP7_75t_L g1558 ( .A(n_194), .Y(n_1558) );
OAI211xp5_ASAP7_75t_L g1116 ( .A1(n_195), .A2(n_520), .B(n_1117), .C(n_1120), .Y(n_1116) );
INVx1_ASAP7_75t_L g1148 ( .A(n_195), .Y(n_1148) );
AOI22xp33_ASAP7_75t_L g640 ( .A1(n_196), .A2(n_239), .B1(n_458), .B2(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g676 ( .A(n_196), .Y(n_676) );
INVx1_ASAP7_75t_L g658 ( .A(n_197), .Y(n_658) );
INVx1_ASAP7_75t_L g1324 ( .A(n_198), .Y(n_1324) );
CKINVDCx5p33_ASAP7_75t_R g1077 ( .A(n_199), .Y(n_1077) );
INVx1_ASAP7_75t_L g854 ( .A(n_200), .Y(n_854) );
INVx1_ASAP7_75t_L g1283 ( .A(n_201), .Y(n_1283) );
INVxp67_ASAP7_75t_SL g885 ( .A(n_203), .Y(n_885) );
INVx1_ASAP7_75t_L g920 ( .A(n_204), .Y(n_920) );
INVx1_ASAP7_75t_L g802 ( .A(n_206), .Y(n_802) );
INVx1_ASAP7_75t_L g1165 ( .A(n_207), .Y(n_1165) );
CKINVDCx5p33_ASAP7_75t_R g937 ( .A(n_208), .Y(n_937) );
INVx1_ASAP7_75t_L g1261 ( .A(n_209), .Y(n_1261) );
OAI211xp5_ASAP7_75t_L g832 ( .A1(n_210), .A2(n_520), .B(n_833), .C(n_847), .Y(n_832) );
AOI221xp5_ASAP7_75t_L g871 ( .A1(n_210), .A2(n_219), .B1(n_872), .B2(n_874), .C(n_875), .Y(n_871) );
OAI22xp33_ASAP7_75t_L g631 ( .A1(n_211), .A2(n_213), .B1(n_420), .B2(n_632), .Y(n_631) );
OAI221xp5_ASAP7_75t_L g660 ( .A1(n_211), .A2(n_213), .B1(n_661), .B2(n_666), .C(n_669), .Y(n_660) );
CKINVDCx5p33_ASAP7_75t_R g767 ( .A(n_212), .Y(n_767) );
CKINVDCx20_ASAP7_75t_R g1337 ( .A(n_214), .Y(n_1337) );
INVx1_ASAP7_75t_L g302 ( .A(n_215), .Y(n_302) );
INVx2_ASAP7_75t_L g340 ( .A(n_215), .Y(n_340) );
INVx1_ASAP7_75t_L g848 ( .A(n_216), .Y(n_848) );
INVxp33_ASAP7_75t_SL g350 ( .A(n_217), .Y(n_350) );
INVx1_ASAP7_75t_L g973 ( .A(n_218), .Y(n_973) );
OAI221xp5_ASAP7_75t_L g850 ( .A1(n_219), .A2(n_494), .B1(n_851), .B2(n_857), .C(n_861), .Y(n_850) );
OR2x2_ASAP7_75t_L g1063 ( .A(n_220), .B(n_389), .Y(n_1063) );
INVx1_ASAP7_75t_L g1055 ( .A(n_221), .Y(n_1055) );
INVx1_ASAP7_75t_L g1137 ( .A(n_222), .Y(n_1137) );
OAI22xp5_ASAP7_75t_L g1005 ( .A1(n_223), .A2(n_1006), .B1(n_1059), .B2(n_1060), .Y(n_1005) );
INVx1_ASAP7_75t_L g1060 ( .A(n_223), .Y(n_1060) );
INVx1_ASAP7_75t_L g912 ( .A(n_224), .Y(n_912) );
AOI21xp33_ASAP7_75t_L g927 ( .A1(n_224), .A2(n_436), .B(n_624), .Y(n_927) );
INVxp67_ASAP7_75t_SL g319 ( .A(n_225), .Y(n_319) );
AOI221xp5_ASAP7_75t_L g1360 ( .A1(n_228), .A2(n_229), .B1(n_1277), .B2(n_1361), .C(n_1362), .Y(n_1360) );
INVx1_ASAP7_75t_L g1034 ( .A(n_230), .Y(n_1034) );
INVx1_ASAP7_75t_L g1603 ( .A(n_231), .Y(n_1603) );
INVx1_ASAP7_75t_L g1529 ( .A(n_234), .Y(n_1529) );
INVx1_ASAP7_75t_L g1209 ( .A(n_235), .Y(n_1209) );
INVx1_ASAP7_75t_L g1212 ( .A(n_236), .Y(n_1212) );
INVx1_ASAP7_75t_L g648 ( .A(n_237), .Y(n_648) );
INVx1_ASAP7_75t_L g1562 ( .A(n_238), .Y(n_1562) );
INVx1_ASAP7_75t_L g684 ( .A(n_239), .Y(n_684) );
INVx1_ASAP7_75t_L g799 ( .A(n_241), .Y(n_799) );
INVx1_ASAP7_75t_L g913 ( .A(n_242), .Y(n_913) );
INVx1_ASAP7_75t_L g504 ( .A(n_243), .Y(n_504) );
INVx1_ASAP7_75t_L g814 ( .A(n_244), .Y(n_814) );
INVx1_ASAP7_75t_L g1530 ( .A(n_245), .Y(n_1530) );
INVx1_ASAP7_75t_L g1032 ( .A(n_247), .Y(n_1032) );
INVx1_ASAP7_75t_L g1281 ( .A(n_248), .Y(n_1281) );
NAND2xp5_ASAP7_75t_L g1302 ( .A(n_248), .B(n_1297), .Y(n_1302) );
INVx1_ASAP7_75t_L g1020 ( .A(n_249), .Y(n_1020) );
INVx1_ASAP7_75t_L g1216 ( .A(n_250), .Y(n_1216) );
CKINVDCx5p33_ASAP7_75t_R g984 ( .A(n_251), .Y(n_984) );
INVx1_ASAP7_75t_L g1577 ( .A(n_254), .Y(n_1577) );
OAI22xp5_ASAP7_75t_L g1604 ( .A1(n_254), .A2(n_264), .B1(n_1605), .B2(n_1606), .Y(n_1604) );
INVx1_ASAP7_75t_L g1003 ( .A(n_255), .Y(n_1003) );
CKINVDCx5p33_ASAP7_75t_R g647 ( .A(n_256), .Y(n_647) );
CKINVDCx5p33_ASAP7_75t_R g1134 ( .A(n_257), .Y(n_1134) );
INVx2_ASAP7_75t_L g299 ( .A(n_258), .Y(n_299) );
INVx1_ASAP7_75t_L g695 ( .A(n_259), .Y(n_695) );
INVx1_ASAP7_75t_L g1069 ( .A(n_260), .Y(n_1069) );
INVx1_ASAP7_75t_L g1080 ( .A(n_261), .Y(n_1080) );
CKINVDCx5p33_ASAP7_75t_R g1166 ( .A(n_262), .Y(n_1166) );
INVx1_ASAP7_75t_L g1574 ( .A(n_264), .Y(n_1574) );
INVx1_ASAP7_75t_L g849 ( .A(n_265), .Y(n_849) );
INVx1_ASAP7_75t_L g1225 ( .A(n_266), .Y(n_1225) );
INVx1_ASAP7_75t_L g1540 ( .A(n_267), .Y(n_1540) );
INVx1_ASAP7_75t_L g820 ( .A(n_268), .Y(n_820) );
INVx1_ASAP7_75t_L g793 ( .A(n_269), .Y(n_793) );
CKINVDCx5p33_ASAP7_75t_R g646 ( .A(n_271), .Y(n_646) );
AOI21xp33_ASAP7_75t_L g860 ( .A1(n_272), .A2(n_673), .B(n_841), .Y(n_860) );
CKINVDCx5p33_ASAP7_75t_R g1581 ( .A(n_273), .Y(n_1581) );
INVx1_ASAP7_75t_L g1229 ( .A(n_274), .Y(n_1229) );
OAI211xp5_ASAP7_75t_SL g1075 ( .A1(n_275), .A2(n_918), .B(n_1076), .C(n_1079), .Y(n_1075) );
BUFx3_ASAP7_75t_L g402 ( .A(n_276), .Y(n_402) );
INVx1_ASAP7_75t_L g429 ( .A(n_276), .Y(n_429) );
BUFx3_ASAP7_75t_L g404 ( .A(n_277), .Y(n_404) );
INVx1_ASAP7_75t_L g410 ( .A(n_277), .Y(n_410) );
INVx1_ASAP7_75t_L g1010 ( .A(n_278), .Y(n_1010) );
INVx1_ASAP7_75t_L g387 ( .A(n_279), .Y(n_387) );
INVx1_ASAP7_75t_L g1547 ( .A(n_280), .Y(n_1547) );
AOI21xp5_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_303), .B(n_1275), .Y(n_281) );
INVx2_ASAP7_75t_SL g282 ( .A(n_283), .Y(n_282) );
INVx1_ASAP7_75t_SL g283 ( .A(n_284), .Y(n_283) );
AND2x4_ASAP7_75t_L g284 ( .A(n_285), .B(n_290), .Y(n_284) );
AND2x4_ASAP7_75t_L g1567 ( .A(n_285), .B(n_291), .Y(n_1567) );
NOR2xp33_ASAP7_75t_SL g285 ( .A(n_286), .B(n_288), .Y(n_285) );
INVx1_ASAP7_75t_SL g1626 ( .A(n_286), .Y(n_1626) );
NAND2xp5_ASAP7_75t_L g1631 ( .A(n_286), .B(n_288), .Y(n_1631) );
HB1xp67_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g1625 ( .A(n_288), .B(n_1626), .Y(n_1625) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
NOR2xp33_ASAP7_75t_L g291 ( .A(n_292), .B(n_296), .Y(n_291) );
INVxp67_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
HB1xp67_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g361 ( .A(n_294), .B(n_302), .Y(n_361) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
OR2x2_ASAP7_75t_L g673 ( .A(n_295), .B(n_674), .Y(n_673) );
OR2x6_ASAP7_75t_L g296 ( .A(n_297), .B(n_301), .Y(n_296) );
OR2x2_ASAP7_75t_L g390 ( .A(n_297), .B(n_317), .Y(n_390) );
INVx2_ASAP7_75t_SL g512 ( .A(n_297), .Y(n_512) );
INVx1_ASAP7_75t_L g527 ( .A(n_297), .Y(n_527) );
BUFx6f_ASAP7_75t_L g693 ( .A(n_297), .Y(n_693) );
BUFx2_ASAP7_75t_L g810 ( .A(n_297), .Y(n_810) );
INVx2_ASAP7_75t_SL g1046 ( .A(n_297), .Y(n_1046) );
BUFx6f_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_299), .B(n_300), .Y(n_298) );
INVx1_ASAP7_75t_L g323 ( .A(n_299), .Y(n_323) );
INVx1_ASAP7_75t_L g328 ( .A(n_299), .Y(n_328) );
AND2x4_ASAP7_75t_L g336 ( .A(n_299), .B(n_329), .Y(n_336) );
AND2x2_ASAP7_75t_L g349 ( .A(n_299), .B(n_300), .Y(n_349) );
INVx2_ASAP7_75t_L g354 ( .A(n_299), .Y(n_354) );
INVx1_ASAP7_75t_L g315 ( .A(n_300), .Y(n_315) );
INVx2_ASAP7_75t_L g329 ( .A(n_300), .Y(n_329) );
INVx1_ASAP7_75t_L g356 ( .A(n_300), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_300), .B(n_354), .Y(n_501) );
INVx1_ASAP7_75t_L g509 ( .A(n_300), .Y(n_509) );
INVx2_ASAP7_75t_SL g301 ( .A(n_302), .Y(n_301) );
OAI22xp33_ASAP7_75t_L g303 ( .A1(n_304), .A2(n_305), .B1(n_943), .B2(n_944), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
AOI22xp5_ASAP7_75t_L g305 ( .A1(n_306), .A2(n_696), .B1(n_941), .B2(n_942), .Y(n_305) );
INVx1_ASAP7_75t_L g941 ( .A(n_306), .Y(n_941) );
XNOR2xp5_ASAP7_75t_L g306 ( .A(n_307), .B(n_611), .Y(n_306) );
AOI22xp33_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_309), .B1(n_480), .B2(n_610), .Y(n_307) );
INVx2_ASAP7_75t_SL g308 ( .A(n_309), .Y(n_308) );
XNOR2x1_ASAP7_75t_L g309 ( .A(n_310), .B(n_479), .Y(n_309) );
AND2x2_ASAP7_75t_L g310 ( .A(n_311), .B(n_386), .Y(n_310) );
AND4x1_ASAP7_75t_L g311 ( .A(n_312), .B(n_330), .C(n_344), .D(n_357), .Y(n_311) );
AOI221xp5_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_319), .B1(n_320), .B2(n_324), .C(n_325), .Y(n_312) );
AOI221xp5_ASAP7_75t_L g890 ( .A1(n_313), .A2(n_320), .B1(n_325), .B2(n_891), .C(n_892), .Y(n_890) );
AOI221xp5_ASAP7_75t_L g1101 ( .A1(n_313), .A2(n_320), .B1(n_325), .B2(n_1077), .C(n_1078), .Y(n_1101) );
AOI221xp5_ASAP7_75t_L g1210 ( .A1(n_313), .A2(n_320), .B1(n_325), .B2(n_1211), .C(n_1212), .Y(n_1210) );
INVx1_ASAP7_75t_L g1576 ( .A(n_313), .Y(n_1576) );
AND2x4_ASAP7_75t_L g313 ( .A(n_314), .B(n_316), .Y(n_313) );
AND2x2_ASAP7_75t_L g542 ( .A(n_314), .B(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g1267 ( .A(n_314), .B(n_543), .Y(n_1267) );
HB1xp67_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g665 ( .A(n_315), .Y(n_665) );
AND2x4_ASAP7_75t_L g320 ( .A(n_316), .B(n_321), .Y(n_320) );
AND2x4_ASAP7_75t_L g325 ( .A(n_316), .B(n_326), .Y(n_325) );
NAND2x1_ASAP7_75t_SL g663 ( .A(n_316), .B(n_664), .Y(n_663) );
NAND2x1p5_ASAP7_75t_L g667 ( .A(n_316), .B(n_668), .Y(n_667) );
NAND2x1p5_ASAP7_75t_L g670 ( .A(n_316), .B(n_343), .Y(n_670) );
INVx3_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g518 ( .A(n_318), .Y(n_518) );
HB1xp67_ASAP7_75t_L g1573 ( .A(n_320), .Y(n_1573) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g508 ( .A(n_323), .B(n_509), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_323), .B(n_509), .Y(n_681) );
AOI221xp5_ASAP7_75t_L g1572 ( .A1(n_325), .A2(n_1573), .B1(n_1574), .B2(n_1575), .C(n_1577), .Y(n_1572) );
INVx1_ASAP7_75t_L g367 ( .A(n_326), .Y(n_367) );
BUFx2_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
BUFx3_ASAP7_75t_L g343 ( .A(n_327), .Y(n_343) );
BUFx6f_ASAP7_75t_L g379 ( .A(n_327), .Y(n_379) );
BUFx3_ASAP7_75t_L g522 ( .A(n_327), .Y(n_522) );
BUFx6f_ASAP7_75t_L g845 ( .A(n_327), .Y(n_845) );
AND2x4_ASAP7_75t_L g327 ( .A(n_328), .B(n_329), .Y(n_327) );
AOI22xp33_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_332), .B1(n_341), .B2(n_342), .Y(n_330) );
BUFx2_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
BUFx2_ASAP7_75t_L g654 ( .A(n_333), .Y(n_654) );
AOI22xp33_ASAP7_75t_L g797 ( .A1(n_333), .A2(n_342), .B1(n_798), .B2(n_799), .Y(n_797) );
BUFx2_ASAP7_75t_L g909 ( .A(n_333), .Y(n_909) );
BUFx2_ASAP7_75t_L g953 ( .A(n_333), .Y(n_953) );
BUFx2_ASAP7_75t_L g1580 ( .A(n_333), .Y(n_1580) );
AND2x4_ASAP7_75t_L g333 ( .A(n_334), .B(n_337), .Y(n_333) );
BUFx3_ASAP7_75t_L g824 ( .A(n_334), .Y(n_824) );
INVx2_ASAP7_75t_L g855 ( .A(n_334), .Y(n_855) );
INVx1_ASAP7_75t_L g1130 ( .A(n_334), .Y(n_1130) );
INVx3_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
BUFx6f_ASAP7_75t_L g690 ( .A(n_335), .Y(n_690) );
INVx3_ASAP7_75t_L g839 ( .A(n_335), .Y(n_839) );
INVx3_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
BUFx6f_ASAP7_75t_L g372 ( .A(n_336), .Y(n_372) );
INVx1_ASAP7_75t_L g492 ( .A(n_336), .Y(n_492) );
AND2x6_ASAP7_75t_L g342 ( .A(n_337), .B(n_343), .Y(n_342) );
AND2x4_ASAP7_75t_L g346 ( .A(n_337), .B(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g351 ( .A(n_337), .B(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g659 ( .A(n_337), .B(n_352), .Y(n_659) );
AND2x2_ASAP7_75t_L g958 ( .A(n_337), .B(n_352), .Y(n_958) );
AND2x2_ASAP7_75t_L g1033 ( .A(n_337), .B(n_839), .Y(n_1033) );
AND2x2_ASAP7_75t_L g1035 ( .A(n_337), .B(n_379), .Y(n_1035) );
AND2x2_ASAP7_75t_L g1039 ( .A(n_337), .B(n_352), .Y(n_1039) );
AND2x2_ASAP7_75t_L g1179 ( .A(n_337), .B(n_554), .Y(n_1179) );
AND2x2_ASAP7_75t_L g1585 ( .A(n_337), .B(n_352), .Y(n_1585) );
AND2x4_ASAP7_75t_L g337 ( .A(n_338), .B(n_339), .Y(n_337) );
INVx1_ASAP7_75t_L g382 ( .A(n_338), .Y(n_382) );
OR2x2_ASAP7_75t_L g560 ( .A(n_338), .B(n_412), .Y(n_560) );
AND2x2_ASAP7_75t_L g486 ( .A(n_339), .B(n_353), .Y(n_486) );
INVx2_ASAP7_75t_L g490 ( .A(n_339), .Y(n_490) );
AND2x4_ASAP7_75t_L g495 ( .A(n_339), .B(n_365), .Y(n_495) );
INVx1_ASAP7_75t_L g384 ( .A(n_340), .Y(n_384) );
INVx1_ASAP7_75t_L g674 ( .A(n_340), .Y(n_674) );
OAI211xp5_ASAP7_75t_L g424 ( .A1(n_341), .A2(n_425), .B(n_431), .C(n_435), .Y(n_424) );
AOI22xp33_ASAP7_75t_L g652 ( .A1(n_342), .A2(n_653), .B1(n_654), .B2(n_655), .Y(n_652) );
AOI22xp33_ASAP7_75t_L g907 ( .A1(n_342), .A2(n_908), .B1(n_909), .B2(n_910), .Y(n_907) );
AOI22xp33_ASAP7_75t_L g951 ( .A1(n_342), .A2(n_952), .B1(n_953), .B2(n_954), .Y(n_951) );
AOI22xp33_ASAP7_75t_L g1578 ( .A1(n_342), .A2(n_1579), .B1(n_1580), .B2(n_1581), .Y(n_1578) );
AOI22xp33_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_346), .B1(n_350), .B2(n_351), .Y(n_344) );
AOI22xp33_ASAP7_75t_L g656 ( .A1(n_346), .A2(n_657), .B1(n_658), .B2(n_659), .Y(n_656) );
AOI22xp33_ASAP7_75t_L g800 ( .A1(n_346), .A2(n_351), .B1(n_801), .B2(n_802), .Y(n_800) );
AOI22xp33_ASAP7_75t_L g911 ( .A1(n_346), .A2(n_659), .B1(n_912), .B2(n_913), .Y(n_911) );
AOI22xp33_ASAP7_75t_L g955 ( .A1(n_346), .A2(n_956), .B1(n_957), .B2(n_958), .Y(n_955) );
AOI22xp33_ASAP7_75t_L g1036 ( .A1(n_346), .A2(n_1037), .B1(n_1038), .B2(n_1039), .Y(n_1036) );
AOI221xp5_ASAP7_75t_L g1102 ( .A1(n_346), .A2(n_958), .B1(n_1103), .B2(n_1104), .C(n_1105), .Y(n_1102) );
AOI22xp33_ASAP7_75t_L g1582 ( .A1(n_346), .A2(n_1583), .B1(n_1584), .B2(n_1585), .Y(n_1582) );
INVx1_ASAP7_75t_L g842 ( .A(n_347), .Y(n_842) );
INVx1_ASAP7_75t_L g905 ( .A(n_347), .Y(n_905) );
BUFx2_ASAP7_75t_L g1090 ( .A(n_347), .Y(n_1090) );
BUFx3_ASAP7_75t_L g1598 ( .A(n_347), .Y(n_1598) );
INVx2_ASAP7_75t_SL g347 ( .A(n_348), .Y(n_347) );
INVx2_ASAP7_75t_SL g554 ( .A(n_348), .Y(n_554) );
INVx2_ASAP7_75t_L g748 ( .A(n_348), .Y(n_748) );
INVx3_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
BUFx6f_ASAP7_75t_L g365 ( .A(n_349), .Y(n_365) );
INVx2_ASAP7_75t_SL g1595 ( .A(n_352), .Y(n_1595) );
BUFx6f_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
BUFx2_ASAP7_75t_L g369 ( .A(n_353), .Y(n_369) );
BUFx6f_ASAP7_75t_L g737 ( .A(n_353), .Y(n_737) );
INVx1_ASAP7_75t_L g836 ( .A(n_353), .Y(n_836) );
INVx1_ASAP7_75t_L g899 ( .A(n_353), .Y(n_899) );
BUFx6f_ASAP7_75t_L g1122 ( .A(n_353), .Y(n_1122) );
AND2x4_ASAP7_75t_L g353 ( .A(n_354), .B(n_355), .Y(n_353) );
INVx1_ASAP7_75t_L g547 ( .A(n_354), .Y(n_547) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
AOI33xp33_ASAP7_75t_L g357 ( .A1(n_358), .A2(n_362), .A3(n_368), .B1(n_373), .B2(n_374), .B3(n_380), .Y(n_357) );
BUFx2_ASAP7_75t_L g894 ( .A(n_358), .Y(n_894) );
AOI33xp33_ASAP7_75t_L g1088 ( .A1(n_358), .A2(n_1089), .A3(n_1091), .B1(n_1095), .B2(n_1097), .B3(n_1100), .Y(n_1088) );
AND2x4_ASAP7_75t_L g358 ( .A(n_359), .B(n_361), .Y(n_358) );
BUFx2_ASAP7_75t_L g478 ( .A(n_359), .Y(n_478) );
INVx2_ASAP7_75t_L g552 ( .A(n_359), .Y(n_552) );
OR2x6_ASAP7_75t_L g584 ( .A(n_359), .B(n_585), .Y(n_584) );
OR2x2_ASAP7_75t_L g704 ( .A(n_359), .B(n_705), .Y(n_704) );
AND2x2_ASAP7_75t_L g1100 ( .A(n_359), .B(n_531), .Y(n_1100) );
OR2x2_ASAP7_75t_L g1526 ( .A(n_359), .B(n_585), .Y(n_1526) );
AND2x4_ASAP7_75t_L g1588 ( .A(n_359), .B(n_361), .Y(n_1588) );
INVx2_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
BUFx2_ASAP7_75t_L g618 ( .A(n_360), .Y(n_618) );
OR2x6_ASAP7_75t_L g672 ( .A(n_360), .B(n_673), .Y(n_672) );
BUFx2_ASAP7_75t_SL g514 ( .A(n_361), .Y(n_514) );
INVx1_ASAP7_75t_L g1250 ( .A(n_361), .Y(n_1250) );
HB1xp67_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g376 ( .A(n_364), .Y(n_376) );
BUFx6f_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
BUFx2_ASAP7_75t_L g740 ( .A(n_365), .Y(n_740) );
INVx3_ASAP7_75t_L g1099 ( .A(n_365), .Y(n_1099) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx2_ASAP7_75t_SL g371 ( .A(n_372), .Y(n_371) );
INVx2_ASAP7_75t_SL g503 ( .A(n_372), .Y(n_503) );
INVx2_ASAP7_75t_SL g538 ( .A(n_372), .Y(n_538) );
BUFx3_ASAP7_75t_L g686 ( .A(n_372), .Y(n_686) );
INVx4_ASAP7_75t_L g979 ( .A(n_372), .Y(n_979) );
INVx2_ASAP7_75t_SL g1176 ( .A(n_372), .Y(n_1176) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx2_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx2_ASAP7_75t_SL g1591 ( .A(n_378), .Y(n_1591) );
INVx2_ASAP7_75t_SL g378 ( .A(n_379), .Y(n_378) );
BUFx6f_ASAP7_75t_L g896 ( .A(n_379), .Y(n_896) );
INVx2_ASAP7_75t_L g694 ( .A(n_380), .Y(n_694) );
AOI33xp33_ASAP7_75t_L g893 ( .A1(n_380), .A2(n_894), .A3(n_895), .B1(n_897), .B2(n_901), .B3(n_903), .Y(n_893) );
INVx1_ASAP7_75t_L g1177 ( .A(n_380), .Y(n_1177) );
AOI33xp33_ASAP7_75t_L g1586 ( .A1(n_380), .A2(n_1587), .A3(n_1589), .B1(n_1592), .B2(n_1596), .B3(n_1597), .Y(n_1586) );
INVx6_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
OAI33xp33_ASAP7_75t_L g806 ( .A1(n_381), .A2(n_672), .A3(n_807), .B1(n_815), .B2(n_821), .B3(n_825), .Y(n_806) );
INVx5_ASAP7_75t_L g982 ( .A(n_381), .Y(n_982) );
OR2x6_ASAP7_75t_L g381 ( .A(n_382), .B(n_383), .Y(n_381) );
NAND2x1p5_ASAP7_75t_L g578 ( .A(n_382), .B(n_395), .Y(n_578) );
INVx2_ASAP7_75t_L g531 ( .A(n_383), .Y(n_531) );
BUFx2_ASAP7_75t_L g1560 ( .A(n_383), .Y(n_1560) );
NAND2x1p5_ASAP7_75t_L g383 ( .A(n_384), .B(n_385), .Y(n_383) );
AOI21xp5_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_388), .B(n_405), .Y(n_386) );
AOI21xp33_ASAP7_75t_SL g983 ( .A1(n_388), .A2(n_984), .B(n_985), .Y(n_983) );
AOI21xp5_ASAP7_75t_L g1599 ( .A1(n_388), .A2(n_1600), .B(n_1601), .Y(n_1599) );
INVx5_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g649 ( .A(n_389), .Y(n_649) );
INVx2_ASAP7_75t_L g794 ( .A(n_389), .Y(n_794) );
INVx2_ASAP7_75t_SL g1028 ( .A(n_389), .Y(n_1028) );
AND2x4_ASAP7_75t_L g389 ( .A(n_390), .B(n_391), .Y(n_389) );
INVx2_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
OR2x6_ASAP7_75t_L g550 ( .A(n_392), .B(n_551), .Y(n_550) );
AND2x4_ASAP7_75t_L g392 ( .A(n_393), .B(n_394), .Y(n_392) );
AND2x4_ASAP7_75t_L g603 ( .A(n_393), .B(n_439), .Y(n_603) );
AND2x4_ASAP7_75t_L g716 ( .A(n_393), .B(n_439), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g1208 ( .A(n_394), .B(n_1209), .Y(n_1208) );
AND2x2_ASAP7_75t_L g394 ( .A(n_395), .B(n_400), .Y(n_394) );
AND2x4_ASAP7_75t_L g416 ( .A(n_395), .B(n_417), .Y(n_416) );
AND2x2_ASAP7_75t_L g421 ( .A(n_395), .B(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g465 ( .A(n_395), .Y(n_465) );
AND2x4_ASAP7_75t_L g633 ( .A(n_395), .B(n_417), .Y(n_633) );
BUFx2_ASAP7_75t_L g644 ( .A(n_395), .Y(n_644) );
AND2x4_ASAP7_75t_L g779 ( .A(n_395), .B(n_422), .Y(n_779) );
AND2x2_ASAP7_75t_L g1607 ( .A(n_395), .B(n_422), .Y(n_1607) );
AND2x4_ASAP7_75t_L g395 ( .A(n_396), .B(n_398), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
AND2x4_ASAP7_75t_L g439 ( .A(n_398), .B(n_440), .Y(n_439) );
INVx2_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
AND2x2_ASAP7_75t_L g456 ( .A(n_399), .B(n_440), .Y(n_456) );
INVx6_ASAP7_75t_L g437 ( .A(n_400), .Y(n_437) );
INVx2_ASAP7_75t_L g567 ( .A(n_400), .Y(n_567) );
BUFx2_ASAP7_75t_L g788 ( .A(n_400), .Y(n_788) );
AND2x4_ASAP7_75t_L g400 ( .A(n_401), .B(n_403), .Y(n_400) );
INVx1_ASAP7_75t_L g423 ( .A(n_401), .Y(n_423) );
INVx2_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
AND2x4_ASAP7_75t_L g409 ( .A(n_402), .B(n_410), .Y(n_409) );
AND2x2_ASAP7_75t_L g445 ( .A(n_402), .B(n_404), .Y(n_445) );
INVx1_ASAP7_75t_L g419 ( .A(n_403), .Y(n_419) );
INVx2_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
AND2x4_ASAP7_75t_L g434 ( .A(n_404), .B(n_429), .Y(n_434) );
AOI31xp33_ASAP7_75t_L g405 ( .A1(n_406), .A2(n_441), .A3(n_467), .B(n_476), .Y(n_405) );
AOI21xp33_ASAP7_75t_SL g406 ( .A1(n_407), .A2(n_413), .B(n_414), .Y(n_406) );
AOI221xp5_ASAP7_75t_L g620 ( .A1(n_407), .A2(n_621), .B1(n_625), .B2(n_630), .C(n_631), .Y(n_620) );
AOI221xp5_ASAP7_75t_L g766 ( .A1(n_407), .A2(n_767), .B1(n_768), .B2(n_772), .C(n_777), .Y(n_766) );
AOI211xp5_ASAP7_75t_L g986 ( .A1(n_407), .A2(n_973), .B(n_987), .C(n_989), .Y(n_986) );
AOI211xp5_ASAP7_75t_SL g1602 ( .A1(n_407), .A2(n_1603), .B(n_1604), .C(n_1608), .Y(n_1602) );
AND2x4_ASAP7_75t_L g407 ( .A(n_408), .B(n_411), .Y(n_407) );
BUFx3_ASAP7_75t_L g599 ( .A(n_408), .Y(n_599) );
INVx2_ASAP7_75t_SL g997 ( .A(n_408), .Y(n_997) );
BUFx6f_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
BUFx6f_ASAP7_75t_L g432 ( .A(n_409), .Y(n_432) );
BUFx6f_ASAP7_75t_L g450 ( .A(n_409), .Y(n_450) );
INVx2_ASAP7_75t_SL g571 ( .A(n_409), .Y(n_571) );
BUFx3_ASAP7_75t_L g715 ( .A(n_409), .Y(n_715) );
BUFx6f_ASAP7_75t_L g756 ( .A(n_409), .Y(n_756) );
BUFx2_ASAP7_75t_L g773 ( .A(n_409), .Y(n_773) );
HB1xp67_ASAP7_75t_L g1023 ( .A(n_409), .Y(n_1023) );
INVx1_ASAP7_75t_L g430 ( .A(n_410), .Y(n_430) );
AND2x4_ASAP7_75t_L g443 ( .A(n_411), .B(n_444), .Y(n_443) );
AND2x2_ASAP7_75t_L g919 ( .A(n_411), .B(n_756), .Y(n_919) );
INVx2_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
OR2x2_ASAP7_75t_L g470 ( .A(n_412), .B(n_471), .Y(n_470) );
OR2x2_ASAP7_75t_L g474 ( .A(n_412), .B(n_475), .Y(n_474) );
A2O1A1Ixp33_ASAP7_75t_L g1186 ( .A1(n_412), .A2(n_1187), .B(n_1188), .C(n_1190), .Y(n_1186) );
INVx2_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx4_ASAP7_75t_L g922 ( .A(n_416), .Y(n_922) );
INVx1_ASAP7_75t_SL g1026 ( .A(n_416), .Y(n_1026) );
AOI22xp5_ASAP7_75t_L g1076 ( .A1(n_416), .A2(n_779), .B1(n_1077), .B2(n_1078), .Y(n_1076) );
INVx2_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g576 ( .A(n_418), .Y(n_576) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx3_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx2_ASAP7_75t_L g581 ( .A(n_422), .Y(n_581) );
BUFx3_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx2_ASAP7_75t_SL g1072 ( .A(n_426), .Y(n_1072) );
INVx1_ASAP7_75t_L g1081 ( .A(n_426), .Y(n_1081) );
INVx1_ASAP7_75t_L g1201 ( .A(n_426), .Y(n_1201) );
BUFx4f_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx2_ASAP7_75t_L g563 ( .A(n_427), .Y(n_563) );
INVx1_ASAP7_75t_L g925 ( .A(n_427), .Y(n_925) );
INVx1_ASAP7_75t_L g1196 ( .A(n_427), .Y(n_1196) );
INVx1_ASAP7_75t_L g1228 ( .A(n_427), .Y(n_1228) );
AND2x2_ASAP7_75t_L g427 ( .A(n_428), .B(n_430), .Y(n_427) );
OR2x2_ASAP7_75t_L g471 ( .A(n_428), .B(n_430), .Y(n_471) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
BUFx2_ASAP7_75t_L g587 ( .A(n_432), .Y(n_587) );
BUFx3_ASAP7_75t_L g626 ( .A(n_432), .Y(n_626) );
INVx2_ASAP7_75t_L g637 ( .A(n_432), .Y(n_637) );
INVx1_ASAP7_75t_L g1528 ( .A(n_432), .Y(n_1528) );
BUFx6f_ASAP7_75t_L g588 ( .A(n_433), .Y(n_588) );
INVx1_ASAP7_75t_L g601 ( .A(n_433), .Y(n_601) );
BUFx3_ASAP7_75t_L g1610 ( .A(n_433), .Y(n_1610) );
BUFx6f_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g462 ( .A(n_434), .Y(n_462) );
INVx2_ASAP7_75t_L g475 ( .A(n_434), .Y(n_475) );
BUFx6f_ASAP7_75t_L g629 ( .A(n_434), .Y(n_629) );
INVx2_ASAP7_75t_SL g436 ( .A(n_437), .Y(n_436) );
INVx2_ASAP7_75t_L g459 ( .A(n_437), .Y(n_459) );
INVx2_ASAP7_75t_L g596 ( .A(n_437), .Y(n_596) );
BUFx6f_ASAP7_75t_L g623 ( .A(n_437), .Y(n_623) );
INVx1_ASAP7_75t_L g709 ( .A(n_437), .Y(n_709) );
INVx1_ASAP7_75t_L g1203 ( .A(n_437), .Y(n_1203) );
INVx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
CKINVDCx5p33_ASAP7_75t_R g624 ( .A(n_439), .Y(n_624) );
INVx2_ASAP7_75t_SL g771 ( .A(n_439), .Y(n_771) );
HB1xp67_ASAP7_75t_L g993 ( .A(n_439), .Y(n_993) );
AOI221xp5_ASAP7_75t_L g441 ( .A1(n_442), .A2(n_446), .B1(n_447), .B2(n_457), .C(n_463), .Y(n_441) );
AOI221xp5_ASAP7_75t_L g634 ( .A1(n_442), .A2(n_635), .B1(n_640), .B2(n_642), .C(n_643), .Y(n_634) );
AOI221xp5_ASAP7_75t_L g994 ( .A1(n_442), .A2(n_463), .B1(n_975), .B2(n_995), .C(n_1000), .Y(n_994) );
AOI221xp5_ASAP7_75t_L g1612 ( .A1(n_442), .A2(n_463), .B1(n_1613), .B2(n_1614), .C(n_1618), .Y(n_1612) );
BUFx6f_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
HB1xp67_ASAP7_75t_L g781 ( .A(n_443), .Y(n_781) );
HB1xp67_ASAP7_75t_L g929 ( .A(n_443), .Y(n_929) );
INVx2_ASAP7_75t_SL g1014 ( .A(n_443), .Y(n_1014) );
INVx2_ASAP7_75t_SL g592 ( .A(n_444), .Y(n_592) );
BUFx3_ASAP7_75t_L g597 ( .A(n_444), .Y(n_597) );
BUFx6f_ASAP7_75t_L g607 ( .A(n_444), .Y(n_607) );
AND2x4_ASAP7_75t_L g643 ( .A(n_444), .B(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g785 ( .A(n_444), .Y(n_785) );
BUFx4f_ASAP7_75t_L g1189 ( .A(n_444), .Y(n_1189) );
BUFx6f_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
BUFx6f_ASAP7_75t_L g454 ( .A(n_445), .Y(n_454) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx2_ASAP7_75t_SL g990 ( .A(n_449), .Y(n_990) );
INVx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
HB1xp67_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
AND2x2_ASAP7_75t_L g721 ( .A(n_452), .B(n_608), .Y(n_721) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
BUFx6f_ASAP7_75t_L g466 ( .A(n_454), .Y(n_466) );
INVx2_ASAP7_75t_L g713 ( .A(n_454), .Y(n_713) );
BUFx6f_ASAP7_75t_L g999 ( .A(n_454), .Y(n_999) );
INVx2_ASAP7_75t_SL g455 ( .A(n_456), .Y(n_455) );
INVx2_ASAP7_75t_L g585 ( .A(n_456), .Y(n_585) );
BUFx3_ASAP7_75t_L g639 ( .A(n_456), .Y(n_639) );
INVx1_ASAP7_75t_L g705 ( .A(n_456), .Y(n_705) );
INVx1_ASAP7_75t_L g1205 ( .A(n_456), .Y(n_1205) );
BUFx3_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
HB1xp67_ASAP7_75t_L g590 ( .A(n_459), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g1187 ( .A1(n_459), .A2(n_641), .B1(n_1169), .B2(n_1175), .Y(n_1187) );
BUFx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
OR2x6_ASAP7_75t_L g559 ( .A(n_462), .B(n_560), .Y(n_559) );
OR2x2_ASAP7_75t_L g758 ( .A(n_462), .B(n_560), .Y(n_758) );
AND2x4_ASAP7_75t_L g463 ( .A(n_464), .B(n_466), .Y(n_463) );
INVx1_ASAP7_75t_SL g464 ( .A(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g867 ( .A(n_466), .Y(n_867) );
AOI22xp33_ASAP7_75t_L g467 ( .A1(n_468), .A2(n_469), .B1(n_472), .B2(n_473), .Y(n_467) );
AOI22xp33_ASAP7_75t_L g645 ( .A1(n_469), .A2(n_473), .B1(n_646), .B2(n_647), .Y(n_645) );
AOI22xp33_ASAP7_75t_L g790 ( .A1(n_469), .A2(n_473), .B1(n_791), .B2(n_792), .Y(n_790) );
AOI22xp33_ASAP7_75t_L g934 ( .A1(n_469), .A2(n_473), .B1(n_935), .B2(n_936), .Y(n_934) );
AOI22xp33_ASAP7_75t_L g1002 ( .A1(n_469), .A2(n_473), .B1(n_978), .B2(n_980), .Y(n_1002) );
AOI22xp5_ASAP7_75t_L g1009 ( .A1(n_469), .A2(n_473), .B1(n_1010), .B2(n_1011), .Y(n_1009) );
AOI22xp33_ASAP7_75t_L g1620 ( .A1(n_469), .A2(n_473), .B1(n_1621), .B2(n_1622), .Y(n_1620) );
INVx6_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx2_ASAP7_75t_L g753 ( .A(n_471), .Y(n_753) );
INVx1_ASAP7_75t_L g1146 ( .A(n_471), .Y(n_1146) );
BUFx2_ASAP7_75t_L g1224 ( .A(n_471), .Y(n_1224) );
INVx4_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx2_ASAP7_75t_L g776 ( .A(n_475), .Y(n_776) );
INVx1_ASAP7_75t_L g789 ( .A(n_475), .Y(n_789) );
OAI31xp33_ASAP7_75t_L g1548 ( .A1(n_476), .A2(n_1549), .A3(n_1550), .B(n_1554), .Y(n_1548) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
AOI22xp5_ASAP7_75t_L g1007 ( .A1(n_477), .A2(n_1008), .B1(n_1027), .B2(n_1028), .Y(n_1007) );
CKINVDCx8_ASAP7_75t_R g477 ( .A(n_478), .Y(n_477) );
OAI31xp33_ASAP7_75t_L g483 ( .A1(n_478), .A2(n_484), .A3(n_493), .B(n_519), .Y(n_483) );
OAI21xp5_ASAP7_75t_SL g831 ( .A1(n_478), .A2(n_832), .B(n_850), .Y(n_831) );
INVx1_ASAP7_75t_L g610 ( .A(n_480), .Y(n_610) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
NAND3xp33_ASAP7_75t_SL g482 ( .A(n_483), .B(n_548), .C(n_555), .Y(n_482) );
INVx3_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
AOI221x1_ASAP7_75t_L g723 ( .A1(n_486), .A2(n_488), .B1(n_724), .B2(n_725), .C(n_726), .Y(n_723) );
AOI22xp33_ASAP7_75t_L g847 ( .A1(n_486), .A2(n_488), .B1(n_848), .B2(n_849), .Y(n_847) );
AOI22xp33_ASAP7_75t_L g1117 ( .A1(n_486), .A2(n_488), .B1(n_1118), .B2(n_1119), .Y(n_1117) );
INVx3_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
AND2x4_ASAP7_75t_L g488 ( .A(n_489), .B(n_491), .Y(n_488) );
AND2x4_ASAP7_75t_L g521 ( .A(n_489), .B(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx1_ASAP7_75t_L g733 ( .A(n_491), .Y(n_733) );
INVx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g819 ( .A(n_492), .Y(n_819) );
CKINVDCx6p67_ASAP7_75t_R g494 ( .A(n_495), .Y(n_494) );
OAI22xp5_ASAP7_75t_L g496 ( .A1(n_497), .A2(n_502), .B1(n_503), .B2(n_504), .Y(n_496) );
OAI22xp5_ASAP7_75t_SL g682 ( .A1(n_497), .A2(n_683), .B1(n_684), .B2(n_685), .Y(n_682) );
OAI22xp5_ASAP7_75t_L g966 ( .A1(n_497), .A2(n_967), .B1(n_968), .B2(n_970), .Y(n_966) );
OAI221xp5_ASAP7_75t_L g1260 ( .A1(n_497), .A2(n_1176), .B1(n_1261), .B2(n_1262), .C(n_1263), .Y(n_1260) );
INVx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx2_ASAP7_75t_L g816 ( .A(n_498), .Y(n_816) );
INVx1_ASAP7_75t_L g822 ( .A(n_498), .Y(n_822) );
INVx2_ASAP7_75t_L g972 ( .A(n_498), .Y(n_972) );
INVx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
OAI22xp5_ASAP7_75t_L g731 ( .A1(n_499), .A2(n_732), .B1(n_733), .B2(n_734), .Y(n_731) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
BUFx3_ASAP7_75t_L g1053 ( .A(n_500), .Y(n_1053) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g536 ( .A(n_501), .Y(n_536) );
BUFx2_ASAP7_75t_L g1128 ( .A(n_501), .Y(n_1128) );
OAI221xp5_ASAP7_75t_L g505 ( .A1(n_506), .A2(n_510), .B1(n_511), .B2(n_513), .C(n_514), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx2_ASAP7_75t_L g524 ( .A(n_507), .Y(n_524) );
BUFx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx2_ASAP7_75t_L g516 ( .A(n_508), .Y(n_516) );
INVx3_ASAP7_75t_L g728 ( .A(n_508), .Y(n_728) );
INVx2_ASAP7_75t_L g858 ( .A(n_508), .Y(n_858) );
OAI221xp5_ASAP7_75t_L g1132 ( .A1(n_511), .A2(n_514), .B1(n_728), .B2(n_1133), .C(n_1134), .Y(n_1132) );
OAI22xp33_ASAP7_75t_L g1164 ( .A1(n_511), .A2(n_1165), .B1(n_1166), .B2(n_1167), .Y(n_1164) );
OAI221xp5_ASAP7_75t_L g1248 ( .A1(n_511), .A2(n_974), .B1(n_1225), .B2(n_1229), .C(n_1249), .Y(n_1248) );
INVx3_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
OAI21xp5_ASAP7_75t_L g726 ( .A1(n_515), .A2(n_727), .B(n_731), .Y(n_726) );
OR2x6_ASAP7_75t_L g515 ( .A(n_516), .B(n_517), .Y(n_515) );
OAI22xp33_ASAP7_75t_L g825 ( .A1(n_516), .A2(n_782), .B1(n_791), .B2(n_808), .Y(n_825) );
OR2x2_ASAP7_75t_L g861 ( .A(n_516), .B(n_517), .Y(n_861) );
INVx1_ASAP7_75t_L g1049 ( .A(n_516), .Y(n_1049) );
INVx1_ASAP7_75t_L g543 ( .A(n_517), .Y(n_543) );
OR2x6_ASAP7_75t_L g546 ( .A(n_517), .B(n_547), .Y(n_546) );
INVx1_ASAP7_75t_L g745 ( .A(n_517), .Y(n_745) );
INVx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx8_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
AOI221xp5_ASAP7_75t_SL g735 ( .A1(n_521), .A2(n_736), .B1(n_739), .B2(n_742), .C(n_743), .Y(n_735) );
BUFx6f_ASAP7_75t_L g741 ( .A(n_522), .Y(n_741) );
OAI221xp5_ASAP7_75t_L g523 ( .A1(n_524), .A2(n_525), .B1(n_526), .B2(n_528), .C(n_529), .Y(n_523) );
AOI22xp33_ASAP7_75t_L g557 ( .A1(n_525), .A2(n_539), .B1(n_558), .B2(n_561), .Y(n_557) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g677 ( .A(n_527), .Y(n_677) );
INVx2_ASAP7_75t_L g977 ( .A(n_527), .Y(n_977) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_528), .A2(n_537), .B1(n_565), .B2(n_569), .Y(n_564) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx2_ASAP7_75t_SL g530 ( .A(n_531), .Y(n_530) );
INVx1_ASAP7_75t_L g1264 ( .A(n_531), .Y(n_1264) );
OAI22xp5_ASAP7_75t_L g532 ( .A1(n_533), .A2(n_537), .B1(n_538), .B2(n_539), .Y(n_532) );
OAI22xp5_ASAP7_75t_L g687 ( .A1(n_533), .A2(n_630), .B1(n_647), .B2(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
HB1xp67_ASAP7_75t_L g853 ( .A(n_536), .Y(n_853) );
INVx1_ASAP7_75t_L g1174 ( .A(n_536), .Y(n_1174) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_541), .A2(n_542), .B1(n_544), .B2(n_545), .Y(n_540) );
AOI22xp5_ASAP7_75t_L g573 ( .A1(n_541), .A2(n_544), .B1(n_574), .B2(n_579), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_543), .B(n_554), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g1265 ( .A1(n_545), .A2(n_1266), .B1(n_1268), .B2(n_1269), .Y(n_1265) );
AOI22xp33_ASAP7_75t_L g1561 ( .A1(n_545), .A2(n_1267), .B1(n_1562), .B2(n_1563), .Y(n_1561) );
CKINVDCx11_ASAP7_75t_R g545 ( .A(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g668 ( .A(n_547), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_549), .B(n_550), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g862 ( .A(n_550), .B(n_863), .Y(n_862) );
NAND2xp5_ASAP7_75t_L g1136 ( .A(n_550), .B(n_1137), .Y(n_1136) );
NAND2xp5_ASAP7_75t_L g1218 ( .A(n_550), .B(n_1219), .Y(n_1218) );
NAND2xp5_ASAP7_75t_L g1546 ( .A(n_550), .B(n_1547), .Y(n_1546) );
NOR2xp67_ASAP7_75t_L g551 ( .A(n_552), .B(n_553), .Y(n_551) );
INVx2_ASAP7_75t_L g1086 ( .A(n_552), .Y(n_1086) );
NOR2xp33_ASAP7_75t_L g555 ( .A(n_556), .B(n_572), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_557), .B(n_564), .Y(n_556) );
CKINVDCx6p67_ASAP7_75t_R g558 ( .A(n_559), .Y(n_558) );
OR2x6_ASAP7_75t_L g562 ( .A(n_560), .B(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g568 ( .A(n_560), .Y(n_568) );
OR2x2_ASAP7_75t_L g751 ( .A(n_560), .B(n_752), .Y(n_751) );
OR2x2_ASAP7_75t_L g754 ( .A(n_560), .B(n_755), .Y(n_754) );
CKINVDCx6p67_ASAP7_75t_R g561 ( .A(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g1239 ( .A(n_563), .Y(n_1239) );
AOI221xp5_ASAP7_75t_L g883 ( .A1(n_565), .A2(n_569), .B1(n_884), .B2(n_885), .C(n_886), .Y(n_883) );
AOI221xp5_ASAP7_75t_L g1150 ( .A1(n_565), .A2(n_569), .B1(n_1151), .B2(n_1152), .C(n_1153), .Y(n_1150) );
AND2x2_ASAP7_75t_L g565 ( .A(n_566), .B(n_568), .Y(n_565) );
BUFx2_ASAP7_75t_L g874 ( .A(n_566), .Y(n_874) );
INVx2_ASAP7_75t_SL g566 ( .A(n_567), .Y(n_566) );
INVx1_ASAP7_75t_L g1199 ( .A(n_567), .Y(n_1199) );
AND2x2_ASAP7_75t_L g569 ( .A(n_568), .B(n_570), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g1188 ( .A1(n_570), .A2(n_1170), .B1(n_1172), .B2(n_1189), .Y(n_1188) );
INVx2_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx2_ASAP7_75t_SL g707 ( .A(n_571), .Y(n_707) );
OAI22xp5_ASAP7_75t_L g868 ( .A1(n_571), .A2(n_854), .B1(n_856), .B2(n_869), .Y(n_868) );
NAND3xp33_ASAP7_75t_SL g572 ( .A(n_573), .B(n_582), .C(n_604), .Y(n_572) );
INVx1_ASAP7_75t_L g881 ( .A(n_574), .Y(n_881) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx2_ASAP7_75t_L g718 ( .A(n_575), .Y(n_718) );
NAND2x1p5_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
INVx2_ASAP7_75t_SL g577 ( .A(n_578), .Y(n_577) );
OR2x6_ASAP7_75t_L g580 ( .A(n_578), .B(n_581), .Y(n_580) );
INVx1_ASAP7_75t_L g608 ( .A(n_578), .Y(n_608) );
OR2x2_ASAP7_75t_L g882 ( .A(n_578), .B(n_581), .Y(n_882) );
AOI221xp5_ASAP7_75t_L g717 ( .A1(n_579), .A2(n_718), .B1(n_719), .B2(n_720), .C(n_721), .Y(n_717) );
INVx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
AOI33xp33_ASAP7_75t_L g582 ( .A1(n_583), .A2(n_586), .A3(n_589), .B1(n_593), .B2(n_598), .B3(n_602), .Y(n_582) );
CKINVDCx5p33_ASAP7_75t_R g583 ( .A(n_584), .Y(n_583) );
INVx2_ASAP7_75t_L g870 ( .A(n_584), .Y(n_870) );
INVx2_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
INVx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
OAI22xp5_ASAP7_75t_L g1066 ( .A1(n_601), .A2(n_1067), .B1(n_1068), .B2(n_1069), .Y(n_1066) );
OAI22xp33_ASAP7_75t_L g1527 ( .A1(n_601), .A2(n_1528), .B1(n_1529), .B2(n_1530), .Y(n_1527) );
BUFx4f_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
AOI221xp5_ASAP7_75t_L g864 ( .A1(n_603), .A2(n_865), .B1(n_870), .B2(n_871), .C(n_880), .Y(n_864) );
INVx4_ASAP7_75t_L g1143 ( .A(n_603), .Y(n_1143) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .Y(n_606) );
INVx1_ASAP7_75t_L g873 ( .A(n_607), .Y(n_873) );
BUFx2_ASAP7_75t_SL g1617 ( .A(n_607), .Y(n_1617) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx2_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
XNOR2x1_ASAP7_75t_L g613 ( .A(n_614), .B(n_695), .Y(n_613) );
AND2x2_ASAP7_75t_L g614 ( .A(n_615), .B(n_650), .Y(n_614) );
AOI22xp5_ASAP7_75t_L g615 ( .A1(n_616), .A2(n_619), .B1(n_648), .B2(n_649), .Y(n_615) );
INVx2_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
BUFx8_ASAP7_75t_SL g1135 ( .A(n_617), .Y(n_1135) );
INVx2_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
BUFx2_ASAP7_75t_L g749 ( .A(n_618), .Y(n_749) );
NAND3xp33_ASAP7_75t_L g619 ( .A(n_620), .B(n_634), .C(n_645), .Y(n_619) );
INVx4_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx2_ASAP7_75t_L g711 ( .A(n_623), .Y(n_711) );
INVx1_ASAP7_75t_L g769 ( .A(n_623), .Y(n_769) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx2_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
BUFx6f_ASAP7_75t_L g641 ( .A(n_629), .Y(n_641) );
INVx1_ASAP7_75t_L g869 ( .A(n_629), .Y(n_869) );
INVx1_ASAP7_75t_L g879 ( .A(n_629), .Y(n_879) );
HB1xp67_ASAP7_75t_L g1018 ( .A(n_629), .Y(n_1018) );
BUFx6f_ASAP7_75t_L g1234 ( .A(n_629), .Y(n_1234) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g988 ( .A(n_633), .Y(n_988) );
INVx2_ASAP7_75t_SL g1207 ( .A(n_633), .Y(n_1207) );
INVx2_ASAP7_75t_L g1605 ( .A(n_633), .Y(n_1605) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx3_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVxp67_ASAP7_75t_L g932 ( .A(n_639), .Y(n_932) );
INVx2_ASAP7_75t_SL g1539 ( .A(n_641), .Y(n_1539) );
OAI22xp33_ASAP7_75t_L g691 ( .A1(n_642), .A2(n_646), .B1(n_679), .B2(n_692), .Y(n_691) );
AOI221xp5_ASAP7_75t_L g780 ( .A1(n_643), .A2(n_781), .B1(n_782), .B2(n_783), .C(n_787), .Y(n_780) );
AOI221xp5_ASAP7_75t_L g928 ( .A1(n_643), .A2(n_929), .B1(n_930), .B2(n_931), .C(n_933), .Y(n_928) );
AOI221xp5_ASAP7_75t_L g1012 ( .A1(n_643), .A2(n_1013), .B1(n_1015), .B2(n_1016), .C(n_1017), .Y(n_1012) );
INVx1_ASAP7_75t_L g1074 ( .A(n_643), .Y(n_1074) );
INVx1_ASAP7_75t_L g1190 ( .A(n_643), .Y(n_1190) );
NOR3xp33_ASAP7_75t_L g650 ( .A(n_651), .B(n_660), .C(n_671), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_652), .B(n_656), .Y(n_651) );
INVx2_ASAP7_75t_SL g661 ( .A(n_662), .Y(n_661) );
INVx2_ASAP7_75t_L g1041 ( .A(n_662), .Y(n_1041) );
INVx2_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
HB1xp67_ASAP7_75t_L g804 ( .A(n_663), .Y(n_804) );
NAND2x1p5_ASAP7_75t_L g744 ( .A(n_664), .B(n_745), .Y(n_744) );
INVx2_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
BUFx4f_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
BUFx4f_ASAP7_75t_L g805 ( .A(n_667), .Y(n_805) );
BUFx2_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
BUFx3_ASAP7_75t_L g1042 ( .A(n_670), .Y(n_1042) );
OAI33xp33_ASAP7_75t_L g671 ( .A1(n_672), .A2(n_675), .A3(n_682), .B1(n_687), .B2(n_691), .B3(n_694), .Y(n_671) );
OAI33xp33_ASAP7_75t_L g960 ( .A1(n_672), .A2(n_961), .A3(n_966), .B1(n_971), .B2(n_976), .B3(n_981), .Y(n_960) );
OAI33xp33_ASAP7_75t_L g1043 ( .A1(n_672), .A2(n_694), .A3(n_1044), .B1(n_1051), .B2(n_1056), .B3(n_1058), .Y(n_1043) );
OAI22xp33_ASAP7_75t_L g675 ( .A1(n_676), .A2(n_677), .B1(n_678), .B2(n_679), .Y(n_675) );
OAI22xp33_ASAP7_75t_L g1058 ( .A1(n_679), .A2(n_693), .B1(n_1010), .B2(n_1015), .Y(n_1058) );
BUFx3_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx2_ASAP7_75t_L g813 ( .A(n_680), .Y(n_813) );
BUFx3_ASAP7_75t_L g1167 ( .A(n_680), .Y(n_1167) );
OAI22xp33_ASAP7_75t_L g1168 ( .A1(n_680), .A2(n_693), .B1(n_1169), .B2(n_1170), .Y(n_1168) );
BUFx6f_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx3_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx2_ASAP7_75t_L g738 ( .A(n_690), .Y(n_738) );
OAI22xp33_ASAP7_75t_L g961 ( .A1(n_692), .A2(n_962), .B1(n_963), .B2(n_965), .Y(n_961) );
BUFx2_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g942 ( .A(n_696), .Y(n_942) );
XNOR2xp5_ASAP7_75t_L g696 ( .A(n_697), .B(n_828), .Y(n_696) );
AO22x2_ASAP7_75t_L g697 ( .A1(n_698), .A2(n_759), .B1(n_760), .B2(n_827), .Y(n_697) );
INVxp67_ASAP7_75t_SL g827 ( .A(n_698), .Y(n_827) );
INVxp67_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
NOR4xp75_ASAP7_75t_L g700 ( .A(n_701), .B(n_722), .C(n_750), .D(n_757), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_702), .B(n_717), .Y(n_701) );
AOI33xp33_ASAP7_75t_L g702 ( .A1(n_703), .A2(n_706), .A3(n_708), .B1(n_710), .B2(n_714), .B3(n_716), .Y(n_702) );
INVx3_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
OAI22xp5_ASAP7_75t_SL g1140 ( .A1(n_704), .A2(n_1141), .B1(n_1143), .B2(n_1144), .Y(n_1140) );
INVx2_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx3_ASAP7_75t_L g770 ( .A(n_713), .Y(n_770) );
BUFx3_ASAP7_75t_L g1242 ( .A(n_715), .Y(n_1242) );
INVx2_ASAP7_75t_L g1542 ( .A(n_718), .Y(n_1542) );
NOR3xp33_ASAP7_75t_L g1138 ( .A(n_721), .B(n_1139), .C(n_1140), .Y(n_1138) );
BUFx2_ASAP7_75t_L g1243 ( .A(n_721), .Y(n_1243) );
NOR3xp33_ASAP7_75t_SL g1524 ( .A(n_721), .B(n_1525), .C(n_1541), .Y(n_1524) );
AOI21x1_ASAP7_75t_L g722 ( .A1(n_723), .A2(n_735), .B(n_749), .Y(n_722) );
OAI21xp5_ASAP7_75t_SL g727 ( .A1(n_728), .A2(n_729), .B(n_730), .Y(n_727) );
INVx1_ASAP7_75t_L g964 ( .A(n_728), .Y(n_964) );
BUFx2_ASAP7_75t_L g974 ( .A(n_728), .Y(n_974) );
OAI221xp5_ASAP7_75t_L g1553 ( .A1(n_728), .A2(n_808), .B1(n_1249), .B2(n_1532), .C(n_1533), .Y(n_1553) );
INVx1_ASAP7_75t_L g1096 ( .A(n_733), .Y(n_1096) );
HB1xp67_ASAP7_75t_L g969 ( .A(n_738), .Y(n_969) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_747), .B(n_748), .Y(n_746) );
INVx2_ASAP7_75t_L g764 ( .A(n_749), .Y(n_764) );
OAI31xp33_ASAP7_75t_L g1185 ( .A1(n_749), .A2(n_1186), .A3(n_1191), .B(n_1206), .Y(n_1185) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx2_ASAP7_75t_L g992 ( .A(n_753), .Y(n_992) );
INVx2_ASAP7_75t_L g1067 ( .A(n_753), .Y(n_1067) );
INVx2_ASAP7_75t_L g1236 ( .A(n_753), .Y(n_1236) );
INVx1_ASAP7_75t_L g1609 ( .A(n_755), .Y(n_1609) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
BUFx4f_ASAP7_75t_L g786 ( .A(n_756), .Y(n_786) );
INVx1_ASAP7_75t_L g1616 ( .A(n_756), .Y(n_1616) );
INVx2_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
XOR2x2_ASAP7_75t_L g760 ( .A(n_761), .B(n_826), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_762), .B(n_795), .Y(n_761) );
AOI22xp33_ASAP7_75t_L g762 ( .A1(n_763), .A2(n_765), .B1(n_793), .B2(n_794), .Y(n_762) );
AOI22xp5_ASAP7_75t_L g914 ( .A1(n_763), .A2(n_794), .B1(n_915), .B2(n_937), .Y(n_914) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
AOI31xp33_ASAP7_75t_L g985 ( .A1(n_764), .A2(n_986), .A3(n_994), .B(n_1002), .Y(n_985) );
AOI31xp33_ASAP7_75t_L g1601 ( .A1(n_764), .A2(n_1602), .A3(n_1612), .B(n_1620), .Y(n_1601) );
NAND3xp33_ASAP7_75t_L g765 ( .A(n_766), .B(n_780), .C(n_790), .Y(n_765) );
OAI22xp5_ASAP7_75t_L g821 ( .A1(n_767), .A2(n_792), .B1(n_822), .B2(n_823), .Y(n_821) );
INVx1_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
INVx2_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
BUFx2_ASAP7_75t_L g1001 ( .A(n_776), .Y(n_1001) );
INVx2_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
INVx2_ASAP7_75t_SL g923 ( .A(n_779), .Y(n_923) );
INVx1_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
INVx1_ASAP7_75t_L g876 ( .A(n_786), .Y(n_876) );
NOR3xp33_ASAP7_75t_L g795 ( .A(n_796), .B(n_803), .C(n_806), .Y(n_795) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_797), .B(n_800), .Y(n_796) );
OAI22xp33_ASAP7_75t_L g807 ( .A1(n_808), .A2(n_811), .B1(n_812), .B2(n_814), .Y(n_807) );
INVx2_ASAP7_75t_SL g808 ( .A(n_809), .Y(n_808) );
INVx2_ASAP7_75t_SL g809 ( .A(n_810), .Y(n_809) );
INVx2_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
OAI22xp5_ASAP7_75t_L g815 ( .A1(n_816), .A2(n_817), .B1(n_818), .B2(n_820), .Y(n_815) );
INVx1_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
HB1xp67_ASAP7_75t_L g900 ( .A(n_819), .Y(n_900) );
INVx1_ASAP7_75t_L g1057 ( .A(n_819), .Y(n_1057) );
INVx1_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
OAI22xp33_ASAP7_75t_L g1362 ( .A1(n_826), .A2(n_1363), .B1(n_1364), .B2(n_1365), .Y(n_1362) );
AO22x1_ASAP7_75t_SL g828 ( .A1(n_829), .A2(n_887), .B1(n_939), .B2(n_940), .Y(n_828) );
INVx1_ASAP7_75t_L g939 ( .A(n_829), .Y(n_939) );
NAND4xp25_ASAP7_75t_L g830 ( .A(n_831), .B(n_862), .C(n_864), .D(n_883), .Y(n_830) );
AOI21xp5_ASAP7_75t_L g833 ( .A1(n_834), .A2(n_840), .B(n_846), .Y(n_833) );
INVx2_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
INVx2_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
INVx2_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
INVx2_ASAP7_75t_L g1094 ( .A(n_839), .Y(n_1094) );
HB1xp67_ASAP7_75t_L g1163 ( .A(n_839), .Y(n_1163) );
INVx1_ASAP7_75t_L g1257 ( .A(n_839), .Y(n_1257) );
INVx1_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
INVx2_ASAP7_75t_L g843 ( .A(n_844), .Y(n_843) );
INVx2_ASAP7_75t_SL g844 ( .A(n_845), .Y(n_844) );
BUFx2_ASAP7_75t_L g906 ( .A(n_845), .Y(n_906) );
OAI22xp5_ASAP7_75t_L g875 ( .A1(n_848), .A2(n_849), .B1(n_876), .B2(n_877), .Y(n_875) );
OAI22xp5_ASAP7_75t_L g851 ( .A1(n_852), .A2(n_854), .B1(n_855), .B2(n_856), .Y(n_851) );
OAI22xp5_ASAP7_75t_L g1056 ( .A1(n_852), .A2(n_1011), .B1(n_1020), .B2(n_1057), .Y(n_1056) );
INVx1_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
INVx1_ASAP7_75t_L g902 ( .A(n_855), .Y(n_902) );
OAI22xp5_ASAP7_75t_L g1051 ( .A1(n_855), .A2(n_1052), .B1(n_1054), .B2(n_1055), .Y(n_1051) );
OAI21xp5_ASAP7_75t_SL g857 ( .A1(n_858), .A2(n_859), .B(n_860), .Y(n_857) );
INVx1_ASAP7_75t_L g866 ( .A(n_867), .Y(n_866) );
INVx1_ASAP7_75t_L g1024 ( .A(n_869), .Y(n_1024) );
INVx1_ASAP7_75t_L g1222 ( .A(n_870), .Y(n_1222) );
INVx1_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
INVx1_ASAP7_75t_L g877 ( .A(n_878), .Y(n_877) );
INVx1_ASAP7_75t_L g878 ( .A(n_879), .Y(n_878) );
INVx1_ASAP7_75t_L g940 ( .A(n_887), .Y(n_940) );
XNOR2x1_ASAP7_75t_L g887 ( .A(n_888), .B(n_938), .Y(n_887) );
NAND2x1_ASAP7_75t_L g888 ( .A(n_889), .B(n_914), .Y(n_888) );
AND4x1_ASAP7_75t_L g889 ( .A(n_890), .B(n_893), .C(n_907), .D(n_911), .Y(n_889) );
INVx1_ASAP7_75t_L g898 ( .A(n_899), .Y(n_898) );
INVx1_ASAP7_75t_L g1092 ( .A(n_899), .Y(n_1092) );
INVx1_ASAP7_75t_L g904 ( .A(n_905), .Y(n_904) );
OAI211xp5_ASAP7_75t_L g924 ( .A1(n_910), .A2(n_925), .B(n_926), .C(n_927), .Y(n_924) );
NAND3xp33_ASAP7_75t_L g915 ( .A(n_916), .B(n_928), .C(n_934), .Y(n_915) );
AOI21xp5_ASAP7_75t_SL g916 ( .A1(n_917), .A2(n_920), .B(n_921), .Y(n_916) );
INVx1_ASAP7_75t_L g917 ( .A(n_918), .Y(n_917) );
INVx1_ASAP7_75t_L g918 ( .A(n_919), .Y(n_918) );
AOI221xp5_ASAP7_75t_L g1019 ( .A1(n_919), .A2(n_1020), .B1(n_1021), .B2(n_1022), .C(n_1025), .Y(n_1019) );
OAI221xp5_ASAP7_75t_L g991 ( .A1(n_925), .A2(n_954), .B1(n_956), .B2(n_992), .C(n_993), .Y(n_991) );
OAI221xp5_ASAP7_75t_L g1611 ( .A1(n_925), .A2(n_993), .B1(n_1145), .B2(n_1581), .C(n_1583), .Y(n_1611) );
INVx2_ASAP7_75t_L g943 ( .A(n_944), .Y(n_943) );
XNOR2xp5_ASAP7_75t_L g944 ( .A(n_945), .B(n_1111), .Y(n_944) );
OAI22xp5_ASAP7_75t_L g945 ( .A1(n_946), .A2(n_947), .B1(n_1004), .B2(n_1110), .Y(n_945) );
INVx2_ASAP7_75t_L g946 ( .A(n_947), .Y(n_946) );
XNOR2x1_ASAP7_75t_L g947 ( .A(n_948), .B(n_1003), .Y(n_947) );
AND2x2_ASAP7_75t_L g948 ( .A(n_949), .B(n_983), .Y(n_948) );
NOR3xp33_ASAP7_75t_L g949 ( .A(n_950), .B(n_959), .C(n_960), .Y(n_949) );
NAND2xp5_ASAP7_75t_L g950 ( .A(n_951), .B(n_955), .Y(n_950) );
INVx1_ASAP7_75t_L g963 ( .A(n_964), .Y(n_963) );
INVx1_ASAP7_75t_L g968 ( .A(n_969), .Y(n_968) );
OAI22xp5_ASAP7_75t_L g971 ( .A1(n_972), .A2(n_973), .B1(n_974), .B2(n_975), .Y(n_971) );
OAI22xp5_ASAP7_75t_L g976 ( .A1(n_977), .A2(n_978), .B1(n_979), .B2(n_980), .Y(n_976) );
OAI221xp5_ASAP7_75t_L g1555 ( .A1(n_979), .A2(n_1556), .B1(n_1557), .B2(n_1558), .C(n_1559), .Y(n_1555) );
INVx2_ASAP7_75t_SL g1590 ( .A(n_979), .Y(n_1590) );
CKINVDCx8_ASAP7_75t_R g981 ( .A(n_982), .Y(n_981) );
OAI221xp5_ASAP7_75t_L g1141 ( .A1(n_992), .A2(n_1072), .B1(n_1133), .B2(n_1134), .C(n_1142), .Y(n_1141) );
INVx1_ASAP7_75t_L g996 ( .A(n_997), .Y(n_996) );
INVx1_ASAP7_75t_L g1231 ( .A(n_997), .Y(n_1231) );
OAI22xp5_ASAP7_75t_L g1537 ( .A1(n_997), .A2(n_1538), .B1(n_1539), .B2(n_1540), .Y(n_1537) );
HB1xp67_ASAP7_75t_L g998 ( .A(n_999), .Y(n_998) );
INVx2_ASAP7_75t_L g1110 ( .A(n_1004), .Y(n_1110) );
XOR2x2_ASAP7_75t_L g1004 ( .A(n_1005), .B(n_1061), .Y(n_1004) );
INVx1_ASAP7_75t_L g1059 ( .A(n_1006), .Y(n_1059) );
NAND2xp5_ASAP7_75t_L g1006 ( .A(n_1007), .B(n_1029), .Y(n_1006) );
NAND3xp33_ASAP7_75t_L g1008 ( .A(n_1009), .B(n_1012), .C(n_1019), .Y(n_1008) );
INVx1_ASAP7_75t_L g1013 ( .A(n_1014), .Y(n_1013) );
NOR3xp33_ASAP7_75t_L g1029 ( .A(n_1030), .B(n_1040), .C(n_1043), .Y(n_1029) );
NAND2xp5_ASAP7_75t_SL g1030 ( .A(n_1031), .B(n_1036), .Y(n_1030) );
AOI22xp33_ASAP7_75t_L g1031 ( .A1(n_1032), .A2(n_1033), .B1(n_1034), .B2(n_1035), .Y(n_1031) );
INVx2_ASAP7_75t_L g1106 ( .A(n_1033), .Y(n_1106) );
INVx1_ASAP7_75t_L g1107 ( .A(n_1035), .Y(n_1107) );
INVxp67_ASAP7_75t_L g1183 ( .A(n_1035), .Y(n_1183) );
INVx1_ASAP7_75t_L g1182 ( .A(n_1039), .Y(n_1182) );
OAI22xp33_ASAP7_75t_L g1044 ( .A1(n_1045), .A2(n_1047), .B1(n_1048), .B2(n_1050), .Y(n_1044) );
INVx2_ASAP7_75t_L g1045 ( .A(n_1046), .Y(n_1045) );
INVx1_ASAP7_75t_L g1048 ( .A(n_1049), .Y(n_1048) );
OAI22xp5_ASAP7_75t_L g1551 ( .A1(n_1052), .A2(n_1529), .B1(n_1530), .B2(n_1552), .Y(n_1551) );
INVx2_ASAP7_75t_L g1052 ( .A(n_1053), .Y(n_1052) );
INVx2_ASAP7_75t_SL g1253 ( .A(n_1053), .Y(n_1253) );
INVx2_ASAP7_75t_L g1556 ( .A(n_1053), .Y(n_1556) );
INVx1_ASAP7_75t_L g1109 ( .A(n_1062), .Y(n_1109) );
NAND4xp75_ASAP7_75t_L g1062 ( .A(n_1063), .B(n_1064), .C(n_1087), .D(n_1102), .Y(n_1062) );
OAI31xp33_ASAP7_75t_L g1064 ( .A1(n_1065), .A2(n_1075), .A3(n_1084), .B(n_1085), .Y(n_1064) );
OAI21xp33_ASAP7_75t_L g1070 ( .A1(n_1071), .A2(n_1072), .B(n_1073), .Y(n_1070) );
OAI221xp5_ASAP7_75t_L g1144 ( .A1(n_1072), .A2(n_1145), .B1(n_1147), .B2(n_1148), .C(n_1149), .Y(n_1144) );
OAI211xp5_ASAP7_75t_L g1079 ( .A1(n_1080), .A2(n_1081), .B(n_1082), .C(n_1083), .Y(n_1079) );
OAI22xp33_ASAP7_75t_L g1534 ( .A1(n_1081), .A2(n_1236), .B1(n_1535), .B2(n_1536), .Y(n_1534) );
INVx1_ASAP7_75t_L g1085 ( .A(n_1086), .Y(n_1085) );
OAI31xp33_ASAP7_75t_SL g1245 ( .A1(n_1086), .A2(n_1246), .A3(n_1247), .B(n_1259), .Y(n_1245) );
AND2x2_ASAP7_75t_SL g1087 ( .A(n_1088), .B(n_1101), .Y(n_1087) );
INVx1_ASAP7_75t_L g1552 ( .A(n_1093), .Y(n_1552) );
INVx1_ASAP7_75t_L g1093 ( .A(n_1094), .Y(n_1093) );
INVx2_ASAP7_75t_L g1098 ( .A(n_1099), .Y(n_1098) );
INVx2_ASAP7_75t_SL g1593 ( .A(n_1099), .Y(n_1593) );
AOI22xp33_ASAP7_75t_L g1111 ( .A1(n_1112), .A2(n_1215), .B1(n_1273), .B2(n_1274), .Y(n_1111) );
INVx1_ASAP7_75t_L g1273 ( .A(n_1112), .Y(n_1273) );
XNOR2x1_ASAP7_75t_L g1112 ( .A(n_1113), .B(n_1156), .Y(n_1112) );
INVx1_ASAP7_75t_L g1154 ( .A(n_1114), .Y(n_1154) );
NAND4xp25_ASAP7_75t_L g1114 ( .A(n_1115), .B(n_1136), .C(n_1138), .D(n_1150), .Y(n_1114) );
OAI21xp5_ASAP7_75t_L g1115 ( .A1(n_1116), .A2(n_1125), .B(n_1135), .Y(n_1115) );
AOI21xp5_ASAP7_75t_L g1120 ( .A1(n_1121), .A2(n_1123), .B(n_1124), .Y(n_1120) );
OAI22xp5_ASAP7_75t_L g1126 ( .A1(n_1127), .A2(n_1129), .B1(n_1130), .B2(n_1131), .Y(n_1126) );
OAI22xp5_ASAP7_75t_L g1159 ( .A1(n_1127), .A2(n_1160), .B1(n_1161), .B2(n_1162), .Y(n_1159) );
BUFx2_ASAP7_75t_L g1127 ( .A(n_1128), .Y(n_1127) );
OAI22xp33_ASAP7_75t_L g1221 ( .A1(n_1143), .A2(n_1222), .B1(n_1223), .B2(n_1235), .Y(n_1221) );
OAI33xp33_ASAP7_75t_L g1525 ( .A1(n_1143), .A2(n_1526), .A3(n_1527), .B1(n_1531), .B2(n_1534), .B3(n_1537), .Y(n_1525) );
INVx2_ASAP7_75t_L g1145 ( .A(n_1146), .Y(n_1145) );
INVx1_ASAP7_75t_SL g1214 ( .A(n_1157), .Y(n_1214) );
NAND4xp75_ASAP7_75t_L g1157 ( .A(n_1158), .B(n_1180), .C(n_1185), .D(n_1210), .Y(n_1157) );
INVx1_ASAP7_75t_L g1162 ( .A(n_1163), .Y(n_1162) );
OAI211xp5_ASAP7_75t_L g1200 ( .A1(n_1166), .A2(n_1201), .B(n_1202), .C(n_1204), .Y(n_1200) );
OAI22xp5_ASAP7_75t_L g1171 ( .A1(n_1172), .A2(n_1173), .B1(n_1175), .B2(n_1176), .Y(n_1171) );
BUFx2_ASAP7_75t_L g1173 ( .A(n_1174), .Y(n_1173) );
INVx1_ASAP7_75t_L g1178 ( .A(n_1179), .Y(n_1178) );
NOR2x1_ASAP7_75t_L g1180 ( .A(n_1181), .B(n_1184), .Y(n_1180) );
NAND2xp5_ASAP7_75t_L g1191 ( .A(n_1192), .B(n_1200), .Y(n_1191) );
OAI211xp5_ASAP7_75t_L g1192 ( .A1(n_1193), .A2(n_1194), .B(n_1197), .C(n_1198), .Y(n_1192) );
INVx1_ASAP7_75t_L g1194 ( .A(n_1195), .Y(n_1194) );
INVx1_ASAP7_75t_L g1195 ( .A(n_1196), .Y(n_1195) );
INVxp67_ASAP7_75t_SL g1274 ( .A(n_1215), .Y(n_1274) );
XNOR2xp5_ASAP7_75t_L g1215 ( .A(n_1216), .B(n_1217), .Y(n_1215) );
AND4x1_ASAP7_75t_L g1217 ( .A(n_1218), .B(n_1220), .C(n_1245), .D(n_1270), .Y(n_1217) );
NOR3xp33_ASAP7_75t_L g1220 ( .A(n_1221), .B(n_1243), .C(n_1244), .Y(n_1220) );
OAI221xp5_ASAP7_75t_L g1223 ( .A1(n_1224), .A2(n_1225), .B1(n_1226), .B2(n_1229), .C(n_1230), .Y(n_1223) );
OAI22xp33_ASAP7_75t_L g1531 ( .A1(n_1226), .A2(n_1236), .B1(n_1532), .B2(n_1533), .Y(n_1531) );
INVx2_ASAP7_75t_L g1226 ( .A(n_1227), .Y(n_1226) );
INVx1_ASAP7_75t_L g1227 ( .A(n_1228), .Y(n_1227) );
INVx1_ASAP7_75t_L g1232 ( .A(n_1233), .Y(n_1232) );
INVx1_ASAP7_75t_L g1233 ( .A(n_1234), .Y(n_1233) );
HB1xp67_ASAP7_75t_L g1619 ( .A(n_1234), .Y(n_1619) );
OAI221xp5_ASAP7_75t_L g1235 ( .A1(n_1236), .A2(n_1237), .B1(n_1238), .B2(n_1240), .C(n_1241), .Y(n_1235) );
INVx2_ASAP7_75t_L g1238 ( .A(n_1239), .Y(n_1238) );
INVx2_ASAP7_75t_L g1249 ( .A(n_1250), .Y(n_1249) );
OAI22xp5_ASAP7_75t_L g1251 ( .A1(n_1252), .A2(n_1254), .B1(n_1255), .B2(n_1258), .Y(n_1251) );
BUFx2_ASAP7_75t_L g1252 ( .A(n_1253), .Y(n_1252) );
INVx2_ASAP7_75t_SL g1255 ( .A(n_1256), .Y(n_1255) );
INVx1_ASAP7_75t_L g1256 ( .A(n_1257), .Y(n_1256) );
HB1xp67_ASAP7_75t_L g1266 ( .A(n_1267), .Y(n_1266) );
NOR2xp33_ASAP7_75t_L g1270 ( .A(n_1271), .B(n_1272), .Y(n_1270) );
OAI21xp33_ASAP7_75t_L g1275 ( .A1(n_1276), .A2(n_1284), .B(n_1517), .Y(n_1275) );
INVx1_ASAP7_75t_L g1276 ( .A(n_1277), .Y(n_1276) );
BUFx3_ASAP7_75t_L g1277 ( .A(n_1278), .Y(n_1277) );
INVx1_ASAP7_75t_L g1321 ( .A(n_1278), .Y(n_1321) );
AND2x4_ASAP7_75t_L g1278 ( .A(n_1279), .B(n_1282), .Y(n_1278) );
AND2x2_ASAP7_75t_L g1304 ( .A(n_1279), .B(n_1282), .Y(n_1304) );
HB1xp67_ASAP7_75t_L g1630 ( .A(n_1279), .Y(n_1630) );
INVx1_ASAP7_75t_L g1279 ( .A(n_1280), .Y(n_1279) );
AND2x4_ASAP7_75t_L g1305 ( .A(n_1280), .B(n_1282), .Y(n_1305) );
INVx1_ASAP7_75t_L g1280 ( .A(n_1281), .Y(n_1280) );
NAND2xp5_ASAP7_75t_L g1296 ( .A(n_1281), .B(n_1297), .Y(n_1296) );
INVx1_ASAP7_75t_L g1297 ( .A(n_1283), .Y(n_1297) );
NOR2xp33_ASAP7_75t_L g1284 ( .A(n_1285), .B(n_1449), .Y(n_1284) );
OAI211xp5_ASAP7_75t_L g1285 ( .A1(n_1286), .A2(n_1393), .B(n_1420), .C(n_1436), .Y(n_1285) );
AOI21xp33_ASAP7_75t_L g1286 ( .A1(n_1287), .A2(n_1368), .B(n_1369), .Y(n_1286) );
AOI21xp5_ASAP7_75t_L g1393 ( .A1(n_1287), .A2(n_1394), .B(n_1419), .Y(n_1393) );
OAI211xp5_ASAP7_75t_L g1287 ( .A1(n_1288), .A2(n_1309), .B(n_1325), .C(n_1350), .Y(n_1287) );
NOR2xp33_ASAP7_75t_L g1478 ( .A(n_1288), .B(n_1479), .Y(n_1478) );
INVx1_ASAP7_75t_L g1288 ( .A(n_1289), .Y(n_1288) );
AND2x2_ASAP7_75t_L g1289 ( .A(n_1290), .B(n_1306), .Y(n_1289) );
INVx1_ASAP7_75t_L g1376 ( .A(n_1290), .Y(n_1376) );
NOR2xp33_ASAP7_75t_L g1412 ( .A(n_1290), .B(n_1306), .Y(n_1412) );
INVx1_ASAP7_75t_L g1290 ( .A(n_1291), .Y(n_1290) );
AND2x2_ASAP7_75t_L g1327 ( .A(n_1291), .B(n_1328), .Y(n_1327) );
AND2x2_ASAP7_75t_L g1355 ( .A(n_1291), .B(n_1329), .Y(n_1355) );
INVx1_ASAP7_75t_L g1291 ( .A(n_1292), .Y(n_1291) );
AND2x2_ASAP7_75t_L g1346 ( .A(n_1292), .B(n_1347), .Y(n_1346) );
AND2x2_ASAP7_75t_L g1401 ( .A(n_1292), .B(n_1329), .Y(n_1401) );
AND2x2_ASAP7_75t_L g1292 ( .A(n_1293), .B(n_1303), .Y(n_1292) );
AND2x4_ASAP7_75t_L g1294 ( .A(n_1295), .B(n_1298), .Y(n_1294) );
INVx1_ASAP7_75t_L g1295 ( .A(n_1296), .Y(n_1295) );
OR2x2_ASAP7_75t_L g1339 ( .A(n_1296), .B(n_1299), .Y(n_1339) );
HB1xp67_ASAP7_75t_L g1629 ( .A(n_1297), .Y(n_1629) );
AND2x4_ASAP7_75t_L g1300 ( .A(n_1298), .B(n_1301), .Y(n_1300) );
INVx1_ASAP7_75t_L g1298 ( .A(n_1299), .Y(n_1298) );
OR2x2_ASAP7_75t_L g1342 ( .A(n_1299), .B(n_1302), .Y(n_1342) );
INVx1_ASAP7_75t_L g1301 ( .A(n_1302), .Y(n_1301) );
INVx2_ASAP7_75t_L g1323 ( .A(n_1305), .Y(n_1323) );
AND2x2_ASAP7_75t_L g1332 ( .A(n_1306), .B(n_1333), .Y(n_1332) );
AND2x2_ASAP7_75t_L g1345 ( .A(n_1306), .B(n_1346), .Y(n_1345) );
CKINVDCx5p33_ASAP7_75t_R g1357 ( .A(n_1306), .Y(n_1357) );
AND2x2_ASAP7_75t_L g1375 ( .A(n_1306), .B(n_1376), .Y(n_1375) );
OR2x2_ASAP7_75t_L g1385 ( .A(n_1306), .B(n_1376), .Y(n_1385) );
NAND2xp5_ASAP7_75t_L g1390 ( .A(n_1306), .B(n_1329), .Y(n_1390) );
AND2x2_ASAP7_75t_L g1391 ( .A(n_1306), .B(n_1355), .Y(n_1391) );
OR2x2_ASAP7_75t_L g1430 ( .A(n_1306), .B(n_1410), .Y(n_1430) );
NOR2xp33_ASAP7_75t_L g1439 ( .A(n_1306), .B(n_1409), .Y(n_1439) );
AND2x2_ASAP7_75t_L g1484 ( .A(n_1306), .B(n_1327), .Y(n_1484) );
AND2x4_ASAP7_75t_SL g1306 ( .A(n_1307), .B(n_1308), .Y(n_1306) );
INVx1_ASAP7_75t_L g1423 ( .A(n_1309), .Y(n_1423) );
NOR2xp33_ASAP7_75t_L g1447 ( .A(n_1309), .B(n_1448), .Y(n_1447) );
OR2x2_ASAP7_75t_L g1309 ( .A(n_1310), .B(n_1318), .Y(n_1309) );
INVx2_ASAP7_75t_L g1453 ( .A(n_1310), .Y(n_1453) );
INVx1_ASAP7_75t_L g1480 ( .A(n_1310), .Y(n_1480) );
NAND2xp5_ASAP7_75t_L g1310 ( .A(n_1311), .B(n_1315), .Y(n_1310) );
AND2x2_ASAP7_75t_L g1352 ( .A(n_1311), .B(n_1353), .Y(n_1352) );
INVx1_ASAP7_75t_L g1311 ( .A(n_1312), .Y(n_1311) );
INVx1_ASAP7_75t_L g1349 ( .A(n_1312), .Y(n_1349) );
AND2x2_ASAP7_75t_L g1371 ( .A(n_1312), .B(n_1353), .Y(n_1371) );
AND2x2_ASAP7_75t_L g1382 ( .A(n_1312), .B(n_1315), .Y(n_1382) );
AND2x2_ASAP7_75t_L g1418 ( .A(n_1312), .B(n_1318), .Y(n_1418) );
BUFx6f_ASAP7_75t_L g1426 ( .A(n_1312), .Y(n_1426) );
AND2x2_ASAP7_75t_L g1312 ( .A(n_1313), .B(n_1314), .Y(n_1312) );
AND2x2_ASAP7_75t_L g1343 ( .A(n_1315), .B(n_1344), .Y(n_1343) );
INVx1_ASAP7_75t_L g1353 ( .A(n_1315), .Y(n_1353) );
INVx1_ASAP7_75t_L g1392 ( .A(n_1315), .Y(n_1392) );
INVx1_ASAP7_75t_L g1416 ( .A(n_1315), .Y(n_1416) );
AOI321xp33_ASAP7_75t_L g1436 ( .A1(n_1315), .A2(n_1437), .A3(n_1440), .B1(n_1442), .B2(n_1444), .C(n_1447), .Y(n_1436) );
NAND2xp5_ASAP7_75t_SL g1442 ( .A(n_1315), .B(n_1443), .Y(n_1442) );
AND2x2_ASAP7_75t_L g1315 ( .A(n_1316), .B(n_1317), .Y(n_1315) );
CKINVDCx6p67_ASAP7_75t_R g1344 ( .A(n_1318), .Y(n_1344) );
NAND2xp5_ASAP7_75t_L g1367 ( .A(n_1318), .B(n_1359), .Y(n_1367) );
AND2x2_ASAP7_75t_L g1396 ( .A(n_1318), .B(n_1349), .Y(n_1396) );
NAND2xp5_ASAP7_75t_L g1414 ( .A(n_1318), .B(n_1415), .Y(n_1414) );
CKINVDCx5p33_ASAP7_75t_R g1419 ( .A(n_1318), .Y(n_1419) );
OR2x2_ASAP7_75t_L g1494 ( .A(n_1318), .B(n_1349), .Y(n_1494) );
OR2x6_ASAP7_75t_L g1318 ( .A(n_1319), .B(n_1320), .Y(n_1318) );
OR2x2_ASAP7_75t_L g1499 ( .A(n_1319), .B(n_1320), .Y(n_1499) );
OAI22xp5_ASAP7_75t_SL g1320 ( .A1(n_1321), .A2(n_1322), .B1(n_1323), .B2(n_1324), .Y(n_1320) );
INVx2_ASAP7_75t_L g1335 ( .A(n_1323), .Y(n_1335) );
INVx1_ASAP7_75t_L g1361 ( .A(n_1323), .Y(n_1361) );
AOI22xp5_ASAP7_75t_L g1325 ( .A1(n_1326), .A2(n_1343), .B1(n_1345), .B2(n_1348), .Y(n_1325) );
O2A1O1Ixp33_ASAP7_75t_L g1377 ( .A1(n_1326), .A2(n_1378), .B(n_1382), .C(n_1383), .Y(n_1377) );
AND2x2_ASAP7_75t_L g1326 ( .A(n_1327), .B(n_1332), .Y(n_1326) );
AND2x2_ASAP7_75t_L g1454 ( .A(n_1327), .B(n_1455), .Y(n_1454) );
AND2x2_ASAP7_75t_L g1475 ( .A(n_1327), .B(n_1357), .Y(n_1475) );
INVx1_ASAP7_75t_L g1328 ( .A(n_1329), .Y(n_1328) );
INVxp67_ASAP7_75t_SL g1347 ( .A(n_1329), .Y(n_1347) );
INVx1_ASAP7_75t_L g1410 ( .A(n_1329), .Y(n_1410) );
AND2x2_ASAP7_75t_L g1329 ( .A(n_1330), .B(n_1331), .Y(n_1329) );
AOI211xp5_ASAP7_75t_L g1397 ( .A1(n_1332), .A2(n_1384), .B(n_1398), .C(n_1402), .Y(n_1397) );
AND2x2_ASAP7_75t_L g1469 ( .A(n_1332), .B(n_1346), .Y(n_1469) );
AND2x2_ASAP7_75t_L g1482 ( .A(n_1332), .B(n_1355), .Y(n_1482) );
INVx2_ASAP7_75t_SL g1374 ( .A(n_1333), .Y(n_1374) );
BUFx2_ASAP7_75t_L g1380 ( .A(n_1333), .Y(n_1380) );
NOR2xp33_ASAP7_75t_L g1400 ( .A(n_1333), .B(n_1353), .Y(n_1400) );
BUFx3_ASAP7_75t_L g1407 ( .A(n_1333), .Y(n_1407) );
INVx2_ASAP7_75t_SL g1333 ( .A(n_1334), .Y(n_1333) );
AND2x2_ASAP7_75t_L g1356 ( .A(n_1334), .B(n_1357), .Y(n_1356) );
AND2x2_ASAP7_75t_L g1498 ( .A(n_1334), .B(n_1353), .Y(n_1498) );
OAI22xp33_ASAP7_75t_L g1336 ( .A1(n_1337), .A2(n_1338), .B1(n_1340), .B2(n_1341), .Y(n_1336) );
BUFx3_ASAP7_75t_L g1363 ( .A(n_1338), .Y(n_1363) );
BUFx6f_ASAP7_75t_L g1338 ( .A(n_1339), .Y(n_1338) );
HB1xp67_ASAP7_75t_L g1341 ( .A(n_1342), .Y(n_1341) );
INVx1_ASAP7_75t_L g1366 ( .A(n_1342), .Y(n_1366) );
AOI22xp33_ASAP7_75t_L g1490 ( .A1(n_1343), .A2(n_1388), .B1(n_1491), .B2(n_1493), .Y(n_1490) );
AND2x2_ASAP7_75t_L g1348 ( .A(n_1344), .B(n_1349), .Y(n_1348) );
NAND2xp5_ASAP7_75t_L g1368 ( .A(n_1344), .B(n_1358), .Y(n_1368) );
AND2x2_ASAP7_75t_L g1502 ( .A(n_1344), .B(n_1371), .Y(n_1502) );
INVx1_ASAP7_75t_L g1448 ( .A(n_1345), .Y(n_1448) );
INVx1_ASAP7_75t_L g1381 ( .A(n_1346), .Y(n_1381) );
AND2x2_ASAP7_75t_L g1432 ( .A(n_1346), .B(n_1357), .Y(n_1432) );
AND2x2_ASAP7_75t_L g1514 ( .A(n_1346), .B(n_1356), .Y(n_1514) );
INVx1_ASAP7_75t_L g1443 ( .A(n_1348), .Y(n_1443) );
AOI21xp33_ASAP7_75t_SL g1495 ( .A1(n_1348), .A2(n_1391), .B(n_1496), .Y(n_1495) );
NAND2xp5_ASAP7_75t_L g1441 ( .A(n_1349), .B(n_1358), .Y(n_1441) );
INVx1_ASAP7_75t_L g1509 ( .A(n_1349), .Y(n_1509) );
A2O1A1Ixp33_ASAP7_75t_SL g1350 ( .A1(n_1351), .A2(n_1354), .B(n_1358), .C(n_1367), .Y(n_1350) );
NOR2xp33_ASAP7_75t_L g1515 ( .A(n_1351), .B(n_1516), .Y(n_1515) );
INVx1_ASAP7_75t_L g1351 ( .A(n_1352), .Y(n_1351) );
AND2x2_ASAP7_75t_L g1458 ( .A(n_1352), .B(n_1374), .Y(n_1458) );
OAI21xp33_ASAP7_75t_L g1483 ( .A1(n_1352), .A2(n_1421), .B(n_1484), .Y(n_1483) );
OAI21xp5_ASAP7_75t_L g1487 ( .A1(n_1352), .A2(n_1472), .B(n_1488), .Y(n_1487) );
AND2x2_ASAP7_75t_L g1354 ( .A(n_1355), .B(n_1356), .Y(n_1354) );
INVx2_ASAP7_75t_L g1384 ( .A(n_1355), .Y(n_1384) );
OAI21xp5_ASAP7_75t_SL g1431 ( .A1(n_1355), .A2(n_1432), .B(n_1433), .Y(n_1431) );
NAND2xp5_ASAP7_75t_L g1446 ( .A(n_1355), .B(n_1374), .Y(n_1446) );
OR2x2_ASAP7_75t_L g1403 ( .A(n_1357), .B(n_1379), .Y(n_1403) );
AND2x2_ASAP7_75t_L g1421 ( .A(n_1357), .B(n_1422), .Y(n_1421) );
OR2x2_ASAP7_75t_L g1445 ( .A(n_1357), .B(n_1446), .Y(n_1445) );
AND2x2_ASAP7_75t_L g1461 ( .A(n_1357), .B(n_1401), .Y(n_1461) );
INVx2_ASAP7_75t_L g1435 ( .A(n_1358), .Y(n_1435) );
A2O1A1Ixp33_ASAP7_75t_L g1459 ( .A1(n_1358), .A2(n_1425), .B(n_1460), .C(n_1462), .Y(n_1459) );
INVx1_ASAP7_75t_L g1358 ( .A(n_1359), .Y(n_1358) );
INVx1_ASAP7_75t_L g1359 ( .A(n_1360), .Y(n_1359) );
INVx1_ASAP7_75t_L g1365 ( .A(n_1366), .Y(n_1365) );
INVx1_ASAP7_75t_L g1503 ( .A(n_1367), .Y(n_1503) );
OAI211xp5_ASAP7_75t_SL g1369 ( .A1(n_1370), .A2(n_1372), .B(n_1377), .C(n_1387), .Y(n_1369) );
A2O1A1Ixp33_ASAP7_75t_L g1451 ( .A1(n_1370), .A2(n_1372), .B(n_1389), .C(n_1452), .Y(n_1451) );
INVx1_ASAP7_75t_L g1370 ( .A(n_1371), .Y(n_1370) );
NAND2xp5_ASAP7_75t_L g1386 ( .A(n_1371), .B(n_1380), .Y(n_1386) );
INVx1_ASAP7_75t_L g1372 ( .A(n_1373), .Y(n_1372) );
AND2x2_ASAP7_75t_L g1373 ( .A(n_1374), .B(n_1375), .Y(n_1373) );
NOR2xp33_ASAP7_75t_L g1402 ( .A(n_1374), .B(n_1381), .Y(n_1402) );
AND2x2_ASAP7_75t_L g1411 ( .A(n_1374), .B(n_1412), .Y(n_1411) );
NOR2x1p5_ASAP7_75t_L g1422 ( .A(n_1374), .B(n_1384), .Y(n_1422) );
HB1xp67_ASAP7_75t_L g1474 ( .A(n_1374), .Y(n_1474) );
NAND2xp5_ASAP7_75t_L g1489 ( .A(n_1375), .B(n_1407), .Y(n_1489) );
INVx1_ASAP7_75t_L g1378 ( .A(n_1379), .Y(n_1378) );
OR2x2_ASAP7_75t_L g1379 ( .A(n_1380), .B(n_1381), .Y(n_1379) );
OR2x2_ASAP7_75t_L g1389 ( .A(n_1380), .B(n_1390), .Y(n_1389) );
NOR2xp33_ASAP7_75t_L g1429 ( .A(n_1380), .B(n_1430), .Y(n_1429) );
NAND2xp5_ASAP7_75t_L g1438 ( .A(n_1380), .B(n_1439), .Y(n_1438) );
INVx2_ASAP7_75t_L g1464 ( .A(n_1380), .Y(n_1464) );
AND2x2_ASAP7_75t_L g1508 ( .A(n_1380), .B(n_1509), .Y(n_1508) );
NOR2xp33_ASAP7_75t_L g1456 ( .A(n_1381), .B(n_1457), .Y(n_1456) );
INVx1_ASAP7_75t_L g1406 ( .A(n_1382), .Y(n_1406) );
AOI21xp33_ASAP7_75t_SL g1383 ( .A1(n_1384), .A2(n_1385), .B(n_1386), .Y(n_1383) );
OAI21xp33_ASAP7_75t_L g1491 ( .A1(n_1385), .A2(n_1464), .B(n_1492), .Y(n_1491) );
INVx1_ASAP7_75t_L g1433 ( .A(n_1386), .Y(n_1433) );
OAI21xp5_ASAP7_75t_L g1387 ( .A1(n_1388), .A2(n_1391), .B(n_1392), .Y(n_1387) );
INVx1_ASAP7_75t_L g1388 ( .A(n_1389), .Y(n_1388) );
INVx1_ASAP7_75t_L g1506 ( .A(n_1390), .Y(n_1506) );
NAND2xp67_ASAP7_75t_L g1468 ( .A(n_1392), .B(n_1469), .Y(n_1468) );
NAND2xp5_ASAP7_75t_L g1513 ( .A(n_1392), .B(n_1514), .Y(n_1513) );
OAI211xp5_ASAP7_75t_L g1394 ( .A1(n_1395), .A2(n_1397), .B(n_1403), .C(n_1404), .Y(n_1394) );
INVx1_ASAP7_75t_L g1395 ( .A(n_1396), .Y(n_1395) );
INVx1_ASAP7_75t_L g1398 ( .A(n_1399), .Y(n_1398) );
NAND2xp5_ASAP7_75t_L g1399 ( .A(n_1400), .B(n_1401), .Y(n_1399) );
NAND2xp5_ASAP7_75t_L g1477 ( .A(n_1400), .B(n_1475), .Y(n_1477) );
INVx1_ASAP7_75t_L g1500 ( .A(n_1401), .Y(n_1500) );
NAND2xp5_ASAP7_75t_L g1501 ( .A(n_1401), .B(n_1502), .Y(n_1501) );
INVx1_ASAP7_75t_L g1424 ( .A(n_1403), .Y(n_1424) );
A2O1A1Ixp33_ASAP7_75t_L g1404 ( .A1(n_1405), .A2(n_1408), .B(n_1411), .C(n_1413), .Y(n_1404) );
NOR2xp33_ASAP7_75t_L g1405 ( .A(n_1406), .B(n_1407), .Y(n_1405) );
O2A1O1Ixp33_ASAP7_75t_SL g1427 ( .A1(n_1406), .A2(n_1428), .B(n_1431), .C(n_1434), .Y(n_1427) );
INVx1_ASAP7_75t_L g1455 ( .A(n_1407), .Y(n_1455) );
NAND2xp5_ASAP7_75t_L g1460 ( .A(n_1407), .B(n_1461), .Y(n_1460) );
INVx1_ASAP7_75t_L g1408 ( .A(n_1409), .Y(n_1408) );
INVx1_ASAP7_75t_L g1409 ( .A(n_1410), .Y(n_1409) );
NAND2xp5_ASAP7_75t_L g1413 ( .A(n_1414), .B(n_1417), .Y(n_1413) );
INVx1_ASAP7_75t_L g1466 ( .A(n_1415), .Y(n_1466) );
INVx3_ASAP7_75t_L g1415 ( .A(n_1416), .Y(n_1415) );
INVx1_ASAP7_75t_L g1417 ( .A(n_1418), .Y(n_1417) );
AOI31xp33_ASAP7_75t_L g1470 ( .A1(n_1419), .A2(n_1471), .A3(n_1481), .B(n_1483), .Y(n_1470) );
AOI221xp5_ASAP7_75t_L g1420 ( .A1(n_1421), .A2(n_1423), .B1(n_1424), .B2(n_1425), .C(n_1427), .Y(n_1420) );
AOI211xp5_ASAP7_75t_L g1471 ( .A1(n_1425), .A2(n_1472), .B(n_1476), .C(n_1478), .Y(n_1471) );
CKINVDCx14_ASAP7_75t_R g1425 ( .A(n_1426), .Y(n_1425) );
OAI21xp33_ASAP7_75t_L g1481 ( .A1(n_1426), .A2(n_1467), .B(n_1482), .Y(n_1481) );
OAI221xp5_ASAP7_75t_L g1504 ( .A1(n_1426), .A2(n_1460), .B1(n_1505), .B2(n_1507), .C(n_1510), .Y(n_1504) );
INVxp67_ASAP7_75t_SL g1428 ( .A(n_1429), .Y(n_1428) );
INVx1_ASAP7_75t_L g1492 ( .A(n_1432), .Y(n_1492) );
AOI21xp5_ASAP7_75t_L g1452 ( .A1(n_1434), .A2(n_1453), .B(n_1454), .Y(n_1452) );
AOI22xp5_ASAP7_75t_L g1485 ( .A1(n_1434), .A2(n_1486), .B1(n_1503), .B2(n_1504), .Y(n_1485) );
INVx3_ASAP7_75t_L g1434 ( .A(n_1435), .Y(n_1434) );
INVx1_ASAP7_75t_L g1437 ( .A(n_1438), .Y(n_1437) );
AND2x2_ASAP7_75t_L g1463 ( .A(n_1439), .B(n_1464), .Y(n_1463) );
INVx1_ASAP7_75t_L g1440 ( .A(n_1441), .Y(n_1440) );
INVx2_ASAP7_75t_L g1444 ( .A(n_1445), .Y(n_1444) );
NAND2xp5_ASAP7_75t_L g1449 ( .A(n_1450), .B(n_1485), .Y(n_1449) );
O2A1O1Ixp33_ASAP7_75t_L g1450 ( .A1(n_1451), .A2(n_1456), .B(n_1459), .C(n_1470), .Y(n_1450) );
NAND2xp5_ASAP7_75t_L g1479 ( .A(n_1455), .B(n_1480), .Y(n_1479) );
INVx1_ASAP7_75t_L g1457 ( .A(n_1458), .Y(n_1457) );
INVx1_ASAP7_75t_L g1516 ( .A(n_1461), .Y(n_1516) );
AOI21xp5_ASAP7_75t_L g1462 ( .A1(n_1463), .A2(n_1465), .B(n_1467), .Y(n_1462) );
INVx1_ASAP7_75t_L g1465 ( .A(n_1466), .Y(n_1465) );
INVx1_ASAP7_75t_L g1511 ( .A(n_1466), .Y(n_1511) );
INVx1_ASAP7_75t_L g1467 ( .A(n_1468), .Y(n_1467) );
INVx1_ASAP7_75t_L g1472 ( .A(n_1473), .Y(n_1472) );
NAND2xp5_ASAP7_75t_L g1473 ( .A(n_1474), .B(n_1475), .Y(n_1473) );
NOR2xp33_ASAP7_75t_L g1505 ( .A(n_1475), .B(n_1506), .Y(n_1505) );
INVx1_ASAP7_75t_L g1476 ( .A(n_1477), .Y(n_1476) );
AOI211xp5_ASAP7_75t_SL g1510 ( .A1(n_1482), .A2(n_1511), .B(n_1512), .C(n_1515), .Y(n_1510) );
NAND4xp25_ASAP7_75t_L g1486 ( .A(n_1487), .B(n_1490), .C(n_1495), .D(n_1501), .Y(n_1486) );
INVxp67_ASAP7_75t_SL g1488 ( .A(n_1489), .Y(n_1488) );
INVx1_ASAP7_75t_L g1493 ( .A(n_1494), .Y(n_1493) );
NOR3xp33_ASAP7_75t_L g1496 ( .A(n_1497), .B(n_1499), .C(n_1500), .Y(n_1496) );
INVx1_ASAP7_75t_L g1497 ( .A(n_1498), .Y(n_1497) );
INVx1_ASAP7_75t_L g1507 ( .A(n_1508), .Y(n_1507) );
INVx1_ASAP7_75t_L g1512 ( .A(n_1513), .Y(n_1512) );
INVx1_ASAP7_75t_L g1518 ( .A(n_1519), .Y(n_1518) );
INVx1_ASAP7_75t_L g1519 ( .A(n_1520), .Y(n_1519) );
HB1xp67_ASAP7_75t_L g1520 ( .A(n_1521), .Y(n_1520) );
INVx1_ASAP7_75t_L g1521 ( .A(n_1522), .Y(n_1521) );
AND4x1_ASAP7_75t_L g1523 ( .A(n_1524), .B(n_1543), .C(n_1546), .D(n_1548), .Y(n_1523) );
NOR2xp33_ASAP7_75t_L g1543 ( .A(n_1544), .B(n_1545), .Y(n_1543) );
BUFx2_ASAP7_75t_L g1564 ( .A(n_1565), .Y(n_1564) );
INVx1_ASAP7_75t_L g1565 ( .A(n_1566), .Y(n_1565) );
INVx1_ASAP7_75t_L g1566 ( .A(n_1567), .Y(n_1566) );
INVxp67_ASAP7_75t_L g1568 ( .A(n_1569), .Y(n_1568) );
AND2x4_ASAP7_75t_L g1570 ( .A(n_1571), .B(n_1599), .Y(n_1570) );
AND4x1_ASAP7_75t_L g1571 ( .A(n_1572), .B(n_1578), .C(n_1582), .D(n_1586), .Y(n_1571) );
INVx1_ASAP7_75t_L g1575 ( .A(n_1576), .Y(n_1575) );
BUFx3_ASAP7_75t_L g1587 ( .A(n_1588), .Y(n_1587) );
INVx3_ASAP7_75t_L g1594 ( .A(n_1595), .Y(n_1594) );
INVx2_ASAP7_75t_SL g1606 ( .A(n_1607), .Y(n_1606) );
INVx1_ASAP7_75t_L g1615 ( .A(n_1616), .Y(n_1615) );
INVx1_ASAP7_75t_L g1623 ( .A(n_1624), .Y(n_1623) );
CKINVDCx5p33_ASAP7_75t_R g1624 ( .A(n_1625), .Y(n_1624) );
A2O1A1Ixp33_ASAP7_75t_L g1627 ( .A1(n_1626), .A2(n_1628), .B(n_1630), .C(n_1631), .Y(n_1627) );
INVx1_ASAP7_75t_L g1628 ( .A(n_1629), .Y(n_1628) );
endmodule