module fake_jpeg_18832_n_102 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_102);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_102;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

INVx6_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_4),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_2),
.B(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_25),
.B(n_33),
.Y(n_44)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_22),
.B(n_14),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_28),
.B(n_31),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_12),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_30),
.Y(n_37)
);

OAI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_12),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_22),
.B(n_3),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

OAI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_20),
.A2(n_4),
.B1(n_5),
.B2(n_8),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_4),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

CKINVDCx14_ASAP7_75t_R g56 ( 
.A(n_36),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_28),
.B(n_15),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_39),
.B(n_40),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_31),
.B(n_15),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_42),
.A2(n_13),
.B1(n_11),
.B2(n_23),
.Y(n_55)
);

NOR2x1_ASAP7_75t_L g43 ( 
.A(n_29),
.B(n_14),
.Y(n_43)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_32),
.B(n_16),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_46),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_25),
.B(n_16),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_25),
.B(n_17),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_17),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_35),
.A2(n_20),
.B1(n_24),
.B2(n_26),
.Y(n_50)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_54),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

A2O1A1O1Ixp25_ASAP7_75t_L g54 ( 
.A1(n_43),
.A2(n_32),
.B(n_27),
.C(n_33),
.D(n_21),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_58),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_SL g59 ( 
.A1(n_37),
.A2(n_13),
.B(n_11),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_63),
.Y(n_66)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_60),
.Y(n_68)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_62),
.B(n_41),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_43),
.A2(n_21),
.B1(n_23),
.B2(n_33),
.Y(n_63)
);

BUFx24_ASAP7_75t_SL g67 ( 
.A(n_61),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_67),
.B(n_70),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_37),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_69),
.B(n_74),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_57),
.B(n_38),
.Y(n_70)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_71),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_42),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g77 ( 
.A1(n_66),
.A2(n_54),
.B(n_59),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_80),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_72),
.B(n_56),
.C(n_63),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_81),
.C(n_82),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_65),
.B(n_38),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_55),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_66),
.B(n_44),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_74),
.A2(n_40),
.B(n_36),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_83),
.Y(n_84)
);

BUFx12f_ASAP7_75t_SL g85 ( 
.A(n_76),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_85),
.A2(n_84),
.B(n_86),
.Y(n_94)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_82),
.Y(n_87)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_87),
.Y(n_91)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_81),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_88),
.A2(n_68),
.B1(n_49),
.B2(n_41),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_89),
.B(n_72),
.C(n_75),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_90),
.B(n_93),
.C(n_91),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_92),
.B(n_60),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_89),
.B(n_79),
.C(n_73),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_94),
.A2(n_85),
.B(n_64),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_96),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_51),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_98),
.B(n_33),
.C(n_53),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_100),
.A2(n_99),
.B(n_35),
.Y(n_101)
);

BUFx24_ASAP7_75t_SL g102 ( 
.A(n_101),
.Y(n_102)
);


endmodule