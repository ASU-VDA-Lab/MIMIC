module real_aes_993_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_776, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_776;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_766;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_502;
wire n_434;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_753;
wire n_741;
wire n_283;
wire n_252;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_L g520 ( .A(n_0), .B(n_167), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_1), .B(n_771), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_2), .B(n_142), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_3), .B(n_169), .Y(n_181) );
INVx1_ASAP7_75t_L g138 ( .A(n_4), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_5), .B(n_142), .Y(n_480) );
NAND2xp33_ASAP7_75t_SL g539 ( .A(n_6), .B(n_148), .Y(n_539) );
INVx1_ASAP7_75t_L g532 ( .A(n_7), .Y(n_532) );
AOI22xp5_ASAP7_75t_L g751 ( .A1(n_8), .A2(n_60), .B1(n_752), .B2(n_753), .Y(n_751) );
CKINVDCx20_ASAP7_75t_R g752 ( .A(n_8), .Y(n_752) );
CKINVDCx16_ASAP7_75t_R g771 ( .A(n_9), .Y(n_771) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_10), .A2(n_105), .B1(n_766), .B2(n_774), .Y(n_104) );
AND2x2_ASAP7_75t_L g478 ( .A(n_11), .B(n_128), .Y(n_478) );
AND2x2_ASAP7_75t_L g172 ( .A(n_12), .B(n_173), .Y(n_172) );
AND2x2_ASAP7_75t_L g183 ( .A(n_13), .B(n_184), .Y(n_183) );
XNOR2xp5_ASAP7_75t_L g108 ( .A(n_14), .B(n_109), .Y(n_108) );
INVx2_ASAP7_75t_L g129 ( .A(n_15), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_16), .B(n_169), .Y(n_209) );
CKINVDCx16_ASAP7_75t_R g116 ( .A(n_17), .Y(n_116) );
NOR3xp33_ASAP7_75t_L g769 ( .A(n_17), .B(n_770), .C(n_772), .Y(n_769) );
AOI221x1_ASAP7_75t_L g535 ( .A1(n_18), .A2(n_150), .B1(n_173), .B2(n_536), .C(n_538), .Y(n_535) );
NAND2xp5_ASAP7_75t_SL g501 ( .A(n_19), .B(n_142), .Y(n_501) );
OAI22xp5_ASAP7_75t_SL g112 ( .A1(n_20), .A2(n_72), .B1(n_113), .B2(n_114), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g114 ( .A(n_20), .Y(n_114) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_21), .B(n_142), .Y(n_225) );
INVx1_ASAP7_75t_L g743 ( .A(n_22), .Y(n_743) );
AOI22xp5_ASAP7_75t_L g755 ( .A1(n_23), .A2(n_90), .B1(n_756), .B2(n_757), .Y(n_755) );
INVx1_ASAP7_75t_L g756 ( .A(n_23), .Y(n_756) );
AOI22xp33_ASAP7_75t_L g132 ( .A1(n_24), .A2(n_93), .B1(n_133), .B2(n_142), .Y(n_132) );
AOI21xp5_ASAP7_75t_L g481 ( .A1(n_25), .A2(n_150), .B(n_482), .Y(n_481) );
AOI221xp5_ASAP7_75t_SL g510 ( .A1(n_26), .A2(n_40), .B1(n_142), .B2(n_150), .C(n_511), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_27), .B(n_167), .Y(n_483) );
CKINVDCx20_ASAP7_75t_R g764 ( .A(n_28), .Y(n_764) );
OR2x2_ASAP7_75t_L g130 ( .A(n_29), .B(n_92), .Y(n_130) );
OA21x2_ASAP7_75t_L g162 ( .A1(n_29), .A2(n_92), .B(n_129), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_30), .B(n_169), .Y(n_505) );
INVxp67_ASAP7_75t_L g534 ( .A(n_31), .Y(n_534) );
AND2x2_ASAP7_75t_L g475 ( .A(n_32), .B(n_127), .Y(n_475) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_33), .A2(n_150), .B(n_519), .Y(n_518) );
AO21x2_ASAP7_75t_L g204 ( .A1(n_34), .A2(n_173), .B(n_205), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_35), .B(n_169), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g178 ( .A1(n_36), .A2(n_150), .B(n_179), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_37), .B(n_169), .Y(n_239) );
AND2x2_ASAP7_75t_L g140 ( .A(n_38), .B(n_141), .Y(n_140) );
AND2x2_ASAP7_75t_L g148 ( .A(n_38), .B(n_138), .Y(n_148) );
INVx1_ASAP7_75t_L g154 ( .A(n_38), .Y(n_154) );
OR2x6_ASAP7_75t_L g741 ( .A(n_39), .B(n_742), .Y(n_741) );
INVxp67_ASAP7_75t_L g772 ( .A(n_39), .Y(n_772) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_41), .B(n_142), .Y(n_182) );
AOI22xp5_ASAP7_75t_L g456 ( .A1(n_42), .A2(n_85), .B1(n_150), .B2(n_152), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_43), .B(n_169), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_44), .B(n_142), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_45), .B(n_167), .Y(n_473) );
AOI21xp5_ASAP7_75t_L g164 ( .A1(n_46), .A2(n_150), .B(n_165), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_47), .B(n_167), .Y(n_195) );
AND2x2_ASAP7_75t_L g523 ( .A(n_48), .B(n_127), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_49), .B(n_127), .Y(n_514) );
AOI22xp5_ASAP7_75t_SL g109 ( .A1(n_50), .A2(n_110), .B1(n_111), .B2(n_112), .Y(n_109) );
CKINVDCx20_ASAP7_75t_R g110 ( .A(n_50), .Y(n_110) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_51), .B(n_142), .Y(n_206) );
INVx1_ASAP7_75t_L g136 ( .A(n_52), .Y(n_136) );
INVx1_ASAP7_75t_L g145 ( .A(n_52), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_53), .B(n_169), .Y(n_168) );
AND2x2_ASAP7_75t_L g215 ( .A(n_54), .B(n_127), .Y(n_215) );
NAND2xp5_ASAP7_75t_SL g474 ( .A(n_55), .B(n_142), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_56), .B(n_167), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_57), .B(n_167), .Y(n_238) );
AND2x2_ASAP7_75t_L g466 ( .A(n_58), .B(n_127), .Y(n_466) );
NAND2xp5_ASAP7_75t_SL g171 ( .A(n_59), .B(n_142), .Y(n_171) );
CKINVDCx20_ASAP7_75t_R g753 ( .A(n_60), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_61), .B(n_169), .Y(n_521) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_62), .B(n_142), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g236 ( .A1(n_63), .A2(n_150), .B(n_237), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_64), .B(n_167), .Y(n_464) );
AND2x2_ASAP7_75t_SL g506 ( .A(n_65), .B(n_128), .Y(n_506) );
AND2x2_ASAP7_75t_L g231 ( .A(n_66), .B(n_128), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g470 ( .A1(n_67), .A2(n_150), .B(n_471), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_68), .B(n_169), .Y(n_484) );
AND2x2_ASAP7_75t_SL g457 ( .A(n_69), .B(n_184), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_70), .B(n_167), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_71), .B(n_167), .Y(n_210) );
CKINVDCx20_ASAP7_75t_R g113 ( .A(n_72), .Y(n_113) );
AOI22xp5_ASAP7_75t_L g149 ( .A1(n_73), .A2(n_95), .B1(n_150), .B2(n_152), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_74), .B(n_169), .Y(n_228) );
INVx1_ASAP7_75t_L g141 ( .A(n_75), .Y(n_141) );
INVx1_ASAP7_75t_L g147 ( .A(n_75), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_76), .B(n_167), .Y(n_180) );
AOI21xp5_ASAP7_75t_L g218 ( .A1(n_77), .A2(n_150), .B(n_219), .Y(n_218) );
CKINVDCx20_ASAP7_75t_R g745 ( .A(n_78), .Y(n_745) );
AOI21xp5_ASAP7_75t_L g192 ( .A1(n_79), .A2(n_150), .B(n_193), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_80), .A2(n_150), .B(n_208), .Y(n_207) );
AND2x2_ASAP7_75t_L g241 ( .A(n_81), .B(n_128), .Y(n_241) );
NAND2xp5_ASAP7_75t_SL g126 ( .A(n_82), .B(n_127), .Y(n_126) );
AOI22xp5_ASAP7_75t_L g455 ( .A1(n_83), .A2(n_87), .B1(n_133), .B2(n_142), .Y(n_455) );
NAND2xp5_ASAP7_75t_SL g465 ( .A(n_84), .B(n_142), .Y(n_465) );
INVx1_ASAP7_75t_L g744 ( .A(n_86), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_88), .B(n_167), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_89), .B(n_167), .Y(n_513) );
AND2x2_ASAP7_75t_L g196 ( .A(n_90), .B(n_184), .Y(n_196) );
CKINVDCx20_ASAP7_75t_R g757 ( .A(n_90), .Y(n_757) );
AOI21xp5_ASAP7_75t_L g461 ( .A1(n_91), .A2(n_150), .B(n_462), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_94), .B(n_169), .Y(n_463) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_96), .A2(n_150), .B(n_227), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_97), .B(n_169), .Y(n_194) );
BUFx2_ASAP7_75t_L g230 ( .A(n_98), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_99), .B(n_142), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_100), .B(n_169), .Y(n_472) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_101), .A2(n_150), .B(n_503), .Y(n_502) );
INVxp67_ASAP7_75t_L g537 ( .A(n_102), .Y(n_537) );
AO221x2_ASAP7_75t_L g105 ( .A1(n_103), .A2(n_106), .B1(n_749), .B2(n_759), .C(n_763), .Y(n_105) );
BUFx2_ASAP7_75t_L g762 ( .A(n_103), .Y(n_762) );
OAI22x1_ASAP7_75t_L g106 ( .A1(n_107), .A2(n_740), .B1(n_745), .B2(n_746), .Y(n_106) );
XNOR2xp5_ASAP7_75t_L g107 ( .A(n_108), .B(n_115), .Y(n_107) );
INVx1_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
OAI22xp5_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_117), .B1(n_446), .B2(n_739), .Y(n_115) );
CKINVDCx16_ASAP7_75t_R g739 ( .A(n_116), .Y(n_739) );
OR2x2_ASAP7_75t_L g748 ( .A(n_116), .B(n_741), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_116), .B(n_740), .Y(n_761) );
AND2x4_ASAP7_75t_L g117 ( .A(n_118), .B(n_371), .Y(n_117) );
NOR3xp33_ASAP7_75t_L g118 ( .A(n_119), .B(n_307), .C(n_354), .Y(n_118) );
NAND4xp25_ASAP7_75t_SL g119 ( .A(n_120), .B(n_242), .C(n_260), .D(n_286), .Y(n_119) );
OAI21xp33_ASAP7_75t_SL g120 ( .A1(n_121), .A2(n_200), .B(n_201), .Y(n_120) );
NAND2xp5_ASAP7_75t_SL g121 ( .A(n_122), .B(n_185), .Y(n_121) );
INVx1_ASAP7_75t_L g422 ( .A(n_122), .Y(n_422) );
OR2x2_ASAP7_75t_L g122 ( .A(n_123), .B(n_157), .Y(n_122) );
INVx2_ASAP7_75t_L g246 ( .A(n_123), .Y(n_246) );
AND2x2_ASAP7_75t_L g266 ( .A(n_123), .B(n_267), .Y(n_266) );
OR2x2_ASAP7_75t_L g368 ( .A(n_123), .B(n_187), .Y(n_368) );
AND2x2_ASAP7_75t_L g428 ( .A(n_123), .B(n_247), .Y(n_428) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_124), .B(n_281), .Y(n_280) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
OR2x2_ASAP7_75t_L g312 ( .A(n_125), .B(n_160), .Y(n_312) );
BUFx3_ASAP7_75t_L g322 ( .A(n_125), .Y(n_322) );
AND2x2_ASAP7_75t_L g385 ( .A(n_125), .B(n_386), .Y(n_385) );
AND2x4_ASAP7_75t_L g125 ( .A(n_126), .B(n_131), .Y(n_125) );
AND2x4_ASAP7_75t_L g199 ( .A(n_126), .B(n_131), .Y(n_199) );
AO21x2_ASAP7_75t_L g131 ( .A1(n_127), .A2(n_132), .B(n_149), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g176 ( .A(n_127), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g190 ( .A1(n_127), .A2(n_191), .B(n_192), .Y(n_190) );
OA21x2_ASAP7_75t_L g509 ( .A1(n_127), .A2(n_510), .B(n_514), .Y(n_509) );
BUFx6f_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
AND2x2_ASAP7_75t_SL g128 ( .A(n_129), .B(n_130), .Y(n_128) );
AND2x4_ASAP7_75t_L g211 ( .A(n_129), .B(n_130), .Y(n_211) );
AOI22xp5_ASAP7_75t_L g530 ( .A1(n_133), .A2(n_152), .B1(n_531), .B2(n_533), .Y(n_530) );
AND2x4_ASAP7_75t_L g133 ( .A(n_134), .B(n_139), .Y(n_133) );
AND2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_137), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
AND2x2_ASAP7_75t_L g151 ( .A(n_136), .B(n_138), .Y(n_151) );
AND2x4_ASAP7_75t_L g169 ( .A(n_136), .B(n_146), .Y(n_169) );
HB1xp67_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
BUFx3_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
AND2x6_ASAP7_75t_L g150 ( .A(n_140), .B(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g156 ( .A(n_141), .Y(n_156) );
AND2x6_ASAP7_75t_L g167 ( .A(n_141), .B(n_144), .Y(n_167) );
AND2x4_ASAP7_75t_L g142 ( .A(n_143), .B(n_148), .Y(n_142) );
INVx1_ASAP7_75t_L g540 ( .A(n_143), .Y(n_540) );
AND2x4_ASAP7_75t_L g143 ( .A(n_144), .B(n_146), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx5_ASAP7_75t_L g170 ( .A(n_148), .Y(n_170) );
AND2x4_ASAP7_75t_L g152 ( .A(n_151), .B(n_153), .Y(n_152) );
NOR2x1p5_ASAP7_75t_L g153 ( .A(n_154), .B(n_155), .Y(n_153) );
INVx3_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx1_ASAP7_75t_SL g157 ( .A(n_158), .Y(n_157) );
INVx1_ASAP7_75t_L g431 ( .A(n_158), .Y(n_431) );
AND2x2_ASAP7_75t_L g158 ( .A(n_159), .B(n_174), .Y(n_158) );
AND2x2_ASAP7_75t_L g198 ( .A(n_159), .B(n_199), .Y(n_198) );
INVx1_ASAP7_75t_L g386 ( .A(n_159), .Y(n_386) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
AND2x2_ASAP7_75t_L g200 ( .A(n_160), .B(n_189), .Y(n_200) );
AND2x2_ASAP7_75t_L g263 ( .A(n_160), .B(n_174), .Y(n_263) );
INVx2_ASAP7_75t_L g268 ( .A(n_160), .Y(n_268) );
AND2x2_ASAP7_75t_L g270 ( .A(n_160), .B(n_175), .Y(n_270) );
AO21x2_ASAP7_75t_L g160 ( .A1(n_161), .A2(n_163), .B(n_172), .Y(n_160) );
INVx4_ASAP7_75t_L g173 ( .A(n_161), .Y(n_173) );
AOI21x1_ASAP7_75t_L g516 ( .A1(n_161), .A2(n_517), .B(n_523), .Y(n_516) );
INVx3_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
BUFx4f_ASAP7_75t_L g184 ( .A(n_162), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_164), .B(n_171), .Y(n_163) );
AOI21xp5_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_168), .B(n_170), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_167), .B(n_230), .Y(n_229) );
AOI21xp5_ASAP7_75t_L g179 ( .A1(n_170), .A2(n_180), .B(n_181), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g193 ( .A1(n_170), .A2(n_194), .B(n_195), .Y(n_193) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_170), .A2(n_209), .B(n_210), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_170), .A2(n_220), .B(n_221), .Y(n_219) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_170), .A2(n_228), .B(n_229), .Y(n_227) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_170), .A2(n_238), .B(n_239), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g462 ( .A1(n_170), .A2(n_463), .B(n_464), .Y(n_462) );
AOI21xp5_ASAP7_75t_L g471 ( .A1(n_170), .A2(n_472), .B(n_473), .Y(n_471) );
AOI21xp5_ASAP7_75t_L g482 ( .A1(n_170), .A2(n_483), .B(n_484), .Y(n_482) );
AOI21xp5_ASAP7_75t_L g503 ( .A1(n_170), .A2(n_504), .B(n_505), .Y(n_503) );
AOI21xp5_ASAP7_75t_L g511 ( .A1(n_170), .A2(n_512), .B(n_513), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_170), .A2(n_520), .B(n_521), .Y(n_519) );
INVx3_ASAP7_75t_L g234 ( .A(n_173), .Y(n_234) );
INVx1_ASAP7_75t_L g248 ( .A(n_174), .Y(n_248) );
INVx2_ASAP7_75t_L g252 ( .A(n_174), .Y(n_252) );
AND2x4_ASAP7_75t_SL g283 ( .A(n_174), .B(n_189), .Y(n_283) );
HB1xp67_ASAP7_75t_L g315 ( .A(n_174), .Y(n_315) );
INVx3_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
HB1xp67_ASAP7_75t_L g197 ( .A(n_175), .Y(n_197) );
AOI21x1_ASAP7_75t_L g175 ( .A1(n_176), .A2(n_177), .B(n_183), .Y(n_175) );
AO21x2_ASAP7_75t_L g459 ( .A1(n_176), .A2(n_460), .B(n_466), .Y(n_459) );
AO21x2_ASAP7_75t_L g468 ( .A1(n_176), .A2(n_469), .B(n_475), .Y(n_468) );
AO21x2_ASAP7_75t_L g495 ( .A1(n_176), .A2(n_469), .B(n_475), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_178), .B(n_182), .Y(n_177) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_184), .A2(n_225), .B(n_226), .Y(n_224) );
INVx2_ASAP7_75t_SL g453 ( .A(n_184), .Y(n_453) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_184), .A2(n_501), .B(n_502), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_186), .B(n_198), .Y(n_185) );
AND2x2_ASAP7_75t_L g349 ( .A(n_186), .B(n_294), .Y(n_349) );
INVx2_ASAP7_75t_SL g437 ( .A(n_186), .Y(n_437) );
INVx1_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_188), .B(n_197), .Y(n_187) );
NAND2x1p5_ASAP7_75t_L g250 ( .A(n_188), .B(n_251), .Y(n_250) );
AND2x2_ASAP7_75t_L g357 ( .A(n_188), .B(n_270), .Y(n_357) );
INVx4_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
BUFx2_ASAP7_75t_L g245 ( .A(n_189), .Y(n_245) );
AND2x4_ASAP7_75t_L g247 ( .A(n_189), .B(n_248), .Y(n_247) );
NOR2x1_ASAP7_75t_L g267 ( .A(n_189), .B(n_268), .Y(n_267) );
INVx1_ASAP7_75t_L g340 ( .A(n_189), .Y(n_340) );
AND2x2_ASAP7_75t_L g359 ( .A(n_189), .B(n_298), .Y(n_359) );
AND2x2_ASAP7_75t_L g390 ( .A(n_189), .B(n_299), .Y(n_390) );
OR2x6_ASAP7_75t_L g189 ( .A(n_190), .B(n_196), .Y(n_189) );
AND2x2_ASAP7_75t_L g329 ( .A(n_198), .B(n_283), .Y(n_329) );
NAND2xp5_ASAP7_75t_SL g365 ( .A(n_198), .B(n_340), .Y(n_365) );
AOI22xp5_ASAP7_75t_L g439 ( .A1(n_198), .A2(n_440), .B1(n_442), .B2(n_443), .Y(n_439) );
AND2x2_ASAP7_75t_L g442 ( .A(n_198), .B(n_249), .Y(n_442) );
INVx3_ASAP7_75t_L g295 ( .A(n_199), .Y(n_295) );
AND2x2_ASAP7_75t_L g298 ( .A(n_199), .B(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g314 ( .A(n_200), .B(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g323 ( .A(n_200), .Y(n_323) );
AND2x4_ASAP7_75t_SL g201 ( .A(n_202), .B(n_212), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_202), .B(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g374 ( .A(n_202), .B(n_375), .Y(n_374) );
NOR3xp33_ASAP7_75t_L g426 ( .A(n_202), .B(n_336), .C(n_427), .Y(n_426) );
OR2x2_ASAP7_75t_L g444 ( .A(n_202), .B(n_338), .Y(n_444) );
INVx3_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
OR2x2_ASAP7_75t_L g259 ( .A(n_204), .B(n_223), .Y(n_259) );
INVx1_ASAP7_75t_L g276 ( .A(n_204), .Y(n_276) );
INVx2_ASAP7_75t_L g289 ( .A(n_204), .Y(n_289) );
HB1xp67_ASAP7_75t_L g304 ( .A(n_204), .Y(n_304) );
AND2x2_ASAP7_75t_L g318 ( .A(n_204), .B(n_291), .Y(n_318) );
AND2x2_ASAP7_75t_L g397 ( .A(n_204), .B(n_214), .Y(n_397) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_206), .A2(n_207), .B(n_211), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_211), .A2(n_217), .B(n_218), .Y(n_216) );
AOI21xp5_ASAP7_75t_L g479 ( .A1(n_211), .A2(n_480), .B(n_481), .Y(n_479) );
NOR2xp33_ASAP7_75t_L g531 ( .A(n_211), .B(n_532), .Y(n_531) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_211), .B(n_534), .Y(n_533) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_211), .B(n_537), .Y(n_536) );
NOR3xp33_ASAP7_75t_L g538 ( .A(n_211), .B(n_539), .C(n_540), .Y(n_538) );
AOI221xp5_ASAP7_75t_L g260 ( .A1(n_212), .A2(n_261), .B1(n_264), .B2(n_271), .C(n_277), .Y(n_260) );
AOI221xp5_ASAP7_75t_L g389 ( .A1(n_212), .A2(n_390), .B1(n_391), .B2(n_392), .C(n_393), .Y(n_389) );
AND2x2_ASAP7_75t_L g212 ( .A(n_213), .B(n_222), .Y(n_212) );
INVx2_ASAP7_75t_L g331 ( .A(n_213), .Y(n_331) );
AND2x2_ASAP7_75t_L g391 ( .A(n_213), .B(n_275), .Y(n_391) );
AND2x2_ASAP7_75t_L g401 ( .A(n_213), .B(n_287), .Y(n_401) );
OR2x2_ASAP7_75t_L g441 ( .A(n_213), .B(n_325), .Y(n_441) );
INVx2_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
OR2x2_ASAP7_75t_SL g258 ( .A(n_214), .B(n_259), .Y(n_258) );
NAND2x1_ASAP7_75t_L g274 ( .A(n_214), .B(n_223), .Y(n_274) );
INVx4_ASAP7_75t_L g303 ( .A(n_214), .Y(n_303) );
OR2x2_ASAP7_75t_L g345 ( .A(n_214), .B(n_232), .Y(n_345) );
OR2x6_ASAP7_75t_L g214 ( .A(n_215), .B(n_216), .Y(n_214) );
AND2x2_ASAP7_75t_L g396 ( .A(n_222), .B(n_397), .Y(n_396) );
AND2x2_ASAP7_75t_L g222 ( .A(n_223), .B(n_232), .Y(n_222) );
INVx2_ASAP7_75t_SL g284 ( .A(n_223), .Y(n_284) );
NOR2x1_ASAP7_75t_SL g290 ( .A(n_223), .B(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g305 ( .A(n_223), .B(n_306), .Y(n_305) );
OR2x2_ASAP7_75t_L g336 ( .A(n_223), .B(n_303), .Y(n_336) );
AND2x2_ASAP7_75t_L g343 ( .A(n_223), .B(n_289), .Y(n_343) );
BUFx2_ASAP7_75t_L g377 ( .A(n_223), .Y(n_377) );
AND2x2_ASAP7_75t_L g388 ( .A(n_223), .B(n_303), .Y(n_388) );
OR2x6_ASAP7_75t_L g223 ( .A(n_224), .B(n_231), .Y(n_223) );
HB1xp67_ASAP7_75t_L g256 ( .A(n_232), .Y(n_256) );
AND2x2_ASAP7_75t_L g275 ( .A(n_232), .B(n_276), .Y(n_275) );
INVx2_ASAP7_75t_L g306 ( .A(n_232), .Y(n_306) );
AND2x2_ASAP7_75t_L g332 ( .A(n_232), .B(n_288), .Y(n_332) );
INVx3_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
AO21x2_ASAP7_75t_L g233 ( .A1(n_234), .A2(n_235), .B(n_241), .Y(n_233) );
AO21x1_ASAP7_75t_SL g291 ( .A1(n_234), .A2(n_235), .B(n_241), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_236), .B(n_240), .Y(n_235) );
OAI31xp33_ASAP7_75t_L g242 ( .A1(n_243), .A2(n_247), .A3(n_249), .B(n_253), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_245), .B(n_246), .Y(n_244) );
INVx2_ASAP7_75t_L g351 ( .A(n_245), .Y(n_351) );
NOR2xp67_ASAP7_75t_L g261 ( .A(n_246), .B(n_262), .Y(n_261) );
AOI322xp5_ASAP7_75t_L g341 ( .A1(n_246), .A2(n_335), .A3(n_342), .B1(n_346), .B2(n_347), .C1(n_349), .C2(n_350), .Y(n_341) );
AND2x2_ASAP7_75t_L g413 ( .A(n_246), .B(n_390), .Y(n_413) );
AOI221xp5_ASAP7_75t_SL g326 ( .A1(n_247), .A2(n_327), .B1(n_329), .B2(n_330), .C(n_333), .Y(n_326) );
INVx2_ASAP7_75t_L g346 ( .A(n_247), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_249), .B(n_311), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_249), .B(n_342), .Y(n_445) );
INVx1_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
OR2x2_ASAP7_75t_L g320 ( .A(n_250), .B(n_295), .Y(n_320) );
INVx1_ASAP7_75t_SL g251 ( .A(n_252), .Y(n_251) );
AND2x2_ASAP7_75t_L g299 ( .A(n_252), .B(n_268), .Y(n_299) );
AND2x4_ASAP7_75t_L g253 ( .A(n_254), .B(n_257), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
INVx1_ASAP7_75t_L g370 ( .A(n_256), .Y(n_370) );
O2A1O1Ixp5_ASAP7_75t_L g361 ( .A1(n_257), .A2(n_362), .B(n_364), .C(n_366), .Y(n_361) );
INVx2_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
OAI22xp5_ASAP7_75t_L g393 ( .A1(n_258), .A2(n_394), .B1(n_395), .B2(n_398), .Y(n_393) );
OR2x2_ASAP7_75t_L g348 ( .A(n_259), .B(n_345), .Y(n_348) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
NAND2xp5_ASAP7_75t_SL g264 ( .A(n_265), .B(n_269), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
INVx1_ASAP7_75t_L g281 ( .A(n_268), .Y(n_281) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_270), .B(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_273), .B(n_275), .Y(n_272) );
INVx3_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
OR2x2_ASAP7_75t_L g324 ( .A(n_274), .B(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_274), .B(n_275), .Y(n_367) );
OR2x2_ASAP7_75t_L g369 ( .A(n_274), .B(n_370), .Y(n_369) );
NOR2xp33_ASAP7_75t_L g417 ( .A(n_274), .B(n_418), .Y(n_417) );
BUFx2_ASAP7_75t_L g285 ( .A(n_276), .Y(n_285) );
NOR4xp25_ASAP7_75t_L g277 ( .A(n_278), .B(n_282), .C(n_284), .D(n_285), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g405 ( .A(n_279), .B(n_406), .Y(n_405) );
AND2x2_ASAP7_75t_L g433 ( .A(n_279), .B(n_282), .Y(n_433) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
INVx1_ASAP7_75t_L g363 ( .A(n_281), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_282), .B(n_311), .Y(n_398) );
AOI321xp33_ASAP7_75t_L g400 ( .A1(n_282), .A2(n_401), .A3(n_402), .B1(n_403), .B2(n_405), .C(n_408), .Y(n_400) );
INVx2_ASAP7_75t_SL g282 ( .A(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_SL g362 ( .A(n_283), .B(n_363), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_283), .B(n_322), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_284), .B(n_306), .Y(n_411) );
OR2x2_ASAP7_75t_L g438 ( .A(n_285), .B(n_322), .Y(n_438) );
AOI21xp5_ASAP7_75t_L g286 ( .A1(n_287), .A2(n_292), .B(n_296), .Y(n_286) );
AND2x2_ASAP7_75t_L g327 ( .A(n_287), .B(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_290), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g353 ( .A(n_289), .B(n_291), .Y(n_353) );
INVx2_ASAP7_75t_L g338 ( .A(n_290), .Y(n_338) );
INVx1_ASAP7_75t_SL g292 ( .A(n_293), .Y(n_292) );
NOR2xp33_ASAP7_75t_L g408 ( .A(n_293), .B(n_409), .Y(n_408) );
OR2x2_ASAP7_75t_L g394 ( .A(n_294), .B(n_346), .Y(n_394) );
INVx2_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g352 ( .A(n_295), .B(n_353), .Y(n_352) );
NOR2x1_ASAP7_75t_L g430 ( .A(n_295), .B(n_431), .Y(n_430) );
NOR2xp67_ASAP7_75t_L g296 ( .A(n_297), .B(n_300), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g381 ( .A(n_299), .Y(n_381) );
INVx2_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g301 ( .A(n_302), .B(n_305), .Y(n_301) );
NOR2xp67_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_303), .B(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g328 ( .A(n_303), .Y(n_328) );
BUFx2_ASAP7_75t_L g410 ( .A(n_303), .Y(n_410) );
INVxp67_ASAP7_75t_L g418 ( .A(n_306), .Y(n_418) );
NAND3xp33_ASAP7_75t_L g307 ( .A(n_308), .B(n_326), .C(n_341), .Y(n_307) );
AOI21xp5_ASAP7_75t_L g308 ( .A1(n_309), .A2(n_316), .B(n_319), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_310), .B(n_313), .Y(n_309) );
INVx2_ASAP7_75t_SL g311 ( .A(n_312), .Y(n_311) );
OR2x2_ASAP7_75t_L g339 ( .A(n_312), .B(n_340), .Y(n_339) );
INVx2_ASAP7_75t_L g392 ( .A(n_313), .Y(n_392) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx2_ASAP7_75t_L g407 ( .A(n_315), .Y(n_407) );
AOI21xp5_ASAP7_75t_L g412 ( .A1(n_316), .A2(n_413), .B(n_414), .Y(n_412) );
INVx1_ASAP7_75t_SL g316 ( .A(n_317), .Y(n_316) );
INVx2_ASAP7_75t_SL g325 ( .A(n_318), .Y(n_325) );
AND2x2_ASAP7_75t_L g387 ( .A(n_318), .B(n_388), .Y(n_387) );
AOI21xp33_ASAP7_75t_L g319 ( .A1(n_320), .A2(n_321), .B(n_324), .Y(n_319) );
OAI22xp5_ASAP7_75t_L g366 ( .A1(n_320), .A2(n_367), .B1(n_368), .B2(n_369), .Y(n_366) );
OR2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
INVx1_ASAP7_75t_L g356 ( .A(n_322), .Y(n_356) );
OR2x2_ASAP7_75t_L g404 ( .A(n_325), .B(n_336), .Y(n_404) );
NOR4xp25_ASAP7_75t_L g436 ( .A(n_328), .B(n_377), .C(n_437), .D(n_438), .Y(n_436) );
AND2x2_ASAP7_75t_L g330 ( .A(n_331), .B(n_332), .Y(n_330) );
OR2x2_ASAP7_75t_L g337 ( .A(n_331), .B(n_338), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_331), .B(n_353), .Y(n_435) );
AOI21xp33_ASAP7_75t_SL g333 ( .A1(n_334), .A2(n_337), .B(n_339), .Y(n_333) );
INVx2_ASAP7_75t_SL g335 ( .A(n_336), .Y(n_335) );
OR2x2_ASAP7_75t_L g424 ( .A(n_336), .B(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g432 ( .A(n_338), .Y(n_432) );
AND2x4_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
INVxp67_ASAP7_75t_L g360 ( .A(n_343), .Y(n_360) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
OR2x2_ASAP7_75t_L g376 ( .A(n_345), .B(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g350 ( .A(n_351), .B(n_352), .Y(n_350) );
AND2x2_ASAP7_75t_L g379 ( .A(n_351), .B(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g425 ( .A(n_353), .Y(n_425) );
A2O1A1Ixp33_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_358), .B(n_360), .C(n_361), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_356), .B(n_357), .Y(n_355) );
INVx1_ASAP7_75t_L g415 ( .A(n_357), .Y(n_415) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVxp67_ASAP7_75t_L g419 ( .A(n_362), .Y(n_419) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
NOR3xp33_ASAP7_75t_L g371 ( .A(n_372), .B(n_399), .C(n_420), .Y(n_371) );
OAI211xp5_ASAP7_75t_SL g372 ( .A1(n_373), .A2(n_378), .B(n_382), .C(n_389), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_SL g375 ( .A(n_376), .Y(n_375) );
INVxp67_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx2_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
OAI21xp5_ASAP7_75t_SL g382 ( .A1(n_383), .A2(n_385), .B(n_387), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
O2A1O1Ixp33_ASAP7_75t_L g421 ( .A1(n_385), .A2(n_422), .B(n_423), .C(n_426), .Y(n_421) );
BUFx2_ASAP7_75t_L g402 ( .A(n_386), .Y(n_402) );
INVx2_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_400), .B(n_412), .Y(n_399) );
INVx2_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx2_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
OAI22xp5_ASAP7_75t_L g414 ( .A1(n_409), .A2(n_415), .B1(n_416), .B2(n_419), .Y(n_414) );
OR2x2_ASAP7_75t_L g409 ( .A(n_410), .B(n_411), .Y(n_409) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
NAND4xp25_ASAP7_75t_L g420 ( .A(n_421), .B(n_429), .C(n_439), .D(n_445), .Y(n_420) );
INVx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
AOI221xp5_ASAP7_75t_L g429 ( .A1(n_430), .A2(n_432), .B1(n_433), .B2(n_434), .C(n_436), .Y(n_429) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
XNOR2x1_ASAP7_75t_L g750 ( .A(n_446), .B(n_751), .Y(n_750) );
AND3x4_ASAP7_75t_L g446 ( .A(n_447), .B(n_610), .C(n_684), .Y(n_446) );
NOR3xp33_ASAP7_75t_L g447 ( .A(n_448), .B(n_552), .C(n_583), .Y(n_447) );
A2O1A1Ixp33_ASAP7_75t_L g448 ( .A1(n_449), .A2(n_487), .B(n_496), .C(n_524), .Y(n_448) );
AOI21x1_ASAP7_75t_SL g449 ( .A1(n_450), .A2(n_467), .B(n_485), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g585 ( .A1(n_450), .A2(n_586), .B1(n_592), .B2(n_595), .Y(n_585) );
AND2x2_ASAP7_75t_L g719 ( .A(n_450), .B(n_489), .Y(n_719) );
AND2x2_ASAP7_75t_L g450 ( .A(n_451), .B(n_458), .Y(n_450) );
BUFx2_ASAP7_75t_L g492 ( .A(n_451), .Y(n_492) );
AND2x2_ASAP7_75t_L g578 ( .A(n_451), .B(n_459), .Y(n_578) );
AND2x2_ASAP7_75t_L g649 ( .A(n_451), .B(n_495), .Y(n_649) );
INVx2_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
BUFx6f_ASAP7_75t_L g543 ( .A(n_452), .Y(n_543) );
AOI21x1_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_454), .B(n_457), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_455), .B(n_456), .Y(n_454) );
AND2x4_ASAP7_75t_L g542 ( .A(n_458), .B(n_543), .Y(n_542) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
AND2x2_ASAP7_75t_L g486 ( .A(n_459), .B(n_477), .Y(n_486) );
OR2x2_ASAP7_75t_L g494 ( .A(n_459), .B(n_495), .Y(n_494) );
AND2x4_ASAP7_75t_L g547 ( .A(n_459), .B(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g594 ( .A(n_459), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_459), .B(n_495), .Y(n_602) );
AND2x2_ASAP7_75t_L g639 ( .A(n_459), .B(n_543), .Y(n_639) );
HB1xp67_ASAP7_75t_L g648 ( .A(n_459), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_459), .B(n_476), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_461), .B(n_465), .Y(n_460) );
INVx2_ASAP7_75t_L g581 ( .A(n_467), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_467), .B(n_542), .Y(n_637) );
HB1xp67_ASAP7_75t_L g738 ( .A(n_467), .Y(n_738) );
AND2x4_ASAP7_75t_L g467 ( .A(n_468), .B(n_476), .Y(n_467) );
AND2x2_ASAP7_75t_L g485 ( .A(n_468), .B(n_486), .Y(n_485) );
OR2x2_ASAP7_75t_L g563 ( .A(n_468), .B(n_477), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_468), .B(n_594), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_470), .B(n_474), .Y(n_469) );
AND2x2_ASAP7_75t_L g630 ( .A(n_476), .B(n_547), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_476), .B(n_542), .Y(n_686) );
INVx5_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx2_ASAP7_75t_L g490 ( .A(n_477), .Y(n_490) );
AND2x2_ASAP7_75t_L g557 ( .A(n_477), .B(n_548), .Y(n_557) );
HB1xp67_ASAP7_75t_L g577 ( .A(n_477), .Y(n_577) );
AND2x4_ASAP7_75t_L g584 ( .A(n_477), .B(n_495), .Y(n_584) );
AND2x2_ASAP7_75t_SL g731 ( .A(n_477), .B(n_543), .Y(n_731) );
OR2x6_ASAP7_75t_L g477 ( .A(n_478), .B(n_479), .Y(n_477) );
INVx1_ASAP7_75t_L g710 ( .A(n_485), .Y(n_710) );
INVx1_ASAP7_75t_L g652 ( .A(n_486), .Y(n_652) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_489), .B(n_491), .Y(n_488) );
INVx2_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
OR2x2_ASAP7_75t_L g574 ( .A(n_490), .B(n_494), .Y(n_574) );
NOR2xp33_ASAP7_75t_L g667 ( .A(n_490), .B(n_543), .Y(n_667) );
AND2x2_ASAP7_75t_L g669 ( .A(n_490), .B(n_493), .Y(n_669) );
AOI32xp33_ASAP7_75t_L g735 ( .A1(n_490), .A2(n_551), .A3(n_706), .B1(n_736), .B2(n_738), .Y(n_735) );
AND2x2_ASAP7_75t_L g491 ( .A(n_492), .B(n_493), .Y(n_491) );
AND2x2_ASAP7_75t_L g561 ( .A(n_492), .B(n_562), .Y(n_561) );
OR2x2_ASAP7_75t_L g679 ( .A(n_492), .B(n_680), .Y(n_679) );
OR2x2_ASAP7_75t_L g702 ( .A(n_492), .B(n_563), .Y(n_702) );
AND2x2_ASAP7_75t_L g729 ( .A(n_492), .B(n_630), .Y(n_729) );
AND2x2_ASAP7_75t_L g655 ( .A(n_493), .B(n_543), .Y(n_655) );
AND2x2_ASAP7_75t_L g730 ( .A(n_493), .B(n_731), .Y(n_730) );
INVx2_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx2_ASAP7_75t_L g548 ( .A(n_495), .Y(n_548) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_498), .B(n_507), .Y(n_497) );
NOR2x1p5_ASAP7_75t_L g588 ( .A(n_498), .B(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g606 ( .A(n_498), .Y(n_606) );
OR2x2_ASAP7_75t_L g634 ( .A(n_498), .B(n_635), .Y(n_634) );
INVx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
AND2x4_ASAP7_75t_SL g551 ( .A(n_499), .B(n_529), .Y(n_551) );
AND2x4_ASAP7_75t_L g567 ( .A(n_499), .B(n_568), .Y(n_567) );
OR2x2_ASAP7_75t_L g570 ( .A(n_499), .B(n_571), .Y(n_570) );
OR2x2_ASAP7_75t_L g598 ( .A(n_499), .B(n_509), .Y(n_598) );
OR2x2_ASAP7_75t_L g623 ( .A(n_499), .B(n_572), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_499), .B(n_628), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_499), .B(n_509), .Y(n_658) );
INVx2_ASAP7_75t_L g674 ( .A(n_499), .Y(n_674) );
AND2x2_ASAP7_75t_L g689 ( .A(n_499), .B(n_528), .Y(n_689) );
HB1xp67_ASAP7_75t_L g713 ( .A(n_499), .Y(n_713) );
INVx1_ASAP7_75t_L g718 ( .A(n_499), .Y(n_718) );
OR2x6_ASAP7_75t_L g499 ( .A(n_500), .B(n_506), .Y(n_499) );
AND2x2_ASAP7_75t_L g582 ( .A(n_507), .B(n_567), .Y(n_582) );
AND2x2_ASAP7_75t_L g603 ( .A(n_507), .B(n_551), .Y(n_603) );
INVx1_ASAP7_75t_L g635 ( .A(n_507), .Y(n_635) );
AND2x2_ASAP7_75t_L g507 ( .A(n_508), .B(n_515), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx1_ASAP7_75t_L g527 ( .A(n_509), .Y(n_527) );
INVx2_ASAP7_75t_L g572 ( .A(n_509), .Y(n_572) );
BUFx3_ASAP7_75t_L g589 ( .A(n_509), .Y(n_589) );
AND2x2_ASAP7_75t_L g628 ( .A(n_509), .B(n_515), .Y(n_628) );
HB1xp67_ASAP7_75t_L g726 ( .A(n_509), .Y(n_726) );
INVx2_ASAP7_75t_L g541 ( .A(n_515), .Y(n_541) );
HB1xp67_ASAP7_75t_L g550 ( .A(n_515), .Y(n_550) );
INVx1_ASAP7_75t_L g566 ( .A(n_515), .Y(n_566) );
OR2x2_ASAP7_75t_L g571 ( .A(n_515), .B(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g591 ( .A(n_515), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_515), .B(n_568), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_515), .B(n_674), .Y(n_673) );
INVx3_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_518), .B(n_522), .Y(n_517) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_525), .A2(n_542), .B(n_544), .Y(n_524) );
AND2x2_ASAP7_75t_SL g525 ( .A(n_526), .B(n_528), .Y(n_525) );
HB1xp67_ASAP7_75t_L g734 ( .A(n_526), .Y(n_734) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVxp67_ASAP7_75t_SL g560 ( .A(n_527), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_527), .B(n_566), .Y(n_608) );
HB1xp67_ASAP7_75t_L g723 ( .A(n_527), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_528), .B(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g613 ( .A(n_528), .B(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g664 ( .A(n_528), .Y(n_664) );
AOI221xp5_ASAP7_75t_L g668 ( .A1(n_528), .A2(n_669), .B1(n_670), .B2(n_675), .C(n_678), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_528), .B(n_718), .Y(n_717) );
AND2x4_ASAP7_75t_L g528 ( .A(n_529), .B(n_541), .Y(n_528) );
INVx3_ASAP7_75t_L g568 ( .A(n_529), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_529), .B(n_572), .Y(n_672) );
AND2x2_ASAP7_75t_L g701 ( .A(n_529), .B(n_674), .Y(n_701) );
NOR2xp33_ASAP7_75t_L g732 ( .A(n_529), .B(n_733), .Y(n_732) );
AND2x4_ASAP7_75t_L g529 ( .A(n_530), .B(n_535), .Y(n_529) );
AND2x2_ASAP7_75t_L g609 ( .A(n_542), .B(n_584), .Y(n_609) );
AOI21xp5_ASAP7_75t_L g645 ( .A1(n_542), .A2(n_562), .B(n_646), .Y(n_645) );
AND2x2_ASAP7_75t_L g546 ( .A(n_543), .B(n_547), .Y(n_546) );
INVx2_ASAP7_75t_L g555 ( .A(n_543), .Y(n_555) );
OR2x2_ASAP7_75t_L g601 ( .A(n_543), .B(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_SL g693 ( .A(n_543), .B(n_584), .Y(n_693) );
OR2x2_ASAP7_75t_L g725 ( .A(n_543), .B(n_726), .Y(n_725) );
OR2x2_ASAP7_75t_L g737 ( .A(n_543), .B(n_643), .Y(n_737) );
INVxp67_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_546), .B(n_549), .Y(n_545) );
INVx2_ASAP7_75t_L g615 ( .A(n_546), .Y(n_615) );
INVx3_ASAP7_75t_SL g681 ( .A(n_547), .Y(n_681) );
INVxp67_ASAP7_75t_L g631 ( .A(n_549), .Y(n_631) );
AND2x2_ASAP7_75t_L g549 ( .A(n_550), .B(n_551), .Y(n_549) );
AOI322xp5_ASAP7_75t_L g553 ( .A1(n_551), .A2(n_554), .A3(n_558), .B1(n_561), .B2(n_564), .C1(n_569), .C2(n_573), .Y(n_553) );
INVx1_ASAP7_75t_SL g642 ( .A(n_551), .Y(n_642) );
AND2x4_ASAP7_75t_L g727 ( .A(n_551), .B(n_614), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_553), .B(n_575), .Y(n_552) );
NOR2x1_ASAP7_75t_L g554 ( .A(n_555), .B(n_556), .Y(n_554) );
OR2x2_ASAP7_75t_L g580 ( .A(n_555), .B(n_581), .Y(n_580) );
OR2x2_ASAP7_75t_L g676 ( .A(n_555), .B(n_677), .Y(n_676) );
AND2x2_ASAP7_75t_L g704 ( .A(n_555), .B(n_557), .Y(n_704) );
AOI32xp33_ASAP7_75t_L g705 ( .A1(n_555), .A2(n_556), .A3(n_706), .B1(n_708), .B2(n_711), .Y(n_705) );
OR2x2_ASAP7_75t_L g709 ( .A(n_555), .B(n_602), .Y(n_709) );
NAND3xp33_ASAP7_75t_L g665 ( .A(n_556), .B(n_581), .C(n_666), .Y(n_665) );
OAI22xp33_ASAP7_75t_SL g685 ( .A1(n_556), .A2(n_622), .B1(n_686), .B2(n_687), .Y(n_685) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVxp67_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g688 ( .A(n_559), .B(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx1_ASAP7_75t_SL g562 ( .A(n_563), .Y(n_562) );
NOR2xp33_ASAP7_75t_L g724 ( .A(n_563), .B(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_566), .B(n_567), .Y(n_565) );
OAI322xp33_ASAP7_75t_L g611 ( .A1(n_567), .A2(n_571), .A3(n_580), .B1(n_612), .B2(n_615), .C1(n_616), .C2(n_617), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_567), .B(n_620), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_567), .B(n_683), .Y(n_682) );
AND2x2_ASAP7_75t_L g590 ( .A(n_568), .B(n_591), .Y(n_590) );
OR2x2_ASAP7_75t_L g622 ( .A(n_568), .B(n_623), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_568), .B(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx1_ASAP7_75t_L g683 ( .A(n_571), .Y(n_683) );
HB1xp67_ASAP7_75t_L g614 ( .A(n_572), .Y(n_614) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
OAI21xp5_ASAP7_75t_L g575 ( .A1(n_576), .A2(n_579), .B(n_582), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_577), .B(n_578), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_578), .B(n_626), .Y(n_625) );
AOI322xp5_ASAP7_75t_SL g720 ( .A1(n_578), .A2(n_584), .A3(n_701), .B1(n_719), .B2(n_721), .C1(n_724), .C2(n_727), .Y(n_720) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
OAI21xp33_ASAP7_75t_L g583 ( .A1(n_584), .A2(n_585), .B(n_599), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_584), .B(n_594), .Y(n_616) );
INVx2_ASAP7_75t_SL g626 ( .A(n_584), .Y(n_626) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_588), .B(n_590), .Y(n_587) );
INVx1_ASAP7_75t_SL g651 ( .A(n_590), .Y(n_651) );
HB1xp67_ASAP7_75t_L g621 ( .A(n_591), .Y(n_621) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
HB1xp67_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
AND2x2_ASAP7_75t_L g696 ( .A(n_597), .B(n_697), .Y(n_696) );
INVx1_ASAP7_75t_SL g597 ( .A(n_598), .Y(n_597) );
OR2x2_ASAP7_75t_L g650 ( .A(n_598), .B(n_651), .Y(n_650) );
AOI22xp33_ASAP7_75t_L g599 ( .A1(n_600), .A2(n_603), .B1(n_604), .B2(n_609), .Y(n_599) );
INVx1_ASAP7_75t_SL g600 ( .A(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_606), .B(n_607), .Y(n_605) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
NOR4xp75_ASAP7_75t_L g610 ( .A(n_611), .B(n_624), .C(n_644), .D(n_660), .Y(n_610) );
INVx1_ASAP7_75t_SL g612 ( .A(n_613), .Y(n_612) );
INVxp67_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
NAND2xp5_ASAP7_75t_SL g618 ( .A(n_619), .B(n_622), .Y(n_618) );
INVxp67_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
OAI22xp5_ASAP7_75t_L g698 ( .A1(n_622), .A2(n_699), .B1(n_702), .B2(n_703), .Y(n_698) );
OR2x2_ASAP7_75t_L g663 ( .A(n_623), .B(n_664), .Y(n_663) );
INVx2_ASAP7_75t_L g707 ( .A(n_623), .Y(n_707) );
OAI221xp5_ASAP7_75t_L g624 ( .A1(n_625), .A2(n_627), .B1(n_629), .B2(n_631), .C(n_632), .Y(n_624) );
INVx2_ASAP7_75t_L g643 ( .A(n_628), .Y(n_643) );
AND2x2_ASAP7_75t_L g700 ( .A(n_628), .B(n_701), .Y(n_700) );
INVx2_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
AOI22xp5_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_636), .B1(n_638), .B2(n_640), .Y(n_632) );
INVx1_ASAP7_75t_SL g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
BUFx2_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g695 ( .A(n_639), .Y(n_695) );
AOI22xp5_ASAP7_75t_L g661 ( .A1(n_640), .A2(n_646), .B1(n_662), .B2(n_665), .Y(n_661) );
INVx1_ASAP7_75t_SL g640 ( .A(n_641), .Y(n_640) );
OR2x2_ASAP7_75t_L g641 ( .A(n_642), .B(n_643), .Y(n_641) );
OAI221xp5_ASAP7_75t_L g644 ( .A1(n_645), .A2(n_650), .B1(n_652), .B2(n_653), .C(n_776), .Y(n_644) );
AND2x2_ASAP7_75t_SL g646 ( .A(n_647), .B(n_649), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
OR2x2_ASAP7_75t_L g712 ( .A(n_651), .B(n_713), .Y(n_712) );
INVxp67_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
AND2x2_ASAP7_75t_L g654 ( .A(n_655), .B(n_656), .Y(n_654) );
INVx2_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
OR2x2_ASAP7_75t_L g657 ( .A(n_658), .B(n_659), .Y(n_657) );
INVx1_ASAP7_75t_L g697 ( .A(n_659), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_661), .B(n_668), .Y(n_660) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx2_ASAP7_75t_SL g670 ( .A(n_671), .Y(n_670) );
OR2x2_ASAP7_75t_L g671 ( .A(n_672), .B(n_673), .Y(n_671) );
INVx1_ASAP7_75t_SL g675 ( .A(n_676), .Y(n_675) );
AOI21xp33_ASAP7_75t_L g678 ( .A1(n_679), .A2(n_681), .B(n_682), .Y(n_678) );
NOR3xp33_ASAP7_75t_SL g684 ( .A(n_685), .B(n_690), .C(n_714), .Y(n_684) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_691), .B(n_705), .Y(n_690) );
O2A1O1Ixp33_ASAP7_75t_L g691 ( .A1(n_692), .A2(n_694), .B(n_696), .C(n_698), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
AND2x4_ASAP7_75t_L g706 ( .A(n_697), .B(n_707), .Y(n_706) );
INVx1_ASAP7_75t_SL g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_SL g703 ( .A(n_704), .Y(n_703) );
NAND2xp5_ASAP7_75t_SL g708 ( .A(n_709), .B(n_710), .Y(n_708) );
INVx1_ASAP7_75t_SL g711 ( .A(n_712), .Y(n_711) );
NAND4xp25_ASAP7_75t_SL g714 ( .A(n_715), .B(n_720), .C(n_728), .D(n_735), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_716), .B(n_719), .Y(n_715) );
INVx1_ASAP7_75t_SL g716 ( .A(n_717), .Y(n_716) );
INVxp67_ASAP7_75t_SL g721 ( .A(n_722), .Y(n_721) );
OAI21xp5_ASAP7_75t_SL g728 ( .A1(n_729), .A2(n_730), .B(n_732), .Y(n_728) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx3_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
CKINVDCx5p33_ASAP7_75t_R g740 ( .A(n_741), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_743), .B(n_744), .Y(n_742) );
NOR2xp33_ASAP7_75t_L g773 ( .A(n_743), .B(n_744), .Y(n_773) );
CKINVDCx5p33_ASAP7_75t_R g746 ( .A(n_747), .Y(n_746) );
INVx3_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
OAI22xp5_ASAP7_75t_L g749 ( .A1(n_750), .A2(n_754), .B1(n_755), .B2(n_758), .Y(n_749) );
INVx2_ASAP7_75t_L g758 ( .A(n_750), .Y(n_758) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
NOR2x1_ASAP7_75t_R g759 ( .A(n_760), .B(n_762), .Y(n_759) );
INVxp67_ASAP7_75t_SL g760 ( .A(n_761), .Y(n_760) );
BUFx3_ASAP7_75t_L g765 ( .A(n_761), .Y(n_765) );
NOR2xp33_ASAP7_75t_L g763 ( .A(n_764), .B(n_765), .Y(n_763) );
BUFx2_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
CKINVDCx20_ASAP7_75t_R g774 ( .A(n_767), .Y(n_774) );
INVx3_ASAP7_75t_SL g767 ( .A(n_768), .Y(n_767) );
NAND2xp5_ASAP7_75t_SL g768 ( .A(n_769), .B(n_773), .Y(n_768) );
endmodule