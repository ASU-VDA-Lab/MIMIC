module fake_netlist_1_11115_n_657 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_74, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_657);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_74;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_657;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_446;
wire n_342;
wire n_423;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx16_ASAP7_75t_R g75 ( .A(n_14), .Y(n_75) );
CKINVDCx20_ASAP7_75t_R g76 ( .A(n_51), .Y(n_76) );
CKINVDCx20_ASAP7_75t_R g77 ( .A(n_24), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_55), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_32), .Y(n_79) );
BUFx2_ASAP7_75t_L g80 ( .A(n_34), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_53), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_40), .Y(n_82) );
BUFx6f_ASAP7_75t_L g83 ( .A(n_1), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_22), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_2), .Y(n_85) );
INVx2_ASAP7_75t_L g86 ( .A(n_8), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_6), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_8), .Y(n_88) );
CKINVDCx16_ASAP7_75t_R g89 ( .A(n_52), .Y(n_89) );
INVx2_ASAP7_75t_L g90 ( .A(n_0), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_54), .Y(n_91) );
INVx1_ASAP7_75t_SL g92 ( .A(n_31), .Y(n_92) );
BUFx2_ASAP7_75t_L g93 ( .A(n_30), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_6), .Y(n_94) );
BUFx3_ASAP7_75t_L g95 ( .A(n_46), .Y(n_95) );
HB1xp67_ASAP7_75t_L g96 ( .A(n_35), .Y(n_96) );
INVxp33_ASAP7_75t_SL g97 ( .A(n_20), .Y(n_97) );
CKINVDCx16_ASAP7_75t_R g98 ( .A(n_44), .Y(n_98) );
INVx3_ASAP7_75t_L g99 ( .A(n_71), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_25), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_26), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_36), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_49), .Y(n_103) );
INVx2_ASAP7_75t_SL g104 ( .A(n_50), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_74), .Y(n_105) );
INVx2_ASAP7_75t_L g106 ( .A(n_73), .Y(n_106) );
INVx2_ASAP7_75t_L g107 ( .A(n_10), .Y(n_107) );
INVx1_ASAP7_75t_SL g108 ( .A(n_10), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_5), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_60), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_47), .Y(n_111) );
BUFx2_ASAP7_75t_L g112 ( .A(n_57), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_15), .Y(n_113) );
HB1xp67_ASAP7_75t_L g114 ( .A(n_14), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_56), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_23), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_70), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_59), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_68), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_43), .Y(n_120) );
AND2x4_ASAP7_75t_L g121 ( .A(n_80), .B(n_0), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_78), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_99), .Y(n_123) );
BUFx6f_ASAP7_75t_L g124 ( .A(n_99), .Y(n_124) );
BUFx6f_ASAP7_75t_L g125 ( .A(n_99), .Y(n_125) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_95), .Y(n_126) );
AOI22xp5_ASAP7_75t_L g127 ( .A1(n_75), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_127) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_95), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_106), .Y(n_129) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_83), .Y(n_130) );
OA21x2_ASAP7_75t_L g131 ( .A1(n_78), .A2(n_33), .B(n_69), .Y(n_131) );
OAI21x1_ASAP7_75t_L g132 ( .A1(n_106), .A2(n_29), .B(n_67), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_79), .Y(n_133) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_83), .Y(n_134) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_83), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_80), .B(n_3), .Y(n_136) );
INVx3_ASAP7_75t_L g137 ( .A(n_83), .Y(n_137) );
AND2x2_ASAP7_75t_L g138 ( .A(n_93), .B(n_4), .Y(n_138) );
INVx3_ASAP7_75t_L g139 ( .A(n_83), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_79), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_81), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_81), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_104), .Y(n_143) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_104), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_82), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_82), .Y(n_146) );
AOI22xp5_ASAP7_75t_L g147 ( .A1(n_114), .A2(n_4), .B1(n_5), .B2(n_7), .Y(n_147) );
AOI22x1_ASAP7_75t_SL g148 ( .A1(n_76), .A2(n_7), .B1(n_9), .B2(n_11), .Y(n_148) );
AND2x6_ASAP7_75t_L g149 ( .A(n_84), .B(n_38), .Y(n_149) );
HB1xp67_ASAP7_75t_L g150 ( .A(n_85), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_84), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_91), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_91), .Y(n_153) );
AND2x4_ASAP7_75t_L g154 ( .A(n_93), .B(n_9), .Y(n_154) );
AND2x2_ASAP7_75t_SL g155 ( .A(n_112), .B(n_72), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_101), .Y(n_156) );
AND2x4_ASAP7_75t_L g157 ( .A(n_112), .B(n_11), .Y(n_157) );
AND2x2_ASAP7_75t_L g158 ( .A(n_89), .B(n_12), .Y(n_158) );
AOI22xp5_ASAP7_75t_SL g159 ( .A1(n_77), .A2(n_12), .B1(n_13), .B2(n_15), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_101), .Y(n_160) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_102), .Y(n_161) );
OAI22xp5_ASAP7_75t_L g162 ( .A1(n_85), .A2(n_13), .B1(n_16), .B2(n_17), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_124), .Y(n_163) );
INVx3_ASAP7_75t_L g164 ( .A(n_144), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_143), .B(n_98), .Y(n_165) );
NAND2xp33_ASAP7_75t_L g166 ( .A(n_149), .B(n_96), .Y(n_166) );
OR2x6_ASAP7_75t_L g167 ( .A(n_121), .B(n_88), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_143), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_124), .Y(n_169) );
AND2x2_ASAP7_75t_L g170 ( .A(n_138), .B(n_86), .Y(n_170) );
CKINVDCx5p33_ASAP7_75t_R g171 ( .A(n_158), .Y(n_171) );
INVx2_ASAP7_75t_SL g172 ( .A(n_121), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_124), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_124), .Y(n_174) );
AND2x6_ASAP7_75t_L g175 ( .A(n_121), .B(n_105), .Y(n_175) );
BUFx6f_ASAP7_75t_SL g176 ( .A(n_155), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_124), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_123), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_122), .B(n_103), .Y(n_179) );
INVx1_ASAP7_75t_SL g180 ( .A(n_158), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_123), .Y(n_181) );
AOI22xp5_ASAP7_75t_L g182 ( .A1(n_155), .A2(n_87), .B1(n_113), .B2(n_109), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_122), .B(n_115), .Y(n_183) );
NAND3xp33_ASAP7_75t_L g184 ( .A(n_150), .B(n_87), .C(n_88), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_133), .B(n_110), .Y(n_185) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_133), .B(n_105), .Y(n_186) );
NAND2xp5_ASAP7_75t_SL g187 ( .A(n_141), .B(n_116), .Y(n_187) );
INVx2_ASAP7_75t_SL g188 ( .A(n_121), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_140), .Y(n_189) );
INVx5_ASAP7_75t_L g190 ( .A(n_149), .Y(n_190) );
NAND2xp5_ASAP7_75t_SL g191 ( .A(n_141), .B(n_116), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_145), .B(n_97), .Y(n_192) );
NOR2x1p5_ASAP7_75t_L g193 ( .A(n_136), .B(n_109), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_125), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_125), .Y(n_195) );
BUFx3_ASAP7_75t_L g196 ( .A(n_144), .Y(n_196) );
BUFx6f_ASAP7_75t_L g197 ( .A(n_132), .Y(n_197) );
INVx1_ASAP7_75t_SL g198 ( .A(n_138), .Y(n_198) );
OR2x2_ASAP7_75t_L g199 ( .A(n_154), .B(n_108), .Y(n_199) );
INVx2_ASAP7_75t_L g200 ( .A(n_125), .Y(n_200) );
BUFx10_ASAP7_75t_L g201 ( .A(n_154), .Y(n_201) );
INVx5_ASAP7_75t_L g202 ( .A(n_149), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_140), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_145), .B(n_117), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_125), .Y(n_205) );
AOI22xp33_ASAP7_75t_L g206 ( .A1(n_154), .A2(n_94), .B1(n_113), .B2(n_86), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_152), .B(n_100), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_152), .B(n_119), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_140), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_142), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_142), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_142), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g213 ( .A(n_153), .B(n_119), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_146), .Y(n_214) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_153), .B(n_102), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g216 ( .A(n_165), .B(n_154), .Y(n_216) );
AOI22xp33_ASAP7_75t_SL g217 ( .A1(n_176), .A2(n_155), .B1(n_159), .B2(n_148), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_168), .Y(n_218) );
INVx3_ASAP7_75t_L g219 ( .A(n_201), .Y(n_219) );
NAND2xp33_ASAP7_75t_L g220 ( .A(n_175), .B(n_149), .Y(n_220) );
A2O1A1Ixp33_ASAP7_75t_L g221 ( .A1(n_213), .A2(n_157), .B(n_156), .C(n_160), .Y(n_221) );
AOI22xp5_ASAP7_75t_L g222 ( .A1(n_182), .A2(n_157), .B1(n_127), .B2(n_120), .Y(n_222) );
AOI22xp33_ASAP7_75t_L g223 ( .A1(n_176), .A2(n_156), .B1(n_160), .B2(n_149), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_192), .B(n_157), .Y(n_224) );
INVx8_ASAP7_75t_L g225 ( .A(n_167), .Y(n_225) );
INVx2_ASAP7_75t_SL g226 ( .A(n_167), .Y(n_226) );
AOI22xp5_ASAP7_75t_L g227 ( .A1(n_176), .A2(n_157), .B1(n_127), .B2(n_147), .Y(n_227) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_190), .B(n_144), .Y(n_228) );
BUFx3_ASAP7_75t_L g229 ( .A(n_175), .Y(n_229) );
AND2x4_ASAP7_75t_L g230 ( .A(n_167), .B(n_147), .Y(n_230) );
CKINVDCx5p33_ASAP7_75t_R g231 ( .A(n_171), .Y(n_231) );
NAND2xp5_ASAP7_75t_SL g232 ( .A(n_201), .B(n_144), .Y(n_232) );
NOR2x2_ASAP7_75t_L g233 ( .A(n_167), .B(n_148), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_198), .B(n_146), .Y(n_234) );
CKINVDCx5p33_ASAP7_75t_R g235 ( .A(n_171), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_170), .B(n_151), .Y(n_236) );
INVx1_ASAP7_75t_SL g237 ( .A(n_180), .Y(n_237) );
A2O1A1Ixp33_ASAP7_75t_L g238 ( .A1(n_172), .A2(n_151), .B(n_129), .C(n_132), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_170), .B(n_149), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_178), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_179), .B(n_149), .Y(n_241) );
BUFx4f_ASAP7_75t_L g242 ( .A(n_175), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_183), .B(n_144), .Y(n_243) );
NAND2xp5_ASAP7_75t_SL g244 ( .A(n_201), .B(n_92), .Y(n_244) );
NAND2xp5_ASAP7_75t_SL g245 ( .A(n_190), .B(n_125), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_185), .B(n_129), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_204), .B(n_129), .Y(n_247) );
BUFx2_ASAP7_75t_L g248 ( .A(n_175), .Y(n_248) );
INVx2_ASAP7_75t_L g249 ( .A(n_189), .Y(n_249) );
NOR2xp33_ASAP7_75t_L g250 ( .A(n_199), .B(n_111), .Y(n_250) );
NOR2xp33_ASAP7_75t_SL g251 ( .A(n_190), .B(n_162), .Y(n_251) );
AND2x2_ASAP7_75t_SL g252 ( .A(n_166), .B(n_131), .Y(n_252) );
NAND2x1p5_ASAP7_75t_L g253 ( .A(n_199), .B(n_94), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_203), .Y(n_254) );
AOI22xp33_ASAP7_75t_L g255 ( .A1(n_175), .A2(n_161), .B1(n_90), .B2(n_107), .Y(n_255) );
INVxp67_ASAP7_75t_SL g256 ( .A(n_172), .Y(n_256) );
AO22x1_ASAP7_75t_L g257 ( .A1(n_175), .A2(n_159), .B1(n_111), .B2(n_118), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_209), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_206), .B(n_118), .Y(n_259) );
NAND2xp33_ASAP7_75t_L g260 ( .A(n_190), .B(n_202), .Y(n_260) );
AOI21xp5_ASAP7_75t_L g261 ( .A1(n_166), .A2(n_131), .B(n_126), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_181), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_193), .B(n_161), .Y(n_263) );
INVx2_ASAP7_75t_SL g264 ( .A(n_188), .Y(n_264) );
INVx3_ASAP7_75t_L g265 ( .A(n_188), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_207), .B(n_161), .Y(n_266) );
NAND2xp5_ASAP7_75t_SL g267 ( .A(n_190), .B(n_161), .Y(n_267) );
AOI22xp33_ASAP7_75t_L g268 ( .A1(n_214), .A2(n_161), .B1(n_90), .B2(n_107), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_208), .B(n_126), .Y(n_269) );
OAI22xp5_ASAP7_75t_L g270 ( .A1(n_184), .A2(n_126), .B1(n_128), .B2(n_139), .Y(n_270) );
AOI22xp5_ASAP7_75t_L g271 ( .A1(n_186), .A2(n_126), .B1(n_128), .B2(n_131), .Y(n_271) );
NAND2xp5_ASAP7_75t_SL g272 ( .A(n_202), .B(n_126), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_210), .B(n_128), .Y(n_273) );
NAND2xp5_ASAP7_75t_SL g274 ( .A(n_202), .B(n_128), .Y(n_274) );
OAI22xp5_ASAP7_75t_L g275 ( .A1(n_227), .A2(n_212), .B1(n_211), .B2(n_187), .Y(n_275) );
BUFx6f_ASAP7_75t_L g276 ( .A(n_225), .Y(n_276) );
AOI21xp5_ASAP7_75t_L g277 ( .A1(n_241), .A2(n_202), .B(n_197), .Y(n_277) );
AOI21xp5_ASAP7_75t_L g278 ( .A1(n_220), .A2(n_202), .B(n_197), .Y(n_278) );
O2A1O1Ixp5_ASAP7_75t_L g279 ( .A1(n_261), .A2(n_215), .B(n_186), .C(n_187), .Y(n_279) );
BUFx2_ASAP7_75t_L g280 ( .A(n_237), .Y(n_280) );
OAI22xp5_ASAP7_75t_SL g281 ( .A1(n_217), .A2(n_131), .B1(n_197), .B2(n_16), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_253), .B(n_215), .Y(n_282) );
NOR2xp33_ASAP7_75t_L g283 ( .A(n_253), .B(n_191), .Y(n_283) );
AOI21xp5_ASAP7_75t_L g284 ( .A1(n_239), .A2(n_197), .B(n_191), .Y(n_284) );
NAND2xp5_ASAP7_75t_SL g285 ( .A(n_226), .B(n_197), .Y(n_285) );
CKINVDCx11_ASAP7_75t_R g286 ( .A(n_225), .Y(n_286) );
AOI22xp5_ASAP7_75t_L g287 ( .A1(n_225), .A2(n_164), .B1(n_196), .B2(n_128), .Y(n_287) );
INVx4_ASAP7_75t_L g288 ( .A(n_242), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_216), .B(n_164), .Y(n_289) );
NAND3xp33_ASAP7_75t_SL g290 ( .A(n_231), .B(n_205), .C(n_200), .Y(n_290) );
O2A1O1Ixp33_ASAP7_75t_L g291 ( .A1(n_221), .A2(n_164), .B(n_139), .C(n_137), .Y(n_291) );
BUFx2_ASAP7_75t_SL g292 ( .A(n_229), .Y(n_292) );
NAND2xp5_ASAP7_75t_SL g293 ( .A(n_242), .B(n_196), .Y(n_293) );
AOI21xp5_ASAP7_75t_L g294 ( .A1(n_238), .A2(n_205), .B(n_200), .Y(n_294) );
BUFx8_ASAP7_75t_L g295 ( .A(n_230), .Y(n_295) );
NOR2xp33_ASAP7_75t_R g296 ( .A(n_235), .B(n_18), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_236), .Y(n_297) );
AND2x2_ASAP7_75t_L g298 ( .A(n_230), .B(n_137), .Y(n_298) );
AND2x2_ASAP7_75t_L g299 ( .A(n_222), .B(n_137), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_216), .B(n_195), .Y(n_300) );
NAND2x1p5_ASAP7_75t_L g301 ( .A(n_229), .B(n_163), .Y(n_301) );
AOI21xp5_ASAP7_75t_L g302 ( .A1(n_260), .A2(n_163), .B(n_194), .Y(n_302) );
BUFx6f_ASAP7_75t_L g303 ( .A(n_248), .Y(n_303) );
NAND2xp5_ASAP7_75t_SL g304 ( .A(n_219), .B(n_195), .Y(n_304) );
INVx2_ASAP7_75t_SL g305 ( .A(n_234), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_250), .B(n_194), .Y(n_306) );
CKINVDCx20_ASAP7_75t_R g307 ( .A(n_250), .Y(n_307) );
O2A1O1Ixp33_ASAP7_75t_L g308 ( .A1(n_259), .A2(n_139), .B(n_137), .C(n_173), .Y(n_308) );
NOR2xp33_ASAP7_75t_L g309 ( .A(n_224), .B(n_177), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_218), .B(n_177), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_249), .B(n_174), .Y(n_311) );
BUFx6f_ASAP7_75t_L g312 ( .A(n_219), .Y(n_312) );
OAI21xp33_ASAP7_75t_SL g313 ( .A1(n_223), .A2(n_174), .B(n_173), .Y(n_313) );
OAI22xp5_ASAP7_75t_L g314 ( .A1(n_223), .A2(n_139), .B1(n_169), .B2(n_135), .Y(n_314) );
BUFx6f_ASAP7_75t_L g315 ( .A(n_249), .Y(n_315) );
NOR3xp33_ASAP7_75t_SL g316 ( .A(n_233), .B(n_19), .C(n_21), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_254), .B(n_169), .Y(n_317) );
OAI21xp33_ASAP7_75t_SL g318 ( .A1(n_252), .A2(n_27), .B(n_28), .Y(n_318) );
NAND2xp5_ASAP7_75t_SL g319 ( .A(n_265), .B(n_135), .Y(n_319) );
BUFx12f_ASAP7_75t_L g320 ( .A(n_264), .Y(n_320) );
INVx3_ASAP7_75t_L g321 ( .A(n_254), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_258), .B(n_135), .Y(n_322) );
OAI21x1_ASAP7_75t_L g323 ( .A1(n_271), .A2(n_37), .B(n_39), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_321), .Y(n_324) );
AO31x2_ASAP7_75t_L g325 ( .A1(n_275), .A2(n_269), .A3(n_246), .B(n_247), .Y(n_325) );
A2O1A1Ixp33_ASAP7_75t_L g326 ( .A1(n_318), .A2(n_258), .B(n_266), .C(n_243), .Y(n_326) );
A2O1A1Ixp33_ASAP7_75t_L g327 ( .A1(n_291), .A2(n_240), .B(n_262), .C(n_252), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_321), .Y(n_328) );
OAI22xp5_ASAP7_75t_L g329 ( .A1(n_307), .A2(n_255), .B1(n_256), .B2(n_265), .Y(n_329) );
AOI221xp5_ASAP7_75t_L g330 ( .A1(n_275), .A2(n_257), .B1(n_251), .B2(n_263), .C(n_244), .Y(n_330) );
AO31x2_ASAP7_75t_L g331 ( .A1(n_314), .A2(n_273), .A3(n_270), .B(n_268), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_297), .Y(n_332) );
BUFx2_ASAP7_75t_SL g333 ( .A(n_276), .Y(n_333) );
A2O1A1Ixp33_ASAP7_75t_L g334 ( .A1(n_309), .A2(n_268), .B(n_255), .C(n_232), .Y(n_334) );
OAI21x1_ASAP7_75t_L g335 ( .A1(n_294), .A2(n_274), .B(n_272), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_305), .B(n_245), .Y(n_336) );
NAND3xp33_ASAP7_75t_L g337 ( .A(n_313), .B(n_314), .C(n_308), .Y(n_337) );
AOI21xp5_ASAP7_75t_L g338 ( .A1(n_277), .A2(n_245), .B(n_228), .Y(n_338) );
O2A1O1Ixp33_ASAP7_75t_SL g339 ( .A1(n_285), .A2(n_228), .B(n_272), .C(n_274), .Y(n_339) );
BUFx6f_ASAP7_75t_L g340 ( .A(n_276), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_299), .B(n_267), .Y(n_341) );
INVx3_ASAP7_75t_SL g342 ( .A(n_276), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_315), .Y(n_343) );
AOI21xp5_ASAP7_75t_L g344 ( .A1(n_284), .A2(n_135), .B(n_134), .Y(n_344) );
AO31x2_ASAP7_75t_L g345 ( .A1(n_278), .A2(n_135), .A3(n_134), .B(n_130), .Y(n_345) );
BUFx10_ASAP7_75t_L g346 ( .A(n_283), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_280), .B(n_134), .Y(n_347) );
OAI22xp5_ASAP7_75t_L g348 ( .A1(n_282), .A2(n_130), .B1(n_134), .B2(n_45), .Y(n_348) );
A2O1A1Ixp33_ASAP7_75t_L g349 ( .A1(n_279), .A2(n_134), .B(n_130), .C(n_48), .Y(n_349) );
BUFx6f_ASAP7_75t_SL g350 ( .A(n_286), .Y(n_350) );
OA21x2_ASAP7_75t_L g351 ( .A1(n_323), .A2(n_130), .B(n_42), .Y(n_351) );
AOI21xp5_ASAP7_75t_L g352 ( .A1(n_300), .A2(n_130), .B(n_58), .Y(n_352) );
CKINVDCx20_ASAP7_75t_R g353 ( .A(n_295), .Y(n_353) );
OA21x2_ASAP7_75t_L g354 ( .A1(n_322), .A2(n_41), .B(n_61), .Y(n_354) );
NOR2xp33_ASAP7_75t_L g355 ( .A(n_332), .B(n_295), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_346), .B(n_298), .Y(n_356) );
INVxp67_ASAP7_75t_L g357 ( .A(n_350), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_346), .B(n_316), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_342), .B(n_315), .Y(n_359) );
NAND2x1p5_ASAP7_75t_L g360 ( .A(n_340), .B(n_312), .Y(n_360) );
AOI221xp5_ASAP7_75t_L g361 ( .A1(n_330), .A2(n_281), .B1(n_289), .B2(n_306), .C(n_296), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_347), .Y(n_362) );
OAI221xp5_ASAP7_75t_L g363 ( .A1(n_326), .A2(n_289), .B1(n_287), .B2(n_310), .C(n_288), .Y(n_363) );
AOI21xp5_ASAP7_75t_L g364 ( .A1(n_326), .A2(n_290), .B(n_304), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_336), .Y(n_365) );
OAI221xp5_ASAP7_75t_L g366 ( .A1(n_327), .A2(n_288), .B1(n_315), .B2(n_317), .C(n_311), .Y(n_366) );
AOI22xp5_ASAP7_75t_L g367 ( .A1(n_329), .A2(n_320), .B1(n_312), .B2(n_292), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_341), .Y(n_368) );
INVx4_ASAP7_75t_L g369 ( .A(n_340), .Y(n_369) );
OAI21x1_ASAP7_75t_SL g370 ( .A1(n_354), .A2(n_302), .B(n_312), .Y(n_370) );
AOI22xp33_ASAP7_75t_L g371 ( .A1(n_337), .A2(n_303), .B1(n_293), .B2(n_301), .Y(n_371) );
OAI21x1_ASAP7_75t_L g372 ( .A1(n_351), .A2(n_301), .B(n_319), .Y(n_372) );
AOI21xp5_ASAP7_75t_L g373 ( .A1(n_344), .A2(n_303), .B(n_63), .Y(n_373) );
AOI221xp5_ASAP7_75t_L g374 ( .A1(n_327), .A2(n_303), .B1(n_64), .B2(n_65), .C(n_66), .Y(n_374) );
OAI21x1_ASAP7_75t_L g375 ( .A1(n_351), .A2(n_62), .B(n_352), .Y(n_375) );
OA21x2_ASAP7_75t_L g376 ( .A1(n_349), .A2(n_335), .B(n_338), .Y(n_376) );
AND2x2_ASAP7_75t_L g377 ( .A(n_325), .B(n_342), .Y(n_377) );
HB1xp67_ASAP7_75t_L g378 ( .A(n_340), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_324), .Y(n_379) );
AOI21xp5_ASAP7_75t_L g380 ( .A1(n_349), .A2(n_339), .B(n_334), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_328), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_376), .Y(n_382) );
OA21x2_ASAP7_75t_L g383 ( .A1(n_380), .A2(n_348), .B(n_334), .Y(n_383) );
OA21x2_ASAP7_75t_L g384 ( .A1(n_370), .A2(n_343), .B(n_325), .Y(n_384) );
OA21x2_ASAP7_75t_L g385 ( .A1(n_370), .A2(n_325), .B(n_345), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_377), .B(n_325), .Y(n_386) );
AO21x2_ASAP7_75t_L g387 ( .A1(n_364), .A2(n_339), .B(n_354), .Y(n_387) );
OAI21xp5_ASAP7_75t_L g388 ( .A1(n_361), .A2(n_354), .B(n_331), .Y(n_388) );
BUFx2_ASAP7_75t_L g389 ( .A(n_377), .Y(n_389) );
BUFx2_ASAP7_75t_L g390 ( .A(n_369), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_368), .B(n_340), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_365), .B(n_331), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_362), .B(n_331), .Y(n_393) );
HB1xp67_ASAP7_75t_L g394 ( .A(n_378), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_369), .B(n_331), .Y(n_395) );
OR2x6_ASAP7_75t_L g396 ( .A(n_369), .B(n_333), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_381), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_379), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_376), .Y(n_399) );
BUFx2_ASAP7_75t_L g400 ( .A(n_360), .Y(n_400) );
OAI22xp5_ASAP7_75t_L g401 ( .A1(n_367), .A2(n_353), .B1(n_350), .B2(n_345), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_376), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_375), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_360), .Y(n_404) );
INVx1_ASAP7_75t_SL g405 ( .A(n_359), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_375), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_372), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_372), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_366), .Y(n_409) );
OR2x6_ASAP7_75t_L g410 ( .A(n_373), .B(n_345), .Y(n_410) );
BUFx3_ASAP7_75t_L g411 ( .A(n_356), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_371), .B(n_345), .Y(n_412) );
INVx3_ASAP7_75t_L g413 ( .A(n_358), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_363), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_393), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_382), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_393), .B(n_371), .Y(n_417) );
NOR2xp33_ASAP7_75t_L g418 ( .A(n_411), .B(n_355), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_393), .B(n_374), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_392), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_386), .B(n_355), .Y(n_421) );
OR2x2_ASAP7_75t_L g422 ( .A(n_389), .B(n_357), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_382), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_386), .B(n_389), .Y(n_424) );
NOR2xp33_ASAP7_75t_L g425 ( .A(n_411), .B(n_413), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_386), .B(n_395), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_395), .B(n_392), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_395), .Y(n_428) );
NOR3xp33_ASAP7_75t_L g429 ( .A(n_401), .B(n_413), .C(n_414), .Y(n_429) );
OR2x2_ASAP7_75t_L g430 ( .A(n_405), .B(n_394), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_397), .B(n_398), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_397), .B(n_398), .Y(n_432) );
INVx4_ASAP7_75t_L g433 ( .A(n_396), .Y(n_433) );
OR2x6_ASAP7_75t_L g434 ( .A(n_396), .B(n_401), .Y(n_434) );
BUFx3_ASAP7_75t_L g435 ( .A(n_390), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_384), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_382), .Y(n_437) );
HB1xp67_ASAP7_75t_L g438 ( .A(n_405), .Y(n_438) );
AND2x4_ASAP7_75t_L g439 ( .A(n_412), .B(n_402), .Y(n_439) );
AOI211xp5_ASAP7_75t_L g440 ( .A1(n_411), .A2(n_413), .B(n_414), .C(n_388), .Y(n_440) );
HB1xp67_ASAP7_75t_L g441 ( .A(n_394), .Y(n_441) );
INVxp67_ASAP7_75t_L g442 ( .A(n_390), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_391), .B(n_413), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_384), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_391), .B(n_412), .Y(n_445) );
AND2x4_ASAP7_75t_L g446 ( .A(n_412), .B(n_402), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_391), .B(n_388), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_399), .Y(n_448) );
HB1xp67_ASAP7_75t_L g449 ( .A(n_396), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_413), .B(n_385), .Y(n_450) );
OR2x2_ASAP7_75t_L g451 ( .A(n_385), .B(n_404), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_384), .Y(n_452) );
HB1xp67_ASAP7_75t_L g453 ( .A(n_396), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_384), .Y(n_454) );
BUFx3_ASAP7_75t_L g455 ( .A(n_396), .Y(n_455) );
BUFx3_ASAP7_75t_L g456 ( .A(n_396), .Y(n_456) );
AOI21xp33_ASAP7_75t_SL g457 ( .A1(n_404), .A2(n_385), .B(n_400), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_409), .B(n_400), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_385), .B(n_384), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_385), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_426), .B(n_399), .Y(n_461) );
NAND4xp25_ASAP7_75t_L g462 ( .A(n_429), .B(n_409), .C(n_399), .D(n_407), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_431), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_431), .B(n_409), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_432), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_426), .B(n_407), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_432), .Y(n_467) );
OR2x2_ASAP7_75t_L g468 ( .A(n_428), .B(n_408), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_427), .B(n_408), .Y(n_469) );
AND2x4_ASAP7_75t_L g470 ( .A(n_434), .B(n_410), .Y(n_470) );
INVx3_ASAP7_75t_L g471 ( .A(n_433), .Y(n_471) );
AOI22xp33_ASAP7_75t_L g472 ( .A1(n_429), .A2(n_383), .B1(n_410), .B2(n_387), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_427), .B(n_408), .Y(n_473) );
INVxp67_ASAP7_75t_L g474 ( .A(n_438), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_416), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_420), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_445), .B(n_387), .Y(n_477) );
INVx2_ASAP7_75t_L g478 ( .A(n_416), .Y(n_478) );
NOR2xp33_ASAP7_75t_R g479 ( .A(n_435), .B(n_403), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_445), .B(n_387), .Y(n_480) );
AOI22xp33_ASAP7_75t_L g481 ( .A1(n_434), .A2(n_383), .B1(n_410), .B2(n_387), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_428), .B(n_403), .Y(n_482) );
OR2x2_ASAP7_75t_L g483 ( .A(n_424), .B(n_403), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_424), .B(n_406), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_415), .B(n_406), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_420), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_415), .B(n_406), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_436), .Y(n_488) );
OR2x2_ASAP7_75t_L g489 ( .A(n_430), .B(n_410), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_447), .B(n_410), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_447), .B(n_410), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_421), .B(n_383), .Y(n_492) );
BUFx2_ASAP7_75t_SL g493 ( .A(n_433), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_439), .B(n_383), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_439), .B(n_383), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_416), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_421), .B(n_441), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_436), .Y(n_498) );
OR2x2_ASAP7_75t_L g499 ( .A(n_430), .B(n_417), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_439), .B(n_446), .Y(n_500) );
OR2x2_ASAP7_75t_L g501 ( .A(n_417), .B(n_443), .Y(n_501) );
BUFx2_ASAP7_75t_L g502 ( .A(n_435), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_444), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_439), .B(n_446), .Y(n_504) );
OR2x2_ASAP7_75t_L g505 ( .A(n_443), .B(n_446), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_444), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_452), .Y(n_507) );
HB1xp67_ASAP7_75t_L g508 ( .A(n_435), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_452), .Y(n_509) );
INVx2_ASAP7_75t_L g510 ( .A(n_423), .Y(n_510) );
NAND2x1p5_ASAP7_75t_L g511 ( .A(n_433), .B(n_456), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_446), .B(n_450), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_454), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_422), .B(n_418), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_422), .B(n_425), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_463), .Y(n_516) );
NAND2x1p5_ASAP7_75t_L g517 ( .A(n_502), .B(n_433), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_500), .B(n_434), .Y(n_518) );
OR2x2_ASAP7_75t_L g519 ( .A(n_497), .B(n_451), .Y(n_519) );
INVx2_ASAP7_75t_L g520 ( .A(n_475), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_463), .B(n_442), .Y(n_521) );
OAI21xp33_ASAP7_75t_L g522 ( .A1(n_490), .A2(n_440), .B(n_434), .Y(n_522) );
NOR2xp67_ASAP7_75t_L g523 ( .A(n_462), .B(n_457), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_465), .B(n_442), .Y(n_524) );
NAND3xp33_ASAP7_75t_L g525 ( .A(n_474), .B(n_457), .C(n_440), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_512), .B(n_450), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_465), .Y(n_527) );
INVxp67_ASAP7_75t_SL g528 ( .A(n_475), .Y(n_528) );
NAND2x1p5_ASAP7_75t_L g529 ( .A(n_502), .B(n_456), .Y(n_529) );
AND2x4_ASAP7_75t_SL g530 ( .A(n_508), .B(n_434), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_512), .B(n_459), .Y(n_531) );
INVx2_ASAP7_75t_L g532 ( .A(n_478), .Y(n_532) );
OR2x2_ASAP7_75t_L g533 ( .A(n_499), .B(n_451), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_467), .B(n_458), .Y(n_534) );
OR2x2_ASAP7_75t_L g535 ( .A(n_499), .B(n_458), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_500), .B(n_453), .Y(n_536) );
AND2x4_ASAP7_75t_L g537 ( .A(n_470), .B(n_456), .Y(n_537) );
HB1xp67_ASAP7_75t_L g538 ( .A(n_478), .Y(n_538) );
OR2x2_ASAP7_75t_L g539 ( .A(n_501), .B(n_449), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_494), .B(n_459), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_494), .B(n_454), .Y(n_541) );
INVx2_ASAP7_75t_L g542 ( .A(n_496), .Y(n_542) );
NAND2x1_ASAP7_75t_SL g543 ( .A(n_471), .B(n_460), .Y(n_543) );
NAND3xp33_ASAP7_75t_L g544 ( .A(n_472), .B(n_481), .C(n_489), .Y(n_544) );
NOR2xp67_ASAP7_75t_L g545 ( .A(n_471), .B(n_460), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_467), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_501), .B(n_419), .Y(n_547) );
OR2x2_ASAP7_75t_L g548 ( .A(n_505), .B(n_423), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_476), .Y(n_549) );
INVx2_ASAP7_75t_L g550 ( .A(n_496), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_504), .B(n_455), .Y(n_551) );
NAND2xp5_ASAP7_75t_SL g552 ( .A(n_479), .B(n_455), .Y(n_552) );
OR2x2_ASAP7_75t_L g553 ( .A(n_505), .B(n_423), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_476), .Y(n_554) );
INVxp67_ASAP7_75t_L g555 ( .A(n_514), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_495), .B(n_437), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_486), .B(n_419), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_486), .B(n_437), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_488), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_495), .B(n_437), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_466), .B(n_448), .Y(n_561) );
NAND3xp33_ASAP7_75t_L g562 ( .A(n_489), .B(n_455), .C(n_448), .Y(n_562) );
NOR2xp33_ASAP7_75t_L g563 ( .A(n_515), .B(n_448), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_466), .B(n_464), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_461), .B(n_480), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_547), .B(n_480), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_539), .Y(n_567) );
OR2x2_ASAP7_75t_L g568 ( .A(n_533), .B(n_461), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_531), .B(n_504), .Y(n_569) );
OR2x2_ASAP7_75t_L g570 ( .A(n_519), .B(n_483), .Y(n_570) );
INVx2_ASAP7_75t_SL g571 ( .A(n_543), .Y(n_571) );
INVx2_ASAP7_75t_L g572 ( .A(n_520), .Y(n_572) );
OR2x2_ASAP7_75t_L g573 ( .A(n_565), .B(n_483), .Y(n_573) );
NOR3xp33_ASAP7_75t_L g574 ( .A(n_525), .B(n_471), .C(n_509), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_555), .B(n_477), .Y(n_575) );
OR2x2_ASAP7_75t_L g576 ( .A(n_565), .B(n_469), .Y(n_576) );
OAI332xp33_ASAP7_75t_L g577 ( .A1(n_557), .A2(n_492), .A3(n_509), .B1(n_507), .B2(n_506), .B3(n_503), .C1(n_498), .C2(n_513), .Y(n_577) );
AOI22xp5_ASAP7_75t_L g578 ( .A1(n_522), .A2(n_490), .B1(n_491), .B2(n_470), .Y(n_578) );
AND2x4_ASAP7_75t_L g579 ( .A(n_545), .B(n_470), .Y(n_579) );
INVx2_ASAP7_75t_L g580 ( .A(n_520), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_516), .Y(n_581) );
INVx2_ASAP7_75t_L g582 ( .A(n_532), .Y(n_582) );
OAI22xp5_ASAP7_75t_L g583 ( .A1(n_517), .A2(n_493), .B1(n_511), .B2(n_470), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_563), .B(n_477), .Y(n_584) );
AOI22xp5_ASAP7_75t_L g585 ( .A1(n_544), .A2(n_491), .B1(n_493), .B2(n_473), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_563), .B(n_473), .Y(n_586) );
OR2x2_ASAP7_75t_L g587 ( .A(n_564), .B(n_469), .Y(n_587) );
INVx1_ASAP7_75t_SL g588 ( .A(n_548), .Y(n_588) );
AOI31xp33_ASAP7_75t_SL g589 ( .A1(n_535), .A2(n_468), .A3(n_511), .B(n_510), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_527), .B(n_498), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_531), .B(n_484), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_526), .B(n_484), .Y(n_592) );
AND2x2_ASAP7_75t_L g593 ( .A(n_526), .B(n_482), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_546), .Y(n_594) );
OAI21xp5_ASAP7_75t_L g595 ( .A1(n_523), .A2(n_511), .B(n_513), .Y(n_595) );
AND2x2_ASAP7_75t_L g596 ( .A(n_540), .B(n_482), .Y(n_596) );
NOR2xp33_ASAP7_75t_L g597 ( .A(n_540), .B(n_503), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_541), .B(n_488), .Y(n_598) );
OR2x2_ASAP7_75t_L g599 ( .A(n_553), .B(n_561), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_559), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_577), .B(n_541), .Y(n_601) );
BUFx2_ASAP7_75t_L g602 ( .A(n_579), .Y(n_602) );
NAND2xp5_ASAP7_75t_SL g603 ( .A(n_574), .B(n_552), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_597), .B(n_556), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_597), .B(n_556), .Y(n_605) );
AOI222xp33_ASAP7_75t_L g606 ( .A1(n_595), .A2(n_521), .B1(n_524), .B2(n_534), .C1(n_530), .C2(n_518), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_566), .B(n_560), .Y(n_607) );
OAI21xp33_ASAP7_75t_L g608 ( .A1(n_585), .A2(n_530), .B(n_536), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_598), .Y(n_609) );
AOI221xp5_ASAP7_75t_L g610 ( .A1(n_574), .A2(n_554), .B1(n_549), .B2(n_562), .C(n_537), .Y(n_610) );
OAI22xp5_ASAP7_75t_L g611 ( .A1(n_578), .A2(n_517), .B1(n_552), .B2(n_537), .Y(n_611) );
INVx2_ASAP7_75t_L g612 ( .A(n_572), .Y(n_612) );
NOR2xp33_ASAP7_75t_L g613 ( .A(n_567), .B(n_551), .Y(n_613) );
OAI21xp5_ASAP7_75t_SL g614 ( .A1(n_583), .A2(n_529), .B(n_537), .Y(n_614) );
AOI22xp5_ASAP7_75t_L g615 ( .A1(n_575), .A2(n_560), .B1(n_507), .B2(n_506), .Y(n_615) );
OAI22xp33_ASAP7_75t_L g616 ( .A1(n_571), .A2(n_529), .B1(n_589), .B2(n_586), .Y(n_616) );
OAI21xp5_ASAP7_75t_L g617 ( .A1(n_571), .A2(n_528), .B(n_538), .Y(n_617) );
AOI22xp33_ASAP7_75t_L g618 ( .A1(n_584), .A2(n_485), .B1(n_487), .B2(n_538), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_596), .B(n_528), .Y(n_619) );
INVxp67_ASAP7_75t_L g620 ( .A(n_600), .Y(n_620) );
INVx2_ASAP7_75t_L g621 ( .A(n_572), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_581), .Y(n_622) );
A2O1A1Ixp33_ASAP7_75t_L g623 ( .A1(n_614), .A2(n_579), .B(n_588), .C(n_596), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_620), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_620), .Y(n_625) );
NAND2xp5_ASAP7_75t_SL g626 ( .A(n_616), .B(n_579), .Y(n_626) );
AND2x2_ASAP7_75t_L g627 ( .A(n_602), .B(n_569), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_622), .Y(n_628) );
OAI21xp5_ASAP7_75t_L g629 ( .A1(n_603), .A2(n_592), .B(n_593), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_619), .Y(n_630) );
AND2x2_ASAP7_75t_L g631 ( .A(n_618), .B(n_592), .Y(n_631) );
AOI21xp5_ASAP7_75t_L g632 ( .A1(n_616), .A2(n_590), .B(n_558), .Y(n_632) );
OAI221xp5_ASAP7_75t_L g633 ( .A1(n_608), .A2(n_594), .B1(n_570), .B2(n_573), .C(n_587), .Y(n_633) );
INVxp67_ASAP7_75t_L g634 ( .A(n_601), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_615), .B(n_593), .Y(n_635) );
OAI211xp5_ASAP7_75t_L g636 ( .A1(n_634), .A2(n_606), .B(n_610), .C(n_611), .Y(n_636) );
AOI221xp5_ASAP7_75t_L g637 ( .A1(n_626), .A2(n_618), .B1(n_609), .B2(n_617), .C(n_613), .Y(n_637) );
NAND2xp33_ASAP7_75t_R g638 ( .A(n_632), .B(n_604), .Y(n_638) );
OAI211xp5_ASAP7_75t_L g639 ( .A1(n_626), .A2(n_605), .B(n_607), .C(n_621), .Y(n_639) );
OAI221xp5_ASAP7_75t_L g640 ( .A1(n_623), .A2(n_612), .B1(n_568), .B2(n_576), .C(n_599), .Y(n_640) );
AOI221xp5_ASAP7_75t_L g641 ( .A1(n_623), .A2(n_591), .B1(n_582), .B2(n_580), .C(n_485), .Y(n_641) );
INVx2_ASAP7_75t_L g642 ( .A(n_627), .Y(n_642) );
AOI21xp5_ASAP7_75t_L g643 ( .A1(n_636), .A2(n_629), .B(n_633), .Y(n_643) );
NOR2xp33_ASAP7_75t_L g644 ( .A(n_639), .B(n_625), .Y(n_644) );
AOI221xp5_ASAP7_75t_SL g645 ( .A1(n_637), .A2(n_631), .B1(n_624), .B2(n_635), .C(n_630), .Y(n_645) );
NOR2xp33_ASAP7_75t_L g646 ( .A(n_640), .B(n_628), .Y(n_646) );
NOR3xp33_ASAP7_75t_SL g647 ( .A(n_643), .B(n_638), .C(n_641), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_644), .Y(n_648) );
NOR3xp33_ASAP7_75t_SL g649 ( .A(n_646), .B(n_642), .C(n_627), .Y(n_649) );
NOR4xp25_ASAP7_75t_L g650 ( .A(n_648), .B(n_645), .C(n_582), .D(n_580), .Y(n_650) );
INVx2_ASAP7_75t_L g651 ( .A(n_647), .Y(n_651) );
BUFx3_ASAP7_75t_L g652 ( .A(n_651), .Y(n_652) );
AOI22xp5_ASAP7_75t_L g653 ( .A1(n_652), .A2(n_649), .B1(n_650), .B2(n_542), .Y(n_653) );
OAI22xp5_ASAP7_75t_L g654 ( .A1(n_653), .A2(n_652), .B1(n_532), .B2(n_542), .Y(n_654) );
INVxp67_ASAP7_75t_SL g655 ( .A(n_654), .Y(n_655) );
NAND3xp33_ASAP7_75t_SL g656 ( .A(n_655), .B(n_550), .C(n_468), .Y(n_656) );
AOI211xp5_ASAP7_75t_L g657 ( .A1(n_656), .A2(n_550), .B(n_487), .C(n_510), .Y(n_657) );
endmodule