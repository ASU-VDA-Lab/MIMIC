module fake_jpeg_30290_n_182 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_182);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_182;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx4f_ASAP7_75t_L g53 ( 
.A(n_52),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_11),
.Y(n_55)
);

CKINVDCx9p33_ASAP7_75t_R g56 ( 
.A(n_49),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_43),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_0),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_6),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_9),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_10),
.Y(n_63)
);

BUFx24_ASAP7_75t_L g64 ( 
.A(n_4),
.Y(n_64)
);

CKINVDCx14_ASAP7_75t_R g65 ( 
.A(n_25),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_24),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_18),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_26),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_13),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_28),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_48),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_19),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_27),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_3),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_37),
.Y(n_76)
);

BUFx16f_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_56),
.B(n_0),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_86),
.Y(n_94)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_77),
.Y(n_82)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_78),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_68),
.Y(n_91)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_60),
.B(n_75),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_78),
.Y(n_87)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_63),
.B(n_55),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_88),
.B(n_58),
.Y(n_97)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_89),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_91),
.B(n_66),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_62),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_98),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_83),
.A2(n_58),
.B1(n_53),
.B2(n_61),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_96),
.A2(n_102),
.B1(n_103),
.B2(n_54),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_73),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_87),
.B(n_65),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_89),
.A2(n_53),
.B1(n_79),
.B2(n_65),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_82),
.A2(n_70),
.B1(n_69),
.B2(n_71),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_103),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_104),
.B(n_107),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_101),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_105),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_106),
.A2(n_111),
.B1(n_114),
.B2(n_118),
.Y(n_140)
);

A2O1A1Ixp33_ASAP7_75t_L g107 ( 
.A1(n_94),
.A2(n_72),
.B(n_64),
.C(n_3),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_95),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_108),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_101),
.Y(n_110)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_110),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_100),
.A2(n_57),
.B1(n_76),
.B2(n_74),
.Y(n_111)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_99),
.Y(n_112)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_112),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_82),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_113),
.B(n_116),
.Y(n_128)
);

OAI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_100),
.A2(n_72),
.B1(n_64),
.B2(n_73),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_115),
.B(n_16),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_92),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_117),
.B(n_122),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_95),
.A2(n_22),
.B1(n_50),
.B2(n_45),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_99),
.Y(n_119)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_119),
.Y(n_138)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_90),
.Y(n_120)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_120),
.Y(n_142)
);

OAI21xp33_ASAP7_75t_L g121 ( 
.A1(n_90),
.A2(n_21),
.B(n_42),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_121),
.A2(n_14),
.B(n_35),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_93),
.B(n_1),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_93),
.B(n_1),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_123),
.B(n_2),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_126),
.B(n_131),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_113),
.A2(n_17),
.B1(n_41),
.B2(n_40),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_129),
.B(n_134),
.Y(n_152)
);

OA22x2_ASAP7_75t_L g132 ( 
.A1(n_114),
.A2(n_15),
.B1(n_38),
.B2(n_36),
.Y(n_132)
);

O2A1O1Ixp33_ASAP7_75t_L g157 ( 
.A1(n_132),
.A2(n_30),
.B(n_31),
.C(n_33),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_133),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_117),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_109),
.B(n_5),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_135),
.B(n_137),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_108),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_121),
.B(n_7),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_141),
.B(n_145),
.Y(n_158)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_105),
.Y(n_143)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_143),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_110),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_144),
.B(n_138),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_104),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_128),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_146),
.B(n_148),
.Y(n_164)
);

AND2x4_ASAP7_75t_L g149 ( 
.A(n_125),
.B(n_12),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_149),
.Y(n_168)
);

MAJx2_ASAP7_75t_L g150 ( 
.A(n_124),
.B(n_32),
.C(n_29),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_150),
.A2(n_151),
.B(n_51),
.Y(n_169)
);

NAND2x1_ASAP7_75t_L g151 ( 
.A(n_132),
.B(n_12),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g153 ( 
.A(n_127),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_153),
.B(n_155),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_129),
.Y(n_155)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_157),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_140),
.B(n_34),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_160),
.B(n_140),
.Y(n_163)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_130),
.Y(n_161)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_161),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_163),
.B(n_169),
.Y(n_172)
);

AO221x1_ASAP7_75t_L g166 ( 
.A1(n_147),
.A2(n_127),
.B1(n_139),
.B2(n_142),
.C(n_136),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_166),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_164),
.B(n_154),
.C(n_150),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_170),
.B(n_158),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_165),
.B(n_159),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_173),
.A2(n_162),
.B1(n_152),
.B2(n_154),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_174),
.B(n_175),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_176),
.B(n_174),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_177),
.A2(n_172),
.B1(n_168),
.B2(n_151),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_168),
.C(n_171),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_179),
.A2(n_157),
.B(n_156),
.Y(n_180)
);

O2A1O1Ixp33_ASAP7_75t_SL g181 ( 
.A1(n_180),
.A2(n_149),
.B(n_132),
.C(n_167),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_181),
.B(n_149),
.Y(n_182)
);


endmodule