module fake_jpeg_21527_n_172 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_172);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_172;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVxp67_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_17),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_35),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_1),
.Y(n_58)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_29),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_8),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_47),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_14),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_4),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_18),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_20),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_4),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_7),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_44),
.Y(n_73)
);

INVx6_ASAP7_75t_SL g74 ( 
.A(n_45),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_11),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_0),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_38),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

BUFx8_ASAP7_75t_L g79 ( 
.A(n_28),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_84),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_81),
.Y(n_89)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

INVx2_ASAP7_75t_SL g84 ( 
.A(n_75),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

INVx2_ASAP7_75t_SL g88 ( 
.A(n_86),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_86),
.B(n_51),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_87),
.B(n_72),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_67),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_90),
.B(n_95),
.Y(n_100)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_97),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_85),
.B(n_64),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_84),
.A2(n_59),
.B1(n_62),
.B2(n_70),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_94),
.Y(n_98)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_98),
.Y(n_119)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_89),
.Y(n_99)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_99),
.Y(n_118)
);

INVx13_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_101),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_102),
.Y(n_124)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_94),
.Y(n_103)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_103),
.Y(n_122)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_89),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_104),
.Y(n_111)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_105),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_92),
.A2(n_96),
.B1(n_93),
.B2(n_61),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_106),
.A2(n_79),
.B1(n_77),
.B2(n_68),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_110),
.Y(n_125)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_97),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_108),
.A2(n_58),
.B(n_76),
.Y(n_116)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_91),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_109),
.A2(n_57),
.B1(n_71),
.B2(n_60),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_112),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_100),
.A2(n_66),
.B1(n_78),
.B2(n_56),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_113),
.A2(n_117),
.B1(n_120),
.B2(n_126),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_114),
.A2(n_115),
.B1(n_123),
.B2(n_2),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_99),
.A2(n_71),
.B1(n_55),
.B2(n_54),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_116),
.B(n_128),
.Y(n_135)
);

O2A1O1Ixp33_ASAP7_75t_L g117 ( 
.A1(n_106),
.A2(n_48),
.B(n_69),
.C(n_65),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_101),
.A2(n_77),
.B1(n_73),
.B2(n_49),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_109),
.A2(n_63),
.B1(n_30),
.B2(n_42),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_109),
.A2(n_74),
.B1(n_79),
.B2(n_53),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_100),
.B(n_76),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_125),
.B(n_0),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_129),
.B(n_132),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_130),
.A2(n_138),
.B1(n_141),
.B2(n_9),
.Y(n_151)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_119),
.Y(n_131)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_131),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_121),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_118),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_133),
.B(n_134),
.Y(n_150)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_122),
.Y(n_134)
);

XNOR2x1_ASAP7_75t_L g136 ( 
.A(n_112),
.B(n_2),
.Y(n_136)
);

XOR2x2_ASAP7_75t_L g149 ( 
.A(n_136),
.B(n_9),
.Y(n_149)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_119),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_127),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_139),
.A2(n_111),
.B(n_6),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_123),
.B(n_3),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_140),
.B(n_142),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_114),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_117),
.B(n_26),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_135),
.B(n_124),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_144),
.B(n_142),
.C(n_137),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_146),
.B(n_149),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_143),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_147),
.A2(n_151),
.B1(n_136),
.B2(n_143),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_150),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_153),
.B(n_154),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_148),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_156),
.A2(n_157),
.B1(n_149),
.B2(n_145),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_158),
.B(n_155),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_160),
.B(n_158),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_159),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_162),
.Y(n_163)
);

AOI21x1_ASAP7_75t_L g164 ( 
.A1(n_163),
.A2(n_153),
.B(n_152),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_150),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_10),
.C(n_12),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_15),
.Y(n_167)
);

AO21x1_ASAP7_75t_L g168 ( 
.A1(n_167),
.A2(n_22),
.B(n_23),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_168),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_169),
.B(n_27),
.C(n_31),
.Y(n_170)
);

OAI21xp33_ASAP7_75t_L g171 ( 
.A1(n_170),
.A2(n_41),
.B(n_33),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_171),
.B(n_40),
.Y(n_172)
);


endmodule