module fake_jpeg_8777_n_78 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_78);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_78;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

INVx1_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_9),
.B(n_4),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_3),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_5),
.B(n_8),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_1),
.B(n_2),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_15),
.B(n_0),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_22),
.B(n_23),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_15),
.B(n_0),
.Y(n_23)
);

A2O1A1Ixp33_ASAP7_75t_L g24 ( 
.A1(n_18),
.A2(n_0),
.B(n_1),
.C(n_3),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_24),
.B(n_27),
.Y(n_34)
);

HAxp5_ASAP7_75t_SL g25 ( 
.A(n_13),
.B(n_1),
.CON(n_25),
.SN(n_25)
);

O2A1O1Ixp33_ASAP7_75t_L g32 ( 
.A1(n_25),
.A2(n_10),
.B(n_17),
.C(n_14),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_28),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_20),
.B(n_3),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_22),
.B(n_10),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_36),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_32),
.A2(n_13),
.B1(n_21),
.B2(n_6),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_22),
.B(n_20),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_16),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_37),
.B(n_19),
.Y(n_41)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_24),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_39),
.A2(n_24),
.B1(n_29),
.B2(n_23),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_40),
.B(n_41),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_45),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_34),
.A2(n_29),
.B1(n_32),
.B2(n_38),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_28),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_16),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_46),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_SL g47 ( 
.A(n_34),
.B(n_25),
.Y(n_47)
);

AO22x1_ASAP7_75t_L g58 ( 
.A1(n_47),
.A2(n_50),
.B1(n_31),
.B2(n_30),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_36),
.A2(n_29),
.B1(n_14),
.B2(n_17),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_49),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_30),
.B(n_19),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_50),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_51),
.B(n_52),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g59 ( 
.A(n_58),
.B(n_42),
.Y(n_59)
);

AOI322xp5_ASAP7_75t_L g67 ( 
.A1(n_59),
.A2(n_40),
.A3(n_58),
.B1(n_51),
.B2(n_54),
.C1(n_46),
.C2(n_38),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_55),
.B(n_42),
.Y(n_60)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_56),
.B(n_43),
.C(n_47),
.Y(n_61)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_57),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_62),
.A2(n_35),
.B1(n_12),
.B2(n_21),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_67),
.B(n_68),
.C(n_61),
.Y(n_69)
);

AOI222xp33_ASAP7_75t_L g73 ( 
.A1(n_69),
.A2(n_21),
.B1(n_26),
.B2(n_28),
.C1(n_8),
.C2(n_5),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_66),
.B(n_63),
.C(n_64),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_70),
.B(n_71),
.C(n_65),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_66),
.A2(n_65),
.B(n_64),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_72),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_73),
.A2(n_28),
.B1(n_26),
.B2(n_5),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_74),
.B(n_4),
.Y(n_76)
);

AOI322xp5_ASAP7_75t_L g77 ( 
.A1(n_76),
.A2(n_4),
.A3(n_26),
.B1(n_28),
.B2(n_75),
.C1(n_68),
.C2(n_71),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_28),
.Y(n_78)
);


endmodule