module fake_jpeg_29007_n_317 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_317);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_317;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx4f_ASAP7_75t_SL g33 ( 
.A(n_17),
.Y(n_33)
);

BUFx8_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_10),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_7),
.B(n_15),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_41),
.Y(n_88)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_9),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_47),
.Y(n_59)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_46),
.Y(n_95)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx6_ASAP7_75t_SL g49 ( 
.A(n_20),
.Y(n_49)
);

INVx5_ASAP7_75t_SL g99 ( 
.A(n_49),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_51),
.B(n_53),
.Y(n_87)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_39),
.B(n_0),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_54),
.B(n_34),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_41),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_55),
.B(n_80),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_40),
.C(n_36),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_56),
.B(n_69),
.Y(n_123)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_57),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_45),
.B(n_24),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_58),
.B(n_62),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_52),
.A2(n_40),
.B1(n_31),
.B2(n_35),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_61),
.A2(n_78),
.B1(n_83),
.B2(n_89),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_18),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_42),
.B(n_24),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_63),
.B(n_68),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_48),
.A2(n_40),
.B1(n_31),
.B2(n_35),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_65),
.A2(n_85),
.B1(n_102),
.B2(n_1),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_18),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_67),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_28),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_28),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_51),
.B(n_21),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_70),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_49),
.A2(n_29),
.B1(n_35),
.B2(n_26),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_71),
.A2(n_72),
.B1(n_77),
.B2(n_82),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_53),
.A2(n_29),
.B1(n_35),
.B2(n_26),
.Y(n_72)
);

BUFx12_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

INVx13_ASAP7_75t_L g124 ( 
.A(n_73),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_53),
.A2(n_29),
.B1(n_26),
.B2(n_22),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_46),
.A2(n_26),
.B1(n_29),
.B2(n_23),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_51),
.A2(n_38),
.B1(n_30),
.B2(n_32),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_79),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_50),
.B(n_23),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_50),
.B(n_32),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_81),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_49),
.A2(n_22),
.B1(n_30),
.B2(n_27),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_44),
.A2(n_27),
.B1(n_25),
.B2(n_38),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_49),
.A2(n_25),
.B1(n_34),
.B2(n_33),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_84),
.A2(n_91),
.B1(n_96),
.B2(n_97),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_L g85 ( 
.A1(n_48),
.A2(n_34),
.B1(n_33),
.B2(n_2),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_44),
.A2(n_34),
.B1(n_33),
.B2(n_11),
.Y(n_89)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_90),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_49),
.A2(n_34),
.B1(n_33),
.B2(n_11),
.Y(n_91)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_41),
.Y(n_92)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_92),
.Y(n_120)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_93),
.Y(n_108)
);

OR2x4_ASAP7_75t_L g126 ( 
.A(n_94),
.B(n_1),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_49),
.A2(n_33),
.B1(n_9),
.B2(n_11),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_49),
.A2(n_8),
.B1(n_16),
.B2(n_15),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_44),
.Y(n_98)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_98),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_45),
.B(n_6),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_100),
.A2(n_101),
.B(n_13),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_45),
.B(n_6),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_L g102 ( 
.A1(n_48),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_102)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_60),
.Y(n_106)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_106),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g111 ( 
.A(n_73),
.Y(n_111)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_111),
.Y(n_167)
);

BUFx12f_ASAP7_75t_L g113 ( 
.A(n_60),
.Y(n_113)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_113),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_75),
.A2(n_76),
.B1(n_99),
.B2(n_95),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_115),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_116),
.B(n_130),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_75),
.A2(n_13),
.B1(n_16),
.B2(n_4),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_117),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_118),
.B(n_125),
.Y(n_163)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_93),
.Y(n_121)
);

INVx1_ASAP7_75t_SL g152 ( 
.A(n_121),
.Y(n_152)
);

NOR2x1_ASAP7_75t_R g156 ( 
.A(n_126),
.B(n_17),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_56),
.A2(n_5),
.B1(n_12),
.B2(n_14),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_128),
.A2(n_132),
.B1(n_3),
.B2(n_99),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_87),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_76),
.A2(n_5),
.B1(n_12),
.B2(n_14),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_131),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_68),
.A2(n_12),
.B1(n_15),
.B2(n_16),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_99),
.A2(n_3),
.B1(n_17),
.B2(n_95),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_134),
.Y(n_165)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_64),
.Y(n_135)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_135),
.Y(n_139)
);

FAx1_ASAP7_75t_SL g137 ( 
.A(n_123),
.B(n_69),
.CI(n_80),
.CON(n_137),
.SN(n_137)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_137),
.B(n_164),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_114),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_138),
.B(n_142),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_103),
.B(n_59),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_140),
.B(n_145),
.Y(n_175)
);

OA21x2_ASAP7_75t_L g141 ( 
.A1(n_109),
.A2(n_87),
.B(n_79),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_141),
.Y(n_176)
);

A2O1A1Ixp33_ASAP7_75t_L g142 ( 
.A1(n_133),
.A2(n_94),
.B(n_59),
.C(n_101),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_118),
.A2(n_78),
.B1(n_86),
.B2(n_74),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_143),
.A2(n_158),
.B1(n_163),
.B2(n_90),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_123),
.B(n_63),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_123),
.B(n_74),
.C(n_98),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_146),
.B(n_161),
.C(n_125),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_114),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_148),
.B(n_162),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_119),
.A2(n_81),
.B(n_65),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_149),
.A2(n_66),
.B(n_120),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_133),
.B(n_64),
.Y(n_150)
);

A2O1A1O1Ixp25_ASAP7_75t_L g202 ( 
.A1(n_150),
.A2(n_153),
.B(n_155),
.C(n_168),
.D(n_113),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_122),
.B(n_58),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_122),
.B(n_100),
.Y(n_155)
);

OAI21xp33_ASAP7_75t_SL g189 ( 
.A1(n_156),
.A2(n_73),
.B(n_107),
.Y(n_189)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_105),
.Y(n_157)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_157),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_119),
.A2(n_55),
.B1(n_57),
.B2(n_92),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_105),
.Y(n_159)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_159),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_130),
.B(n_66),
.C(n_57),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_111),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_127),
.B(n_104),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_104),
.B(n_116),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_166),
.B(n_170),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_128),
.B(n_92),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_169),
.A2(n_148),
.B1(n_151),
.B2(n_147),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_124),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_171),
.B(n_190),
.C(n_191),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_163),
.A2(n_112),
.B1(n_126),
.B2(n_135),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_174),
.A2(n_179),
.B1(n_198),
.B2(n_201),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_163),
.A2(n_110),
.B1(n_132),
.B2(n_120),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_180),
.A2(n_192),
.B1(n_170),
.B2(n_152),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_136),
.A2(n_110),
.B(n_108),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_181),
.A2(n_188),
.B(n_200),
.Y(n_215)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_139),
.Y(n_182)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_182),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_164),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_185),
.B(n_187),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_137),
.B(n_121),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_186),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_140),
.B(n_108),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_189),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_146),
.B(n_107),
.C(n_129),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_145),
.B(n_73),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_143),
.A2(n_107),
.B1(n_88),
.B2(n_106),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_162),
.B(n_124),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_193),
.B(n_194),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_167),
.B(n_124),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_167),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_195),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_160),
.Y(n_196)
);

BUFx12f_ASAP7_75t_L g211 ( 
.A(n_196),
.Y(n_211)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_139),
.Y(n_197)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_197),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_138),
.A2(n_88),
.B1(n_129),
.B2(n_60),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_157),
.Y(n_199)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_199),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_144),
.A2(n_129),
.B(n_90),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_202),
.B(n_137),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_176),
.A2(n_168),
.B1(n_136),
.B2(n_141),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_204),
.A2(n_206),
.B1(n_174),
.B2(n_202),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_176),
.A2(n_158),
.B1(n_149),
.B2(n_141),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_209),
.B(n_220),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_173),
.Y(n_214)
);

INVx13_ASAP7_75t_L g233 ( 
.A(n_214),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_217),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_171),
.B(n_150),
.C(n_161),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_219),
.B(n_221),
.C(n_222),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_184),
.B(n_155),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_190),
.B(n_142),
.C(n_166),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_191),
.B(n_153),
.C(n_141),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_180),
.A2(n_169),
.B1(n_165),
.B2(n_156),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_223),
.B(n_179),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_188),
.A2(n_152),
.B(n_154),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_224),
.A2(n_200),
.B(n_181),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_183),
.B(n_154),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_226),
.B(n_178),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_228),
.A2(n_230),
.B(n_205),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_229),
.A2(n_243),
.B1(n_245),
.B2(n_204),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_215),
.A2(n_195),
.B(n_186),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_213),
.B(n_186),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_232),
.B(n_246),
.Y(n_259)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_210),
.Y(n_234)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_234),
.Y(n_255)
);

BUFx12_ASAP7_75t_L g235 ( 
.A(n_211),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_235),
.B(n_241),
.Y(n_257)
);

NOR3xp33_ASAP7_75t_SL g236 ( 
.A(n_220),
.B(n_175),
.C(n_172),
.Y(n_236)
);

NAND3xp33_ASAP7_75t_SL g253 ( 
.A(n_236),
.B(n_217),
.C(n_216),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_213),
.B(n_175),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_237),
.B(n_219),
.C(n_215),
.Y(n_256)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_210),
.Y(n_238)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_238),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_239),
.A2(n_208),
.B1(n_203),
.B2(n_221),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_207),
.B(n_185),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_212),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_242),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_207),
.B(n_172),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_244),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_225),
.B(n_198),
.Y(n_245)
);

FAx1_ASAP7_75t_SL g246 ( 
.A(n_222),
.B(n_192),
.CI(n_199),
.CON(n_246),
.SN(n_246)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_226),
.B(n_182),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_247),
.B(n_218),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_248),
.A2(n_230),
.B1(n_240),
.B2(n_232),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_249),
.A2(n_239),
.B1(n_227),
.B2(n_241),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_250),
.A2(n_228),
.B(n_247),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_229),
.A2(n_223),
.B1(n_209),
.B2(n_208),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_252),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_253),
.B(n_236),
.Y(n_274)
);

BUFx2_ASAP7_75t_L g254 ( 
.A(n_235),
.Y(n_254)
);

INVx13_ASAP7_75t_L g276 ( 
.A(n_254),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_256),
.B(n_260),
.C(n_261),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_231),
.B(n_224),
.C(n_212),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_231),
.B(n_218),
.C(n_197),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g277 ( 
.A(n_262),
.B(n_259),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_237),
.B(n_177),
.C(n_178),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_263),
.B(n_227),
.C(n_246),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_265),
.B(n_266),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_259),
.B(n_244),
.Y(n_266)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_257),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_268),
.B(n_278),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_269),
.A2(n_250),
.B(n_260),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_270),
.A2(n_245),
.B1(n_258),
.B2(n_255),
.Y(n_279)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_251),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_271),
.B(n_272),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_256),
.B(n_246),
.C(n_243),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_273),
.B(n_274),
.Y(n_286)
);

FAx1_ASAP7_75t_SL g287 ( 
.A(n_277),
.B(n_266),
.CI(n_273),
.CON(n_287),
.SN(n_287)
);

HB1xp67_ASAP7_75t_L g278 ( 
.A(n_262),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_279),
.B(n_287),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_L g281 ( 
.A1(n_268),
.A2(n_225),
.B1(n_254),
.B2(n_264),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_281),
.B(n_242),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_282),
.A2(n_283),
.B(n_265),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_269),
.A2(n_252),
.B(n_246),
.Y(n_283)
);

INVx6_ASAP7_75t_L g284 ( 
.A(n_276),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_284),
.B(n_289),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_275),
.B(n_234),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_286),
.B(n_261),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_291),
.B(n_293),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_292),
.B(n_279),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_280),
.B(n_267),
.C(n_272),
.Y(n_293)
);

OA21x2_ASAP7_75t_SL g294 ( 
.A1(n_285),
.A2(n_236),
.B(n_267),
.Y(n_294)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_294),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_295),
.B(n_285),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_282),
.A2(n_275),
.B(n_238),
.Y(n_296)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_296),
.Y(n_302)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_299),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_290),
.B(n_284),
.Y(n_301)
);

NAND3xp33_ASAP7_75t_L g309 ( 
.A(n_301),
.B(n_233),
.C(n_276),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_292),
.A2(n_289),
.B(n_283),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_303),
.A2(n_304),
.B(n_297),
.Y(n_305)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_305),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_298),
.B(n_293),
.C(n_297),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_306),
.A2(n_307),
.B(n_303),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_300),
.A2(n_288),
.B(n_287),
.Y(n_307)
);

AOI21x1_ASAP7_75t_L g312 ( 
.A1(n_309),
.A2(n_233),
.B(n_235),
.Y(n_312)
);

AO21x1_ASAP7_75t_L g313 ( 
.A1(n_311),
.A2(n_312),
.B(n_302),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_313),
.A2(n_314),
.B(n_263),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_310),
.B(n_308),
.C(n_304),
.Y(n_314)
);

BUFx24_ASAP7_75t_SL g316 ( 
.A(n_315),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_316),
.B(n_287),
.Y(n_317)
);


endmodule