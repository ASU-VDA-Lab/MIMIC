module real_jpeg_32640_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_661;
wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_630;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_663;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_648;
wire n_541;
wire n_441;
wire n_657;
wire n_643;
wire n_656;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_669;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_640;
wire n_666;
wire n_160;
wire n_211;
wire n_574;
wire n_627;
wire n_595;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_578;
wire n_456;
wire n_620;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_668;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_605;
wire n_483;
wire n_367;
wire n_639;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_658;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_516;
wire n_348;
wire n_473;
wire n_252;
wire n_601;
wire n_655;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_611;
wire n_104;
wire n_153;
wire n_634;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_646;
wire n_214;
wire n_671;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_631;
wire n_338;
wire n_175;
wire n_653;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_650;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_262;
wire n_652;
wire n_334;
wire n_647;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_651;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_615;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_672;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_670;
wire n_524;
wire n_589;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_644;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_632;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_633;
wire n_497;
wire n_638;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_596;
wire n_617;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_594;
wire n_161;
wire n_207;
wire n_526;
wire n_604;
wire n_420;
wire n_357;
wire n_431;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_572;
wire n_586;
wire n_548;
wire n_319;
wire n_664;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_637;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_613;
wire n_231;
wire n_44;
wire n_635;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_642;
wire n_172;
wire n_546;
wire n_285;
wire n_531;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_654;
wire n_616;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_667;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_628;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_662;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_649;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_636;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_597;
wire n_618;
wire n_609;
wire n_94;
wire n_645;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_641;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_629;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_659;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_660;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_625;
wire n_96;
wire n_665;
wire n_308;
wire n_433;
wire n_364;

BUFx3_ASAP7_75t_L g223 ( 
.A(n_0),
.Y(n_223)
);

BUFx12f_ASAP7_75t_L g233 ( 
.A(n_0),
.Y(n_233)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_0),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_0),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_1),
.A2(n_339),
.B(n_342),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_1),
.B(n_343),
.Y(n_342)
);

INVx2_ASAP7_75t_SL g397 ( 
.A(n_1),
.Y(n_397)
);

OAI32xp33_ASAP7_75t_L g500 ( 
.A1(n_1),
.A2(n_162),
.A3(n_501),
.B1(n_505),
.B2(n_508),
.Y(n_500)
);

AOI22xp33_ASAP7_75t_L g541 ( 
.A1(n_1),
.A2(n_397),
.B1(n_542),
.B2(n_543),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_1),
.B(n_134),
.Y(n_595)
);

OAI22xp33_ASAP7_75t_SL g629 ( 
.A1(n_1),
.A2(n_222),
.B1(n_616),
.B2(n_630),
.Y(n_629)
);

AO22x1_ASAP7_75t_L g265 ( 
.A1(n_2),
.A2(n_266),
.B1(n_268),
.B2(n_269),
.Y(n_265)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_2),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_2),
.A2(n_76),
.B1(n_268),
.B2(n_276),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_2),
.A2(n_268),
.B1(n_357),
.B2(n_360),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_2),
.A2(n_268),
.B1(n_379),
.B2(n_383),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_4),
.A2(n_76),
.B1(n_346),
.B2(n_347),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_4),
.Y(n_346)
);

AOI22xp33_ASAP7_75t_SL g368 ( 
.A1(n_4),
.A2(n_346),
.B1(n_369),
.B2(n_372),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g572 ( 
.A1(n_4),
.A2(n_346),
.B1(n_573),
.B2(n_575),
.Y(n_572)
);

AOI22xp5_ASAP7_75t_SL g616 ( 
.A1(n_4),
.A2(n_346),
.B1(n_617),
.B2(n_619),
.Y(n_616)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_5),
.A2(n_75),
.B1(n_79),
.B2(n_80),
.Y(n_74)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_5),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_5),
.A2(n_79),
.B1(n_211),
.B2(n_214),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_5),
.A2(n_79),
.B1(n_197),
.B2(n_241),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_5),
.A2(n_79),
.B1(n_227),
.B2(n_392),
.Y(n_391)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_6),
.A2(n_61),
.B1(n_65),
.B2(n_68),
.Y(n_60)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_6),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_6),
.A2(n_68),
.B1(n_123),
.B2(n_127),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_6),
.A2(n_68),
.B1(n_146),
.B2(n_151),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_6),
.A2(n_68),
.B1(n_235),
.B2(n_236),
.Y(n_234)
);

OAI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_7),
.A2(n_257),
.B1(n_259),
.B2(n_260),
.Y(n_256)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_7),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g351 ( 
.A1(n_7),
.A2(n_259),
.B1(n_352),
.B2(n_355),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_7),
.A2(n_259),
.B1(n_445),
.B2(n_446),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_SL g516 ( 
.A1(n_7),
.A2(n_259),
.B1(n_517),
.B2(n_520),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_8),
.A2(n_249),
.B1(n_251),
.B2(n_252),
.Y(n_248)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_8),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_8),
.A2(n_251),
.B1(n_329),
.B2(n_333),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g497 ( 
.A1(n_8),
.A2(n_251),
.B1(n_355),
.B2(n_498),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g584 ( 
.A1(n_8),
.A2(n_226),
.B1(n_251),
.B2(n_585),
.Y(n_584)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_9),
.A2(n_61),
.B1(n_83),
.B2(n_88),
.Y(n_82)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_9),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_9),
.A2(n_88),
.B1(n_205),
.B2(n_207),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g242 ( 
.A1(n_9),
.A2(n_88),
.B1(n_241),
.B2(n_243),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_9),
.A2(n_88),
.B1(n_236),
.B2(n_421),
.Y(n_420)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_10),
.A2(n_50),
.B1(n_54),
.B2(n_58),
.Y(n_49)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_10),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_10),
.A2(n_58),
.B1(n_170),
.B2(n_174),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g193 ( 
.A1(n_10),
.A2(n_58),
.B1(n_194),
.B2(n_197),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_10),
.A2(n_58),
.B1(n_226),
.B2(n_231),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_11),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_12),
.Y(n_139)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_12),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_13),
.Y(n_96)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_13),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_13),
.Y(n_386)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_13),
.Y(n_589)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_14),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_15),
.A2(n_21),
.B(n_671),
.Y(n_20)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_15),
.Y(n_672)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_16),
.A2(n_320),
.B1(n_324),
.B2(n_325),
.Y(n_319)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_16),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_16),
.A2(n_76),
.B1(n_324),
.B2(n_437),
.Y(n_436)
);

AOI22xp33_ASAP7_75t_L g547 ( 
.A1(n_16),
.A2(n_197),
.B1(n_324),
.B2(n_548),
.Y(n_547)
);

AOI22xp33_ASAP7_75t_SL g603 ( 
.A1(n_16),
.A2(n_324),
.B1(n_604),
.B2(n_607),
.Y(n_603)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_17),
.Y(n_110)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_17),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_17),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_18),
.B(n_672),
.Y(n_671)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_19),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_19),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_19),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_183),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_182),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_69),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_25),
.B(n_69),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_49),
.B1(n_59),
.B2(n_60),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_26),
.A2(n_59),
.B1(n_73),
.B2(n_82),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_26),
.A2(n_49),
.B1(n_59),
.B2(n_82),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_26),
.A2(n_59),
.B1(n_248),
.B2(n_255),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_26),
.A2(n_59),
.B1(n_338),
.B2(n_345),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g456 ( 
.A1(n_26),
.A2(n_59),
.B1(n_248),
.B2(n_436),
.Y(n_456)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AO22x1_ASAP7_75t_L g274 ( 
.A1(n_27),
.A2(n_256),
.B1(n_275),
.B2(n_279),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_27),
.A2(n_74),
.B1(n_275),
.B2(n_279),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_27),
.A2(n_279),
.B1(n_435),
.B2(n_441),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_39),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_32),
.B1(n_35),
.B2(n_37),
.Y(n_28)
);

INVx3_ASAP7_75t_SL g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_31),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_31),
.Y(n_250)
);

INVx3_ASAP7_75t_L g440 ( 
.A(n_31),
.Y(n_440)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_34),
.Y(n_404)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_35),
.Y(n_341)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_36),
.Y(n_344)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

HB1xp67_ASAP7_75t_L g411 ( 
.A(n_38),
.Y(n_411)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_42),
.B1(n_45),
.B2(n_47),
.Y(n_39)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_40),
.Y(n_206)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_41),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_41),
.Y(n_271)
);

INVx4_ASAP7_75t_SL g42 ( 
.A(n_43),
.Y(n_42)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_46),
.Y(n_161)
);

INVx2_ASAP7_75t_SL g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx4_ASAP7_75t_SL g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_53),
.Y(n_254)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_59),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_59),
.B(n_397),
.Y(n_396)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_63),
.Y(n_349)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_64),
.Y(n_408)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_178),
.C(n_179),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g661 ( 
.A1(n_70),
.A2(n_71),
.B1(n_662),
.B2(n_663),
.Y(n_661)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_89),
.C(n_131),
.Y(n_71)
);

XNOR2x1_ASAP7_75t_L g310 ( 
.A(n_72),
.B(n_311),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_78),
.Y(n_278)
);

INVx4_ASAP7_75t_SL g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_SL g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx6_ASAP7_75t_L g262 ( 
.A(n_87),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_89),
.A2(n_297),
.B(n_299),
.Y(n_296)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_90),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_90),
.B(n_307),
.C(n_308),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_SL g311 ( 
.A(n_90),
.B(n_132),
.Y(n_311)
);

AOI21x1_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_104),
.B(n_122),
.Y(n_90)
);

INVx2_ASAP7_75t_SL g202 ( 
.A(n_91),
.Y(n_202)
);

OAI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_91),
.A2(n_200),
.B1(n_240),
.B2(n_242),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_91),
.A2(n_193),
.B1(n_200),
.B2(n_242),
.Y(n_285)
);

OAI22xp33_ASAP7_75t_SL g350 ( 
.A1(n_91),
.A2(n_200),
.B1(n_351),
.B2(n_356),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g427 ( 
.A1(n_91),
.A2(n_200),
.B1(n_240),
.B2(n_356),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_L g596 ( 
.A1(n_91),
.A2(n_200),
.B1(n_547),
.B2(n_571),
.Y(n_596)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVxp33_ASAP7_75t_SL g121 ( 
.A(n_93),
.Y(n_121)
);

AO21x2_ASAP7_75t_L g200 ( 
.A1(n_93),
.A2(n_106),
.B(n_115),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_97),
.B1(n_100),
.B2(n_102),
.Y(n_93)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_94),
.Y(n_224)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_96),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_96),
.Y(n_382)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_96),
.Y(n_395)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_97),
.Y(n_116)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_98),
.Y(n_564)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_99),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_99),
.Y(n_113)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_101),
.Y(n_231)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_114),
.B(n_121),
.Y(n_104)
);

AO21x1_ASAP7_75t_L g556 ( 
.A1(n_105),
.A2(n_557),
.B(n_559),
.Y(n_556)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_111),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_109),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_110),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_110),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_110),
.Y(n_354)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVxp33_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

NAND2xp67_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_117),
.Y(n_115)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx5_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g513 ( 
.A(n_120),
.Y(n_513)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_122),
.Y(n_201)
);

INVx2_ASAP7_75t_SL g123 ( 
.A(n_124),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx4_ASAP7_75t_L g362 ( 
.A(n_125),
.Y(n_362)
);

INVx4_ASAP7_75t_L g575 ( 
.A(n_125),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_126),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_126),
.Y(n_141)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_126),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_126),
.Y(n_359)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

BUFx4f_ASAP7_75t_L g574 ( 
.A(n_128),
.Y(n_574)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_130),
.Y(n_581)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

OA22x2_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_145),
.B1(n_155),
.B2(n_169),
.Y(n_132)
);

OA22x2_ASAP7_75t_L g297 ( 
.A1(n_133),
.A2(n_155),
.B1(n_169),
.B2(n_298),
.Y(n_297)
);

OAI22xp33_ASAP7_75t_L g367 ( 
.A1(n_133),
.A2(n_155),
.B1(n_319),
.B2(n_368),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g443 ( 
.A1(n_133),
.A2(n_155),
.B1(n_328),
.B2(n_444),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g540 ( 
.A1(n_133),
.A2(n_155),
.B1(n_368),
.B2(n_541),
.Y(n_540)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_134),
.A2(n_180),
.B(n_181),
.Y(n_179)
);

AOI22x1_ASAP7_75t_L g203 ( 
.A1(n_134),
.A2(n_180),
.B1(n_204),
.B2(n_210),
.Y(n_203)
);

AOI22x1_ASAP7_75t_L g264 ( 
.A1(n_134),
.A2(n_180),
.B1(n_210),
.B2(n_265),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_134),
.A2(n_180),
.B1(n_318),
.B2(n_327),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_134),
.A2(n_180),
.B1(n_265),
.B2(n_458),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_134),
.A2(n_180),
.B1(n_265),
.B2(n_458),
.Y(n_468)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

AO21x2_ASAP7_75t_L g155 ( 
.A1(n_135),
.A2(n_156),
.B(n_162),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_137),
.B1(n_140),
.B2(n_142),
.Y(n_135)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_139),
.Y(n_159)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

HB1xp67_ASAP7_75t_L g507 ( 
.A(n_141),
.Y(n_507)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_144),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_145),
.Y(n_181)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_150),
.Y(n_213)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_150),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_150),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_150),
.Y(n_375)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx8_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx8_ASAP7_75t_L g209 ( 
.A(n_154),
.Y(n_209)
);

INVx3_ASAP7_75t_SL g180 ( 
.A(n_155),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_160),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_166),
.Y(n_162)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_163),
.Y(n_445)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_164),
.Y(n_173)
);

BUFx2_ASAP7_75t_L g401 ( 
.A(n_164),
.Y(n_401)
);

INVx8_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

HB1xp67_ASAP7_75t_L g371 ( 
.A(n_165),
.Y(n_371)
);

INVx3_ASAP7_75t_L g414 ( 
.A(n_165),
.Y(n_414)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_171),
.Y(n_170)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_174),
.Y(n_542)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g663 ( 
.A(n_178),
.B(n_179),
.Y(n_663)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_660),
.B(n_665),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_312),
.Y(n_184)
);

NOR2xp67_ASAP7_75t_SL g185 ( 
.A(n_186),
.B(n_301),
.Y(n_185)
);

NOR2xp67_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_286),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_187),
.B(n_286),
.Y(n_668)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_218),
.C(n_272),
.Y(n_187)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g479 ( 
.A1(n_189),
.A2(n_190),
.B1(n_273),
.B2(n_480),
.Y(n_479)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_203),
.B(n_217),
.Y(n_190)
);

NAND2x1p5_ASAP7_75t_L g217 ( 
.A(n_191),
.B(n_203),
.Y(n_217)
);

AOI22x1_ASAP7_75t_SL g191 ( 
.A1(n_192),
.A2(n_199),
.B1(n_201),
.B2(n_202),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_194),
.Y(n_355)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_196),
.Y(n_198)
);

BUFx6f_ASAP7_75t_SL g197 ( 
.A(n_198),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g545 ( 
.A1(n_199),
.A2(n_202),
.B1(n_497),
.B2(n_546),
.Y(n_545)
);

INVx1_ASAP7_75t_SL g576 ( 
.A(n_199),
.Y(n_576)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g494 ( 
.A1(n_200),
.A2(n_351),
.B1(n_495),
.B2(n_496),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_202),
.Y(n_495)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_204),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx5_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_209),
.Y(n_216)
);

INVx5_ASAP7_75t_L g267 ( 
.A(n_209),
.Y(n_267)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_213),
.Y(n_326)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_216),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_217),
.B(n_293),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_217),
.B(n_287),
.C(n_304),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_218),
.B(n_479),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_246),
.C(n_263),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g472 ( 
.A1(n_219),
.A2(n_220),
.B1(n_473),
.B2(n_475),
.Y(n_472)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_239),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_SL g463 ( 
.A(n_221),
.B(n_239),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_225),
.B1(n_232),
.B2(n_234),
.Y(n_221)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_222),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_222),
.A2(n_225),
.B1(n_420),
.B2(n_429),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_L g583 ( 
.A1(n_222),
.A2(n_584),
.B1(n_590),
.B2(n_593),
.Y(n_583)
);

OAI22xp5_ASAP7_75t_SL g615 ( 
.A1(n_222),
.A2(n_603),
.B1(n_616),
.B2(n_623),
.Y(n_615)
);

OR2x2_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx5_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_228),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_229),
.Y(n_618)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_230),
.Y(n_238)
);

INVx3_ASAP7_75t_L g519 ( 
.A(n_230),
.Y(n_519)
);

INVx3_ASAP7_75t_L g523 ( 
.A(n_230),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g606 ( 
.A(n_230),
.Y(n_606)
);

INVx4_ASAP7_75t_L g283 ( 
.A(n_232),
.Y(n_283)
);

INVx8_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx8_ASAP7_75t_L g418 ( 
.A(n_233),
.Y(n_418)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_234),
.Y(n_284)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

BUFx2_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_247),
.A2(n_263),
.B1(n_264),
.B2(n_474),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_247),
.Y(n_474)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx4_ASAP7_75t_L g258 ( 
.A(n_250),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx5_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx4_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_273),
.Y(n_480)
);

XNOR2x1_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_280),
.Y(n_273)
);

INVxp67_ASAP7_75t_SL g291 ( 
.A(n_274),
.Y(n_291)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

BUFx3_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

OAI21x1_ASAP7_75t_L g469 ( 
.A1(n_280),
.A2(n_290),
.B(n_470),
.Y(n_469)
);

OR2x2_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_285),
.Y(n_280)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_281),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_282),
.A2(n_283),
.B(n_284),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_282),
.A2(n_378),
.B1(n_387),
.B2(n_391),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_282),
.A2(n_391),
.B1(n_417),
.B2(n_419),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_282),
.A2(n_378),
.B1(n_516),
.B2(n_524),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_SL g601 ( 
.A1(n_282),
.A2(n_602),
.B1(n_608),
.B2(n_609),
.Y(n_601)
);

HB1xp67_ASAP7_75t_L g289 ( 
.A(n_285),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_292),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_288),
.A2(n_290),
.B(n_291),
.Y(n_287)
);

NAND2xp33_ASAP7_75t_SL g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_289),
.Y(n_470)
);

HB1xp67_ASAP7_75t_L g304 ( 
.A(n_293),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_296),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_295),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_297),
.B(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_297),
.Y(n_308)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

AOI21x1_ASAP7_75t_SL g667 ( 
.A1(n_302),
.A2(n_668),
.B(n_669),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_305),
.Y(n_302)
);

NOR2xp67_ASAP7_75t_SL g669 ( 
.A(n_303),
.B(n_305),
.Y(n_669)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_309),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g664 ( 
.A(n_306),
.B(n_307),
.C(n_310),
.Y(n_664)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_307),
.B(n_310),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_313),
.A2(n_489),
.B(n_651),
.Y(n_312)
);

NAND4xp25_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_450),
.C(n_476),
.D(n_481),
.Y(n_313)
);

OR2x2_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_424),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_315),
.B(n_424),
.Y(n_653)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_365),
.C(n_398),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g647 ( 
.A(n_316),
.B(n_648),
.Y(n_647)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_336),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_317),
.B(n_363),
.C(n_364),
.Y(n_430)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

BUFx3_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_332),
.Y(n_335)
);

INVx2_ASAP7_75t_SL g544 ( 
.A(n_332),
.Y(n_544)
);

INVx1_ASAP7_75t_SL g333 ( 
.A(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_337),
.A2(n_350),
.B1(n_363),
.B2(n_364),
.Y(n_336)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_337),
.Y(n_363)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g415 ( 
.A(n_342),
.Y(n_415)
);

INVx4_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_345),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_350),
.Y(n_364)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

BUFx2_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_359),
.Y(n_498)
);

INVx2_ASAP7_75t_SL g360 ( 
.A(n_361),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

HB1xp67_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g648 ( 
.A(n_366),
.B(n_398),
.Y(n_648)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_376),
.C(n_396),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g532 ( 
.A(n_367),
.B(n_533),
.Y(n_532)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

BUFx3_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx3_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

BUFx3_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_375),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_L g533 ( 
.A1(n_376),
.A2(n_377),
.B1(n_396),
.B2(n_534),
.Y(n_533)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

BUFx3_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

HB1xp67_ASAP7_75t_L g558 ( 
.A(n_382),
.Y(n_558)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

BUFx2_ASAP7_75t_SL g384 ( 
.A(n_385),
.Y(n_384)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_385),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g562 ( 
.A(n_386),
.Y(n_562)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_386),
.Y(n_622)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

BUFx2_ASAP7_75t_L g634 ( 
.A(n_389),
.Y(n_634)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_390),
.Y(n_626)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_396),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_397),
.B(n_509),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_397),
.B(n_566),
.Y(n_565)
);

OA21x2_ASAP7_75t_SL g577 ( 
.A1(n_397),
.A2(n_565),
.B(n_578),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_SL g627 ( 
.A(n_397),
.B(n_495),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_397),
.B(n_633),
.Y(n_632)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_399),
.A2(n_416),
.B1(n_422),
.B2(n_423),
.Y(n_398)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_399),
.Y(n_422)
);

OAI32xp33_ASAP7_75t_L g399 ( 
.A1(n_400),
.A2(n_402),
.A3(n_405),
.B1(n_409),
.B2(n_415),
.Y(n_399)
);

OAI32xp33_ASAP7_75t_L g449 ( 
.A1(n_400),
.A2(n_402),
.A3(n_405),
.B1(n_409),
.B2(n_415),
.Y(n_449)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

BUFx2_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_SL g409 ( 
.A(n_410),
.B(n_412),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx3_ASAP7_75t_SL g413 ( 
.A(n_414),
.Y(n_413)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_416),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_417),
.Y(n_429)
);

INVx5_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_421),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_423),
.B(n_449),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_423),
.B(n_449),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_425),
.B(n_431),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_430),
.Y(n_425)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_426),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_428),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_427),
.B(n_428),
.Y(n_454)
);

HB1xp67_ASAP7_75t_L g485 ( 
.A(n_430),
.Y(n_485)
);

INVxp67_ASAP7_75t_L g483 ( 
.A(n_431),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_432),
.B(n_448),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_433),
.A2(n_434),
.B1(n_442),
.B2(n_443),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

HB1xp67_ASAP7_75t_L g461 ( 
.A(n_434),
.Y(n_461)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_442),
.B(n_460),
.C(n_461),
.Y(n_459)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_444),
.Y(n_458)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_451),
.B(n_464),
.Y(n_450)
);

AOI22xp33_ASAP7_75t_L g654 ( 
.A1(n_451),
.A2(n_464),
.B1(n_482),
.B2(n_653),
.Y(n_654)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_451),
.Y(n_657)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_452),
.B(n_459),
.C(n_462),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_452),
.B(n_463),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_453),
.B(n_455),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_454),
.B(n_467),
.C(n_468),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_456),
.B(n_457),
.Y(n_455)
);

INVxp67_ASAP7_75t_SL g467 ( 
.A(n_456),
.Y(n_467)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_459),
.Y(n_487)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_464),
.Y(n_658)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_465),
.B(n_471),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_466),
.B(n_469),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_466),
.B(n_469),
.C(n_472),
.Y(n_477)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_473),
.Y(n_475)
);

A2O1A1Ixp33_ASAP7_75t_L g651 ( 
.A1(n_476),
.A2(n_652),
.B(n_654),
.C(n_655),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_477),
.B(n_478),
.Y(n_476)
);

OR2x2_ASAP7_75t_L g659 ( 
.A(n_477),
.B(n_478),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_482),
.B(n_486),
.Y(n_481)
);

OAI21xp33_ASAP7_75t_L g652 ( 
.A1(n_482),
.A2(n_486),
.B(n_653),
.Y(n_652)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_483),
.B(n_484),
.C(n_485),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_487),
.B(n_488),
.Y(n_486)
);

AOI21x1_ASAP7_75t_L g489 ( 
.A1(n_490),
.A2(n_646),
.B(n_650),
.Y(n_489)
);

OAI21x1_ASAP7_75t_SL g490 ( 
.A1(n_491),
.A2(n_552),
.B(n_645),
.Y(n_490)
);

AOI211xp5_ASAP7_75t_L g491 ( 
.A1(n_492),
.A2(n_530),
.B(n_535),
.C(n_536),
.Y(n_491)
);

A2O1A1Ixp33_ASAP7_75t_L g645 ( 
.A1(n_492),
.A2(n_530),
.B(n_535),
.C(n_536),
.Y(n_645)
);

HB1xp67_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_493),
.B(n_532),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_L g493 ( 
.A1(n_494),
.A2(n_499),
.B1(n_528),
.B2(n_529),
.Y(n_493)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_494),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g649 ( 
.A(n_494),
.B(n_528),
.C(n_531),
.Y(n_649)
);

OAI22x1_ASAP7_75t_L g570 ( 
.A1(n_495),
.A2(n_571),
.B1(n_576),
.B2(n_577),
.Y(n_570)
);

INVxp67_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_499),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_500),
.B(n_514),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g537 ( 
.A1(n_500),
.A2(n_514),
.B1(n_515),
.B2(n_538),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_500),
.Y(n_538)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

BUFx2_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_507),
.Y(n_506)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_512),
.Y(n_569)
);

INVx5_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_513),
.Y(n_551)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

INVxp67_ASAP7_75t_L g593 ( 
.A(n_516),
.Y(n_593)
);

INVx3_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

INVx4_ASAP7_75t_L g518 ( 
.A(n_519),
.Y(n_518)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);

HB1xp67_ASAP7_75t_L g521 ( 
.A(n_522),
.Y(n_521)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_522),
.Y(n_635)
);

BUFx12f_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

INVx3_ASAP7_75t_L g524 ( 
.A(n_525),
.Y(n_524)
);

INVx3_ASAP7_75t_L g525 ( 
.A(n_526),
.Y(n_525)
);

BUFx3_ASAP7_75t_L g526 ( 
.A(n_527),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g592 ( 
.A(n_527),
.Y(n_592)
);

BUFx6f_ASAP7_75t_L g611 ( 
.A(n_527),
.Y(n_611)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_531),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_532),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_537),
.B(n_539),
.C(n_545),
.Y(n_536)
);

XNOR2xp5_ASAP7_75t_L g641 ( 
.A(n_537),
.B(n_642),
.Y(n_641)
);

AOI22xp5_ASAP7_75t_L g642 ( 
.A1(n_539),
.A2(n_540),
.B1(n_545),
.B2(n_643),
.Y(n_642)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_540),
.Y(n_539)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_544),
.Y(n_543)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_545),
.Y(n_643)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_547),
.Y(n_546)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_549),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_550),
.Y(n_549)
);

INVx2_ASAP7_75t_SL g550 ( 
.A(n_551),
.Y(n_550)
);

AOI21x1_ASAP7_75t_L g552 ( 
.A1(n_553),
.A2(n_639),
.B(n_644),
.Y(n_552)
);

OAI21x1_ASAP7_75t_SL g553 ( 
.A1(n_554),
.A2(n_599),
.B(n_638),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_555),
.B(n_582),
.Y(n_554)
);

OR2x2_ASAP7_75t_L g638 ( 
.A(n_555),
.B(n_582),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_556),
.B(n_570),
.Y(n_555)
);

XNOR2xp5_ASAP7_75t_SL g612 ( 
.A(n_556),
.B(n_570),
.Y(n_612)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_558),
.Y(n_557)
);

AOI21xp5_ASAP7_75t_L g559 ( 
.A1(n_560),
.A2(n_563),
.B(n_565),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_561),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_562),
.Y(n_561)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_564),
.Y(n_563)
);

INVx3_ASAP7_75t_L g566 ( 
.A(n_567),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_568),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_569),
.Y(n_568)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_572),
.Y(n_571)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_574),
.Y(n_573)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_579),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_580),
.Y(n_579)
);

BUFx3_ASAP7_75t_L g580 ( 
.A(n_581),
.Y(n_580)
);

XNOR2xp5_ASAP7_75t_L g582 ( 
.A(n_583),
.B(n_594),
.Y(n_582)
);

MAJIxp5_ASAP7_75t_L g640 ( 
.A(n_583),
.B(n_596),
.C(n_597),
.Y(n_640)
);

INVxp67_ASAP7_75t_L g608 ( 
.A(n_584),
.Y(n_608)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_586),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_587),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_588),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_589),
.Y(n_588)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_591),
.Y(n_590)
);

HB1xp67_ASAP7_75t_L g591 ( 
.A(n_592),
.Y(n_591)
);

OAI22xp5_ASAP7_75t_L g594 ( 
.A1(n_595),
.A2(n_596),
.B1(n_597),
.B2(n_598),
.Y(n_594)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_595),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_596),
.Y(n_598)
);

AOI21x1_ASAP7_75t_L g599 ( 
.A1(n_600),
.A2(n_613),
.B(n_637),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_601),
.B(n_612),
.Y(n_600)
);

NOR2xp67_ASAP7_75t_L g637 ( 
.A(n_601),
.B(n_612),
.Y(n_637)
);

INVxp67_ASAP7_75t_L g602 ( 
.A(n_603),
.Y(n_602)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_605),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_606),
.Y(n_605)
);

INVx3_ASAP7_75t_SL g609 ( 
.A(n_610),
.Y(n_609)
);

INVx8_ASAP7_75t_L g610 ( 
.A(n_611),
.Y(n_610)
);

OAI21xp5_ASAP7_75t_SL g613 ( 
.A1(n_614),
.A2(n_628),
.B(n_636),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_615),
.B(n_627),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_615),
.B(n_627),
.Y(n_636)
);

BUFx2_ASAP7_75t_L g617 ( 
.A(n_618),
.Y(n_617)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_620),
.Y(n_619)
);

INVx4_ASAP7_75t_L g620 ( 
.A(n_621),
.Y(n_620)
);

INVx4_ASAP7_75t_L g621 ( 
.A(n_622),
.Y(n_621)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_624),
.Y(n_623)
);

INVx4_ASAP7_75t_L g630 ( 
.A(n_624),
.Y(n_630)
);

INVx4_ASAP7_75t_L g624 ( 
.A(n_625),
.Y(n_624)
);

INVx2_ASAP7_75t_SL g625 ( 
.A(n_626),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_629),
.B(n_631),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_SL g631 ( 
.A(n_632),
.B(n_635),
.Y(n_631)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_634),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_640),
.B(n_641),
.Y(n_639)
);

NOR2xp67_ASAP7_75t_SL g644 ( 
.A(n_640),
.B(n_641),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_647),
.B(n_649),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_647),
.B(n_649),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_656),
.B(n_659),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_657),
.B(n_658),
.Y(n_656)
);

OAI21xp5_ASAP7_75t_SL g666 ( 
.A1(n_660),
.A2(n_667),
.B(n_670),
.Y(n_666)
);

NOR2x1_ASAP7_75t_R g660 ( 
.A(n_661),
.B(n_664),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_661),
.B(n_664),
.Y(n_670)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_663),
.Y(n_662)
);

INVxp33_ASAP7_75t_L g665 ( 
.A(n_666),
.Y(n_665)
);


endmodule