module fake_jpeg_24294_n_283 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_283);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_283;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_16),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_37),
.B(n_40),
.Y(n_48)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_42),
.Y(n_47)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_17),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_31),
.Y(n_51)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_50),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_43),
.A2(n_31),
.B1(n_26),
.B2(n_32),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_45),
.A2(n_58),
.B1(n_32),
.B2(n_21),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_42),
.B(n_24),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_49),
.B(n_20),
.Y(n_89)
);

INVx2_ASAP7_75t_SL g50 ( 
.A(n_36),
.Y(n_50)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_42),
.B(n_34),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_63),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_43),
.A2(n_31),
.B1(n_25),
.B2(n_39),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_53),
.A2(n_62),
.B1(n_33),
.B2(n_23),
.Y(n_77)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_28),
.Y(n_55)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_28),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_56),
.B(n_55),
.Y(n_78)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_61),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_39),
.A2(n_26),
.B1(n_32),
.B2(n_21),
.Y(n_58)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_37),
.A2(n_28),
.B1(n_25),
.B2(n_17),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_35),
.B(n_34),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_63),
.B(n_0),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_65),
.B(n_78),
.Y(n_120)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_64),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_67),
.B(n_75),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_69),
.A2(n_92),
.B1(n_95),
.B2(n_67),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_51),
.A2(n_25),
.B1(n_33),
.B2(n_21),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_70),
.A2(n_91),
.B1(n_29),
.B2(n_27),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_46),
.A2(n_33),
.B1(n_23),
.B2(n_22),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_71),
.Y(n_111)
);

CKINVDCx12_ASAP7_75t_R g74 ( 
.A(n_50),
.Y(n_74)
);

CKINVDCx14_ASAP7_75t_R g105 ( 
.A(n_74),
.Y(n_105)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_48),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_48),
.B(n_40),
.C(n_37),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_76),
.B(n_82),
.C(n_86),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_77),
.A2(n_60),
.B1(n_18),
.B2(n_29),
.Y(n_114)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_79),
.B(n_81),
.Y(n_112)
);

A2O1A1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_47),
.A2(n_27),
.B(n_29),
.C(n_33),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_80),
.B(n_29),
.Y(n_101)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_47),
.B(n_40),
.C(n_38),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_61),
.B(n_24),
.Y(n_83)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_83),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_84),
.B(n_2),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_52),
.B(n_41),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_86),
.B(n_99),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_49),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_87),
.B(n_90),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

INVx13_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_89),
.B(n_93),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_46),
.A2(n_38),
.B1(n_22),
.B2(n_19),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_46),
.A2(n_20),
.B1(n_19),
.B2(n_18),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_61),
.B(n_0),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_59),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_94),
.B(n_96),
.Y(n_122)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_64),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_60),
.B(n_2),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_64),
.Y(n_97)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_97),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_54),
.Y(n_98)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_98),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_54),
.B(n_41),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_44),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_100),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_101),
.A2(n_85),
.B(n_66),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_82),
.A2(n_53),
.B1(n_57),
.B2(n_60),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_102),
.A2(n_123),
.B1(n_111),
.B2(n_77),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_104),
.B(n_121),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_73),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_108),
.B(n_128),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_109),
.B(n_84),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_114),
.A2(n_127),
.B1(n_111),
.B2(n_95),
.Y(n_142)
);

AND2x6_ASAP7_75t_L g116 ( 
.A(n_78),
.B(n_2),
.Y(n_116)
);

AND2x6_ASAP7_75t_L g136 ( 
.A(n_116),
.B(n_117),
.Y(n_136)
);

AND2x6_ASAP7_75t_L g117 ( 
.A(n_90),
.B(n_3),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_65),
.B(n_29),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_119),
.B(n_84),
.Y(n_135)
);

AND2x6_ASAP7_75t_L g121 ( 
.A(n_76),
.B(n_3),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_99),
.B(n_3),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_124),
.A2(n_72),
.B(n_88),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_68),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_129),
.A2(n_149),
.B1(n_158),
.B2(n_154),
.Y(n_178)
);

AND2x2_ASAP7_75t_SL g130 ( 
.A(n_125),
.B(n_75),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_130),
.A2(n_144),
.B(n_153),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_132),
.B(n_29),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_106),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_133),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_104),
.A2(n_80),
.B1(n_66),
.B2(n_85),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_134),
.A2(n_142),
.B1(n_143),
.B2(n_152),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_135),
.B(n_140),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_138),
.B(n_139),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_112),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_125),
.B(n_119),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_103),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_141),
.B(n_146),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_114),
.A2(n_72),
.B1(n_97),
.B2(n_100),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_102),
.B(n_88),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_145),
.B(n_106),
.C(n_115),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_122),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_118),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_147),
.B(n_157),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_128),
.B(n_88),
.Y(n_148)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_148),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_101),
.A2(n_123),
.B1(n_120),
.B2(n_121),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_120),
.B(n_98),
.Y(n_150)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_150),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_124),
.B(n_41),
.Y(n_151)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_151),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_116),
.A2(n_94),
.B1(n_81),
.B2(n_79),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_117),
.A2(n_41),
.B(n_35),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_124),
.B(n_35),
.Y(n_154)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_154),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_108),
.B(n_4),
.Y(n_155)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_155),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_113),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_156),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g157 ( 
.A(n_107),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_113),
.A2(n_35),
.B1(n_18),
.B2(n_27),
.Y(n_158)
);

MAJx2_ASAP7_75t_L g160 ( 
.A(n_132),
.B(n_109),
.C(n_126),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_160),
.B(n_5),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_157),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_163),
.B(n_144),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_134),
.A2(n_129),
.B1(n_145),
.B2(n_152),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_165),
.A2(n_130),
.B1(n_136),
.B2(n_156),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_149),
.B(n_109),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_166),
.B(n_176),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_133),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_168),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_131),
.B(n_126),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_170),
.B(n_177),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_173),
.B(n_182),
.C(n_15),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_147),
.B(n_115),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_178),
.A2(n_181),
.B1(n_186),
.B2(n_139),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_141),
.B(n_107),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_179),
.B(n_158),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_153),
.A2(n_110),
.B1(n_107),
.B2(n_18),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_137),
.B(n_105),
.C(n_110),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_150),
.A2(n_27),
.B(n_6),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_184),
.B(n_15),
.Y(n_205)
);

AO21x2_ASAP7_75t_L g186 ( 
.A1(n_156),
.A2(n_27),
.B(n_6),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_187),
.A2(n_196),
.B1(n_203),
.B2(n_204),
.Y(n_214)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_188),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_164),
.B(n_140),
.Y(n_191)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_191),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_192),
.B(n_193),
.Y(n_226)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_171),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_163),
.B(n_137),
.Y(n_194)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_194),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_162),
.B(n_151),
.Y(n_195)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_195),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_178),
.A2(n_136),
.B1(n_130),
.B2(n_135),
.Y(n_196)
);

INVxp33_ASAP7_75t_SL g197 ( 
.A(n_186),
.Y(n_197)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_197),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_164),
.B(n_167),
.Y(n_198)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_198),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_199),
.A2(n_182),
.B1(n_173),
.B2(n_174),
.Y(n_210)
);

NOR3xp33_ASAP7_75t_L g200 ( 
.A(n_184),
.B(n_5),
.C(n_7),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_200),
.B(n_201),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_172),
.B(n_5),
.Y(n_201)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_181),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_167),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_205),
.B(n_207),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_206),
.B(n_166),
.C(n_174),
.Y(n_212)
);

BUFx2_ASAP7_75t_L g208 ( 
.A(n_186),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_208),
.A2(n_209),
.B(n_186),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_175),
.B(n_8),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_210),
.A2(n_222),
.B(n_9),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_212),
.B(n_9),
.C(n_11),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_206),
.B(n_165),
.C(n_180),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_213),
.B(n_220),
.C(n_227),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_196),
.B(n_180),
.C(n_175),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_199),
.A2(n_161),
.B1(n_159),
.B2(n_186),
.Y(n_221)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_221),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_187),
.A2(n_161),
.B1(n_185),
.B2(n_160),
.Y(n_224)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_224),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_191),
.B(n_176),
.C(n_183),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_217),
.B(n_189),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_228),
.B(n_235),
.Y(n_249)
);

BUFx12f_ASAP7_75t_L g229 ( 
.A(n_223),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_229),
.Y(n_246)
);

NAND3xp33_ASAP7_75t_L g231 ( 
.A(n_219),
.B(n_209),
.C(n_207),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_231),
.B(n_218),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_222),
.A2(n_198),
.B(n_208),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_232),
.A2(n_241),
.B(n_225),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_219),
.B(n_169),
.Y(n_235)
);

MAJx2_ASAP7_75t_L g236 ( 
.A(n_210),
.B(n_202),
.C(n_205),
.Y(n_236)
);

HB1xp67_ASAP7_75t_SL g248 ( 
.A(n_236),
.Y(n_248)
);

INVx13_ASAP7_75t_L g237 ( 
.A(n_226),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_237),
.B(n_238),
.Y(n_254)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_214),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_220),
.A2(n_202),
.B1(n_190),
.B2(n_10),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_239),
.A2(n_227),
.B1(n_216),
.B2(n_212),
.Y(n_253)
);

AO22x1_ASAP7_75t_L g240 ( 
.A1(n_221),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_240)
);

AO21x1_ASAP7_75t_L g251 ( 
.A1(n_240),
.A2(n_211),
.B(n_215),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_242),
.B(n_218),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_243),
.A2(n_230),
.B(n_240),
.Y(n_259)
);

XNOR2x1_ASAP7_75t_L g244 ( 
.A(n_241),
.B(n_224),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_244),
.A2(n_245),
.B(n_239),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_247),
.B(n_252),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_233),
.B(n_213),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_250),
.B(n_233),
.Y(n_260)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_251),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_229),
.Y(n_252)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_253),
.Y(n_258)
);

AOI322xp5_ASAP7_75t_L g257 ( 
.A1(n_244),
.A2(n_230),
.A3(n_234),
.B1(n_232),
.B2(n_237),
.C1(n_229),
.C2(n_236),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_257),
.B(n_262),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_259),
.A2(n_251),
.B(n_249),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_260),
.B(n_261),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_254),
.B(n_242),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_248),
.B(n_12),
.C(n_13),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_263),
.B(n_12),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_255),
.B(n_246),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_266),
.B(n_268),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_267),
.A2(n_257),
.B(n_250),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_262),
.B(n_253),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_269),
.B(n_270),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_256),
.B(n_247),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_265),
.B(n_263),
.Y(n_272)
);

OR2x2_ASAP7_75t_L g276 ( 
.A(n_272),
.B(n_267),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_264),
.B(n_258),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_274),
.B(n_275),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_276),
.B(n_13),
.Y(n_280)
);

AO21x1_ASAP7_75t_L g278 ( 
.A1(n_271),
.A2(n_273),
.B(n_13),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_278),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_280),
.B(n_277),
.C(n_14),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_281),
.B(n_14),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_282),
.B(n_279),
.Y(n_283)
);


endmodule