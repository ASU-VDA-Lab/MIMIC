module fake_ibex_1204_n_4966 (n_151, n_85, n_599, n_778, n_822, n_507, n_743, n_540, n_754, n_395, n_84, n_64, n_171, n_756, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_766, n_688, n_130, n_177, n_946, n_707, n_76, n_273, n_309, n_330, n_926, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_845, n_947, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_956, n_790, n_920, n_452, n_86, n_70, n_664, n_255, n_175, n_586, n_773, n_638, n_398, n_59, n_28, n_125, n_304, n_821, n_191, n_873, n_593, n_5, n_62, n_71, n_153, n_862, n_545, n_909, n_583, n_887, n_957, n_678, n_663, n_194, n_249, n_334, n_634, n_733, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_872, n_423, n_608, n_864, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_930, n_336, n_258, n_861, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_727, n_58, n_43, n_216, n_915, n_911, n_33, n_652, n_781, n_421, n_828, n_738, n_475, n_802, n_166, n_163, n_753, n_645, n_500, n_747, n_542, n_114, n_236, n_900, n_34, n_376, n_377, n_584, n_531, n_647, n_15, n_761, n_556, n_748, n_24, n_189, n_498, n_698, n_280, n_317, n_340, n_375, n_708, n_901, n_105, n_187, n_667, n_884, n_1, n_154, n_682, n_850, n_182, n_196, n_326, n_327, n_879, n_89, n_50, n_723, n_144, n_170, n_270, n_346, n_383, n_113, n_886, n_840, n_561, n_883, n_117, n_417, n_471, n_846, n_739, n_755, n_265, n_853, n_504, n_948, n_158, n_859, n_259, n_276, n_339, n_470, n_770, n_210, n_348, n_220, n_875, n_941, n_674, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_671, n_228, n_711, n_876, n_147, n_552, n_251, n_384, n_632, n_373, n_854, n_458, n_244, n_73, n_343, n_310, n_714, n_936, n_703, n_426, n_323, n_469, n_829, n_598, n_825, n_143, n_740, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_939, n_67, n_453, n_591, n_898, n_655, n_333, n_928, n_110, n_306, n_400, n_47, n_550, n_736, n_169, n_10, n_673, n_21, n_732, n_798, n_832, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_641, n_7, n_109, n_127, n_121, n_527, n_893, n_590, n_465, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_690, n_914, n_120, n_835, n_168, n_526, n_785, n_155, n_824, n_929, n_315, n_441, n_604, n_13, n_637, n_122, n_523, n_116, n_694, n_787, n_614, n_370, n_431, n_719, n_574, n_0, n_289, n_716, n_865, n_923, n_12, n_515, n_642, n_150, n_286, n_321, n_133, n_569, n_600, n_907, n_51, n_933, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_669, n_838, n_750, n_746, n_22, n_136, n_261, n_742, n_521, n_665, n_459, n_30, n_518, n_367, n_221, n_852, n_789, n_880, n_654, n_656, n_724, n_437, n_731, n_602, n_904, n_842, n_938, n_355, n_767, n_474, n_878, n_758, n_594, n_636, n_710, n_720, n_407, n_102, n_490, n_568, n_813, n_52, n_448, n_646, n_595, n_99, n_466, n_269, n_944, n_156, n_570, n_126, n_623, n_585, n_715, n_791, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_769, n_222, n_660, n_186, n_524, n_349, n_765, n_849, n_857, n_454, n_777, n_295, n_730, n_331, n_576, n_230, n_96, n_759, n_917, n_185, n_388, n_953, n_625, n_619, n_536, n_611, n_352, n_290, n_558, n_931, n_666, n_174, n_467, n_427, n_607, n_827, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_922, n_438, n_851, n_689, n_793, n_167, n_676, n_128, n_937, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_771, n_205, n_618, n_488, n_139, n_514, n_705, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_659, n_267, n_662, n_910, n_635, n_844, n_245, n_589, n_571, n_229, n_209, n_472, n_648, n_783, n_347, n_847, n_830, n_473, n_445, n_629, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_359, n_826, n_299, n_87, n_262, n_433, n_75, n_439, n_704, n_949, n_924, n_643, n_137, n_679, n_841, n_772, n_810, n_768, n_839, n_338, n_173, n_696, n_796, n_797, n_837, n_477, n_640, n_954, n_363, n_402, n_725, n_180, n_369, n_596, n_201, n_699, n_14, n_351, n_368, n_456, n_834, n_257, n_77, n_935, n_869, n_925, n_718, n_801, n_918, n_44, n_672, n_722, n_401, n_553, n_554, n_66, n_735, n_305, n_882, n_942, n_713, n_307, n_192, n_804, n_140, n_484, n_566, n_480, n_416, n_581, n_651, n_365, n_721, n_4, n_814, n_955, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_630, n_516, n_548, n_567, n_943, n_763, n_745, n_329, n_447, n_940, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_868, n_546, n_199, n_788, n_795, n_592, n_495, n_762, n_410, n_905, n_308, n_675, n_800, n_463, n_624, n_706, n_411, n_135, n_520, n_784, n_684, n_775, n_927, n_934, n_658, n_512, n_615, n_950, n_685, n_283, n_366, n_397, n_111, n_803, n_894, n_692, n_36, n_627, n_18, n_709, n_322, n_53, n_227, n_499, n_115, n_888, n_757, n_11, n_248, n_92, n_702, n_451, n_712, n_101, n_190, n_906, n_138, n_650, n_776, n_409, n_582, n_818, n_653, n_214, n_238, n_579, n_843, n_899, n_902, n_332, n_799, n_517, n_211, n_744, n_817, n_218, n_314, n_691, n_563, n_132, n_277, n_555, n_337, n_522, n_700, n_479, n_534, n_225, n_360, n_881, n_272, n_951, n_511, n_23, n_734, n_468, n_223, n_381, n_525, n_815, n_919, n_780, n_535, n_382, n_502, n_681, n_633, n_532, n_726, n_95, n_405, n_863, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_819, n_161, n_237, n_29, n_203, n_268, n_440, n_858, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_729, n_741, n_603, n_378, n_486, n_952, n_422, n_164, n_38, n_198, n_264, n_616, n_782, n_833, n_217, n_324, n_391, n_831, n_537, n_728, n_78, n_805, n_670, n_820, n_20, n_69, n_892, n_390, n_544, n_891, n_913, n_39, n_178, n_509, n_695, n_786, n_639, n_303, n_362, n_717, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_680, n_501, n_809, n_752, n_856, n_668, n_779, n_871, n_266, n_42, n_294, n_112, n_485, n_870, n_46, n_284, n_811, n_808, n_80, n_172, n_250, n_945, n_493, n_460, n_609, n_476, n_792, n_461, n_575, n_313, n_903, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_774, n_72, n_319, n_195, n_885, n_513, n_212, n_588, n_877, n_693, n_311, n_860, n_661, n_848, n_406, n_606, n_737, n_896, n_97, n_197, n_528, n_181, n_131, n_123, n_631, n_683, n_260, n_620, n_794, n_836, n_462, n_302, n_450, n_443, n_686, n_572, n_867, n_644, n_577, n_344, n_393, n_889, n_897, n_436, n_428, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_697, n_816, n_874, n_890, n_912, n_921, n_83, n_32, n_107, n_149, n_489, n_677, n_399, n_254, n_908, n_213, n_424, n_565, n_916, n_823, n_701, n_271, n_241, n_68, n_503, n_292, n_807, n_394, n_79, n_81, n_35, n_364, n_687, n_895, n_159, n_202, n_231, n_298, n_587, n_760, n_751, n_806, n_932, n_160, n_657, n_764, n_184, n_56, n_492, n_649, n_812, n_855, n_232, n_380, n_749, n_281, n_866, n_559, n_425, n_4966);

input n_151;
input n_85;
input n_599;
input n_778;
input n_822;
input n_507;
input n_743;
input n_540;
input n_754;
input n_395;
input n_84;
input n_64;
input n_171;
input n_756;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_766;
input n_688;
input n_130;
input n_177;
input n_946;
input n_707;
input n_76;
input n_273;
input n_309;
input n_330;
input n_926;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_845;
input n_947;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_956;
input n_790;
input n_920;
input n_452;
input n_86;
input n_70;
input n_664;
input n_255;
input n_175;
input n_586;
input n_773;
input n_638;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_821;
input n_191;
input n_873;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_862;
input n_545;
input n_909;
input n_583;
input n_887;
input n_957;
input n_678;
input n_663;
input n_194;
input n_249;
input n_334;
input n_634;
input n_733;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_872;
input n_423;
input n_608;
input n_864;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_930;
input n_336;
input n_258;
input n_861;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_727;
input n_58;
input n_43;
input n_216;
input n_915;
input n_911;
input n_33;
input n_652;
input n_781;
input n_421;
input n_828;
input n_738;
input n_475;
input n_802;
input n_166;
input n_163;
input n_753;
input n_645;
input n_500;
input n_747;
input n_542;
input n_114;
input n_236;
input n_900;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_647;
input n_15;
input n_761;
input n_556;
input n_748;
input n_24;
input n_189;
input n_498;
input n_698;
input n_280;
input n_317;
input n_340;
input n_375;
input n_708;
input n_901;
input n_105;
input n_187;
input n_667;
input n_884;
input n_1;
input n_154;
input n_682;
input n_850;
input n_182;
input n_196;
input n_326;
input n_327;
input n_879;
input n_89;
input n_50;
input n_723;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_886;
input n_840;
input n_561;
input n_883;
input n_117;
input n_417;
input n_471;
input n_846;
input n_739;
input n_755;
input n_265;
input n_853;
input n_504;
input n_948;
input n_158;
input n_859;
input n_259;
input n_276;
input n_339;
input n_470;
input n_770;
input n_210;
input n_348;
input n_220;
input n_875;
input n_941;
input n_674;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_671;
input n_228;
input n_711;
input n_876;
input n_147;
input n_552;
input n_251;
input n_384;
input n_632;
input n_373;
input n_854;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_714;
input n_936;
input n_703;
input n_426;
input n_323;
input n_469;
input n_829;
input n_598;
input n_825;
input n_143;
input n_740;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_939;
input n_67;
input n_453;
input n_591;
input n_898;
input n_655;
input n_333;
input n_928;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_736;
input n_169;
input n_10;
input n_673;
input n_21;
input n_732;
input n_798;
input n_832;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_641;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_893;
input n_590;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_690;
input n_914;
input n_120;
input n_835;
input n_168;
input n_526;
input n_785;
input n_155;
input n_824;
input n_929;
input n_315;
input n_441;
input n_604;
input n_13;
input n_637;
input n_122;
input n_523;
input n_116;
input n_694;
input n_787;
input n_614;
input n_370;
input n_431;
input n_719;
input n_574;
input n_0;
input n_289;
input n_716;
input n_865;
input n_923;
input n_12;
input n_515;
input n_642;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_907;
input n_51;
input n_933;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_669;
input n_838;
input n_750;
input n_746;
input n_22;
input n_136;
input n_261;
input n_742;
input n_521;
input n_665;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_852;
input n_789;
input n_880;
input n_654;
input n_656;
input n_724;
input n_437;
input n_731;
input n_602;
input n_904;
input n_842;
input n_938;
input n_355;
input n_767;
input n_474;
input n_878;
input n_758;
input n_594;
input n_636;
input n_710;
input n_720;
input n_407;
input n_102;
input n_490;
input n_568;
input n_813;
input n_52;
input n_448;
input n_646;
input n_595;
input n_99;
input n_466;
input n_269;
input n_944;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_715;
input n_791;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_769;
input n_222;
input n_660;
input n_186;
input n_524;
input n_349;
input n_765;
input n_849;
input n_857;
input n_454;
input n_777;
input n_295;
input n_730;
input n_331;
input n_576;
input n_230;
input n_96;
input n_759;
input n_917;
input n_185;
input n_388;
input n_953;
input n_625;
input n_619;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_931;
input n_666;
input n_174;
input n_467;
input n_427;
input n_607;
input n_827;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_922;
input n_438;
input n_851;
input n_689;
input n_793;
input n_167;
input n_676;
input n_128;
input n_937;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_771;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_705;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_659;
input n_267;
input n_662;
input n_910;
input n_635;
input n_844;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_648;
input n_783;
input n_347;
input n_847;
input n_830;
input n_473;
input n_445;
input n_629;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_359;
input n_826;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_704;
input n_949;
input n_924;
input n_643;
input n_137;
input n_679;
input n_841;
input n_772;
input n_810;
input n_768;
input n_839;
input n_338;
input n_173;
input n_696;
input n_796;
input n_797;
input n_837;
input n_477;
input n_640;
input n_954;
input n_363;
input n_402;
input n_725;
input n_180;
input n_369;
input n_596;
input n_201;
input n_699;
input n_14;
input n_351;
input n_368;
input n_456;
input n_834;
input n_257;
input n_77;
input n_935;
input n_869;
input n_925;
input n_718;
input n_801;
input n_918;
input n_44;
input n_672;
input n_722;
input n_401;
input n_553;
input n_554;
input n_66;
input n_735;
input n_305;
input n_882;
input n_942;
input n_713;
input n_307;
input n_192;
input n_804;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_651;
input n_365;
input n_721;
input n_4;
input n_814;
input n_955;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_630;
input n_516;
input n_548;
input n_567;
input n_943;
input n_763;
input n_745;
input n_329;
input n_447;
input n_940;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_868;
input n_546;
input n_199;
input n_788;
input n_795;
input n_592;
input n_495;
input n_762;
input n_410;
input n_905;
input n_308;
input n_675;
input n_800;
input n_463;
input n_624;
input n_706;
input n_411;
input n_135;
input n_520;
input n_784;
input n_684;
input n_775;
input n_927;
input n_934;
input n_658;
input n_512;
input n_615;
input n_950;
input n_685;
input n_283;
input n_366;
input n_397;
input n_111;
input n_803;
input n_894;
input n_692;
input n_36;
input n_627;
input n_18;
input n_709;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_888;
input n_757;
input n_11;
input n_248;
input n_92;
input n_702;
input n_451;
input n_712;
input n_101;
input n_190;
input n_906;
input n_138;
input n_650;
input n_776;
input n_409;
input n_582;
input n_818;
input n_653;
input n_214;
input n_238;
input n_579;
input n_843;
input n_899;
input n_902;
input n_332;
input n_799;
input n_517;
input n_211;
input n_744;
input n_817;
input n_218;
input n_314;
input n_691;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_700;
input n_479;
input n_534;
input n_225;
input n_360;
input n_881;
input n_272;
input n_951;
input n_511;
input n_23;
input n_734;
input n_468;
input n_223;
input n_381;
input n_525;
input n_815;
input n_919;
input n_780;
input n_535;
input n_382;
input n_502;
input n_681;
input n_633;
input n_532;
input n_726;
input n_95;
input n_405;
input n_863;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_819;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_858;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_729;
input n_741;
input n_603;
input n_378;
input n_486;
input n_952;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_782;
input n_833;
input n_217;
input n_324;
input n_391;
input n_831;
input n_537;
input n_728;
input n_78;
input n_805;
input n_670;
input n_820;
input n_20;
input n_69;
input n_892;
input n_390;
input n_544;
input n_891;
input n_913;
input n_39;
input n_178;
input n_509;
input n_695;
input n_786;
input n_639;
input n_303;
input n_362;
input n_717;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_680;
input n_501;
input n_809;
input n_752;
input n_856;
input n_668;
input n_779;
input n_871;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_870;
input n_46;
input n_284;
input n_811;
input n_808;
input n_80;
input n_172;
input n_250;
input n_945;
input n_493;
input n_460;
input n_609;
input n_476;
input n_792;
input n_461;
input n_575;
input n_313;
input n_903;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_774;
input n_72;
input n_319;
input n_195;
input n_885;
input n_513;
input n_212;
input n_588;
input n_877;
input n_693;
input n_311;
input n_860;
input n_661;
input n_848;
input n_406;
input n_606;
input n_737;
input n_896;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_631;
input n_683;
input n_260;
input n_620;
input n_794;
input n_836;
input n_462;
input n_302;
input n_450;
input n_443;
input n_686;
input n_572;
input n_867;
input n_644;
input n_577;
input n_344;
input n_393;
input n_889;
input n_897;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_697;
input n_816;
input n_874;
input n_890;
input n_912;
input n_921;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_677;
input n_399;
input n_254;
input n_908;
input n_213;
input n_424;
input n_565;
input n_916;
input n_823;
input n_701;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_807;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_687;
input n_895;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_760;
input n_751;
input n_806;
input n_932;
input n_160;
input n_657;
input n_764;
input n_184;
input n_56;
input n_492;
input n_649;
input n_812;
input n_855;
input n_232;
input n_380;
input n_749;
input n_281;
input n_866;
input n_559;
input n_425;

output n_4966;

wire n_4557;
wire n_3590;
wire n_4056;
wire n_2960;
wire n_3548;
wire n_1382;
wire n_2949;
wire n_2840;
wire n_3319;
wire n_3915;
wire n_4204;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_1802;
wire n_3817;
wire n_2038;
wire n_2504;
wire n_962;
wire n_4607;
wire n_4514;
wire n_3674;
wire n_4249;
wire n_4931;
wire n_1859;
wire n_4805;
wire n_1034;
wire n_1765;
wire n_2392;
wire n_3280;
wire n_4371;
wire n_4601;
wire n_3458;
wire n_3519;
wire n_2276;
wire n_1782;
wire n_2889;
wire n_2391;
wire n_4585;
wire n_1391;
wire n_3338;
wire n_3168;
wire n_2396;
wire n_3440;
wire n_4169;
wire n_3570;
wire n_4875;
wire n_1957;
wire n_4197;
wire n_2188;
wire n_1144;
wire n_2506;
wire n_3598;
wire n_1752;
wire n_4172;
wire n_1730;
wire n_3479;
wire n_3751;
wire n_3262;
wire n_4673;
wire n_3537;
wire n_2343;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_4781;
wire n_4423;
wire n_1766;
wire n_4065;
wire n_3469;
wire n_3170;
wire n_1922;
wire n_3347;
wire n_3395;
wire n_4808;
wire n_4507;
wire n_3577;
wire n_2995;
wire n_4526;
wire n_3472;
wire n_1981;
wire n_3976;
wire n_4348;
wire n_3807;
wire n_2998;
wire n_3845;
wire n_2163;
wire n_4450;
wire n_4467;
wire n_4801;
wire n_3639;
wire n_1664;
wire n_4144;
wire n_3298;
wire n_1427;
wire n_4447;
wire n_4955;
wire n_3208;
wire n_4569;
wire n_3671;
wire n_1778;
wire n_2839;
wire n_1698;
wire n_1496;
wire n_2333;
wire n_2705;
wire n_1214;
wire n_1274;
wire n_1595;
wire n_1070;
wire n_4510;
wire n_4567;
wire n_2362;
wire n_968;
wire n_2822;
wire n_1306;
wire n_1493;
wire n_2597;
wire n_2774;
wire n_3681;
wire n_2753;
wire n_3603;
wire n_1960;
wire n_3979;
wire n_3714;
wire n_2844;
wire n_3565;
wire n_3883;
wire n_3943;
wire n_4563;
wire n_1309;
wire n_1316;
wire n_1562;
wire n_4854;
wire n_3769;
wire n_1445;
wire n_2147;
wire n_2253;
wire n_4479;
wire n_3858;
wire n_4173;
wire n_1078;
wire n_4422;
wire n_1865;
wire n_4786;
wire n_4842;
wire n_1170;
wire n_3842;
wire n_2980;
wire n_1322;
wire n_4457;
wire n_4060;
wire n_1305;
wire n_2088;
wire n_1248;
wire n_2171;
wire n_3307;
wire n_1388;
wire n_3780;
wire n_1653;
wire n_1375;
wire n_1118;
wire n_1881;
wire n_3798;
wire n_4809;
wire n_3060;
wire n_4124;
wire n_971;
wire n_4499;
wire n_1350;
wire n_3627;
wire n_2957;
wire n_2586;
wire n_3958;
wire n_1093;
wire n_2412;
wire n_2783;
wire n_3293;
wire n_2550;
wire n_3381;
wire n_2750;
wire n_1650;
wire n_1453;
wire n_1108;
wire n_1423;
wire n_3836;
wire n_1239;
wire n_4714;
wire n_1209;
wire n_3732;
wire n_3295;
wire n_3199;
wire n_1616;
wire n_2389;
wire n_2107;
wire n_3435;
wire n_4828;
wire n_4480;
wire n_1613;
wire n_3874;
wire n_2782;
wire n_4258;
wire n_4290;
wire n_1549;
wire n_1531;
wire n_2919;
wire n_4577;
wire n_1424;
wire n_2444;
wire n_2625;
wire n_3652;
wire n_4913;
wire n_2199;
wire n_1610;
wire n_4398;
wire n_1298;
wire n_1844;
wire n_4055;
wire n_3194;
wire n_4692;
wire n_2431;
wire n_2084;
wire n_1243;
wire n_3572;
wire n_1121;
wire n_4823;
wire n_3951;
wire n_4927;
wire n_3355;
wire n_2019;
wire n_1407;
wire n_4680;
wire n_1821;
wire n_4757;
wire n_3698;
wire n_2731;
wire n_4451;
wire n_4653;
wire n_3466;
wire n_3370;
wire n_1504;
wire n_1781;
wire n_4331;
wire n_2028;
wire n_3678;
wire n_4216;
wire n_2856;
wire n_1921;
wire n_1293;
wire n_3968;
wire n_4825;
wire n_3950;
wire n_1042;
wire n_1319;
wire n_4376;
wire n_4050;
wire n_4623;
wire n_1041;
wire n_4523;
wire n_4411;
wire n_3811;
wire n_1271;
wire n_3416;
wire n_3147;
wire n_3628;
wire n_3983;
wire n_2425;
wire n_2800;
wire n_4225;
wire n_3859;
wire n_4489;
wire n_3455;
wire n_1591;
wire n_2289;
wire n_2841;
wire n_4271;
wire n_1409;
wire n_1015;
wire n_2744;
wire n_3524;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_4404;
wire n_1521;
wire n_3054;
wire n_2456;
wire n_2924;
wire n_2264;
wire n_1987;
wire n_1129;
wire n_1244;
wire n_3365;
wire n_4725;
wire n_1932;
wire n_3775;
wire n_3741;
wire n_3854;
wire n_1217;
wire n_4658;
wire n_2655;
wire n_3487;
wire n_1715;
wire n_3300;
wire n_1713;
wire n_3621;
wire n_2036;
wire n_1255;
wire n_2740;
wire n_2622;
wire n_4250;
wire n_1218;
wire n_4572;
wire n_4374;
wire n_3708;
wire n_2626;
wire n_1446;
wire n_3218;
wire n_2880;
wire n_2423;
wire n_3849;
wire n_3490;
wire n_3055;
wire n_1633;
wire n_4469;
wire n_2580;
wire n_3222;
wire n_3529;
wire n_3352;
wire n_1051;
wire n_4180;
wire n_1008;
wire n_2964;
wire n_4062;
wire n_1498;
wire n_1207;
wire n_1735;
wire n_1032;
wire n_3813;
wire n_1825;
wire n_4232;
wire n_4199;
wire n_1210;
wire n_4033;
wire n_2522;
wire n_4608;
wire n_1201;
wire n_1246;
wire n_4231;
wire n_1724;
wire n_2838;
wire n_1540;
wire n_3243;
wire n_3214;
wire n_1890;
wire n_3128;
wire n_4073;
wire n_2549;
wire n_4325;
wire n_2440;
wire n_4113;
wire n_1440;
wire n_4646;
wire n_1751;
wire n_2146;
wire n_2341;
wire n_1737;
wire n_4819;
wire n_4261;
wire n_4884;
wire n_1083;
wire n_3205;
wire n_4490;
wire n_2358;
wire n_2361;
wire n_4128;
wire n_2062;
wire n_3932;
wire n_2339;
wire n_1963;
wire n_1418;
wire n_1137;
wire n_2552;
wire n_3119;
wire n_2590;
wire n_1977;
wire n_3345;
wire n_4114;
wire n_1776;
wire n_3544;
wire n_1279;
wire n_4209;
wire n_3692;
wire n_1064;
wire n_1408;
wire n_3913;
wire n_3535;
wire n_2287;
wire n_3597;
wire n_4190;
wire n_2954;
wire n_2046;
wire n_4443;
wire n_4151;
wire n_4625;
wire n_4170;
wire n_4424;
wire n_1465;
wire n_4674;
wire n_1232;
wire n_2715;
wire n_4679;
wire n_1345;
wire n_4456;
wire n_1590;
wire n_2133;
wire n_3553;
wire n_1471;
wire n_3441;
wire n_4559;
wire n_2551;
wire n_4641;
wire n_4064;
wire n_4110;
wire n_4379;
wire n_3397;
wire n_4145;
wire n_1627;
wire n_3880;
wire n_4664;
wire n_3829;
wire n_1864;
wire n_2010;
wire n_2733;
wire n_3796;
wire n_1836;
wire n_4753;
wire n_1420;
wire n_2651;
wire n_1699;
wire n_4894;
wire n_4115;
wire n_2905;
wire n_3460;
wire n_3978;
wire n_3954;
wire n_4321;
wire n_2418;
wire n_1087;
wire n_1599;
wire n_3070;
wire n_3477;
wire n_1575;
wire n_4416;
wire n_4024;
wire n_3975;
wire n_3164;
wire n_1448;
wire n_3034;
wire n_2628;
wire n_4361;
wire n_1705;
wire n_4237;
wire n_2263;
wire n_3495;
wire n_3169;
wire n_3759;
wire n_4777;
wire n_4800;
wire n_3629;
wire n_4117;
wire n_2884;
wire n_3383;
wire n_3687;
wire n_4154;
wire n_3459;
wire n_2691;
wire n_2243;
wire n_3092;
wire n_4385;
wire n_2759;
wire n_3434;
wire n_2654;
wire n_2975;
wire n_2503;
wire n_4072;
wire n_1512;
wire n_4908;
wire n_3885;
wire n_1426;
wire n_2365;
wire n_2245;
wire n_3877;
wire n_3260;
wire n_2776;
wire n_2630;
wire n_1967;
wire n_1095;
wire n_3834;
wire n_1378;
wire n_3257;
wire n_2459;
wire n_2439;
wire n_1430;
wire n_2450;
wire n_4195;
wire n_1475;
wire n_3337;
wire n_4851;
wire n_4963;
wire n_1122;
wire n_3387;
wire n_4495;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_1514;
wire n_2728;
wire n_4685;
wire n_3428;
wire n_2427;
wire n_1127;
wire n_1004;
wire n_1845;
wire n_3835;
wire n_3723;
wire n_3389;
wire n_2422;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1578;
wire n_2712;
wire n_972;
wire n_4314;
wire n_2788;
wire n_2089;
wire n_1857;
wire n_1997;
wire n_3314;
wire n_1349;
wire n_3891;
wire n_4704;
wire n_1777;
wire n_3409;
wire n_1546;
wire n_4003;
wire n_4775;
wire n_3420;
wire n_4192;
wire n_4633;
wire n_1950;
wire n_4593;
wire n_3914;
wire n_3289;
wire n_1834;
wire n_3372;
wire n_4121;
wire n_2862;
wire n_3850;
wire n_4488;
wire n_3405;
wire n_1657;
wire n_1741;
wire n_4264;
wire n_4183;
wire n_4118;
wire n_4302;
wire n_2138;
wire n_4916;
wire n_4858;
wire n_1914;
wire n_3833;
wire n_3339;
wire n_3673;
wire n_2620;
wire n_1826;
wire n_1855;
wire n_4241;
wire n_3556;
wire n_1340;
wire n_2562;
wire n_3269;
wire n_2223;
wire n_3876;
wire n_1267;
wire n_2683;
wire n_3432;
wire n_1816;
wire n_4645;
wire n_4619;
wire n_2318;
wire n_2141;
wire n_1422;
wire n_4339;
wire n_4085;
wire n_3190;
wire n_1055;
wire n_3878;
wire n_4661;
wire n_2947;
wire n_4080;
wire n_1754;
wire n_3686;
wire n_1025;
wire n_2679;
wire n_4028;
wire n_1517;
wire n_3670;
wire n_3002;
wire n_2087;
wire n_2920;
wire n_4289;
wire n_977;
wire n_1895;
wire n_1860;
wire n_1763;
wire n_3912;
wire n_1607;
wire n_2959;
wire n_2420;
wire n_2380;
wire n_3265;
wire n_2221;
wire n_1774;
wire n_2516;
wire n_2031;
wire n_1348;
wire n_1021;
wire n_1191;
wire n_4099;
wire n_3899;
wire n_4729;
wire n_1617;
wire n_2639;
wire n_3099;
wire n_1001;
wire n_4745;
wire n_4057;
wire n_2410;
wire n_3206;
wire n_2633;
wire n_1017;
wire n_2049;
wire n_2113;
wire n_1690;
wire n_4466;
wire n_4132;
wire n_3361;
wire n_4603;
wire n_1135;
wire n_4300;
wire n_3277;
wire n_2758;
wire n_4417;
wire n_1550;
wire n_1169;
wire n_1938;
wire n_3452;
wire n_4022;
wire n_1072;
wire n_2194;
wire n_4320;
wire n_1173;
wire n_2736;
wire n_2845;
wire n_3886;
wire n_1901;
wire n_3096;
wire n_2059;
wire n_1278;
wire n_4730;
wire n_4616;
wire n_4760;
wire n_1710;
wire n_3021;
wire n_1603;
wire n_3404;
wire n_2072;
wire n_2963;
wire n_1489;
wire n_1993;
wire n_4859;
wire n_1455;
wire n_2182;
wire n_3115;
wire n_1057;
wire n_4583;
wire n_1502;
wire n_4923;
wire n_3920;
wire n_4082;
wire n_3273;
wire n_4367;
wire n_4282;
wire n_4475;
wire n_2286;
wire n_2563;
wire n_4893;
wire n_3650;
wire n_3513;
wire n_2677;
wire n_2531;
wire n_4029;
wire n_3212;
wire n_1321;
wire n_1779;
wire n_2489;
wire n_2950;
wire n_2272;
wire n_3574;
wire n_2608;
wire n_3739;
wire n_2825;
wire n_4338;
wire n_2742;
wire n_3604;
wire n_1740;
wire n_3540;
wire n_2680;
wire n_1343;
wire n_1371;
wire n_4198;
wire n_4529;
wire n_2861;
wire n_2976;
wire n_2366;
wire n_4919;
wire n_4200;
wire n_4111;
wire n_1659;
wire n_4575;
wire n_4847;
wire n_4803;
wire n_1047;
wire n_1878;
wire n_1374;
wire n_2851;
wire n_2973;
wire n_3651;
wire n_4666;
wire n_1242;
wire n_2810;
wire n_1119;
wire n_3027;
wire n_4189;
wire n_4076;
wire n_3438;
wire n_4835;
wire n_3464;
wire n_4390;
wire n_4722;
wire n_1530;
wire n_3215;
wire n_2871;
wire n_2764;
wire n_3648;
wire n_3234;
wire n_4058;
wire n_985;
wire n_4611;
wire n_2714;
wire n_2669;
wire n_4081;
wire n_4391;
wire n_1459;
wire n_4032;
wire n_2232;
wire n_4541;
wire n_4530;
wire n_1570;
wire n_995;
wire n_1303;
wire n_1994;
wire n_1526;
wire n_4268;
wire n_2367;
wire n_3236;
wire n_1961;
wire n_3013;
wire n_4265;
wire n_1050;
wire n_3062;
wire n_3806;
wire n_3256;
wire n_3126;
wire n_1257;
wire n_2864;
wire n_1632;
wire n_3104;
wire n_4895;
wire n_3354;
wire n_4069;
wire n_3373;
wire n_2784;
wire n_4140;
wire n_1909;
wire n_4125;
wire n_2495;
wire n_4531;
wire n_4778;
wire n_4789;
wire n_2703;
wire n_2574;
wire n_1887;
wire n_3504;
wire n_3511;
wire n_2428;
wire n_3159;
wire n_1768;
wire n_3697;
wire n_2068;
wire n_2636;
wire n_3101;
wire n_2364;
wire n_2641;
wire n_1077;
wire n_4751;
wire n_3774;
wire n_2494;
wire n_3863;
wire n_2228;
wire n_4474;
wire n_1518;
wire n_4350;
wire n_4478;
wire n_2872;
wire n_2411;
wire n_3539;
wire n_1061;
wire n_2266;
wire n_4473;
wire n_3761;
wire n_2830;
wire n_4675;
wire n_3083;
wire n_1010;
wire n_3844;
wire n_4049;
wire n_2044;
wire n_2091;
wire n_4945;
wire n_3362;
wire n_3035;
wire n_4165;
wire n_4891;
wire n_2394;
wire n_1572;
wire n_1245;
wire n_4867;
wire n_2929;
wire n_4911;
wire n_1329;
wire n_2409;
wire n_2405;
wire n_2601;
wire n_4405;
wire n_3118;
wire n_3742;
wire n_3532;
wire n_4686;
wire n_4682;
wire n_2914;
wire n_1833;
wire n_1986;
wire n_2882;
wire n_4301;
wire n_2493;
wire n_2115;
wire n_2013;
wire n_1556;
wire n_3547;
wire n_4898;
wire n_3700;
wire n_4733;
wire n_987;
wire n_3947;
wire n_4684;
wire n_3663;
wire n_2129;
wire n_3230;
wire n_2532;
wire n_3782;
wire n_1720;
wire n_3831;
wire n_2293;
wire n_3068;
wire n_3071;
wire n_3683;
wire n_3919;
wire n_2734;
wire n_1166;
wire n_2310;
wire n_2674;
wire n_1284;
wire n_2689;
wire n_1992;
wire n_4493;
wire n_4797;
wire n_1082;
wire n_4962;
wire n_2596;
wire n_1488;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_3606;
wire n_1866;
wire n_2169;
wire n_2111;
wire n_1262;
wire n_4644;
wire n_1012;
wire n_960;
wire n_4412;
wire n_4266;
wire n_2982;
wire n_3124;
wire n_2634;
wire n_3015;
wire n_3321;
wire n_3081;
wire n_4639;
wire n_2291;
wire n_4102;
wire n_3612;
wire n_2172;
wire n_1728;
wire n_1230;
wire n_3622;
wire n_3857;
wire n_2357;
wire n_4354;
wire n_2937;
wire n_3728;
wire n_4401;
wire n_4727;
wire n_4296;
wire n_2967;
wire n_3005;
wire n_4627;
wire n_4309;
wire n_4027;
wire n_2056;
wire n_2054;
wire n_2226;
wire n_1402;
wire n_3267;
wire n_3008;
wire n_2802;
wire n_4728;
wire n_2279;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_4046;
wire n_2961;
wire n_3689;
wire n_4631;
wire n_3283;
wire n_1736;
wire n_2907;
wire n_1948;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1033;
wire n_990;
wire n_3675;
wire n_2378;
wire n_2749;
wire n_3658;
wire n_4901;
wire n_3133;
wire n_3527;
wire n_2014;
wire n_3901;
wire n_4539;
wire n_1205;
wire n_2969;
wire n_3550;
wire n_3287;
wire n_3534;
wire n_1837;
wire n_1414;
wire n_1002;
wire n_2195;
wire n_2940;
wire n_4150;
wire n_3275;
wire n_2645;
wire n_1714;
wire n_1958;
wire n_1611;
wire n_1675;
wire n_1551;
wire n_1533;
wire n_3792;
wire n_2515;
wire n_3089;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_3406;
wire n_3988;
wire n_3758;
wire n_2353;
wire n_4106;
wire n_4251;
wire n_3662;
wire n_1354;
wire n_3329;
wire n_1277;
wire n_3233;
wire n_3193;
wire n_2582;
wire n_3789;
wire n_2174;
wire n_2510;
wire n_2435;
wire n_3934;
wire n_2583;
wire n_1678;
wire n_4606;
wire n_1287;
wire n_1525;
wire n_1150;
wire n_1674;
wire n_3980;
wire n_2912;
wire n_2710;
wire n_2970;
wire n_1393;
wire n_4691;
wire n_984;
wire n_2978;
wire n_3502;
wire n_3935;
wire n_1854;
wire n_1084;
wire n_2804;
wire n_4926;
wire n_4688;
wire n_3144;
wire n_4234;
wire n_4146;
wire n_2835;
wire n_4656;
wire n_4932;
wire n_1930;
wire n_1234;
wire n_4881;
wire n_3755;
wire n_1469;
wire n_4632;
wire n_3255;
wire n_1652;
wire n_969;
wire n_2183;
wire n_1883;
wire n_2037;
wire n_4550;
wire n_1226;
wire n_4651;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2682;
wire n_3605;
wire n_3105;
wire n_3146;
wire n_4892;
wire n_4343;
wire n_3931;
wire n_4421;
wire n_2322;
wire n_3025;
wire n_3411;
wire n_2955;
wire n_1045;
wire n_3235;
wire n_2989;
wire n_1856;
wire n_3843;
wire n_2847;
wire n_4399;
wire n_1308;
wire n_3904;
wire n_4378;
wire n_3729;
wire n_3484;
wire n_2485;
wire n_4477;
wire n_2179;
wire n_4654;
wire n_3984;
wire n_4233;
wire n_4765;
wire n_3086;
wire n_2475;
wire n_3721;
wire n_3726;
wire n_4277;
wire n_4431;
wire n_4771;
wire n_4652;
wire n_3804;
wire n_1908;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_4285;
wire n_4928;
wire n_3251;
wire n_2921;
wire n_3724;
wire n_3192;
wire n_3753;
wire n_3566;
wire n_2820;
wire n_2311;
wire n_4403;
wire n_3242;
wire n_1654;
wire n_3330;
wire n_2707;
wire n_4746;
wire n_4382;
wire n_4002;
wire n_3631;
wire n_2537;
wire n_1130;
wire n_4246;
wire n_2643;
wire n_4545;
wire n_2336;
wire n_3987;
wire n_3969;
wire n_1081;
wire n_4437;
wire n_3856;
wire n_1155;
wire n_1292;
wire n_2432;
wire n_3043;
wire n_2273;
wire n_4491;
wire n_4672;
wire n_2421;
wire n_3237;
wire n_1970;
wire n_3946;
wire n_2953;
wire n_3949;
wire n_3507;
wire n_3926;
wire n_3688;
wire n_1094;
wire n_2462;
wire n_2436;
wire n_1663;
wire n_4267;
wire n_4723;
wire n_2269;
wire n_2472;
wire n_2846;
wire n_3699;
wire n_4312;
wire n_2249;
wire n_3022;
wire n_4014;
wire n_3766;
wire n_3707;
wire n_4217;
wire n_3973;
wire n_4769;
wire n_4724;
wire n_2260;
wire n_4721;
wire n_1071;
wire n_2663;
wire n_3882;
wire n_2595;
wire n_4433;
wire n_3030;
wire n_4503;
wire n_3917;
wire n_3679;
wire n_4517;
wire n_3221;
wire n_3210;
wire n_4511;
wire n_1672;
wire n_4171;
wire n_3764;
wire n_3795;
wire n_4788;
wire n_4754;
wire n_1817;
wire n_1301;
wire n_4166;
wire n_2242;
wire n_4845;
wire n_1561;
wire n_2247;
wire n_3177;
wire n_3399;
wire n_4850;
wire n_1869;
wire n_2189;
wire n_2482;
wire n_3799;
wire n_3676;
wire n_1753;
wire n_4610;
wire n_4067;
wire n_4393;
wire n_3777;
wire n_4553;
wire n_3961;
wire n_1520;
wire n_2509;
wire n_4283;
wire n_4174;
wire n_4870;
wire n_2399;
wire n_1370;
wire n_1708;
wire n_3038;
wire n_4804;
wire n_3716;
wire n_1649;
wire n_3450;
wire n_4518;
wire n_4732;
wire n_1936;
wire n_1717;
wire n_2257;
wire n_4856;
wire n_1467;
wire n_3217;
wire n_2511;
wire n_3909;
wire n_3971;
wire n_1332;
wire n_2661;
wire n_4079;
wire n_3573;
wire n_3563;
wire n_3510;
wire n_4248;
wire n_2334;
wire n_2350;
wire n_1709;
wire n_2649;
wire n_3607;
wire n_4476;
wire n_3241;
wire n_2746;
wire n_2256;
wire n_2445;
wire n_1980;
wire n_3583;
wire n_3832;
wire n_4649;
wire n_3508;
wire n_1862;
wire n_4693;
wire n_3415;
wire n_2355;
wire n_1543;
wire n_3386;
wire n_4568;
wire n_4359;
wire n_3814;
wire n_1441;
wire n_4573;
wire n_4105;
wire n_4206;
wire n_4177;
wire n_1888;
wire n_3320;
wire n_1786;
wire n_2033;
wire n_4700;
wire n_2828;
wire n_1964;
wire n_3720;
wire n_1196;
wire n_1182;
wire n_4074;
wire n_3633;
wire n_1731;
wire n_2879;
wire n_3514;
wire n_3091;
wire n_4037;
wire n_4582;
wire n_3426;
wire n_4308;
wire n_2288;
wire n_3075;
wire n_1671;
wire n_3448;
wire n_3788;
wire n_2076;
wire n_974;
wire n_3733;
wire n_1831;
wire n_4853;
wire n_959;
wire n_1312;
wire n_3684;
wire n_1318;
wire n_4006;
wire n_1508;
wire n_3970;
wire n_3291;
wire n_2454;
wire n_4008;
wire n_2829;
wire n_2968;
wire n_4494;
wire n_3473;
wire n_3263;
wire n_4501;
wire n_1772;
wire n_2858;
wire n_1283;
wire n_1421;
wire n_4922;
wire n_2424;
wire n_1793;
wire n_2573;
wire n_2390;
wire n_965;
wire n_4402;
wire n_2793;
wire n_4813;
wire n_3098;
wire n_1711;
wire n_3069;
wire n_3107;
wire n_4134;
wire n_4131;
wire n_4330;
wire n_1053;
wire n_2176;
wire n_2805;
wire n_2319;
wire n_3757;
wire n_1933;
wire n_1842;
wire n_3364;
wire n_3429;
wire n_3306;
wire n_3787;
wire n_3445;
wire n_2080;
wire n_2554;
wire n_1676;
wire n_1013;
wire n_1136;
wire n_1918;
wire n_3642;
wire n_2461;
wire n_1229;
wire n_1490;
wire n_1179;
wire n_4818;
wire n_4462;
wire n_1153;
wire n_2787;
wire n_4540;
wire n_4187;
wire n_1273;
wire n_3821;
wire n_2930;
wire n_2616;
wire n_1014;
wire n_3503;
wire n_2441;
wire n_4063;
wire n_4362;
wire n_3312;
wire n_1848;
wire n_4009;
wire n_2650;
wire n_2888;
wire n_3614;
wire n_3394;
wire n_2530;
wire n_2792;
wire n_2372;
wire n_4191;
wire n_4965;
wire n_1522;
wire n_2523;
wire n_3488;
wire n_2832;
wire n_1028;
wire n_4525;
wire n_4011;
wire n_3526;
wire n_2142;
wire n_3703;
wire n_4554;
wire n_1260;
wire n_4097;
wire n_4861;
wire n_3239;
wire n_2600;
wire n_1069;
wire n_3952;
wire n_1171;
wire n_1126;
wire n_4596;
wire n_2434;
wire n_3578;
wire n_4734;
wire n_4492;
wire n_3470;
wire n_1738;
wire n_998;
wire n_1729;
wire n_2094;
wire n_1479;
wire n_2306;
wire n_4579;
wire n_2568;
wire n_2629;
wire n_3587;
wire n_4936;
wire n_2097;
wire n_2109;
wire n_2648;
wire n_2398;
wire n_1593;
wire n_986;
wire n_1775;
wire n_2570;
wire n_4025;
wire n_2184;
wire n_3948;
wire n_2842;
wire n_1400;
wire n_2469;
wire n_3074;
wire n_4640;
wire n_3136;
wire n_3108;
wire n_2395;
wire n_4059;
wire n_4130;
wire n_2752;
wire n_2124;
wire n_3991;
wire n_3974;
wire n_4642;
wire n_3625;
wire n_1746;
wire n_2716;
wire n_2212;
wire n_4878;
wire n_3718;
wire n_1832;
wire n_1128;
wire n_2376;
wire n_3398;
wire n_2170;
wire n_4904;
wire n_1785;
wire n_3999;
wire n_1405;
wire n_4087;
wire n_997;
wire n_3238;
wire n_4318;
wire n_3731;
wire n_3555;
wire n_3254;
wire n_4717;
wire n_4052;
wire n_2463;
wire n_2478;
wire n_3178;
wire n_4245;
wire n_3378;
wire n_3350;
wire n_4873;
wire n_3936;
wire n_1560;
wire n_3166;
wire n_3953;
wire n_3385;
wire n_1265;
wire n_2488;
wire n_2042;
wire n_1925;
wire n_1251;
wire n_3090;
wire n_1247;
wire n_3816;
wire n_4636;
wire n_4256;
wire n_1185;
wire n_3575;
wire n_2765;
wire n_4278;
wire n_4609;
wire n_4822;
wire n_2936;
wire n_2985;
wire n_3106;
wire n_4030;
wire n_4276;
wire n_4612;
wire n_1148;
wire n_1667;
wire n_1011;
wire n_3902;
wire n_1707;
wire n_4203;
wire n_2055;
wire n_4866;
wire n_2385;
wire n_3864;
wire n_3026;
wire n_3294;
wire n_4831;
wire n_1143;
wire n_2584;
wire n_4381;
wire n_2442;
wire n_1067;
wire n_4441;
wire n_2000;
wire n_4083;
wire n_2696;
wire n_4960;
wire n_1894;
wire n_2904;
wire n_3064;
wire n_2896;
wire n_4228;
wire n_4699;
wire n_1331;
wire n_1223;
wire n_1739;
wire n_3130;
wire n_1353;
wire n_2386;
wire n_3324;
wire n_3073;
wire n_2029;
wire n_4254;
wire n_4536;
wire n_1320;
wire n_4247;
wire n_4071;
wire n_2238;
wire n_4924;
wire n_4138;
wire n_3100;
wire n_1727;
wire n_1294;
wire n_1351;
wire n_1380;
wire n_3336;
wire n_1291;
wire n_3763;
wire n_4284;
wire n_4370;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_1830;
wire n_3476;
wire n_3990;
wire n_2011;
wire n_4044;
wire n_1662;
wire n_3443;
wire n_3029;
wire n_4135;
wire n_1626;
wire n_3995;
wire n_4104;
wire n_1660;
wire n_4000;
wire n_2556;
wire n_1537;
wire n_3908;
wire n_3696;
wire n_2902;
wire n_3608;
wire n_4269;
wire n_4016;
wire n_4915;
wire n_4286;
wire n_3048;
wire n_1962;
wire n_1624;
wire n_1952;
wire n_4795;
wire n_1598;
wire n_2952;
wire n_2250;
wire n_1491;
wire n_3778;
wire n_2075;
wire n_4816;
wire n_3335;
wire n_4846;
wire n_3669;
wire n_1899;
wire n_4001;
wire n_2892;
wire n_3356;
wire n_4377;
wire n_3220;
wire n_3422;
wire n_1052;
wire n_2309;
wire n_2274;
wire n_3712;
wire n_2143;
wire n_4637;
wire n_4021;
wire n_2739;
wire n_2528;
wire n_2548;
wire n_3216;
wire n_3061;
wire n_3717;
wire n_3424;
wire n_3745;
wire n_3245;
wire n_4855;
wire n_4643;
wire n_4736;
wire n_2817;
wire n_1790;
wire n_4202;
wire n_3196;
wire n_4287;
wire n_2809;
wire n_3921;
wire n_3480;
wire n_1494;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_1726;
wire n_1241;
wire n_2589;
wire n_1231;
wire n_1208;
wire n_1604;
wire n_4947;
wire n_3506;
wire n_1976;
wire n_1337;
wire n_2984;
wire n_4890;
wire n_4538;
wire n_4023;
wire n_3031;
wire n_4920;
wire n_1238;
wire n_3959;
wire n_976;
wire n_1063;
wire n_4288;
wire n_2452;
wire n_2144;
wire n_4763;
wire n_2592;
wire n_2251;
wire n_1644;
wire n_4586;
wire n_3860;
wire n_1871;
wire n_3044;
wire n_2868;
wire n_3493;
wire n_2818;
wire n_3486;
wire n_2426;
wire n_1403;
wire n_2181;
wire n_3253;
wire n_4034;
wire n_1149;
wire n_4905;
wire n_1457;
wire n_3172;
wire n_2159;
wire n_2700;
wire n_1222;
wire n_1630;
wire n_1959;
wire n_1198;
wire n_3637;
wire n_3393;
wire n_1261;
wire n_3327;
wire n_1114;
wire n_3647;
wire n_3619;
wire n_3928;
wire n_4043;
wire n_1846;
wire n_1573;
wire n_1956;
wire n_4270;
wire n_2983;
wire n_4273;
wire n_1018;
wire n_1669;
wire n_1885;
wire n_1989;
wire n_1801;
wire n_3740;
wire n_3001;
wire n_4181;
wire n_2161;
wire n_2191;
wire n_2329;
wire n_2576;
wire n_4344;
wire n_1342;
wire n_2756;
wire n_4408;
wire n_1175;
wire n_1221;
wire n_3875;
wire n_4341;
wire n_4759;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_2567;
wire n_1085;
wire n_2981;
wire n_2222;
wire n_4439;
wire n_4565;
wire n_1451;
wire n_4663;
wire n_2471;
wire n_1288;
wire n_1275;
wire n_4519;
wire n_1622;
wire n_2757;
wire n_3121;
wire n_2121;
wire n_4515;
wire n_1893;
wire n_2278;
wire n_2433;
wire n_2798;
wire n_3425;
wire n_1771;
wire n_3308;
wire n_1507;
wire n_1206;
wire n_3576;
wire n_3109;
wire n_4838;
wire n_2553;
wire n_4524;
wire n_2218;
wire n_2130;
wire n_4862;
wire n_4260;
wire n_4628;
wire n_4696;
wire n_1097;
wire n_3122;
wire n_3012;
wire n_3368;
wire n_3586;
wire n_2381;
wire n_2313;
wire n_4597;
wire n_1812;
wire n_4574;
wire n_4242;
wire n_4949;
wire n_4748;
wire n_4959;
wire n_1747;
wire n_3400;
wire n_2508;
wire n_4243;
wire n_2540;
wire n_3820;
wire n_2672;
wire n_3360;
wire n_1585;
wire n_2316;
wire n_1995;
wire n_4677;
wire n_1631;
wire n_2911;
wire n_1828;
wire n_1389;
wire n_1798;
wire n_4562;
wire n_1584;
wire n_1438;
wire n_1973;
wire n_2156;
wire n_4453;
wire n_1366;
wire n_1187;
wire n_3173;
wire n_4281;
wire n_4332;
wire n_3433;
wire n_3998;
wire n_1686;
wire n_4464;
wire n_3017;
wire n_4605;
wire n_4737;
wire n_2542;
wire n_2843;
wire n_3305;
wire n_1635;
wire n_4310;
wire n_3752;
wire n_2637;
wire n_3543;
wire n_3655;
wire n_3791;
wire n_3050;
wire n_2666;
wire n_4091;
wire n_4906;
wire n_4257;
wire n_4516;
wire n_2913;
wire n_1381;
wire n_2254;
wire n_1597;
wire n_1486;
wire n_1068;
wire n_4196;
wire n_2371;
wire n_3898;
wire n_3366;
wire n_1024;
wire n_3453;
wire n_4107;
wire n_1949;
wire n_1197;
wire n_2408;
wire n_4961;
wire n_2140;
wire n_2134;
wire n_2483;
wire n_2466;
wire n_3661;
wire n_2048;
wire n_2760;
wire n_1299;
wire n_2942;
wire n_4420;
wire n_4964;
wire n_3665;
wire n_2079;
wire n_4807;
wire n_4886;
wire n_4342;
wire n_2671;
wire n_3296;
wire n_1390;
wire n_2775;
wire n_1023;
wire n_3223;
wire n_2005;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_2848;
wire n_1784;
wire n_3200;
wire n_1213;
wire n_3483;
wire n_3207;
wire n_1180;
wire n_4657;
wire n_3869;
wire n_3852;
wire n_1220;
wire n_3036;
wire n_4207;
wire n_1022;
wire n_1760;
wire n_2173;
wire n_2824;
wire n_4038;
wire n_4793;
wire n_4472;
wire n_2588;
wire n_3046;
wire n_1020;
wire n_1142;
wire n_1385;
wire n_4395;
wire n_4274;
wire n_1062;
wire n_2533;
wire n_1500;
wire n_2706;
wire n_1868;
wire n_2303;
wire n_4532;
wire n_3332;
wire n_4413;
wire n_4743;
wire n_2403;
wire n_2702;
wire n_3922;
wire n_2791;
wire n_1450;
wire n_2092;
wire n_3189;
wire n_2797;
wire n_1089;
wire n_4275;
wire n_2988;
wire n_3945;
wire n_1882;
wire n_2996;
wire n_2836;
wire n_1404;
wire n_3582;
wire n_4830;
wire n_4442;
wire n_1442;
wire n_2168;
wire n_4689;
wire n_2886;
wire n_1968;
wire n_4018;
wire n_2609;
wire n_4613;
wire n_1483;
wire n_1703;
wire n_1953;
wire n_3715;
wire n_1059;
wire n_3261;
wire n_3861;
wire n_3161;
wire n_3313;
wire n_1807;
wire n_1310;
wire n_3198;
wire n_3463;
wire n_2559;
wire n_4188;
wire n_2619;
wire n_2726;
wire n_2917;
wire n_3738;
wire n_1640;
wire n_1145;
wire n_2307;
wire n_3546;
wire n_1511;
wire n_1651;
wire n_3944;
wire n_3595;
wire n_1732;
wire n_2167;
wire n_3079;
wire n_1696;
wire n_1355;
wire n_4534;
wire n_3635;
wire n_3270;
wire n_4590;
wire n_4602;
wire n_1335;
wire n_3213;
wire n_4394;
wire n_1900;
wire n_3418;
wire n_2614;
wire n_1091;
wire n_1780;
wire n_3865;
wire n_2769;
wire n_4220;
wire n_3244;
wire n_3195;
wire n_3997;
wire n_4742;
wire n_2100;
wire n_4948;
wire n_3903;
wire n_3895;
wire n_1194;
wire n_4508;
wire n_3851;
wire n_4934;
wire n_3482;
wire n_2282;
wire n_970;
wire n_3654;
wire n_4939;
wire n_4213;
wire n_2430;
wire n_2673;
wire n_2926;
wire n_1534;
wire n_3268;
wire n_4703;
wire n_1655;
wire n_3494;
wire n_3615;
wire n_3363;
wire n_1186;
wire n_3180;
wire n_1743;
wire n_1506;
wire n_2594;
wire n_1474;
wire n_3150;
wire n_4773;
wire n_3853;
wire n_2512;
wire n_4449;
wire n_2607;
wire n_4615;
wire n_3911;
wire n_4883;
wire n_1079;
wire n_3559;
wire n_4943;
wire n_2498;
wire n_4630;
wire n_3812;
wire n_2017;
wire n_1227;
wire n_3750;
wire n_3838;
wire n_1954;
wire n_4749;
wire n_1125;
wire n_2687;
wire n_3456;
wire n_3132;
wire n_4159;
wire n_4372;
wire n_1044;
wire n_4731;
wire n_4004;
wire n_1134;
wire n_1684;
wire n_4353;
wire n_3334;
wire n_3819;
wire n_2023;
wire n_2720;
wire n_3870;
wire n_1233;
wire n_3653;
wire n_4360;
wire n_4897;
wire n_963;
wire n_2139;
wire n_3693;
wire n_1138;
wire n_2943;
wire n_1096;
wire n_3135;
wire n_4239;
wire n_3175;
wire n_1268;
wire n_3187;
wire n_3830;
wire n_2724;
wire n_1829;
wire n_1338;
wire n_1327;
wire n_3407;
wire n_3315;
wire n_4470;
wire n_4690;
wire n_3982;
wire n_2565;
wire n_4201;
wire n_1636;
wire n_1687;
wire n_4584;
wire n_3184;
wire n_4155;
wire n_3890;
wire n_2032;
wire n_3392;
wire n_4802;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_1680;
wire n_1195;
wire n_4304;
wire n_4821;
wire n_4160;
wire n_2860;
wire n_2448;
wire n_2015;
wire n_4910;
wire n_3641;
wire n_4887;
wire n_3996;
wire n_2873;
wire n_1576;
wire n_3049;
wire n_4015;
wire n_4211;
wire n_4119;
wire n_3620;
wire n_2558;
wire n_2347;
wire n_3884;
wire n_3103;
wire n_3770;
wire n_4591;
wire n_2527;
wire n_1509;
wire n_1648;
wire n_2944;
wire n_4349;
wire n_1886;
wire n_1841;
wire n_2685;
wire n_1313;
wire n_4223;
wire n_2090;
wire n_3722;
wire n_3802;
wire n_2215;
wire n_1449;
wire n_1723;
wire n_3129;
wire n_4806;
wire n_2116;
wire n_3592;
wire n_1645;
wire n_3186;
wire n_973;
wire n_1943;
wire n_3541;
wire n_1863;
wire n_1269;
wire n_2773;
wire n_2906;
wire n_3097;
wire n_3910;
wire n_4238;
wire n_1466;
wire n_3667;
wire n_1007;
wire n_3822;
wire n_1276;
wire n_1637;
wire n_2900;
wire n_3765;
wire n_2216;
wire n_4259;
wire n_1620;
wire n_3518;
wire n_2022;
wire n_3967;
wire n_2373;
wire n_1853;
wire n_2275;
wire n_2899;
wire n_3351;
wire n_2008;
wire n_2859;
wire n_2564;
wire n_4799;
wire n_1356;
wire n_2591;
wire n_3965;
wire n_1969;
wire n_1296;
wire n_4444;
wire n_4676;
wire n_1764;
wire n_1019;
wire n_1250;
wire n_1190;
wire n_4598;
wire n_3259;
wire n_4533;
wire n_4078;
wire n_1794;
wire n_3779;
wire n_3203;
wire n_3923;
wire n_4392;
wire n_3808;
wire n_4455;
wire n_3093;
wire n_2664;
wire n_1434;
wire n_4129;
wire n_2114;
wire n_1609;
wire n_3530;
wire n_1132;
wire n_4548;
wire n_1803;
wire n_1281;
wire n_4535;
wire n_1447;
wire n_2150;
wire n_2660;
wire n_4604;
wire n_3467;
wire n_4240;
wire n_2219;
wire n_4522;
wire n_1387;
wire n_1040;
wire n_3371;
wire n_4713;
wire n_1368;
wire n_1154;
wire n_2539;
wire n_1701;
wire n_2387;
wire n_3375;
wire n_2397;
wire n_3317;
wire n_3963;
wire n_3461;
wire n_2729;
wire n_1571;
wire n_2529;
wire n_4103;
wire n_4126;
wire n_4710;
wire n_3282;
wire n_1003;
wire n_2708;
wire n_2748;
wire n_2224;
wire n_2233;
wire n_2499;
wire n_3888;
wire n_4549;
wire n_3309;
wire n_1924;
wire n_3024;
wire n_4767;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_1553;
wire n_3542;
wire n_1090;
wire n_3374;
wire n_3704;
wire n_2786;
wire n_1905;
wire n_4355;
wire n_2958;
wire n_981;
wire n_2118;
wire n_2259;
wire n_2162;
wire n_4834;
wire n_3660;
wire n_2718;
wire n_4712;
wire n_1795;
wire n_3634;
wire n_4096;
wire n_2101;
wire n_1152;
wire n_3626;
wire n_2599;
wire n_4571;
wire n_3171;
wire n_1733;
wire n_3986;
wire n_2853;
wire n_1552;
wire n_4930;
wire n_2217;
wire n_3594;
wire n_2866;
wire n_3153;
wire n_1189;
wire n_4039;
wire n_4253;
wire n_4681;
wire n_2623;
wire n_3232;
wire n_2178;
wire n_1181;
wire n_3815;
wire n_4375;
wire n_4205;
wire n_3790;
wire n_2404;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_1203;
wire n_3640;
wire n_2821;
wire n_4768;
wire n_3299;
wire n_4070;
wire n_4558;
wire n_3065;
wire n_2375;
wire n_2572;
wire n_1656;
wire n_1076;
wire n_2063;
wire n_3082;
wire n_4504;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_4864;
wire n_3855;
wire n_3357;
wire n_4485;
wire n_1510;
wire n_2852;
wire n_2132;
wire n_1236;
wire n_3412;
wire n_1712;
wire n_4537;
wire n_1184;
wire n_2585;
wire n_2220;
wire n_4005;
wire n_1364;
wire n_3183;
wire n_4323;
wire n_4184;
wire n_2468;
wire n_3248;
wire n_2606;
wire n_4337;
wire n_4826;
wire n_2152;
wire n_4952;
wire n_3785;
wire n_3525;
wire n_2779;
wire n_1117;
wire n_2547;
wire n_1748;
wire n_2935;
wire n_2490;
wire n_3127;
wire n_3496;
wire n_3568;
wire n_4876;
wire n_3841;
wire n_4626;
wire n_1334;
wire n_3879;
wire n_2402;
wire n_1200;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_4747;
wire n_3341;
wire n_4347;
wire n_1852;
wire n_3868;
wire n_4791;
wire n_2481;
wire n_4409;
wire n_1264;
wire n_2808;
wire n_3396;
wire n_2102;
wire n_3492;
wire n_3558;
wire n_2751;
wire n_1548;
wire n_4824;
wire n_2977;
wire n_1682;
wire n_3599;
wire n_1896;
wire n_1704;
wire n_2234;
wire n_4152;
wire n_1352;
wire n_2328;
wire n_4587;
wire n_2332;
wire n_1628;
wire n_1773;
wire n_3580;
wire n_2369;
wire n_3584;
wire n_4500;
wire n_1115;
wire n_1395;
wire n_4660;
wire n_2823;
wire n_3274;
wire n_2613;
wire n_1046;
wire n_2419;
wire n_2807;
wire n_4047;
wire n_4157;
wire n_3956;
wire n_1431;
wire n_1086;
wire n_1523;
wire n_1756;
wire n_2241;
wire n_2458;
wire n_3032;
wire n_3401;
wire n_1750;
wire n_2833;
wire n_3179;
wire n_1563;
wire n_4051;
wire n_3123;
wire n_1875;
wire n_1615;
wire n_3719;
wire n_2635;
wire n_4077;
wire n_3897;
wire n_3475;
wire n_2077;
wire n_2520;
wire n_2193;
wire n_4010;
wire n_4942;
wire n_4255;
wire n_2908;
wire n_4561;
wire n_4957;
wire n_2053;
wire n_1580;
wire n_2200;
wire n_2304;
wire n_4683;
wire n_1439;
wire n_2352;
wire n_4839;
wire n_2185;
wire n_2476;
wire n_1266;
wire n_4814;
wire n_2781;
wire n_2460;
wire n_4694;
wire n_3600;
wire n_4109;
wire n_1870;
wire n_2484;
wire n_2721;
wire n_2308;
wire n_3498;
wire n_4520;
wire n_1428;
wire n_4026;
wire n_2903;
wire n_3659;
wire n_4496;
wire n_1528;
wire n_3840;
wire n_3481;
wire n_4719;
wire n_4100;
wire n_3517;
wire n_1413;
wire n_2464;
wire n_2925;
wire n_2270;
wire n_1706;
wire n_1592;
wire n_1461;
wire n_2695;
wire n_3656;
wire n_3137;
wire n_3116;
wire n_4426;
wire n_2414;
wire n_3316;
wire n_2465;
wire n_3925;
wire n_4089;
wire n_1683;
wire n_4175;
wire n_4458;
wire n_3955;
wire n_1035;
wire n_3158;
wire n_3657;
wire n_2684;
wire n_1104;
wire n_2205;
wire n_2875;
wire n_3284;
wire n_1437;
wire n_2747;
wire n_4185;
wire n_2064;
wire n_3088;
wire n_1497;
wire n_2002;
wire n_4815;
wire n_2545;
wire n_2050;
wire n_3695;
wire n_2500;
wire n_1917;
wire n_1444;
wire n_4316;
wire n_3328;
wire n_2763;
wire n_994;
wire n_2761;
wire n_4020;
wire n_1920;
wire n_4306;
wire n_2997;
wire n_961;
wire n_3735;
wire n_2127;
wire n_3028;
wire n_3228;
wire n_3706;
wire n_1432;
wire n_3322;
wire n_996;
wire n_1174;
wire n_4512;
wire n_4483;
wire n_3499;
wire n_3552;
wire n_4164;
wire n_1286;
wire n_3784;
wire n_4142;
wire n_4621;
wire n_3016;
wire n_1629;
wire n_2694;
wire n_3609;
wire n_3447;
wire n_3771;
wire n_4678;
wire n_2647;
wire n_1850;
wire n_1670;
wire n_4123;
wire n_2317;
wire n_1384;
wire n_1612;
wire n_1099;
wire n_3113;
wire n_4305;
wire n_2909;
wire n_4007;
wire n_3960;
wire n_1524;
wire n_4707;
wire n_4429;
wire n_1991;
wire n_2566;
wire n_2210;
wire n_1225;
wire n_2346;
wire n_4695;
wire n_982;
wire n_2180;
wire n_3376;
wire n_2617;
wire n_4163;
wire n_2831;
wire n_2865;
wire n_1625;
wire n_4638;
wire n_4498;
wire n_2240;
wire n_1797;
wire n_4750;
wire n_3993;
wire n_2120;
wire n_1289;
wire n_1557;
wire n_1567;
wire n_2007;
wire n_2004;
wire n_2086;
wire n_4832;
wire n_3666;
wire n_1839;
wire n_1587;
wire n_2330;
wire n_2555;
wire n_2108;
wire n_2535;
wire n_2945;
wire n_3057;
wire n_4319;
wire n_3760;
wire n_1396;
wire n_1224;
wire n_1923;
wire n_2196;
wire n_1538;
wire n_3773;
wire n_2604;
wire n_3462;
wire n_4373;
wire n_2437;
wire n_2351;
wire n_1889;
wire n_1124;
wire n_2688;
wire n_3302;
wire n_1673;
wire n_2085;
wire n_3304;
wire n_1725;
wire n_2149;
wire n_2001;
wire n_1800;
wire n_3746;
wire n_3645;
wire n_4262;
wire n_4019;
wire n_2735;
wire n_2035;
wire n_4436;
wire n_4697;
wire n_1906;
wire n_1647;
wire n_4357;
wire n_4849;
wire n_4366;
wire n_4139;
wire n_1270;
wire n_4340;
wire n_1476;
wire n_1054;
wire n_2027;
wire n_2012;
wire n_3512;
wire n_4720;
wire n_3892;
wire n_1880;
wire n_1642;
wire n_2447;
wire n_3358;
wire n_2894;
wire n_2587;
wire n_1605;
wire n_2099;
wire n_1202;
wire n_3410;
wire n_975;
wire n_4900;
wire n_3408;
wire n_3182;
wire n_1879;
wire n_4941;
wire n_1311;
wire n_2299;
wire n_2078;
wire n_3709;
wire n_3011;
wire n_2315;
wire n_3623;
wire n_2157;
wire n_3446;
wire n_1770;
wire n_1107;
wire n_4167;
wire n_3058;
wire n_4334;
wire n_2211;
wire n_3384;
wire n_4698;
wire n_2225;
wire n_1411;
wire n_1501;
wire n_4397;
wire n_3611;
wire n_4186;
wire n_2093;
wire n_2675;
wire n_4229;
wire n_4294;
wire n_1919;
wire n_4351;
wire n_2893;
wire n_2009;
wire n_4162;
wire n_1416;
wire n_3465;
wire n_1515;
wire n_4127;
wire n_4620;
wire n_1314;
wire n_3059;
wire n_3085;
wire n_2867;
wire n_2229;
wire n_4770;
wire n_3871;
wire n_2388;
wire n_3112;
wire n_3413;
wire n_4580;
wire n_2624;
wire n_1813;
wire n_1005;
wire n_4581;
wire n_4618;
wire n_1105;
wire n_2898;
wire n_2519;
wire n_2231;
wire n_1000;
wire n_2816;
wire n_2803;
wire n_3402;
wire n_1256;
wire n_4670;
wire n_1769;
wire n_1060;
wire n_1372;
wire n_1847;
wire n_3805;
wire n_2406;
wire n_4017;
wire n_1586;
wire n_3497;
wire n_3382;
wire n_4236;
wire n_4313;
wire n_3561;
wire n_2543;
wire n_2992;
wire n_1541;
wire n_4907;
wire n_4659;
wire n_1697;
wire n_2128;
wire n_1872;
wire n_2690;
wire n_3942;
wire n_2020;
wire n_1939;
wire n_4053;
wire n_4279;
wire n_3937;
wire n_3303;
wire n_4555;
wire n_3549;
wire n_1481;
wire n_1928;
wire n_4235;
wire n_3972;
wire n_2314;
wire n_2126;
wire n_3403;
wire n_1363;
wire n_1691;
wire n_1098;
wire n_1361;
wire n_1693;
wire n_2081;
wire n_2993;
wire n_3018;
wire n_4820;
wire n_2449;
wire n_2131;
wire n_2526;
wire n_4794;
wire n_1302;
wire n_3989;
wire n_4752;
wire n_4546;
wire n_3918;
wire n_3191;
wire n_1029;
wire n_3051;
wire n_1317;
wire n_3643;
wire n_2615;
wire n_2487;
wire n_3343;
wire n_4415;
wire n_3163;
wire n_3786;
wire n_4061;
wire n_4432;
wire n_1912;
wire n_4552;
wire n_3143;
wire n_1876;
wire n_4790;
wire n_1811;
wire n_1285;
wire n_967;
wire n_4263;
wire n_3725;
wire n_1529;
wire n_1824;
wire n_3522;
wire n_4528;
wire n_4888;
wire n_4502;
wire n_4335;
wire n_3444;
wire n_4218;
wire n_4705;
wire n_3009;
wire n_1141;
wire n_4471;
wire n_3297;
wire n_1168;
wire n_3000;
wire n_2305;
wire n_1192;
wire n_1290;
wire n_2514;
wire n_4386;
wire n_4547;
wire n_4836;
wire n_3545;
wire n_1101;
wire n_4193;
wire n_1336;
wire n_1358;
wire n_3318;
wire n_1397;
wire n_1359;
wire n_3226;
wire n_3702;
wire n_3981;
wire n_1532;
wire n_3430;
wire n_1685;
wire n_2801;
wire n_3225;
wire n_3067;
wire n_1074;
wire n_1462;
wire n_3823;
wire n_4718;
wire n_3185;
wire n_2326;
wire n_1398;
wire n_1904;
wire n_2966;
wire n_3084;
wire n_4634;
wire n_1692;
wire n_4796;
wire n_4560;
wire n_1240;
wire n_3285;
wire n_1814;
wire n_4882;
wire n_1808;
wire n_2768;
wire n_1658;
wire n_3837;
wire n_4841;
wire n_3076;
wire n_4954;
wire n_4635;
wire n_4521;
wire n_1027;
wire n_3893;
wire n_4272;
wire n_2148;
wire n_2104;
wire n_2653;
wire n_2855;
wire n_2618;
wire n_4448;
wire n_3359;
wire n_2331;
wire n_1600;
wire n_4701;
wire n_4088;
wire n_2136;
wire n_1913;
wire n_1043;
wire n_3056;
wire n_4208;
wire n_1472;
wire n_1365;
wire n_2443;
wire n_3052;
wire n_4865;
wire n_2066;
wire n_1974;
wire n_1158;
wire n_4589;
wire n_3924;
wire n_1915;
wire n_2534;
wire n_4617;
wire n_3311;
wire n_1160;
wire n_4094;
wire n_4772;
wire n_4857;
wire n_3613;
wire n_1383;
wire n_2057;
wire n_1822;
wire n_1804;
wire n_1581;
wire n_4776;
wire n_1975;
wire n_3437;
wire n_3744;
wire n_2246;
wire n_2738;
wire n_1851;
wire n_1755;
wire n_4702;
wire n_1341;
wire n_4486;
wire n_4946;
wire n_2202;
wire n_2262;
wire n_1333;
wire n_4506;
wire n_3157;
wire n_4669;
wire n_4226;
wire n_4153;
wire n_4329;
wire n_4877;
wire n_3442;
wire n_2327;
wire n_4780;
wire n_4327;
wire n_2656;
wire n_4168;
wire n_2258;
wire n_4396;
wire n_2039;
wire n_1016;
wire n_4465;
wire n_2544;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_3266;
wire n_1843;
wire n_2030;
wire n_4576;
wire n_4075;
wire n_3593;
wire n_2536;
wire n_1399;
wire n_3685;
wire n_4833;
wire n_1903;
wire n_1849;
wire n_3768;
wire n_983;
wire n_4224;
wire n_4868;
wire n_2676;
wire n_3515;
wire n_3489;
wire n_3181;
wire n_3644;
wire n_4387;
wire n_2368;
wire n_4896;
wire n_1157;
wire n_2065;
wire n_2901;
wire n_3818;
wire n_4368;
wire n_1295;
wire n_1983;
wire n_992;
wire n_4798;
wire n_1582;
wire n_2201;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_3610;
wire n_2569;
wire n_1998;
wire n_1596;
wire n_3077;
wire n_1100;
wire n_4158;
wire n_4687;
wire n_4756;
wire n_4095;
wire n_2177;
wire n_2123;
wire n_4364;
wire n_3019;
wire n_2235;
wire n_1080;
wire n_2290;
wire n_3272;
wire n_4346;
wire n_2074;
wire n_2897;
wire n_4668;
wire n_2383;
wire n_2640;
wire n_1492;
wire n_1478;
wire n_1796;
wire n_3569;
wire n_1614;
wire n_2374;
wire n_4648;
wire n_2598;
wire n_1722;
wire n_4179;
wire n_3340;
wire n_2335;
wire n_4785;
wire n_2230;
wire n_3033;
wire n_2151;
wire n_4912;
wire n_1971;
wire n_2479;
wire n_4914;
wire n_2359;
wire n_2360;
wire n_4902;
wire n_4369;
wire n_1392;
wire n_2158;
wire n_2571;
wire n_2799;
wire n_4708;
wire n_4592;
wire n_1307;
wire n_2644;
wire n_4445;
wire n_3211;
wire n_1840;
wire n_2837;
wire n_989;
wire n_1668;
wire n_1681;
wire n_4031;
wire n_4120;
wire n_3896;
wire n_3533;
wire n_2192;
wire n_4578;
wire n_3323;
wire n_1937;
wire n_3839;
wire n_3509;
wire n_1749;
wire n_2918;
wire n_3353;
wire n_1945;
wire n_2638;
wire n_3939;
wire n_4874;
wire n_1228;
wire n_4840;
wire n_2354;
wire n_4311;
wire n_1133;
wire n_1926;
wire n_2363;
wire n_2814;
wire n_3264;
wire n_3204;
wire n_2003;
wire n_3727;
wire n_2621;
wire n_2922;
wire n_3881;
wire n_1030;
wire n_1910;
wire n_1606;
wire n_3711;
wire n_2164;
wire n_1618;
wire n_3748;
wire n_4389;
wire n_3668;
wire n_3197;
wire n_1955;
wire n_4556;
wire n_2413;
wire n_3148;
wire n_4779;
wire n_1253;
wire n_1484;
wire n_2686;
wire n_4214;
wire n_4430;
wire n_3151;
wire n_3977;
wire n_3125;
wire n_2812;
wire n_4889;
wire n_4221;
wire n_1638;
wire n_4650;
wire n_1038;
wire n_2280;
wire n_4428;
wire n_4784;
wire n_2393;
wire n_4766;
wire n_3809;
wire n_979;
wire n_1999;
wire n_3810;
wire n_1215;
wire n_3579;
wire n_2777;
wire n_2480;
wire n_2283;
wire n_2806;
wire n_2813;
wire n_4295;
wire n_1716;
wire n_1412;
wire n_3310;
wire n_4182;
wire n_1401;
wire n_2951;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_2579;
wire n_2876;
wire n_3301;
wire n_2370;
wire n_4600;
wire n_2025;
wire n_3451;
wire n_1219;
wire n_4513;
wire n_1252;
wire n_2730;
wire n_1927;
wire n_4735;
wire n_2767;
wire n_4667;
wire n_2826;
wire n_2112;
wire n_2762;
wire n_4774;
wire n_4711;
wire n_3023;
wire n_3224;
wire n_4481;
wire n_3762;
wire n_4671;
wire n_1326;
wire n_978;
wire n_1799;
wire n_1689;
wire n_1304;
wire n_2541;
wire n_4879;
wire n_2987;
wire n_1702;
wire n_3916;
wire n_3630;
wire n_1558;
wire n_1073;
wire n_2722;
wire n_3618;
wire n_2727;
wire n_2719;
wire n_2213;
wire n_3521;
wire n_2723;
wire n_4054;
wire n_1569;
wire n_4012;
wire n_3567;
wire n_4352;
wire n_1988;
wire n_2401;
wire n_1787;
wire n_3094;
wire n_2166;
wire n_2451;
wire n_4665;
wire n_2631;
wire n_1867;
wire n_4252;
wire n_4505;
wire n_4219;
wire n_2292;
wire n_3560;
wire n_1742;
wire n_1818;
wire n_3847;
wire n_2203;
wire n_4909;
wire n_2693;
wire n_1159;
wire n_2281;
wire n_3202;
wire n_2646;
wire n_3887;
wire n_3800;
wire n_4435;
wire n_1235;
wire n_4755;
wire n_3827;
wire n_3156;
wire n_4303;
wire n_3457;
wire n_1058;
wire n_1835;
wire n_2697;
wire n_3531;
wire n_2470;
wire n_2890;
wire n_4400;
wire n_1519;
wire n_1425;
wire n_4812;
wire n_2069;
wire n_2602;
wire n_4090;
wire n_4136;
wire n_1156;
wire n_4358;
wire n_2857;
wire n_1360;
wire n_2070;
wire n_3471;
wire n_4098;
wire n_3117;
wire n_3039;
wire n_3900;
wire n_3478;
wire n_3701;
wire n_2766;
wire n_3756;
wire n_3754;
wire n_4156;
wire n_2416;
wire n_2962;
wire n_1031;
wire n_3694;
wire n_2052;
wire n_3690;
wire n_3006;
wire n_3348;
wire n_4758;
wire n_2236;
wire n_3957;
wire n_2377;
wire n_2577;
wire n_3165;
wire n_4419;
wire n_2795;
wire n_3520;
wire n_2632;
wire n_4406;
wire n_1036;
wire n_1106;
wire n_4655;
wire n_1634;
wire n_1452;
wire n_4953;
wire n_4570;
wire n_3966;
wire n_4293;
wire n_1577;
wire n_1700;
wire n_4542;
wire n_4122;
wire n_2819;
wire n_1140;
wire n_1985;
wire n_4740;
wire n_1056;
wire n_3007;
wire n_1487;
wire n_1237;
wire n_4230;
wire n_1109;
wire n_2741;
wire n_4333;
wire n_3436;
wire n_4460;
wire n_2312;
wire n_2946;
wire n_4040;
wire n_1884;
wire n_1589;
wire n_2717;
wire n_4527;
wire n_2877;
wire n_1996;
wire n_3964;
wire n_3110;
wire n_1677;
wire n_4384;
wire n_2297;
wire n_3037;
wire n_3188;
wire n_2780;
wire n_1792;
wire n_3250;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_4762;
wire n_1877;
wire n_1477;
wire n_3155;
wire n_4938;
wire n_4407;
wire n_1075;
wire n_1249;
wire n_3468;
wire n_2006;
wire n_1990;
wire n_3680;
wire n_3624;
wire n_2467;
wire n_4292;
wire n_3145;
wire n_2662;
wire n_3872;
wire n_3801;
wire n_2883;
wire n_1178;
wire n_1566;
wire n_1464;
wire n_4092;
wire n_3003;
wire n_4244;
wire n_2277;
wire n_1982;
wire n_2252;
wire n_1695;
wire n_2999;
wire n_3331;
wire n_2910;
wire n_4414;
wire n_2294;
wire n_2295;
wire n_4706;
wire n_1602;
wire n_2965;
wire n_2382;
wire n_2557;
wire n_2505;
wire n_3554;
wire n_3730;
wire n_4307;
wire n_4356;
wire n_1935;
wire n_3367;
wire n_1146;
wire n_2785;
wire n_4929;
wire n_1608;
wire n_3776;
wire n_4951;
wire n_1009;
wire n_2160;
wire n_2991;
wire n_2699;
wire n_1436;
wire n_4137;
wire n_1485;
wire n_2239;
wire n_3826;
wire n_4365;
wire n_1979;
wire n_3781;
wire n_4215;
wire n_4315;
wire n_2971;
wire n_3072;
wire n_1545;
wire n_3249;
wire n_3797;
wire n_3281;
wire n_3505;
wire n_4427;
wire n_4564;
wire n_2934;
wire n_4042;
wire n_2525;
wire n_4624;
wire n_4317;
wire n_3087;
wire n_4925;
wire n_2197;
wire n_1470;
wire n_2098;
wire n_1761;
wire n_4041;
wire n_4958;
wire n_4297;
wire n_4709;
wire n_3379;
wire n_4425;
wire n_3390;
wire n_1539;
wire n_1806;
wire n_2711;
wire n_3646;
wire n_2209;
wire n_3020;
wire n_3142;
wire n_2612;
wire n_2095;
wire n_2486;
wire n_2521;
wire n_1574;
wire n_4764;
wire n_4899;
wire n_4141;
wire n_4614;
wire n_2979;
wire n_4739;
wire n_1300;
wire n_4035;
wire n_4291;
wire n_3419;
wire n_4935;
wire n_4880;
wire n_3167;
wire n_2986;
wire n_2400;
wire n_2507;
wire n_3682;
wire n_3131;
wire n_1495;
wire n_1357;
wire n_4566;
wire n_2794;
wire n_3672;
wire n_2496;
wire n_4918;
wire n_2974;
wire n_2990;
wire n_2923;
wire n_3449;
wire n_1339;
wire n_1544;
wire n_4933;
wire n_4872;
wire n_1315;
wire n_4647;
wire n_2340;
wire n_2117;
wire n_1328;
wire n_4837;
wire n_1048;
wire n_3638;
wire n_2106;
wire n_1263;
wire n_4940;
wire n_4176;
wire n_4454;
wire n_964;
wire n_3772;
wire n_2948;
wire n_4322;
wire n_2298;
wire n_2771;
wire n_4336;
wire n_3219;
wire n_3867;
wire n_4956;
wire n_2045;
wire n_1535;
wire n_4227;
wire n_2190;
wire n_1972;
wire n_3080;
wire n_2772;
wire n_2778;
wire n_3929;
wire n_1898;
wire n_1254;
wire n_2524;
wire n_3927;
wire n_1941;
wire n_3564;
wire n_3095;
wire n_1783;
wire n_3279;
wire n_1815;
wire n_3344;
wire n_4133;
wire n_3985;
wire n_3252;
wire n_1162;
wire n_2578;
wire n_2745;
wire n_2110;
wire n_3747;
wire n_991;
wire n_1323;
wire n_3710;
wire n_1429;
wire n_3209;
wire n_2026;
wire n_3588;
wire n_2103;
wire n_4497;
wire n_4388;
wire n_3632;
wire n_1874;
wire n_4116;
wire n_3377;
wire n_1601;
wire n_3414;
wire n_2933;
wire n_3828;
wire n_1367;
wire n_3240;
wire n_2895;
wire n_1694;
wire n_1458;
wire n_2271;
wire n_2356;
wire n_2261;
wire n_4066;
wire n_2994;
wire n_2105;
wire n_2187;
wire n_2642;
wire n_1643;
wire n_1789;
wire n_2415;
wire n_3152;
wire n_3154;
wire n_2344;
wire n_3589;
wire n_1112;
wire n_2384;
wire n_1376;
wire n_1858;
wire n_3523;
wire n_2815;
wire n_2446;
wire n_3388;
wire n_1172;
wire n_2659;
wire n_3616;
wire n_4048;
wire n_4084;
wire n_1527;
wire n_3174;
wire n_4848;
wire n_2849;
wire n_1177;
wire n_3292;
wire n_3940;
wire n_2502;
wire n_4860;
wire n_4438;
wire n_3290;
wire n_3585;
wire n_2878;
wire n_1810;
wire n_3047;
wire n_2610;
wire n_1037;
wire n_3427;
wire n_1188;
wire n_3431;
wire n_2024;
wire n_3783;
wire n_1503;
wire n_1942;
wire n_4326;
wire n_3141;
wire n_2698;
wire n_3930;
wire n_4149;
wire n_1259;
wire n_4101;
wire n_4792;
wire n_2916;
wire n_3736;
wire n_2611;
wire n_4383;
wire n_2709;
wire n_2244;
wire n_3664;
wire n_1456;
wire n_3907;
wire n_2665;
wire n_3063;
wire n_4543;
wire n_2881;
wire n_3862;
wire n_2018;
wire n_3134;
wire n_993;
wire n_2581;
wire n_2268;
wire n_2237;
wire n_2320;
wire n_2255;
wire n_1820;
wire n_3906;
wire n_3474;
wire n_1946;
wire n_3111;
wire n_4212;
wire n_4827;
wire n_1639;
wire n_2154;
wire n_3162;
wire n_4599;
wire n_2732;
wire n_3004;
wire n_3333;
wire n_4509;
wire n_3705;
wire n_4783;
wire n_3276;
wire n_1006;
wire n_2956;
wire n_1415;
wire n_3743;
wire n_4068;
wire n_2153;
wire n_2891;
wire n_2457;
wire n_3825;
wire n_4434;
wire n_2737;
wire n_1406;
wire n_3591;
wire n_2137;
wire n_1473;
wire n_3140;
wire n_2125;
wire n_1176;
wire n_3848;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_4622;
wire n_3139;
wire n_4715;
wire n_4222;
wire n_2206;
wire n_3734;
wire n_3538;
wire n_4716;
wire n_4588;
wire n_2265;
wire n_1167;
wire n_3231;
wire n_3138;
wire n_1282;
wire n_2067;
wire n_2517;
wire n_3349;
wire n_3454;
wire n_4143;
wire n_4410;
wire n_1718;
wire n_3229;
wire n_2546;
wire n_4741;
wire n_1139;
wire n_2345;
wire n_1324;
wire n_4440;
wire n_3649;
wire n_1838;
wire n_3824;
wire n_3439;
wire n_1513;
wire n_1788;
wire n_2348;
wire n_2417;
wire n_2043;
wire n_3601;
wire n_1621;
wire n_2338;
wire n_3571;
wire n_2248;
wire n_958;
wire n_3500;
wire n_2850;
wire n_3962;
wire n_3846;
wire n_4328;
wire n_1433;
wire n_1907;
wire n_3994;
wire n_2135;
wire n_1088;
wire n_1102;
wire n_4487;
wire n_1165;
wire n_4148;
wire n_3066;
wire n_2869;
wire n_4829;
wire n_2455;
wire n_2874;
wire n_4937;
wire n_4463;
wire n_2284;
wire n_1931;
wire n_1809;
wire n_3491;
wire n_4844;
wire n_3271;
wire n_2667;
wire n_1565;
wire n_2325;
wire n_3346;
wire n_3391;
wire n_1542;
wire n_1547;
wire n_1362;
wire n_4178;
wire n_4324;
wire n_3288;
wire n_2518;
wire n_3045;
wire n_3014;
wire n_1951;
wire n_1330;
wire n_1940;
wire n_3767;
wire n_1212;
wire n_1199;
wire n_4852;
wire n_1978;
wire n_1767;
wire n_1443;
wire n_1861;
wire n_1564;
wire n_2593;
wire n_1623;
wire n_1131;
wire n_3120;
wire n_1554;
wire n_4843;
wire n_4761;
wire n_2021;
wire n_2713;
wire n_2938;
wire n_3227;
wire n_3342;
wire n_2939;
wire n_4036;
wire n_1147;
wire n_4380;
wire n_2790;
wire n_2034;
wire n_3102;
wire n_4345;
wire n_1892;
wire n_2061;
wire n_1373;
wire n_3866;
wire n_3803;
wire n_2083;
wire n_2119;
wire n_2207;
wire n_4210;
wire n_3485;
wire n_4810;
wire n_3149;
wire n_2827;
wire n_3278;
wire n_2701;
wire n_2337;
wire n_4045;
wire n_4871;
wire n_2513;
wire n_1369;
wire n_1297;
wire n_1734;
wire n_4461;
wire n_2323;
wire n_3042;
wire n_2561;
wire n_2491;
wire n_1161;
wire n_1103;
wire n_4363;
wire n_3551;
wire n_3992;
wire n_4147;
wire n_4811;
wire n_3176;
wire n_2429;
wire n_3326;
wire n_3581;
wire n_3423;
wire n_1646;
wire n_4161;
wire n_1759;
wire n_2096;
wire n_2296;
wire n_1911;
wire n_2870;
wire n_4869;
wire n_4013;
wire n_1211;
wire n_4482;
wire n_3794;
wire n_1419;
wire n_4738;
wire n_1193;
wire n_980;
wire n_3557;
wire n_2928;
wire n_3380;
wire n_2227;
wire n_2652;
wire n_3596;
wire n_2627;
wire n_1827;
wire n_3369;
wire n_4086;
wire n_4112;
wire n_2501;
wire n_2051;
wire n_1805;
wire n_3737;
wire n_1183;
wire n_3160;
wire n_4744;
wire n_1204;
wire n_1151;
wire n_3286;
wire n_999;
wire n_1092;
wire n_2668;
wire n_1386;
wire n_2931;
wire n_2492;
wire n_3636;
wire n_4787;
wire n_4885;
wire n_2927;
wire n_4459;
wire n_1516;
wire n_4551;
wire n_4484;
wire n_1499;
wire n_2155;
wire n_966;
wire n_3938;
wire n_3114;
wire n_3905;
wire n_1661;
wire n_1965;
wire n_1757;
wire n_4726;
wire n_3617;
wire n_3602;
wire n_4298;
wire n_3053;
wire n_1039;
wire n_3894;
wire n_2407;
wire n_2267;
wire n_2302;
wire n_2082;
wire n_2453;
wire n_2560;
wire n_4544;
wire n_4418;
wire n_4595;
wire n_2770;
wire n_2704;
wire n_1762;
wire n_4944;
wire n_4468;
wire n_3421;
wire n_4950;
wire n_3247;
wire n_1026;
wire n_1454;
wire n_4108;
wire n_4594;
wire n_1325;
wire n_2754;
wire n_4629;
wire n_4903;
wire n_3041;
wire n_4194;
wire n_3713;
wire n_2692;
wire n_3889;
wire n_3325;
wire n_4299;
wire n_1744;
wire n_2324;
wire n_4921;
wire n_1111;
wire n_1819;
wire n_4863;
wire n_2670;
wire n_1745;
wire n_3941;
wire n_3516;
wire n_3933;
wire n_3562;
wire n_1916;
wire n_3873;
wire n_2073;
wire n_4093;
wire n_1947;
wire n_2165;
wire n_2016;
wire n_3793;
wire n_1791;
wire n_1113;
wire n_4817;
wire n_1468;
wire n_4917;
wire n_1164;
wire n_3749;
wire n_3691;
wire n_4452;
wire n_3501;
wire n_2538;
wire n_1559;
wire n_4446;
wire n_1280;
wire n_2854;
wire n_2932;
wire n_3258;
wire n_4280;
wire n_2285;
wire n_1934;
wire n_2040;
wire n_3246;
wire n_2186;
wire n_1665;
wire n_3417;
wire n_2725;
wire n_1482;
wire n_4782;
wire n_2349;
wire n_1902;
wire n_2474;
wire n_1417;
wire n_3536;
wire n_1346;
wire n_2834;
wire n_1123;
wire n_1272;
wire n_2497;
wire n_3040;
wire n_1410;
wire n_988;
wire n_3528;
wire n_3677;
wire n_2657;
wire n_2743;
wire n_4662;
wire n_2658;

INVx1_ASAP7_75t_L g958 ( 
.A(n_327),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_947),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_370),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_870),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_495),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_873),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_541),
.Y(n_964)
);

INVx1_ASAP7_75t_SL g965 ( 
.A(n_0),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_917),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_756),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_850),
.Y(n_968)
);

INVx2_ASAP7_75t_SL g969 ( 
.A(n_804),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_122),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_794),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_161),
.Y(n_972)
);

BUFx3_ASAP7_75t_L g973 ( 
.A(n_686),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_950),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_928),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_544),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_475),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_299),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_809),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_918),
.Y(n_980)
);

BUFx6f_ASAP7_75t_L g981 ( 
.A(n_289),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_422),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_882),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_826),
.Y(n_984)
);

INVx1_ASAP7_75t_SL g985 ( 
.A(n_853),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_912),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_609),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_405),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_857),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_392),
.Y(n_990)
);

BUFx5_ASAP7_75t_L g991 ( 
.A(n_250),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_926),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_944),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_732),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_340),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_228),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_455),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_667),
.Y(n_998)
);

INVx1_ASAP7_75t_SL g999 ( 
.A(n_284),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_721),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_933),
.Y(n_1001)
);

BUFx2_ASAP7_75t_L g1002 ( 
.A(n_818),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_825),
.Y(n_1003)
);

INVxp67_ASAP7_75t_SL g1004 ( 
.A(n_896),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_531),
.Y(n_1005)
);

INVxp33_ASAP7_75t_L g1006 ( 
.A(n_327),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_908),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_845),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_363),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_516),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_815),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_69),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_30),
.Y(n_1013)
);

CKINVDCx20_ASAP7_75t_R g1014 ( 
.A(n_784),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_571),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_794),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_84),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_817),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_136),
.Y(n_1019)
);

BUFx10_ASAP7_75t_L g1020 ( 
.A(n_949),
.Y(n_1020)
);

INVxp67_ASAP7_75t_L g1021 ( 
.A(n_455),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_416),
.Y(n_1022)
);

CKINVDCx20_ASAP7_75t_R g1023 ( 
.A(n_252),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_715),
.Y(n_1024)
);

BUFx3_ASAP7_75t_L g1025 ( 
.A(n_322),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_859),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_893),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_366),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_406),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_933),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_776),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_762),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_443),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_948),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_430),
.Y(n_1035)
);

INVxp67_ASAP7_75t_SL g1036 ( 
.A(n_869),
.Y(n_1036)
);

BUFx10_ASAP7_75t_L g1037 ( 
.A(n_334),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_386),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_901),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_575),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_421),
.Y(n_1041)
);

INVx2_ASAP7_75t_SL g1042 ( 
.A(n_194),
.Y(n_1042)
);

INVx1_ASAP7_75t_SL g1043 ( 
.A(n_868),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_927),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_575),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_749),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_5),
.Y(n_1047)
);

INVx1_ASAP7_75t_SL g1048 ( 
.A(n_709),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_382),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_832),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_762),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_872),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_607),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_462),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_907),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_891),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_233),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_748),
.Y(n_1058)
);

BUFx6f_ASAP7_75t_L g1059 ( 
.A(n_696),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_71),
.Y(n_1060)
);

HB1xp67_ASAP7_75t_L g1061 ( 
.A(n_502),
.Y(n_1061)
);

BUFx10_ASAP7_75t_L g1062 ( 
.A(n_954),
.Y(n_1062)
);

INVx1_ASAP7_75t_SL g1063 ( 
.A(n_176),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_108),
.Y(n_1064)
);

INVx2_ASAP7_75t_SL g1065 ( 
.A(n_570),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_214),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_525),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_619),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_850),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_692),
.Y(n_1070)
);

BUFx10_ASAP7_75t_L g1071 ( 
.A(n_708),
.Y(n_1071)
);

BUFx10_ASAP7_75t_L g1072 ( 
.A(n_657),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_222),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_708),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_246),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_353),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_373),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_847),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_531),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_85),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_503),
.Y(n_1081)
);

BUFx2_ASAP7_75t_R g1082 ( 
.A(n_795),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_830),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_795),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_472),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_165),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_627),
.Y(n_1087)
);

CKINVDCx20_ASAP7_75t_R g1088 ( 
.A(n_771),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_9),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_68),
.Y(n_1090)
);

CKINVDCx20_ASAP7_75t_R g1091 ( 
.A(n_50),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_289),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_615),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_250),
.Y(n_1094)
);

BUFx3_ASAP7_75t_L g1095 ( 
.A(n_403),
.Y(n_1095)
);

BUFx3_ASAP7_75t_L g1096 ( 
.A(n_640),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_767),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_772),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_440),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_926),
.Y(n_1100)
);

CKINVDCx16_ASAP7_75t_R g1101 ( 
.A(n_740),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_856),
.Y(n_1102)
);

INVx1_ASAP7_75t_SL g1103 ( 
.A(n_668),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_8),
.Y(n_1104)
);

BUFx8_ASAP7_75t_SL g1105 ( 
.A(n_537),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_469),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_834),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_482),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_226),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_250),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_322),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_216),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_943),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_665),
.Y(n_1114)
);

CKINVDCx20_ASAP7_75t_R g1115 ( 
.A(n_725),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_865),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_932),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_727),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_557),
.Y(n_1119)
);

CKINVDCx20_ASAP7_75t_R g1120 ( 
.A(n_130),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_889),
.Y(n_1121)
);

INVx2_ASAP7_75t_SL g1122 ( 
.A(n_557),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_493),
.Y(n_1123)
);

CKINVDCx20_ASAP7_75t_R g1124 ( 
.A(n_504),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_217),
.Y(n_1125)
);

CKINVDCx20_ASAP7_75t_R g1126 ( 
.A(n_328),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_841),
.Y(n_1127)
);

INVxp67_ASAP7_75t_L g1128 ( 
.A(n_259),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_643),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_349),
.Y(n_1130)
);

BUFx3_ASAP7_75t_L g1131 ( 
.A(n_860),
.Y(n_1131)
);

CKINVDCx16_ASAP7_75t_R g1132 ( 
.A(n_716),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_941),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_670),
.Y(n_1134)
);

BUFx5_ASAP7_75t_L g1135 ( 
.A(n_225),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_904),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_103),
.Y(n_1137)
);

CKINVDCx20_ASAP7_75t_R g1138 ( 
.A(n_166),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_331),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_391),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_831),
.Y(n_1141)
);

BUFx5_ASAP7_75t_L g1142 ( 
.A(n_275),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_483),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_230),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_662),
.Y(n_1145)
);

INVx1_ASAP7_75t_SL g1146 ( 
.A(n_895),
.Y(n_1146)
);

BUFx10_ASAP7_75t_L g1147 ( 
.A(n_863),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_528),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_31),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_716),
.Y(n_1150)
);

CKINVDCx20_ASAP7_75t_R g1151 ( 
.A(n_878),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_682),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_324),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_495),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_942),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_956),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_939),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_234),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_589),
.Y(n_1159)
);

CKINVDCx20_ASAP7_75t_R g1160 ( 
.A(n_818),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_365),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_945),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_846),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_697),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_486),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_664),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_441),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_920),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_836),
.Y(n_1169)
);

BUFx2_ASAP7_75t_L g1170 ( 
.A(n_912),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_217),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_833),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_247),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_770),
.Y(n_1174)
);

BUFx3_ASAP7_75t_L g1175 ( 
.A(n_411),
.Y(n_1175)
);

CKINVDCx20_ASAP7_75t_R g1176 ( 
.A(n_880),
.Y(n_1176)
);

BUFx3_ASAP7_75t_L g1177 ( 
.A(n_66),
.Y(n_1177)
);

BUFx2_ASAP7_75t_L g1178 ( 
.A(n_155),
.Y(n_1178)
);

BUFx3_ASAP7_75t_L g1179 ( 
.A(n_444),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_822),
.Y(n_1180)
);

CKINVDCx20_ASAP7_75t_R g1181 ( 
.A(n_890),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_86),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_887),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_98),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_384),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_311),
.Y(n_1186)
);

CKINVDCx20_ASAP7_75t_R g1187 ( 
.A(n_340),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_542),
.Y(n_1188)
);

BUFx5_ASAP7_75t_L g1189 ( 
.A(n_304),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_381),
.Y(n_1190)
);

CKINVDCx20_ASAP7_75t_R g1191 ( 
.A(n_130),
.Y(n_1191)
);

BUFx10_ASAP7_75t_L g1192 ( 
.A(n_866),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_216),
.Y(n_1193)
);

INVx2_ASAP7_75t_SL g1194 ( 
.A(n_390),
.Y(n_1194)
);

INVx3_ASAP7_75t_L g1195 ( 
.A(n_539),
.Y(n_1195)
);

INVx1_ASAP7_75t_SL g1196 ( 
.A(n_953),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_879),
.Y(n_1197)
);

CKINVDCx20_ASAP7_75t_R g1198 ( 
.A(n_427),
.Y(n_1198)
);

BUFx8_ASAP7_75t_SL g1199 ( 
.A(n_120),
.Y(n_1199)
);

CKINVDCx20_ASAP7_75t_R g1200 ( 
.A(n_905),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_269),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_399),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_289),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_733),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_872),
.Y(n_1205)
);

CKINVDCx20_ASAP7_75t_R g1206 ( 
.A(n_773),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_496),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_511),
.Y(n_1208)
);

CKINVDCx14_ASAP7_75t_R g1209 ( 
.A(n_419),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_204),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_806),
.Y(n_1211)
);

BUFx2_ASAP7_75t_L g1212 ( 
.A(n_377),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_864),
.Y(n_1213)
);

BUFx5_ASAP7_75t_L g1214 ( 
.A(n_922),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_404),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_562),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_824),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_586),
.Y(n_1218)
);

BUFx3_ASAP7_75t_L g1219 ( 
.A(n_202),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_55),
.Y(n_1220)
);

BUFx10_ASAP7_75t_L g1221 ( 
.A(n_931),
.Y(n_1221)
);

CKINVDCx20_ASAP7_75t_R g1222 ( 
.A(n_197),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_637),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_284),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_72),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_315),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_855),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_594),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_957),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_946),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_902),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_262),
.Y(n_1232)
);

BUFx10_ASAP7_75t_L g1233 ( 
.A(n_287),
.Y(n_1233)
);

CKINVDCx20_ASAP7_75t_R g1234 ( 
.A(n_808),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_885),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_929),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_128),
.Y(n_1237)
);

HB1xp67_ASAP7_75t_L g1238 ( 
.A(n_413),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_293),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_910),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_663),
.Y(n_1241)
);

CKINVDCx5p33_ASAP7_75t_R g1242 ( 
.A(n_742),
.Y(n_1242)
);

CKINVDCx20_ASAP7_75t_R g1243 ( 
.A(n_911),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_923),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_839),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_266),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_915),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_249),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_104),
.Y(n_1249)
);

CKINVDCx5p33_ASAP7_75t_R g1250 ( 
.A(n_433),
.Y(n_1250)
);

INVx1_ASAP7_75t_SL g1251 ( 
.A(n_918),
.Y(n_1251)
);

CKINVDCx20_ASAP7_75t_R g1252 ( 
.A(n_625),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_239),
.Y(n_1253)
);

HB1xp67_ASAP7_75t_L g1254 ( 
.A(n_483),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_292),
.Y(n_1255)
);

CKINVDCx20_ASAP7_75t_R g1256 ( 
.A(n_843),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_538),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_296),
.Y(n_1258)
);

CKINVDCx20_ASAP7_75t_R g1259 ( 
.A(n_596),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_290),
.Y(n_1260)
);

CKINVDCx5p33_ASAP7_75t_R g1261 ( 
.A(n_387),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_657),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_915),
.Y(n_1263)
);

INVx2_ASAP7_75t_L g1264 ( 
.A(n_789),
.Y(n_1264)
);

CKINVDCx20_ASAP7_75t_R g1265 ( 
.A(n_17),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_899),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_420),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_258),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_56),
.Y(n_1269)
);

CKINVDCx5p33_ASAP7_75t_R g1270 ( 
.A(n_691),
.Y(n_1270)
);

BUFx10_ASAP7_75t_L g1271 ( 
.A(n_295),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_512),
.Y(n_1272)
);

INVx2_ASAP7_75t_SL g1273 ( 
.A(n_919),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_582),
.Y(n_1274)
);

CKINVDCx5p33_ASAP7_75t_R g1275 ( 
.A(n_951),
.Y(n_1275)
);

CKINVDCx5p33_ASAP7_75t_R g1276 ( 
.A(n_684),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_488),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_898),
.Y(n_1278)
);

CKINVDCx5p33_ASAP7_75t_R g1279 ( 
.A(n_832),
.Y(n_1279)
);

CKINVDCx20_ASAP7_75t_R g1280 ( 
.A(n_565),
.Y(n_1280)
);

BUFx6f_ASAP7_75t_L g1281 ( 
.A(n_813),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_168),
.Y(n_1282)
);

CKINVDCx5p33_ASAP7_75t_R g1283 ( 
.A(n_77),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_938),
.Y(n_1284)
);

CKINVDCx5p33_ASAP7_75t_R g1285 ( 
.A(n_852),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_86),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_26),
.Y(n_1287)
);

BUFx6f_ASAP7_75t_L g1288 ( 
.A(n_890),
.Y(n_1288)
);

BUFx10_ASAP7_75t_L g1289 ( 
.A(n_921),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_51),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_315),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_292),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_929),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_848),
.Y(n_1294)
);

CKINVDCx20_ASAP7_75t_R g1295 ( 
.A(n_952),
.Y(n_1295)
);

CKINVDCx20_ASAP7_75t_R g1296 ( 
.A(n_940),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_874),
.Y(n_1297)
);

INVx2_ASAP7_75t_L g1298 ( 
.A(n_819),
.Y(n_1298)
);

CKINVDCx20_ASAP7_75t_R g1299 ( 
.A(n_580),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_388),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_630),
.Y(n_1301)
);

CKINVDCx20_ASAP7_75t_R g1302 ( 
.A(n_499),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_411),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_690),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_702),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_445),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_837),
.Y(n_1307)
);

BUFx2_ASAP7_75t_L g1308 ( 
.A(n_9),
.Y(n_1308)
);

CKINVDCx5p33_ASAP7_75t_R g1309 ( 
.A(n_84),
.Y(n_1309)
);

CKINVDCx20_ASAP7_75t_R g1310 ( 
.A(n_879),
.Y(n_1310)
);

INVx2_ASAP7_75t_SL g1311 ( 
.A(n_31),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_130),
.Y(n_1312)
);

CKINVDCx5p33_ASAP7_75t_R g1313 ( 
.A(n_496),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_863),
.Y(n_1314)
);

CKINVDCx20_ASAP7_75t_R g1315 ( 
.A(n_105),
.Y(n_1315)
);

CKINVDCx20_ASAP7_75t_R g1316 ( 
.A(n_594),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_387),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_196),
.Y(n_1318)
);

CKINVDCx5p33_ASAP7_75t_R g1319 ( 
.A(n_849),
.Y(n_1319)
);

CKINVDCx5p33_ASAP7_75t_R g1320 ( 
.A(n_89),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_432),
.Y(n_1321)
);

CKINVDCx5p33_ASAP7_75t_R g1322 ( 
.A(n_585),
.Y(n_1322)
);

CKINVDCx20_ASAP7_75t_R g1323 ( 
.A(n_814),
.Y(n_1323)
);

CKINVDCx5p33_ASAP7_75t_R g1324 ( 
.A(n_26),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_578),
.Y(n_1325)
);

CKINVDCx5p33_ASAP7_75t_R g1326 ( 
.A(n_597),
.Y(n_1326)
);

CKINVDCx5p33_ASAP7_75t_R g1327 ( 
.A(n_284),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_838),
.Y(n_1328)
);

CKINVDCx14_ASAP7_75t_R g1329 ( 
.A(n_537),
.Y(n_1329)
);

CKINVDCx5p33_ASAP7_75t_R g1330 ( 
.A(n_808),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_628),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_509),
.Y(n_1332)
);

CKINVDCx5p33_ASAP7_75t_R g1333 ( 
.A(n_169),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_557),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_513),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_406),
.Y(n_1336)
);

CKINVDCx5p33_ASAP7_75t_R g1337 ( 
.A(n_242),
.Y(n_1337)
);

BUFx10_ASAP7_75t_L g1338 ( 
.A(n_955),
.Y(n_1338)
);

CKINVDCx5p33_ASAP7_75t_R g1339 ( 
.A(n_327),
.Y(n_1339)
);

CKINVDCx5p33_ASAP7_75t_R g1340 ( 
.A(n_346),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_171),
.Y(n_1341)
);

INVx2_ASAP7_75t_L g1342 ( 
.A(n_922),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_632),
.Y(n_1343)
);

BUFx2_ASAP7_75t_L g1344 ( 
.A(n_348),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_92),
.Y(n_1345)
);

CKINVDCx20_ASAP7_75t_R g1346 ( 
.A(n_784),
.Y(n_1346)
);

BUFx3_ASAP7_75t_L g1347 ( 
.A(n_561),
.Y(n_1347)
);

CKINVDCx5p33_ASAP7_75t_R g1348 ( 
.A(n_615),
.Y(n_1348)
);

CKINVDCx5p33_ASAP7_75t_R g1349 ( 
.A(n_934),
.Y(n_1349)
);

CKINVDCx5p33_ASAP7_75t_R g1350 ( 
.A(n_182),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_897),
.Y(n_1351)
);

HB1xp67_ASAP7_75t_L g1352 ( 
.A(n_239),
.Y(n_1352)
);

CKINVDCx5p33_ASAP7_75t_R g1353 ( 
.A(n_87),
.Y(n_1353)
);

CKINVDCx5p33_ASAP7_75t_R g1354 ( 
.A(n_805),
.Y(n_1354)
);

CKINVDCx5p33_ASAP7_75t_R g1355 ( 
.A(n_150),
.Y(n_1355)
);

CKINVDCx5p33_ASAP7_75t_R g1356 ( 
.A(n_855),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1),
.Y(n_1357)
);

CKINVDCx5p33_ASAP7_75t_R g1358 ( 
.A(n_486),
.Y(n_1358)
);

BUFx10_ASAP7_75t_L g1359 ( 
.A(n_614),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_122),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_608),
.Y(n_1361)
);

CKINVDCx20_ASAP7_75t_R g1362 ( 
.A(n_935),
.Y(n_1362)
);

INVx2_ASAP7_75t_SL g1363 ( 
.A(n_778),
.Y(n_1363)
);

CKINVDCx5p33_ASAP7_75t_R g1364 ( 
.A(n_826),
.Y(n_1364)
);

CKINVDCx5p33_ASAP7_75t_R g1365 ( 
.A(n_181),
.Y(n_1365)
);

CKINVDCx5p33_ASAP7_75t_R g1366 ( 
.A(n_658),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_372),
.Y(n_1367)
);

CKINVDCx20_ASAP7_75t_R g1368 ( 
.A(n_416),
.Y(n_1368)
);

CKINVDCx5p33_ASAP7_75t_R g1369 ( 
.A(n_861),
.Y(n_1369)
);

HB1xp67_ASAP7_75t_L g1370 ( 
.A(n_823),
.Y(n_1370)
);

CKINVDCx20_ASAP7_75t_R g1371 ( 
.A(n_173),
.Y(n_1371)
);

BUFx6f_ASAP7_75t_L g1372 ( 
.A(n_19),
.Y(n_1372)
);

CKINVDCx20_ASAP7_75t_R g1373 ( 
.A(n_788),
.Y(n_1373)
);

CKINVDCx5p33_ASAP7_75t_R g1374 ( 
.A(n_205),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_828),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_393),
.Y(n_1376)
);

CKINVDCx5p33_ASAP7_75t_R g1377 ( 
.A(n_532),
.Y(n_1377)
);

CKINVDCx5p33_ASAP7_75t_R g1378 ( 
.A(n_920),
.Y(n_1378)
);

CKINVDCx5p33_ASAP7_75t_R g1379 ( 
.A(n_69),
.Y(n_1379)
);

CKINVDCx5p33_ASAP7_75t_R g1380 ( 
.A(n_924),
.Y(n_1380)
);

CKINVDCx5p33_ASAP7_75t_R g1381 ( 
.A(n_691),
.Y(n_1381)
);

CKINVDCx5p33_ASAP7_75t_R g1382 ( 
.A(n_224),
.Y(n_1382)
);

BUFx6f_ASAP7_75t_L g1383 ( 
.A(n_442),
.Y(n_1383)
);

CKINVDCx5p33_ASAP7_75t_R g1384 ( 
.A(n_900),
.Y(n_1384)
);

CKINVDCx5p33_ASAP7_75t_R g1385 ( 
.A(n_851),
.Y(n_1385)
);

CKINVDCx5p33_ASAP7_75t_R g1386 ( 
.A(n_549),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_432),
.Y(n_1387)
);

CKINVDCx5p33_ASAP7_75t_R g1388 ( 
.A(n_469),
.Y(n_1388)
);

CKINVDCx5p33_ASAP7_75t_R g1389 ( 
.A(n_831),
.Y(n_1389)
);

CKINVDCx20_ASAP7_75t_R g1390 ( 
.A(n_774),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_645),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_709),
.Y(n_1392)
);

CKINVDCx16_ASAP7_75t_R g1393 ( 
.A(n_124),
.Y(n_1393)
);

CKINVDCx5p33_ASAP7_75t_R g1394 ( 
.A(n_498),
.Y(n_1394)
);

CKINVDCx5p33_ASAP7_75t_R g1395 ( 
.A(n_914),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_56),
.Y(n_1396)
);

CKINVDCx5p33_ASAP7_75t_R g1397 ( 
.A(n_740),
.Y(n_1397)
);

CKINVDCx16_ASAP7_75t_R g1398 ( 
.A(n_877),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_854),
.Y(n_1399)
);

CKINVDCx5p33_ASAP7_75t_R g1400 ( 
.A(n_916),
.Y(n_1400)
);

CKINVDCx5p33_ASAP7_75t_R g1401 ( 
.A(n_414),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_704),
.Y(n_1402)
);

BUFx6f_ASAP7_75t_L g1403 ( 
.A(n_73),
.Y(n_1403)
);

CKINVDCx5p33_ASAP7_75t_R g1404 ( 
.A(n_871),
.Y(n_1404)
);

BUFx6f_ASAP7_75t_L g1405 ( 
.A(n_311),
.Y(n_1405)
);

CKINVDCx5p33_ASAP7_75t_R g1406 ( 
.A(n_923),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_841),
.Y(n_1407)
);

CKINVDCx5p33_ASAP7_75t_R g1408 ( 
.A(n_867),
.Y(n_1408)
);

CKINVDCx5p33_ASAP7_75t_R g1409 ( 
.A(n_774),
.Y(n_1409)
);

CKINVDCx5p33_ASAP7_75t_R g1410 ( 
.A(n_159),
.Y(n_1410)
);

CKINVDCx5p33_ASAP7_75t_R g1411 ( 
.A(n_539),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_937),
.Y(n_1412)
);

CKINVDCx5p33_ASAP7_75t_R g1413 ( 
.A(n_815),
.Y(n_1413)
);

CKINVDCx5p33_ASAP7_75t_R g1414 ( 
.A(n_894),
.Y(n_1414)
);

CKINVDCx5p33_ASAP7_75t_R g1415 ( 
.A(n_886),
.Y(n_1415)
);

BUFx10_ASAP7_75t_L g1416 ( 
.A(n_442),
.Y(n_1416)
);

CKINVDCx5p33_ASAP7_75t_R g1417 ( 
.A(n_842),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_159),
.Y(n_1418)
);

CKINVDCx5p33_ASAP7_75t_R g1419 ( 
.A(n_902),
.Y(n_1419)
);

CKINVDCx5p33_ASAP7_75t_R g1420 ( 
.A(n_892),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_542),
.Y(n_1421)
);

CKINVDCx5p33_ASAP7_75t_R g1422 ( 
.A(n_664),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_179),
.Y(n_1423)
);

CKINVDCx5p33_ASAP7_75t_R g1424 ( 
.A(n_508),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_713),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_781),
.Y(n_1426)
);

CKINVDCx5p33_ASAP7_75t_R g1427 ( 
.A(n_593),
.Y(n_1427)
);

CKINVDCx5p33_ASAP7_75t_R g1428 ( 
.A(n_606),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_248),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_711),
.Y(n_1430)
);

CKINVDCx20_ASAP7_75t_R g1431 ( 
.A(n_888),
.Y(n_1431)
);

CKINVDCx20_ASAP7_75t_R g1432 ( 
.A(n_285),
.Y(n_1432)
);

CKINVDCx5p33_ASAP7_75t_R g1433 ( 
.A(n_385),
.Y(n_1433)
);

CKINVDCx5p33_ASAP7_75t_R g1434 ( 
.A(n_544),
.Y(n_1434)
);

CKINVDCx14_ASAP7_75t_R g1435 ( 
.A(n_158),
.Y(n_1435)
);

CKINVDCx5p33_ASAP7_75t_R g1436 ( 
.A(n_909),
.Y(n_1436)
);

CKINVDCx5p33_ASAP7_75t_R g1437 ( 
.A(n_108),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_388),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_79),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_587),
.Y(n_1440)
);

CKINVDCx5p33_ASAP7_75t_R g1441 ( 
.A(n_906),
.Y(n_1441)
);

CKINVDCx16_ASAP7_75t_R g1442 ( 
.A(n_824),
.Y(n_1442)
);

CKINVDCx5p33_ASAP7_75t_R g1443 ( 
.A(n_917),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_769),
.Y(n_1444)
);

CKINVDCx5p33_ASAP7_75t_R g1445 ( 
.A(n_883),
.Y(n_1445)
);

CKINVDCx5p33_ASAP7_75t_R g1446 ( 
.A(n_793),
.Y(n_1446)
);

BUFx3_ASAP7_75t_L g1447 ( 
.A(n_903),
.Y(n_1447)
);

INVxp67_ASAP7_75t_L g1448 ( 
.A(n_946),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_807),
.Y(n_1449)
);

CKINVDCx5p33_ASAP7_75t_R g1450 ( 
.A(n_366),
.Y(n_1450)
);

CKINVDCx5p33_ASAP7_75t_R g1451 ( 
.A(n_812),
.Y(n_1451)
);

CKINVDCx5p33_ASAP7_75t_R g1452 ( 
.A(n_636),
.Y(n_1452)
);

INVxp67_ASAP7_75t_SL g1453 ( 
.A(n_458),
.Y(n_1453)
);

CKINVDCx14_ASAP7_75t_R g1454 ( 
.A(n_862),
.Y(n_1454)
);

CKINVDCx20_ASAP7_75t_R g1455 ( 
.A(n_462),
.Y(n_1455)
);

BUFx6f_ASAP7_75t_L g1456 ( 
.A(n_536),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_925),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_65),
.Y(n_1458)
);

CKINVDCx5p33_ASAP7_75t_R g1459 ( 
.A(n_781),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_156),
.Y(n_1460)
);

INVx1_ASAP7_75t_SL g1461 ( 
.A(n_569),
.Y(n_1461)
);

CKINVDCx5p33_ASAP7_75t_R g1462 ( 
.A(n_658),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_884),
.Y(n_1463)
);

CKINVDCx5p33_ASAP7_75t_R g1464 ( 
.A(n_355),
.Y(n_1464)
);

CKINVDCx5p33_ASAP7_75t_R g1465 ( 
.A(n_811),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_47),
.Y(n_1466)
);

CKINVDCx5p33_ASAP7_75t_R g1467 ( 
.A(n_665),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_844),
.Y(n_1468)
);

CKINVDCx5p33_ASAP7_75t_R g1469 ( 
.A(n_868),
.Y(n_1469)
);

BUFx6f_ASAP7_75t_L g1470 ( 
.A(n_12),
.Y(n_1470)
);

CKINVDCx5p33_ASAP7_75t_R g1471 ( 
.A(n_816),
.Y(n_1471)
);

CKINVDCx5p33_ASAP7_75t_R g1472 ( 
.A(n_770),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_519),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_741),
.Y(n_1474)
);

CKINVDCx5p33_ASAP7_75t_R g1475 ( 
.A(n_514),
.Y(n_1475)
);

CKINVDCx5p33_ASAP7_75t_R g1476 ( 
.A(n_428),
.Y(n_1476)
);

INVx2_ASAP7_75t_SL g1477 ( 
.A(n_426),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_875),
.Y(n_1478)
);

CKINVDCx20_ASAP7_75t_R g1479 ( 
.A(n_141),
.Y(n_1479)
);

BUFx10_ASAP7_75t_L g1480 ( 
.A(n_840),
.Y(n_1480)
);

CKINVDCx5p33_ASAP7_75t_R g1481 ( 
.A(n_313),
.Y(n_1481)
);

CKINVDCx5p33_ASAP7_75t_R g1482 ( 
.A(n_748),
.Y(n_1482)
);

CKINVDCx5p33_ASAP7_75t_R g1483 ( 
.A(n_294),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_876),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_433),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_820),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_347),
.Y(n_1487)
);

CKINVDCx5p33_ASAP7_75t_R g1488 ( 
.A(n_68),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_857),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_532),
.Y(n_1490)
);

CKINVDCx5p33_ASAP7_75t_R g1491 ( 
.A(n_585),
.Y(n_1491)
);

CKINVDCx5p33_ASAP7_75t_R g1492 ( 
.A(n_858),
.Y(n_1492)
);

CKINVDCx5p33_ASAP7_75t_R g1493 ( 
.A(n_821),
.Y(n_1493)
);

CKINVDCx5p33_ASAP7_75t_R g1494 ( 
.A(n_104),
.Y(n_1494)
);

CKINVDCx5p33_ASAP7_75t_R g1495 ( 
.A(n_843),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_711),
.Y(n_1496)
);

CKINVDCx5p33_ASAP7_75t_R g1497 ( 
.A(n_311),
.Y(n_1497)
);

CKINVDCx5p33_ASAP7_75t_R g1498 ( 
.A(n_810),
.Y(n_1498)
);

BUFx5_ASAP7_75t_L g1499 ( 
.A(n_44),
.Y(n_1499)
);

CKINVDCx5p33_ASAP7_75t_R g1500 ( 
.A(n_590),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_729),
.Y(n_1501)
);

CKINVDCx5p33_ASAP7_75t_R g1502 ( 
.A(n_881),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_930),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_764),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_171),
.Y(n_1505)
);

CKINVDCx5p33_ASAP7_75t_R g1506 ( 
.A(n_97),
.Y(n_1506)
);

CKINVDCx5p33_ASAP7_75t_R g1507 ( 
.A(n_742),
.Y(n_1507)
);

CKINVDCx5p33_ASAP7_75t_R g1508 ( 
.A(n_913),
.Y(n_1508)
);

INVx1_ASAP7_75t_SL g1509 ( 
.A(n_827),
.Y(n_1509)
);

CKINVDCx5p33_ASAP7_75t_R g1510 ( 
.A(n_383),
.Y(n_1510)
);

CKINVDCx5p33_ASAP7_75t_R g1511 ( 
.A(n_452),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_928),
.Y(n_1512)
);

CKINVDCx5p33_ASAP7_75t_R g1513 ( 
.A(n_455),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_265),
.Y(n_1514)
);

CKINVDCx20_ASAP7_75t_R g1515 ( 
.A(n_829),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_871),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_75),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_634),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_564),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_884),
.Y(n_1520)
);

CKINVDCx20_ASAP7_75t_R g1521 ( 
.A(n_366),
.Y(n_1521)
);

CKINVDCx20_ASAP7_75t_R g1522 ( 
.A(n_249),
.Y(n_1522)
);

CKINVDCx5p33_ASAP7_75t_R g1523 ( 
.A(n_106),
.Y(n_1523)
);

CKINVDCx5p33_ASAP7_75t_R g1524 ( 
.A(n_313),
.Y(n_1524)
);

CKINVDCx5p33_ASAP7_75t_R g1525 ( 
.A(n_401),
.Y(n_1525)
);

BUFx8_ASAP7_75t_SL g1526 ( 
.A(n_943),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_210),
.Y(n_1527)
);

INVx2_ASAP7_75t_SL g1528 ( 
.A(n_746),
.Y(n_1528)
);

BUFx10_ASAP7_75t_L g1529 ( 
.A(n_835),
.Y(n_1529)
);

CKINVDCx5p33_ASAP7_75t_R g1530 ( 
.A(n_263),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_681),
.Y(n_1531)
);

CKINVDCx5p33_ASAP7_75t_R g1532 ( 
.A(n_936),
.Y(n_1532)
);

CKINVDCx5p33_ASAP7_75t_R g1533 ( 
.A(n_414),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_927),
.Y(n_1534)
);

INVxp67_ASAP7_75t_L g1535 ( 
.A(n_763),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1042),
.Y(n_1536)
);

INVxp67_ASAP7_75t_SL g1537 ( 
.A(n_1006),
.Y(n_1537)
);

INVxp67_ASAP7_75t_SL g1538 ( 
.A(n_1006),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1214),
.Y(n_1539)
);

NOR2xp33_ASAP7_75t_L g1540 ( 
.A(n_1178),
.B(n_0),
.Y(n_1540)
);

INVxp67_ASAP7_75t_L g1541 ( 
.A(n_1212),
.Y(n_1541)
);

CKINVDCx5p33_ASAP7_75t_R g1542 ( 
.A(n_1209),
.Y(n_1542)
);

INVxp67_ASAP7_75t_L g1543 ( 
.A(n_1308),
.Y(n_1543)
);

INVxp33_ASAP7_75t_SL g1544 ( 
.A(n_1061),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1214),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1065),
.Y(n_1546)
);

CKINVDCx20_ASAP7_75t_R g1547 ( 
.A(n_1105),
.Y(n_1547)
);

NOR2xp33_ASAP7_75t_L g1548 ( 
.A(n_1344),
.B(n_1),
.Y(n_1548)
);

CKINVDCx5p33_ASAP7_75t_R g1549 ( 
.A(n_1209),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1122),
.Y(n_1550)
);

CKINVDCx5p33_ASAP7_75t_R g1551 ( 
.A(n_1329),
.Y(n_1551)
);

INVxp67_ASAP7_75t_L g1552 ( 
.A(n_1238),
.Y(n_1552)
);

CKINVDCx5p33_ASAP7_75t_R g1553 ( 
.A(n_1329),
.Y(n_1553)
);

CKINVDCx5p33_ASAP7_75t_R g1554 ( 
.A(n_1435),
.Y(n_1554)
);

CKINVDCx20_ASAP7_75t_R g1555 ( 
.A(n_1105),
.Y(n_1555)
);

NOR2xp33_ASAP7_75t_L g1556 ( 
.A(n_969),
.B(n_1),
.Y(n_1556)
);

CKINVDCx20_ASAP7_75t_R g1557 ( 
.A(n_1199),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1194),
.Y(n_1558)
);

CKINVDCx5p33_ASAP7_75t_R g1559 ( 
.A(n_1435),
.Y(n_1559)
);

CKINVDCx5p33_ASAP7_75t_R g1560 ( 
.A(n_1199),
.Y(n_1560)
);

INVxp33_ASAP7_75t_SL g1561 ( 
.A(n_1254),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1311),
.Y(n_1562)
);

CKINVDCx20_ASAP7_75t_R g1563 ( 
.A(n_1023),
.Y(n_1563)
);

CKINVDCx20_ASAP7_75t_R g1564 ( 
.A(n_1091),
.Y(n_1564)
);

CKINVDCx16_ASAP7_75t_R g1565 ( 
.A(n_1393),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1477),
.Y(n_1566)
);

CKINVDCx20_ASAP7_75t_R g1567 ( 
.A(n_1120),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1195),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1352),
.B(n_2),
.Y(n_1569)
);

CKINVDCx16_ASAP7_75t_R g1570 ( 
.A(n_1037),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1195),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_958),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_964),
.Y(n_1573)
);

CKINVDCx5p33_ASAP7_75t_R g1574 ( 
.A(n_1454),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_970),
.Y(n_1575)
);

CKINVDCx5p33_ASAP7_75t_R g1576 ( 
.A(n_1454),
.Y(n_1576)
);

INVxp67_ASAP7_75t_L g1577 ( 
.A(n_1002),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1170),
.B(n_2),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_972),
.Y(n_1579)
);

CKINVDCx5p33_ASAP7_75t_R g1580 ( 
.A(n_1526),
.Y(n_1580)
);

CKINVDCx20_ASAP7_75t_R g1581 ( 
.A(n_1124),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_987),
.Y(n_1582)
);

CKINVDCx5p33_ASAP7_75t_R g1583 ( 
.A(n_1526),
.Y(n_1583)
);

CKINVDCx20_ASAP7_75t_R g1584 ( 
.A(n_1126),
.Y(n_1584)
);

HB1xp67_ASAP7_75t_L g1585 ( 
.A(n_1370),
.Y(n_1585)
);

CKINVDCx5p33_ASAP7_75t_R g1586 ( 
.A(n_960),
.Y(n_1586)
);

CKINVDCx20_ASAP7_75t_R g1587 ( 
.A(n_1138),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_990),
.Y(n_1588)
);

INVxp67_ASAP7_75t_L g1589 ( 
.A(n_1037),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_998),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1015),
.Y(n_1591)
);

CKINVDCx5p33_ASAP7_75t_R g1592 ( 
.A(n_962),
.Y(n_1592)
);

CKINVDCx20_ASAP7_75t_R g1593 ( 
.A(n_1187),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1019),
.Y(n_1594)
);

BUFx6f_ASAP7_75t_SL g1595 ( 
.A(n_1037),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1040),
.Y(n_1596)
);

CKINVDCx5p33_ASAP7_75t_R g1597 ( 
.A(n_976),
.Y(n_1597)
);

NOR2xp33_ASAP7_75t_L g1598 ( 
.A(n_1273),
.B(n_2),
.Y(n_1598)
);

INVxp33_ASAP7_75t_L g1599 ( 
.A(n_963),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1041),
.Y(n_1600)
);

HB1xp67_ASAP7_75t_L g1601 ( 
.A(n_1021),
.Y(n_1601)
);

CKINVDCx20_ASAP7_75t_R g1602 ( 
.A(n_1191),
.Y(n_1602)
);

CKINVDCx20_ASAP7_75t_R g1603 ( 
.A(n_1198),
.Y(n_1603)
);

CKINVDCx20_ASAP7_75t_R g1604 ( 
.A(n_1222),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1363),
.B(n_3),
.Y(n_1605)
);

INVxp67_ASAP7_75t_SL g1606 ( 
.A(n_973),
.Y(n_1606)
);

CKINVDCx5p33_ASAP7_75t_R g1607 ( 
.A(n_977),
.Y(n_1607)
);

CKINVDCx5p33_ASAP7_75t_R g1608 ( 
.A(n_978),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1045),
.Y(n_1609)
);

CKINVDCx20_ASAP7_75t_R g1610 ( 
.A(n_1252),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1053),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1060),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1068),
.Y(n_1613)
);

CKINVDCx5p33_ASAP7_75t_R g1614 ( 
.A(n_982),
.Y(n_1614)
);

INVxp67_ASAP7_75t_L g1615 ( 
.A(n_1233),
.Y(n_1615)
);

INVxp67_ASAP7_75t_SL g1616 ( 
.A(n_973),
.Y(n_1616)
);

CKINVDCx5p33_ASAP7_75t_R g1617 ( 
.A(n_988),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1070),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1076),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1092),
.Y(n_1620)
);

CKINVDCx16_ASAP7_75t_R g1621 ( 
.A(n_1233),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1099),
.Y(n_1622)
);

CKINVDCx20_ASAP7_75t_R g1623 ( 
.A(n_1259),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1129),
.Y(n_1624)
);

CKINVDCx5p33_ASAP7_75t_R g1625 ( 
.A(n_995),
.Y(n_1625)
);

INVxp33_ASAP7_75t_SL g1626 ( 
.A(n_996),
.Y(n_1626)
);

CKINVDCx20_ASAP7_75t_R g1627 ( 
.A(n_1265),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1134),
.Y(n_1628)
);

INVxp67_ASAP7_75t_L g1629 ( 
.A(n_1233),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1137),
.Y(n_1630)
);

CKINVDCx20_ASAP7_75t_R g1631 ( 
.A(n_1280),
.Y(n_1631)
);

CKINVDCx5p33_ASAP7_75t_R g1632 ( 
.A(n_997),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1528),
.B(n_3),
.Y(n_1633)
);

INVxp67_ASAP7_75t_SL g1634 ( 
.A(n_1025),
.Y(n_1634)
);

CKINVDCx16_ASAP7_75t_R g1635 ( 
.A(n_1271),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1139),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1158),
.Y(n_1637)
);

CKINVDCx5p33_ASAP7_75t_R g1638 ( 
.A(n_1005),
.Y(n_1638)
);

CKINVDCx20_ASAP7_75t_R g1639 ( 
.A(n_1299),
.Y(n_1639)
);

BUFx3_ASAP7_75t_L g1640 ( 
.A(n_1025),
.Y(n_1640)
);

CKINVDCx20_ASAP7_75t_R g1641 ( 
.A(n_1302),
.Y(n_1641)
);

CKINVDCx5p33_ASAP7_75t_R g1642 ( 
.A(n_1009),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1166),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1167),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1173),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1182),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1184),
.Y(n_1647)
);

CKINVDCx5p33_ASAP7_75t_R g1648 ( 
.A(n_1010),
.Y(n_1648)
);

CKINVDCx16_ASAP7_75t_R g1649 ( 
.A(n_1271),
.Y(n_1649)
);

CKINVDCx5p33_ASAP7_75t_R g1650 ( 
.A(n_1012),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1185),
.Y(n_1651)
);

CKINVDCx5p33_ASAP7_75t_R g1652 ( 
.A(n_1013),
.Y(n_1652)
);

CKINVDCx5p33_ASAP7_75t_R g1653 ( 
.A(n_1017),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1214),
.Y(n_1654)
);

INVxp33_ASAP7_75t_SL g1655 ( 
.A(n_1022),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1193),
.Y(n_1656)
);

CKINVDCx5p33_ASAP7_75t_R g1657 ( 
.A(n_1028),
.Y(n_1657)
);

CKINVDCx5p33_ASAP7_75t_R g1658 ( 
.A(n_1029),
.Y(n_1658)
);

CKINVDCx5p33_ASAP7_75t_R g1659 ( 
.A(n_1033),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1201),
.Y(n_1660)
);

CKINVDCx5p33_ASAP7_75t_R g1661 ( 
.A(n_1035),
.Y(n_1661)
);

NOR2xp33_ASAP7_75t_L g1662 ( 
.A(n_1448),
.B(n_3),
.Y(n_1662)
);

CKINVDCx20_ASAP7_75t_R g1663 ( 
.A(n_1315),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1038),
.B(n_4),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1640),
.Y(n_1665)
);

BUFx6f_ASAP7_75t_L g1666 ( 
.A(n_1640),
.Y(n_1666)
);

INVxp67_ASAP7_75t_L g1667 ( 
.A(n_1537),
.Y(n_1667)
);

INVx3_ASAP7_75t_L g1668 ( 
.A(n_1570),
.Y(n_1668)
);

OAI21x1_ASAP7_75t_L g1669 ( 
.A1(n_1539),
.A2(n_1057),
.B(n_1054),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_1545),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_SL g1671 ( 
.A(n_1621),
.B(n_991),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1654),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1568),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1571),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1606),
.Y(n_1675)
);

OA21x2_ASAP7_75t_L g1676 ( 
.A1(n_1572),
.A2(n_1057),
.B(n_1054),
.Y(n_1676)
);

BUFx6f_ASAP7_75t_L g1677 ( 
.A(n_1536),
.Y(n_1677)
);

BUFx3_ASAP7_75t_L g1678 ( 
.A(n_1546),
.Y(n_1678)
);

INVx3_ASAP7_75t_L g1679 ( 
.A(n_1635),
.Y(n_1679)
);

INVx2_ASAP7_75t_L g1680 ( 
.A(n_1550),
.Y(n_1680)
);

CKINVDCx5p33_ASAP7_75t_R g1681 ( 
.A(n_1595),
.Y(n_1681)
);

INVx2_ASAP7_75t_L g1682 ( 
.A(n_1558),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1562),
.Y(n_1683)
);

HB1xp67_ASAP7_75t_L g1684 ( 
.A(n_1649),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1616),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_1566),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1538),
.B(n_1271),
.Y(n_1687)
);

BUFx6f_ASAP7_75t_L g1688 ( 
.A(n_1573),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1552),
.B(n_1047),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1575),
.Y(n_1690)
);

INVx2_ASAP7_75t_L g1691 ( 
.A(n_1579),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1589),
.B(n_1615),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1634),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1605),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1633),
.Y(n_1695)
);

HB1xp67_ASAP7_75t_L g1696 ( 
.A(n_1586),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1582),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1588),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1590),
.Y(n_1699)
);

OA21x2_ASAP7_75t_L g1700 ( 
.A1(n_1591),
.A2(n_1125),
.B(n_1109),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1594),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1596),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1600),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1609),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1611),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1612),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1613),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1618),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1541),
.B(n_1359),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1619),
.Y(n_1710)
);

INVx3_ASAP7_75t_L g1711 ( 
.A(n_1595),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1620),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1622),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_1624),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1628),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1629),
.B(n_1049),
.Y(n_1716)
);

HB1xp67_ASAP7_75t_L g1717 ( 
.A(n_1592),
.Y(n_1717)
);

OA21x2_ASAP7_75t_L g1718 ( 
.A1(n_1630),
.A2(n_1125),
.B(n_1109),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1636),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1543),
.B(n_1064),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1601),
.B(n_1585),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1637),
.Y(n_1722)
);

NOR2xp33_ASAP7_75t_L g1723 ( 
.A(n_1626),
.B(n_1535),
.Y(n_1723)
);

BUFx6f_ASAP7_75t_L g1724 ( 
.A(n_1643),
.Y(n_1724)
);

BUFx6f_ASAP7_75t_L g1725 ( 
.A(n_1644),
.Y(n_1725)
);

BUFx8_ASAP7_75t_L g1726 ( 
.A(n_1569),
.Y(n_1726)
);

BUFx6f_ASAP7_75t_L g1727 ( 
.A(n_1645),
.Y(n_1727)
);

AND2x4_ASAP7_75t_L g1728 ( 
.A(n_1577),
.B(n_1131),
.Y(n_1728)
);

INVx3_ASAP7_75t_L g1729 ( 
.A(n_1646),
.Y(n_1729)
);

INVx2_ASAP7_75t_L g1730 ( 
.A(n_1647),
.Y(n_1730)
);

BUFx6f_ASAP7_75t_L g1731 ( 
.A(n_1651),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1656),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1660),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1556),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1556),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1598),
.Y(n_1736)
);

AND2x4_ASAP7_75t_L g1737 ( 
.A(n_1542),
.B(n_1549),
.Y(n_1737)
);

AND2x4_ASAP7_75t_L g1738 ( 
.A(n_1551),
.B(n_1131),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1544),
.B(n_1066),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1598),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1662),
.Y(n_1741)
);

INVx3_ASAP7_75t_L g1742 ( 
.A(n_1597),
.Y(n_1742)
);

INVxp33_ASAP7_75t_SL g1743 ( 
.A(n_1553),
.Y(n_1743)
);

NAND2xp33_ASAP7_75t_SL g1744 ( 
.A(n_1554),
.B(n_1067),
.Y(n_1744)
);

INVx2_ASAP7_75t_L g1745 ( 
.A(n_1664),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1561),
.B(n_1073),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1662),
.Y(n_1747)
);

INVx3_ASAP7_75t_L g1748 ( 
.A(n_1607),
.Y(n_1748)
);

INVx3_ASAP7_75t_L g1749 ( 
.A(n_1608),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1559),
.B(n_1075),
.Y(n_1750)
);

NOR2xp33_ASAP7_75t_L g1751 ( 
.A(n_1655),
.B(n_1101),
.Y(n_1751)
);

BUFx2_ASAP7_75t_L g1752 ( 
.A(n_1614),
.Y(n_1752)
);

AND2x4_ASAP7_75t_L g1753 ( 
.A(n_1574),
.B(n_1447),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1565),
.B(n_1359),
.Y(n_1754)
);

BUFx6f_ASAP7_75t_L g1755 ( 
.A(n_1578),
.Y(n_1755)
);

AND2x4_ASAP7_75t_L g1756 ( 
.A(n_1576),
.B(n_1447),
.Y(n_1756)
);

BUFx6f_ASAP7_75t_L g1757 ( 
.A(n_1617),
.Y(n_1757)
);

INVx4_ASAP7_75t_L g1758 ( 
.A(n_1625),
.Y(n_1758)
);

INVx4_ASAP7_75t_L g1759 ( 
.A(n_1632),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1540),
.Y(n_1760)
);

HB1xp67_ASAP7_75t_L g1761 ( 
.A(n_1638),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1599),
.B(n_1359),
.Y(n_1762)
);

BUFx6f_ASAP7_75t_L g1763 ( 
.A(n_1642),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1540),
.Y(n_1764)
);

INVx2_ASAP7_75t_L g1765 ( 
.A(n_1548),
.Y(n_1765)
);

BUFx2_ASAP7_75t_L g1766 ( 
.A(n_1648),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1548),
.Y(n_1767)
);

BUFx6f_ASAP7_75t_L g1768 ( 
.A(n_1650),
.Y(n_1768)
);

NOR2xp33_ASAP7_75t_L g1769 ( 
.A(n_1652),
.B(n_1132),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1653),
.Y(n_1770)
);

AND2x4_ASAP7_75t_L g1771 ( 
.A(n_1657),
.B(n_1658),
.Y(n_1771)
);

BUFx6f_ASAP7_75t_L g1772 ( 
.A(n_1659),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1661),
.Y(n_1773)
);

BUFx6f_ASAP7_75t_L g1774 ( 
.A(n_1560),
.Y(n_1774)
);

INVx3_ASAP7_75t_L g1775 ( 
.A(n_1580),
.Y(n_1775)
);

CKINVDCx16_ASAP7_75t_R g1776 ( 
.A(n_1547),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1583),
.Y(n_1777)
);

AND3x2_ASAP7_75t_L g1778 ( 
.A(n_1555),
.B(n_1082),
.C(n_1036),
.Y(n_1778)
);

AND2x4_ASAP7_75t_L g1779 ( 
.A(n_1563),
.B(n_1095),
.Y(n_1779)
);

INVx2_ASAP7_75t_L g1780 ( 
.A(n_1557),
.Y(n_1780)
);

INVx2_ASAP7_75t_L g1781 ( 
.A(n_1564),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1567),
.B(n_1416),
.Y(n_1782)
);

INVx2_ASAP7_75t_L g1783 ( 
.A(n_1581),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1584),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1587),
.B(n_1077),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1593),
.Y(n_1786)
);

AND2x6_ASAP7_75t_L g1787 ( 
.A(n_1602),
.B(n_1095),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1603),
.B(n_1079),
.Y(n_1788)
);

BUFx3_ASAP7_75t_L g1789 ( 
.A(n_1604),
.Y(n_1789)
);

NOR2xp33_ASAP7_75t_L g1790 ( 
.A(n_1610),
.B(n_1398),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1623),
.Y(n_1791)
);

BUFx6f_ASAP7_75t_L g1792 ( 
.A(n_1627),
.Y(n_1792)
);

BUFx6f_ASAP7_75t_L g1793 ( 
.A(n_1631),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1639),
.B(n_1080),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1641),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1663),
.B(n_1081),
.Y(n_1796)
);

INVx2_ASAP7_75t_L g1797 ( 
.A(n_1640),
.Y(n_1797)
);

BUFx6f_ASAP7_75t_L g1798 ( 
.A(n_1640),
.Y(n_1798)
);

BUFx6f_ASAP7_75t_L g1799 ( 
.A(n_1640),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1537),
.B(n_1085),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1539),
.Y(n_1801)
);

INVx2_ASAP7_75t_L g1802 ( 
.A(n_1640),
.Y(n_1802)
);

BUFx6f_ASAP7_75t_L g1803 ( 
.A(n_1640),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1539),
.Y(n_1804)
);

INVx3_ASAP7_75t_L g1805 ( 
.A(n_1570),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1539),
.Y(n_1806)
);

NOR2xp33_ASAP7_75t_L g1807 ( 
.A(n_1536),
.B(n_1442),
.Y(n_1807)
);

INVx3_ASAP7_75t_L g1808 ( 
.A(n_1570),
.Y(n_1808)
);

INVx2_ASAP7_75t_L g1809 ( 
.A(n_1640),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1539),
.Y(n_1810)
);

INVx2_ASAP7_75t_L g1811 ( 
.A(n_1640),
.Y(n_1811)
);

INVx2_ASAP7_75t_L g1812 ( 
.A(n_1640),
.Y(n_1812)
);

BUFx6f_ASAP7_75t_L g1813 ( 
.A(n_1640),
.Y(n_1813)
);

INVx2_ASAP7_75t_L g1814 ( 
.A(n_1640),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1537),
.Y(n_1815)
);

BUFx6f_ASAP7_75t_L g1816 ( 
.A(n_1640),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1537),
.Y(n_1817)
);

BUFx6f_ASAP7_75t_L g1818 ( 
.A(n_1640),
.Y(n_1818)
);

BUFx6f_ASAP7_75t_L g1819 ( 
.A(n_1640),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1537),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_L g1821 ( 
.A(n_1537),
.B(n_1086),
.Y(n_1821)
);

INVx2_ASAP7_75t_L g1822 ( 
.A(n_1640),
.Y(n_1822)
);

BUFx6f_ASAP7_75t_L g1823 ( 
.A(n_1640),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1539),
.Y(n_1824)
);

OAI22xp5_ASAP7_75t_L g1825 ( 
.A1(n_1537),
.A2(n_1089),
.B1(n_1090),
.B2(n_1087),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1640),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1539),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1539),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1539),
.Y(n_1829)
);

NOR2xp33_ASAP7_75t_L g1830 ( 
.A(n_1536),
.B(n_1128),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1537),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1537),
.Y(n_1832)
);

BUFx6f_ASAP7_75t_L g1833 ( 
.A(n_1640),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1537),
.B(n_1093),
.Y(n_1834)
);

BUFx6f_ASAP7_75t_L g1835 ( 
.A(n_1640),
.Y(n_1835)
);

AND2x4_ASAP7_75t_L g1836 ( 
.A(n_1537),
.B(n_1096),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1537),
.Y(n_1837)
);

INVx2_ASAP7_75t_L g1838 ( 
.A(n_1640),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_L g1839 ( 
.A(n_1537),
.B(n_1094),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1537),
.Y(n_1840)
);

OR2x6_ASAP7_75t_L g1841 ( 
.A(n_1541),
.B(n_986),
.Y(n_1841)
);

AND2x4_ASAP7_75t_L g1842 ( 
.A(n_1537),
.B(n_1175),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1537),
.B(n_1104),
.Y(n_1843)
);

INVx4_ASAP7_75t_L g1844 ( 
.A(n_1595),
.Y(n_1844)
);

BUFx2_ASAP7_75t_L g1845 ( 
.A(n_1537),
.Y(n_1845)
);

BUFx3_ASAP7_75t_L g1846 ( 
.A(n_1640),
.Y(n_1846)
);

AND2x4_ASAP7_75t_L g1847 ( 
.A(n_1537),
.B(n_1175),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1537),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1537),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1537),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1537),
.Y(n_1851)
);

INVx2_ASAP7_75t_L g1852 ( 
.A(n_1640),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1537),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1537),
.Y(n_1854)
);

AND2x4_ASAP7_75t_L g1855 ( 
.A(n_1537),
.B(n_1177),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1537),
.Y(n_1856)
);

INVx3_ASAP7_75t_L g1857 ( 
.A(n_1570),
.Y(n_1857)
);

OA21x2_ASAP7_75t_L g1858 ( 
.A1(n_1539),
.A2(n_1239),
.B(n_1159),
.Y(n_1858)
);

BUFx2_ASAP7_75t_L g1859 ( 
.A(n_1537),
.Y(n_1859)
);

INVx2_ASAP7_75t_SL g1860 ( 
.A(n_1570),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_SL g1861 ( 
.A(n_1570),
.B(n_991),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1537),
.B(n_1106),
.Y(n_1862)
);

HB1xp67_ASAP7_75t_L g1863 ( 
.A(n_1570),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1539),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1539),
.Y(n_1865)
);

CKINVDCx5p33_ASAP7_75t_R g1866 ( 
.A(n_1595),
.Y(n_1866)
);

AND2x4_ASAP7_75t_L g1867 ( 
.A(n_1537),
.B(n_1177),
.Y(n_1867)
);

INVx2_ASAP7_75t_L g1868 ( 
.A(n_1640),
.Y(n_1868)
);

INVx2_ASAP7_75t_L g1869 ( 
.A(n_1640),
.Y(n_1869)
);

INVx2_ASAP7_75t_L g1870 ( 
.A(n_1640),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1537),
.B(n_1108),
.Y(n_1871)
);

AND3x2_ASAP7_75t_L g1872 ( 
.A(n_1541),
.B(n_1004),
.C(n_1453),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1537),
.Y(n_1873)
);

CKINVDCx5p33_ASAP7_75t_R g1874 ( 
.A(n_1595),
.Y(n_1874)
);

CKINVDCx20_ASAP7_75t_R g1875 ( 
.A(n_1570),
.Y(n_1875)
);

INVx4_ASAP7_75t_L g1876 ( 
.A(n_1844),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1680),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1682),
.Y(n_1878)
);

OAI22xp33_ASAP7_75t_L g1879 ( 
.A1(n_1752),
.A2(n_1368),
.B1(n_1371),
.B2(n_1316),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1683),
.Y(n_1880)
);

OAI22xp5_ASAP7_75t_L g1881 ( 
.A1(n_1694),
.A2(n_1111),
.B1(n_1112),
.B2(n_1110),
.Y(n_1881)
);

AND2x2_ASAP7_75t_L g1882 ( 
.A(n_1721),
.B(n_1762),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_SL g1883 ( 
.A(n_1695),
.B(n_1416),
.Y(n_1883)
);

INVx4_ASAP7_75t_L g1884 ( 
.A(n_1711),
.Y(n_1884)
);

INVx4_ASAP7_75t_L g1885 ( 
.A(n_1666),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1686),
.Y(n_1886)
);

INVx1_ASAP7_75t_SL g1887 ( 
.A(n_1752),
.Y(n_1887)
);

INVx2_ASAP7_75t_L g1888 ( 
.A(n_1669),
.Y(n_1888)
);

INVx2_ASAP7_75t_L g1889 ( 
.A(n_1676),
.Y(n_1889)
);

INVxp67_ASAP7_75t_L g1890 ( 
.A(n_1684),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1667),
.B(n_991),
.Y(n_1891)
);

OR2x2_ASAP7_75t_L g1892 ( 
.A(n_1863),
.B(n_965),
.Y(n_1892)
);

BUFx6f_ASAP7_75t_SL g1893 ( 
.A(n_1789),
.Y(n_1893)
);

BUFx3_ASAP7_75t_L g1894 ( 
.A(n_1766),
.Y(n_1894)
);

AOI22xp33_ASAP7_75t_L g1895 ( 
.A1(n_1745),
.A2(n_1219),
.B1(n_1347),
.B2(n_1179),
.Y(n_1895)
);

BUFx6f_ASAP7_75t_L g1896 ( 
.A(n_1676),
.Y(n_1896)
);

INVx2_ASAP7_75t_SL g1897 ( 
.A(n_1755),
.Y(n_1897)
);

OR2x2_ASAP7_75t_L g1898 ( 
.A(n_1668),
.B(n_999),
.Y(n_1898)
);

INVx2_ASAP7_75t_L g1899 ( 
.A(n_1700),
.Y(n_1899)
);

NOR2xp33_ASAP7_75t_L g1900 ( 
.A(n_1692),
.B(n_1114),
.Y(n_1900)
);

INVxp67_ASAP7_75t_SL g1901 ( 
.A(n_1729),
.Y(n_1901)
);

INVx2_ASAP7_75t_L g1902 ( 
.A(n_1700),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1718),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_SL g1904 ( 
.A(n_1755),
.B(n_1416),
.Y(n_1904)
);

NOR2xp33_ASAP7_75t_SL g1905 ( 
.A(n_1758),
.B(n_1759),
.Y(n_1905)
);

INVx2_ASAP7_75t_L g1906 ( 
.A(n_1718),
.Y(n_1906)
);

AND3x2_ASAP7_75t_L g1907 ( 
.A(n_1766),
.B(n_1455),
.C(n_1432),
.Y(n_1907)
);

BUFx3_ASAP7_75t_L g1908 ( 
.A(n_1666),
.Y(n_1908)
);

AND2x2_ASAP7_75t_L g1909 ( 
.A(n_1845),
.B(n_1072),
.Y(n_1909)
);

INVx4_ASAP7_75t_L g1910 ( 
.A(n_1798),
.Y(n_1910)
);

NAND3xp33_ASAP7_75t_L g1911 ( 
.A(n_1689),
.B(n_1123),
.C(n_1119),
.Y(n_1911)
);

AOI22xp33_ASAP7_75t_L g1912 ( 
.A1(n_1765),
.A2(n_1219),
.B1(n_1347),
.B2(n_1179),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1677),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_L g1914 ( 
.A(n_1687),
.B(n_991),
.Y(n_1914)
);

INVx4_ASAP7_75t_L g1915 ( 
.A(n_1798),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1677),
.Y(n_1916)
);

AND2x4_ASAP7_75t_L g1917 ( 
.A(n_1770),
.B(n_975),
.Y(n_1917)
);

HB1xp67_ASAP7_75t_L g1918 ( 
.A(n_1679),
.Y(n_1918)
);

INVx2_ASAP7_75t_L g1919 ( 
.A(n_1858),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1836),
.B(n_991),
.Y(n_1920)
);

NOR2xp33_ASAP7_75t_L g1921 ( 
.A(n_1815),
.B(n_1130),
.Y(n_1921)
);

AOI22xp5_ASAP7_75t_L g1922 ( 
.A1(n_1709),
.A2(n_1143),
.B1(n_1144),
.B2(n_1140),
.Y(n_1922)
);

INVx2_ASAP7_75t_L g1923 ( 
.A(n_1858),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_L g1924 ( 
.A(n_1842),
.B(n_1847),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_SL g1925 ( 
.A(n_1855),
.B(n_1867),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1800),
.B(n_1135),
.Y(n_1926)
);

INVx3_ASAP7_75t_L g1927 ( 
.A(n_1805),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1673),
.Y(n_1928)
);

INVx2_ASAP7_75t_L g1929 ( 
.A(n_1799),
.Y(n_1929)
);

BUFx4f_ASAP7_75t_L g1930 ( 
.A(n_1774),
.Y(n_1930)
);

INVxp33_ASAP7_75t_L g1931 ( 
.A(n_1754),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1673),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1674),
.Y(n_1933)
);

INVx3_ASAP7_75t_L g1934 ( 
.A(n_1808),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_SL g1935 ( 
.A(n_1821),
.B(n_1239),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1674),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_SL g1937 ( 
.A(n_1834),
.B(n_1260),
.Y(n_1937)
);

OAI22xp5_ASAP7_75t_SL g1938 ( 
.A1(n_1776),
.A2(n_1521),
.B1(n_1522),
.B2(n_1479),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1688),
.Y(n_1939)
);

HB1xp67_ASAP7_75t_L g1940 ( 
.A(n_1857),
.Y(n_1940)
);

INVx3_ASAP7_75t_L g1941 ( 
.A(n_1678),
.Y(n_1941)
);

INVx2_ASAP7_75t_L g1942 ( 
.A(n_1799),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_SL g1943 ( 
.A(n_1839),
.B(n_1260),
.Y(n_1943)
);

OR2x6_ASAP7_75t_L g1944 ( 
.A(n_1860),
.B(n_986),
.Y(n_1944)
);

INVx2_ASAP7_75t_L g1945 ( 
.A(n_1803),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1688),
.Y(n_1946)
);

INVx4_ASAP7_75t_L g1947 ( 
.A(n_1803),
.Y(n_1947)
);

OR2x2_ASAP7_75t_L g1948 ( 
.A(n_1785),
.B(n_1063),
.Y(n_1948)
);

NOR2xp33_ASAP7_75t_L g1949 ( 
.A(n_1817),
.B(n_1145),
.Y(n_1949)
);

AND2x2_ASAP7_75t_L g1950 ( 
.A(n_1845),
.B(n_1072),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_L g1951 ( 
.A(n_1843),
.B(n_1135),
.Y(n_1951)
);

NAND3xp33_ASAP7_75t_L g1952 ( 
.A(n_1739),
.B(n_1149),
.C(n_1148),
.Y(n_1952)
);

AOI22xp5_ASAP7_75t_L g1953 ( 
.A1(n_1825),
.A2(n_1153),
.B1(n_1154),
.B2(n_1152),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1724),
.Y(n_1954)
);

AND2x2_ASAP7_75t_L g1955 ( 
.A(n_1859),
.B(n_1071),
.Y(n_1955)
);

CKINVDCx5p33_ASAP7_75t_R g1956 ( 
.A(n_1875),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1724),
.Y(n_1957)
);

OR2x6_ASAP7_75t_L g1958 ( 
.A(n_1841),
.B(n_1007),
.Y(n_1958)
);

CKINVDCx5p33_ASAP7_75t_R g1959 ( 
.A(n_1681),
.Y(n_1959)
);

NOR2xp33_ASAP7_75t_L g1960 ( 
.A(n_1820),
.B(n_1161),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1725),
.Y(n_1961)
);

OAI22xp33_ASAP7_75t_SL g1962 ( 
.A1(n_1746),
.A2(n_1165),
.B1(n_1171),
.B2(n_1164),
.Y(n_1962)
);

INVx4_ASAP7_75t_L g1963 ( 
.A(n_1813),
.Y(n_1963)
);

CKINVDCx5p33_ASAP7_75t_R g1964 ( 
.A(n_1866),
.Y(n_1964)
);

INVx2_ASAP7_75t_L g1965 ( 
.A(n_1813),
.Y(n_1965)
);

INVx2_ASAP7_75t_L g1966 ( 
.A(n_1816),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1725),
.Y(n_1967)
);

OR2x2_ASAP7_75t_L g1968 ( 
.A(n_1788),
.B(n_1103),
.Y(n_1968)
);

INVx5_ASAP7_75t_L g1969 ( 
.A(n_1816),
.Y(n_1969)
);

AND2x4_ASAP7_75t_L g1970 ( 
.A(n_1773),
.B(n_1859),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_L g1971 ( 
.A(n_1862),
.B(n_1135),
.Y(n_1971)
);

NOR2xp33_ASAP7_75t_L g1972 ( 
.A(n_1831),
.B(n_1832),
.Y(n_1972)
);

INVx2_ASAP7_75t_L g1973 ( 
.A(n_1818),
.Y(n_1973)
);

INVx2_ASAP7_75t_L g1974 ( 
.A(n_1818),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1727),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1727),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1731),
.Y(n_1977)
);

INVx2_ASAP7_75t_SL g1978 ( 
.A(n_1728),
.Y(n_1978)
);

INVx2_ASAP7_75t_L g1979 ( 
.A(n_1819),
.Y(n_1979)
);

HB1xp67_ASAP7_75t_L g1980 ( 
.A(n_1779),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_SL g1981 ( 
.A(n_1871),
.B(n_1300),
.Y(n_1981)
);

AOI22xp33_ASAP7_75t_L g1982 ( 
.A1(n_1760),
.A2(n_1224),
.B1(n_1225),
.B2(n_1208),
.Y(n_1982)
);

INVx2_ASAP7_75t_SL g1983 ( 
.A(n_1738),
.Y(n_1983)
);

INVx2_ASAP7_75t_L g1984 ( 
.A(n_1819),
.Y(n_1984)
);

AND2x4_ASAP7_75t_L g1985 ( 
.A(n_1837),
.B(n_980),
.Y(n_1985)
);

NAND3xp33_ASAP7_75t_L g1986 ( 
.A(n_1720),
.B(n_1188),
.C(n_1186),
.Y(n_1986)
);

AOI22xp33_ASAP7_75t_L g1987 ( 
.A1(n_1764),
.A2(n_1248),
.B1(n_1249),
.B2(n_1246),
.Y(n_1987)
);

BUFx4f_ASAP7_75t_L g1988 ( 
.A(n_1774),
.Y(n_1988)
);

OR2x6_ASAP7_75t_L g1989 ( 
.A(n_1782),
.B(n_1007),
.Y(n_1989)
);

INVx2_ASAP7_75t_L g1990 ( 
.A(n_1823),
.Y(n_1990)
);

INVxp67_ASAP7_75t_SL g1991 ( 
.A(n_1731),
.Y(n_1991)
);

INVx3_ASAP7_75t_L g1992 ( 
.A(n_1823),
.Y(n_1992)
);

BUFx2_ASAP7_75t_L g1993 ( 
.A(n_1696),
.Y(n_1993)
);

AND2x4_ASAP7_75t_L g1994 ( 
.A(n_1840),
.B(n_989),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_L g1995 ( 
.A(n_1675),
.B(n_1135),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1675),
.Y(n_1996)
);

INVx8_ASAP7_75t_L g1997 ( 
.A(n_1874),
.Y(n_1997)
);

OR2x6_ASAP7_75t_L g1998 ( 
.A(n_1792),
.B(n_1034),
.Y(n_1998)
);

NOR3xp33_ASAP7_75t_L g1999 ( 
.A(n_1794),
.B(n_1461),
.C(n_1043),
.Y(n_1999)
);

CKINVDCx5p33_ASAP7_75t_R g2000 ( 
.A(n_1726),
.Y(n_2000)
);

AND2x2_ASAP7_75t_L g2001 ( 
.A(n_1751),
.B(n_1071),
.Y(n_2001)
);

OAI22xp33_ASAP7_75t_L g2002 ( 
.A1(n_1767),
.A2(n_1202),
.B1(n_1203),
.B2(n_1190),
.Y(n_2002)
);

NOR2xp33_ASAP7_75t_L g2003 ( 
.A(n_1848),
.B(n_1207),
.Y(n_2003)
);

INVx2_ASAP7_75t_L g2004 ( 
.A(n_1833),
.Y(n_2004)
);

BUFx2_ASAP7_75t_L g2005 ( 
.A(n_1717),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1685),
.Y(n_2006)
);

INVx2_ASAP7_75t_L g2007 ( 
.A(n_1833),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1685),
.Y(n_2008)
);

NAND2xp5_ASAP7_75t_SL g2009 ( 
.A(n_1716),
.B(n_1300),
.Y(n_2009)
);

AND2x2_ASAP7_75t_L g2010 ( 
.A(n_1761),
.B(n_1071),
.Y(n_2010)
);

BUFx3_ASAP7_75t_L g2011 ( 
.A(n_1835),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1693),
.Y(n_2012)
);

BUFx2_ASAP7_75t_L g2013 ( 
.A(n_1771),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1849),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_L g2015 ( 
.A(n_1850),
.B(n_1135),
.Y(n_2015)
);

AOI22xp33_ASAP7_75t_L g2016 ( 
.A1(n_1741),
.A2(n_1282),
.B1(n_1287),
.B2(n_1277),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_SL g2017 ( 
.A(n_1734),
.B(n_1317),
.Y(n_2017)
);

AOI21x1_ASAP7_75t_L g2018 ( 
.A1(n_1801),
.A2(n_1301),
.B(n_1290),
.Y(n_2018)
);

INVx1_ASAP7_75t_SL g2019 ( 
.A(n_1796),
.Y(n_2019)
);

INVx2_ASAP7_75t_L g2020 ( 
.A(n_1835),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_SL g2021 ( 
.A(n_1873),
.B(n_1317),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1851),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1853),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1854),
.Y(n_2024)
);

AND2x2_ASAP7_75t_L g2025 ( 
.A(n_1769),
.B(n_1221),
.Y(n_2025)
);

INVx2_ASAP7_75t_L g2026 ( 
.A(n_1665),
.Y(n_2026)
);

NOR2xp33_ASAP7_75t_L g2027 ( 
.A(n_1856),
.B(n_1210),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1690),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1691),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1699),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1704),
.Y(n_2031)
);

INVx4_ASAP7_75t_L g2032 ( 
.A(n_1846),
.Y(n_2032)
);

BUFx6f_ASAP7_75t_L g2033 ( 
.A(n_1797),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_SL g2034 ( 
.A(n_1750),
.B(n_1735),
.Y(n_2034)
);

INVx4_ASAP7_75t_L g2035 ( 
.A(n_1742),
.Y(n_2035)
);

INVxp33_ASAP7_75t_L g2036 ( 
.A(n_1790),
.Y(n_2036)
);

AOI22xp33_ASAP7_75t_L g2037 ( 
.A1(n_1747),
.A2(n_1321),
.B1(n_1331),
.B2(n_1306),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_SL g2038 ( 
.A(n_1736),
.B(n_1335),
.Y(n_2038)
);

AND2x6_ASAP7_75t_L g2039 ( 
.A(n_1740),
.B(n_1335),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_1706),
.Y(n_2040)
);

BUFx6f_ASAP7_75t_L g2041 ( 
.A(n_1802),
.Y(n_2041)
);

INVx2_ASAP7_75t_L g2042 ( 
.A(n_1809),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_1712),
.Y(n_2043)
);

BUFx6f_ASAP7_75t_L g2044 ( 
.A(n_1811),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1714),
.Y(n_2045)
);

NAND2xp5_ASAP7_75t_L g2046 ( 
.A(n_1697),
.B(n_1135),
.Y(n_2046)
);

INVx2_ASAP7_75t_L g2047 ( 
.A(n_1812),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1730),
.Y(n_2048)
);

NOR3xp33_ASAP7_75t_L g2049 ( 
.A(n_1781),
.B(n_1048),
.C(n_985),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_L g2050 ( 
.A(n_1698),
.B(n_1142),
.Y(n_2050)
);

NAND2xp5_ASAP7_75t_L g2051 ( 
.A(n_1701),
.B(n_1142),
.Y(n_2051)
);

AND2x2_ASAP7_75t_L g2052 ( 
.A(n_1748),
.B(n_1221),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1702),
.Y(n_2053)
);

NOR2xp33_ASAP7_75t_L g2054 ( 
.A(n_1753),
.B(n_1215),
.Y(n_2054)
);

INVx2_ASAP7_75t_SL g2055 ( 
.A(n_1756),
.Y(n_2055)
);

INVx2_ASAP7_75t_L g2056 ( 
.A(n_1814),
.Y(n_2056)
);

BUFx6f_ASAP7_75t_L g2057 ( 
.A(n_1822),
.Y(n_2057)
);

AOI22xp33_ASAP7_75t_L g2058 ( 
.A1(n_1703),
.A2(n_1334),
.B1(n_1341),
.B2(n_1332),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_L g2059 ( 
.A(n_1705),
.B(n_1142),
.Y(n_2059)
);

NAND2xp33_ASAP7_75t_L g2060 ( 
.A(n_1707),
.B(n_1142),
.Y(n_2060)
);

NOR2xp33_ASAP7_75t_L g2061 ( 
.A(n_1671),
.B(n_1216),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_1708),
.Y(n_2062)
);

AOI22xp33_ASAP7_75t_L g2063 ( 
.A1(n_1710),
.A2(n_1357),
.B1(n_1360),
.B2(n_1343),
.Y(n_2063)
);

INVx2_ASAP7_75t_L g2064 ( 
.A(n_1826),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_SL g2065 ( 
.A(n_1713),
.B(n_1361),
.Y(n_2065)
);

INVx2_ASAP7_75t_L g2066 ( 
.A(n_1838),
.Y(n_2066)
);

CKINVDCx5p33_ASAP7_75t_R g2067 ( 
.A(n_1792),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_1715),
.Y(n_2068)
);

INVx1_ASAP7_75t_SL g2069 ( 
.A(n_1749),
.Y(n_2069)
);

INVx2_ASAP7_75t_L g2070 ( 
.A(n_1852),
.Y(n_2070)
);

AOI22xp33_ASAP7_75t_L g2071 ( 
.A1(n_1719),
.A2(n_1732),
.B1(n_1733),
.B2(n_1722),
.Y(n_2071)
);

NAND2xp5_ASAP7_75t_L g2072 ( 
.A(n_1830),
.B(n_1142),
.Y(n_2072)
);

BUFx3_ASAP7_75t_L g2073 ( 
.A(n_1757),
.Y(n_2073)
);

NAND2xp5_ASAP7_75t_SL g2074 ( 
.A(n_1723),
.B(n_1361),
.Y(n_2074)
);

NAND2xp33_ASAP7_75t_L g2075 ( 
.A(n_1757),
.B(n_1142),
.Y(n_2075)
);

INVx2_ASAP7_75t_L g2076 ( 
.A(n_1868),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_1869),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_1870),
.Y(n_2078)
);

OAI22xp5_ASAP7_75t_L g2079 ( 
.A1(n_1807),
.A2(n_1524),
.B1(n_1525),
.B2(n_1523),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_1801),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_1804),
.Y(n_2081)
);

NAND2xp5_ASAP7_75t_SL g2082 ( 
.A(n_1737),
.B(n_1439),
.Y(n_2082)
);

NAND3xp33_ASAP7_75t_L g2083 ( 
.A(n_1744),
.B(n_1220),
.C(n_1218),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_1804),
.Y(n_2084)
);

NAND2xp5_ASAP7_75t_L g2085 ( 
.A(n_1861),
.B(n_1806),
.Y(n_2085)
);

OR2x2_ASAP7_75t_L g2086 ( 
.A(n_1783),
.B(n_1795),
.Y(n_2086)
);

INVx3_ASAP7_75t_L g2087 ( 
.A(n_1763),
.Y(n_2087)
);

BUFx10_ASAP7_75t_L g2088 ( 
.A(n_1763),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_1806),
.Y(n_2089)
);

CKINVDCx20_ASAP7_75t_R g2090 ( 
.A(n_1793),
.Y(n_2090)
);

INVx3_ASAP7_75t_L g2091 ( 
.A(n_1768),
.Y(n_2091)
);

AND2x2_ASAP7_75t_L g2092 ( 
.A(n_1768),
.B(n_1221),
.Y(n_2092)
);

INVx4_ASAP7_75t_L g2093 ( 
.A(n_1772),
.Y(n_2093)
);

INVx2_ASAP7_75t_SL g2094 ( 
.A(n_1772),
.Y(n_2094)
);

INVx2_ASAP7_75t_L g2095 ( 
.A(n_1810),
.Y(n_2095)
);

INVx4_ASAP7_75t_L g2096 ( 
.A(n_1670),
.Y(n_2096)
);

AND3x2_ASAP7_75t_L g2097 ( 
.A(n_1784),
.B(n_1088),
.C(n_1014),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_L g2098 ( 
.A(n_1810),
.B(n_1189),
.Y(n_2098)
);

BUFx3_ASAP7_75t_L g2099 ( 
.A(n_1775),
.Y(n_2099)
);

INVx5_ASAP7_75t_L g2100 ( 
.A(n_1672),
.Y(n_2100)
);

BUFx3_ASAP7_75t_L g2101 ( 
.A(n_1787),
.Y(n_2101)
);

AND2x2_ASAP7_75t_L g2102 ( 
.A(n_1787),
.B(n_1529),
.Y(n_2102)
);

INVx2_ASAP7_75t_SL g2103 ( 
.A(n_1872),
.Y(n_2103)
);

INVx2_ASAP7_75t_L g2104 ( 
.A(n_1824),
.Y(n_2104)
);

INVx2_ASAP7_75t_L g2105 ( 
.A(n_1824),
.Y(n_2105)
);

INVx2_ASAP7_75t_L g2106 ( 
.A(n_1827),
.Y(n_2106)
);

NAND2xp5_ASAP7_75t_L g2107 ( 
.A(n_1827),
.B(n_1189),
.Y(n_2107)
);

INVx2_ASAP7_75t_L g2108 ( 
.A(n_1828),
.Y(n_2108)
);

INVx2_ASAP7_75t_L g2109 ( 
.A(n_1828),
.Y(n_2109)
);

NOR2xp33_ASAP7_75t_L g2110 ( 
.A(n_1743),
.B(n_1223),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_1829),
.Y(n_2111)
);

CKINVDCx5p33_ASAP7_75t_R g2112 ( 
.A(n_1793),
.Y(n_2112)
);

BUFx10_ASAP7_75t_L g2113 ( 
.A(n_1787),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_1829),
.Y(n_2114)
);

INVx2_ASAP7_75t_L g2115 ( 
.A(n_1864),
.Y(n_2115)
);

XOR2xp5_ASAP7_75t_L g2116 ( 
.A(n_1786),
.B(n_1176),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_1864),
.Y(n_2117)
);

NOR2xp33_ASAP7_75t_L g2118 ( 
.A(n_1777),
.B(n_1226),
.Y(n_2118)
);

NAND2xp5_ASAP7_75t_SL g2119 ( 
.A(n_1865),
.B(n_1439),
.Y(n_2119)
);

AO22x2_ASAP7_75t_L g2120 ( 
.A1(n_1791),
.A2(n_1196),
.B1(n_1251),
.B2(n_1146),
.Y(n_2120)
);

NAND2xp5_ASAP7_75t_SL g2121 ( 
.A(n_1865),
.B(n_1466),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_L g2122 ( 
.A(n_1780),
.B(n_1189),
.Y(n_2122)
);

NOR2xp33_ASAP7_75t_L g2123 ( 
.A(n_1778),
.B(n_1228),
.Y(n_2123)
);

BUFx4f_ASAP7_75t_L g2124 ( 
.A(n_1774),
.Y(n_2124)
);

INVx3_ASAP7_75t_L g2125 ( 
.A(n_1677),
.Y(n_2125)
);

BUFx6f_ASAP7_75t_L g2126 ( 
.A(n_1676),
.Y(n_2126)
);

INVx2_ASAP7_75t_L g2127 ( 
.A(n_1669),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_1680),
.Y(n_2128)
);

BUFx4f_ASAP7_75t_L g2129 ( 
.A(n_1774),
.Y(n_2129)
);

NAND2xp5_ASAP7_75t_SL g2130 ( 
.A(n_1762),
.B(n_1466),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_1680),
.Y(n_2131)
);

INVx2_ASAP7_75t_L g2132 ( 
.A(n_1669),
.Y(n_2132)
);

INVx2_ASAP7_75t_SL g2133 ( 
.A(n_1762),
.Y(n_2133)
);

NOR2xp33_ASAP7_75t_L g2134 ( 
.A(n_1692),
.B(n_1232),
.Y(n_2134)
);

BUFx3_ASAP7_75t_L g2135 ( 
.A(n_1752),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_1680),
.Y(n_2136)
);

NAND2xp5_ASAP7_75t_SL g2137 ( 
.A(n_1762),
.B(n_1473),
.Y(n_2137)
);

BUFx2_ASAP7_75t_L g2138 ( 
.A(n_1684),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_1680),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_1680),
.Y(n_2140)
);

INVx2_ASAP7_75t_L g2141 ( 
.A(n_1669),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_1680),
.Y(n_2142)
);

INVx2_ASAP7_75t_L g2143 ( 
.A(n_1669),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_1680),
.Y(n_2144)
);

BUFx2_ASAP7_75t_L g2145 ( 
.A(n_1684),
.Y(n_2145)
);

INVx2_ASAP7_75t_L g2146 ( 
.A(n_1669),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_1680),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_1680),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_1680),
.Y(n_2149)
);

INVx3_ASAP7_75t_L g2150 ( 
.A(n_1666),
.Y(n_2150)
);

INVx3_ASAP7_75t_L g2151 ( 
.A(n_1666),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_1680),
.Y(n_2152)
);

INVx2_ASAP7_75t_L g2153 ( 
.A(n_1669),
.Y(n_2153)
);

BUFx2_ASAP7_75t_L g2154 ( 
.A(n_1684),
.Y(n_2154)
);

INVx3_ASAP7_75t_L g2155 ( 
.A(n_1677),
.Y(n_2155)
);

INVx3_ASAP7_75t_L g2156 ( 
.A(n_1677),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_1680),
.Y(n_2157)
);

BUFx3_ASAP7_75t_L g2158 ( 
.A(n_1752),
.Y(n_2158)
);

INVx3_ASAP7_75t_L g2159 ( 
.A(n_1677),
.Y(n_2159)
);

INVx5_ASAP7_75t_L g2160 ( 
.A(n_1666),
.Y(n_2160)
);

NOR2xp33_ASAP7_75t_L g2161 ( 
.A(n_1692),
.B(n_1237),
.Y(n_2161)
);

INVx2_ASAP7_75t_L g2162 ( 
.A(n_1669),
.Y(n_2162)
);

NAND2xp5_ASAP7_75t_SL g2163 ( 
.A(n_1762),
.B(n_1473),
.Y(n_2163)
);

INVx2_ASAP7_75t_L g2164 ( 
.A(n_1669),
.Y(n_2164)
);

NOR2xp33_ASAP7_75t_L g2165 ( 
.A(n_1692),
.B(n_1241),
.Y(n_2165)
);

NOR2xp33_ASAP7_75t_L g2166 ( 
.A(n_1692),
.B(n_1250),
.Y(n_2166)
);

INVx2_ASAP7_75t_L g2167 ( 
.A(n_1896),
.Y(n_2167)
);

INVx2_ASAP7_75t_L g2168 ( 
.A(n_1896),
.Y(n_2168)
);

NAND2xp5_ASAP7_75t_SL g2169 ( 
.A(n_1887),
.B(n_1262),
.Y(n_2169)
);

NAND2xp5_ASAP7_75t_L g2170 ( 
.A(n_1909),
.B(n_1533),
.Y(n_2170)
);

AOI22xp5_ASAP7_75t_L g2171 ( 
.A1(n_2019),
.A2(n_1255),
.B1(n_1257),
.B2(n_1253),
.Y(n_2171)
);

INVx2_ASAP7_75t_L g2172 ( 
.A(n_1896),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_1996),
.Y(n_2173)
);

NAND2xp5_ASAP7_75t_SL g2174 ( 
.A(n_1905),
.B(n_1267),
.Y(n_2174)
);

NAND2xp5_ASAP7_75t_L g2175 ( 
.A(n_1950),
.B(n_1513),
.Y(n_2175)
);

NOR2xp33_ASAP7_75t_L g2176 ( 
.A(n_1931),
.B(n_1258),
.Y(n_2176)
);

INVx2_ASAP7_75t_L g2177 ( 
.A(n_2126),
.Y(n_2177)
);

NAND2xp5_ASAP7_75t_L g2178 ( 
.A(n_1900),
.B(n_1530),
.Y(n_2178)
);

AOI22xp33_ASAP7_75t_L g2179 ( 
.A1(n_2039),
.A2(n_1499),
.B1(n_1189),
.B2(n_1268),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_2006),
.Y(n_2180)
);

NAND2xp5_ASAP7_75t_L g2181 ( 
.A(n_2134),
.B(n_1261),
.Y(n_2181)
);

AOI21xp5_ASAP7_75t_L g2182 ( 
.A1(n_1888),
.A2(n_1531),
.B(n_1367),
.Y(n_2182)
);

NAND2xp5_ASAP7_75t_L g2183 ( 
.A(n_2161),
.B(n_1269),
.Y(n_2183)
);

AND2x2_ASAP7_75t_L g2184 ( 
.A(n_1894),
.B(n_1529),
.Y(n_2184)
);

INVx2_ASAP7_75t_L g2185 ( 
.A(n_2095),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_2008),
.Y(n_2186)
);

AND2x2_ASAP7_75t_L g2187 ( 
.A(n_2135),
.B(n_1529),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_1928),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_1932),
.Y(n_2189)
);

NOR2xp33_ASAP7_75t_L g2190 ( 
.A(n_2133),
.B(n_1270),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_1933),
.Y(n_2191)
);

NAND2xp5_ASAP7_75t_L g2192 ( 
.A(n_2165),
.B(n_1272),
.Y(n_2192)
);

NAND2xp5_ASAP7_75t_L g2193 ( 
.A(n_2166),
.B(n_1274),
.Y(n_2193)
);

AOI22xp5_ASAP7_75t_L g2194 ( 
.A1(n_1882),
.A2(n_1283),
.B1(n_1286),
.B2(n_1276),
.Y(n_2194)
);

INVx2_ASAP7_75t_L g2195 ( 
.A(n_2104),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_1936),
.Y(n_2196)
);

AOI22xp5_ASAP7_75t_L g2197 ( 
.A1(n_1970),
.A2(n_1881),
.B1(n_1922),
.B2(n_1955),
.Y(n_2197)
);

OAI22xp5_ASAP7_75t_L g2198 ( 
.A1(n_2071),
.A2(n_1151),
.B1(n_1160),
.B2(n_1115),
.Y(n_2198)
);

NAND3xp33_ASAP7_75t_L g2199 ( 
.A(n_1999),
.B(n_1292),
.C(n_1291),
.Y(n_2199)
);

NAND2xp33_ASAP7_75t_L g2200 ( 
.A(n_2039),
.B(n_1189),
.Y(n_2200)
);

AND2x4_ASAP7_75t_SL g2201 ( 
.A(n_2088),
.B(n_1181),
.Y(n_2201)
);

INVx2_ASAP7_75t_L g2202 ( 
.A(n_2105),
.Y(n_2202)
);

INVx2_ASAP7_75t_SL g2203 ( 
.A(n_2158),
.Y(n_2203)
);

NAND2xp5_ASAP7_75t_L g2204 ( 
.A(n_1970),
.B(n_1303),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_2012),
.Y(n_2205)
);

NAND3xp33_ASAP7_75t_SL g2206 ( 
.A(n_1956),
.B(n_2112),
.C(n_2067),
.Y(n_2206)
);

BUFx3_ASAP7_75t_L g2207 ( 
.A(n_2090),
.Y(n_2207)
);

NAND2xp5_ASAP7_75t_L g2208 ( 
.A(n_1972),
.B(n_1304),
.Y(n_2208)
);

INVx2_ASAP7_75t_SL g2209 ( 
.A(n_2138),
.Y(n_2209)
);

AND2x2_ASAP7_75t_L g2210 ( 
.A(n_1993),
.B(n_2005),
.Y(n_2210)
);

INVx2_ASAP7_75t_L g2211 ( 
.A(n_2106),
.Y(n_2211)
);

NOR3xp33_ASAP7_75t_L g2212 ( 
.A(n_1879),
.B(n_1509),
.C(n_1309),
.Y(n_2212)
);

NOR2xp33_ASAP7_75t_SL g2213 ( 
.A(n_2145),
.B(n_1200),
.Y(n_2213)
);

AND2x4_ASAP7_75t_L g2214 ( 
.A(n_2035),
.B(n_1000),
.Y(n_2214)
);

OAI22xp5_ASAP7_75t_L g2215 ( 
.A1(n_2014),
.A2(n_1234),
.B1(n_1243),
.B2(n_1206),
.Y(n_2215)
);

NOR3xp33_ASAP7_75t_L g2216 ( 
.A(n_1938),
.B(n_1312),
.C(n_1305),
.Y(n_2216)
);

NAND2xp5_ASAP7_75t_L g2217 ( 
.A(n_1901),
.B(n_1313),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_2053),
.Y(n_2218)
);

NOR2x1p5_ASAP7_75t_L g2219 ( 
.A(n_2000),
.B(n_1318),
.Y(n_2219)
);

INVx2_ASAP7_75t_L g2220 ( 
.A(n_2108),
.Y(n_2220)
);

NOR2xp33_ASAP7_75t_L g2221 ( 
.A(n_2036),
.B(n_1320),
.Y(n_2221)
);

NAND2xp5_ASAP7_75t_SL g2222 ( 
.A(n_2035),
.B(n_1336),
.Y(n_2222)
);

AOI22xp5_ASAP7_75t_L g2223 ( 
.A1(n_2039),
.A2(n_1324),
.B1(n_1325),
.B2(n_1322),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_2062),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_2068),
.Y(n_2225)
);

AND2x2_ASAP7_75t_L g2226 ( 
.A(n_2154),
.B(n_1256),
.Y(n_2226)
);

AND2x6_ASAP7_75t_L g2227 ( 
.A(n_2101),
.B(n_1531),
.Y(n_2227)
);

OR2x2_ASAP7_75t_L g2228 ( 
.A(n_1892),
.B(n_1326),
.Y(n_2228)
);

INVxp67_ASAP7_75t_L g2229 ( 
.A(n_1898),
.Y(n_2229)
);

NAND2xp5_ASAP7_75t_L g2230 ( 
.A(n_2022),
.B(n_1327),
.Y(n_2230)
);

INVx4_ASAP7_75t_L g2231 ( 
.A(n_1876),
.Y(n_2231)
);

BUFx8_ASAP7_75t_L g2232 ( 
.A(n_1893),
.Y(n_2232)
);

BUFx6f_ASAP7_75t_L g2233 ( 
.A(n_1889),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_2023),
.Y(n_2234)
);

AOI22xp33_ASAP7_75t_L g2235 ( 
.A1(n_2039),
.A2(n_1499),
.B1(n_1189),
.B2(n_1337),
.Y(n_2235)
);

INVx2_ASAP7_75t_L g2236 ( 
.A(n_2109),
.Y(n_2236)
);

NAND2xp5_ASAP7_75t_L g2237 ( 
.A(n_2024),
.B(n_1333),
.Y(n_2237)
);

INVx2_ASAP7_75t_L g2238 ( 
.A(n_2115),
.Y(n_2238)
);

OR2x6_ASAP7_75t_L g2239 ( 
.A(n_1997),
.B(n_1034),
.Y(n_2239)
);

NAND2xp5_ASAP7_75t_L g2240 ( 
.A(n_1985),
.B(n_1510),
.Y(n_2240)
);

AND2x2_ASAP7_75t_L g2241 ( 
.A(n_1948),
.B(n_1295),
.Y(n_2241)
);

AOI22xp33_ASAP7_75t_L g2242 ( 
.A1(n_1985),
.A2(n_1499),
.B1(n_1340),
.B2(n_1345),
.Y(n_2242)
);

OR2x2_ASAP7_75t_L g2243 ( 
.A(n_1890),
.B(n_1339),
.Y(n_2243)
);

INVx1_ASAP7_75t_L g2244 ( 
.A(n_1877),
.Y(n_2244)
);

BUFx6f_ASAP7_75t_L g2245 ( 
.A(n_1899),
.Y(n_2245)
);

NAND2xp5_ASAP7_75t_L g2246 ( 
.A(n_1994),
.B(n_1348),
.Y(n_2246)
);

AOI22xp33_ASAP7_75t_L g2247 ( 
.A1(n_1994),
.A2(n_1499),
.B1(n_1353),
.B2(n_1355),
.Y(n_2247)
);

NAND2xp5_ASAP7_75t_L g2248 ( 
.A(n_1921),
.B(n_1949),
.Y(n_2248)
);

BUFx5_ASAP7_75t_L g2249 ( 
.A(n_2080),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_1878),
.Y(n_2250)
);

NAND2xp5_ASAP7_75t_L g2251 ( 
.A(n_1960),
.B(n_1350),
.Y(n_2251)
);

NAND2xp5_ASAP7_75t_L g2252 ( 
.A(n_2003),
.B(n_2027),
.Y(n_2252)
);

AOI22xp5_ASAP7_75t_L g2253 ( 
.A1(n_2002),
.A2(n_1365),
.B1(n_1366),
.B2(n_1358),
.Y(n_2253)
);

INVx2_ASAP7_75t_L g2254 ( 
.A(n_1902),
.Y(n_2254)
);

NAND2xp33_ASAP7_75t_L g2255 ( 
.A(n_1903),
.B(n_1499),
.Y(n_2255)
);

INVx2_ASAP7_75t_SL g2256 ( 
.A(n_1944),
.Y(n_2256)
);

NAND2xp5_ASAP7_75t_L g2257 ( 
.A(n_2034),
.B(n_1374),
.Y(n_2257)
);

BUFx6f_ASAP7_75t_L g2258 ( 
.A(n_1906),
.Y(n_2258)
);

NAND2xp5_ASAP7_75t_L g2259 ( 
.A(n_1968),
.B(n_1377),
.Y(n_2259)
);

BUFx8_ASAP7_75t_L g2260 ( 
.A(n_2013),
.Y(n_2260)
);

INVx2_ASAP7_75t_L g2261 ( 
.A(n_1919),
.Y(n_2261)
);

NAND2x1p5_ASAP7_75t_L g2262 ( 
.A(n_2069),
.B(n_1376),
.Y(n_2262)
);

INVx1_ASAP7_75t_L g2263 ( 
.A(n_1880),
.Y(n_2263)
);

NAND2xp5_ASAP7_75t_L g2264 ( 
.A(n_1982),
.B(n_1987),
.Y(n_2264)
);

OAI22xp5_ASAP7_75t_SL g2265 ( 
.A1(n_2116),
.A2(n_1310),
.B1(n_1323),
.B2(n_1296),
.Y(n_2265)
);

NOR2x1p5_ASAP7_75t_L g2266 ( 
.A(n_1959),
.B(n_1379),
.Y(n_2266)
);

NAND2xp5_ASAP7_75t_L g2267 ( 
.A(n_1886),
.B(n_1381),
.Y(n_2267)
);

AND2x2_ASAP7_75t_L g2268 ( 
.A(n_1944),
.B(n_1346),
.Y(n_2268)
);

INVxp67_ASAP7_75t_L g2269 ( 
.A(n_1958),
.Y(n_2269)
);

INVx2_ASAP7_75t_L g2270 ( 
.A(n_1923),
.Y(n_2270)
);

AO221x1_ASAP7_75t_L g2271 ( 
.A1(n_2120),
.A2(n_1372),
.B1(n_1383),
.B2(n_1059),
.C(n_981),
.Y(n_2271)
);

NAND2xp5_ASAP7_75t_SL g2272 ( 
.A(n_1941),
.B(n_1424),
.Y(n_2272)
);

BUFx6f_ASAP7_75t_L g2273 ( 
.A(n_2033),
.Y(n_2273)
);

NAND2xp5_ASAP7_75t_SL g2274 ( 
.A(n_2100),
.B(n_1434),
.Y(n_2274)
);

NAND2xp5_ASAP7_75t_L g2275 ( 
.A(n_2128),
.B(n_1382),
.Y(n_2275)
);

NOR2xp33_ASAP7_75t_L g2276 ( 
.A(n_2010),
.B(n_1386),
.Y(n_2276)
);

NOR2xp33_ASAP7_75t_L g2277 ( 
.A(n_2001),
.B(n_1388),
.Y(n_2277)
);

NAND2xp5_ASAP7_75t_L g2278 ( 
.A(n_2131),
.B(n_1394),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_2136),
.Y(n_2279)
);

A2O1A1Ixp33_ASAP7_75t_L g2280 ( 
.A1(n_1926),
.A2(n_1391),
.B(n_1402),
.C(n_1387),
.Y(n_2280)
);

INVx8_ASAP7_75t_L g2281 ( 
.A(n_1997),
.Y(n_2281)
);

NAND2xp5_ASAP7_75t_L g2282 ( 
.A(n_2139),
.B(n_1506),
.Y(n_2282)
);

NAND2xp5_ASAP7_75t_L g2283 ( 
.A(n_2140),
.B(n_1511),
.Y(n_2283)
);

NAND2xp5_ASAP7_75t_SL g2284 ( 
.A(n_2100),
.B(n_2096),
.Y(n_2284)
);

INVxp67_ASAP7_75t_L g2285 ( 
.A(n_1958),
.Y(n_2285)
);

NAND2xp5_ASAP7_75t_L g2286 ( 
.A(n_2142),
.B(n_1396),
.Y(n_2286)
);

AND2x2_ASAP7_75t_SL g2287 ( 
.A(n_1930),
.B(n_1362),
.Y(n_2287)
);

NOR2xp33_ASAP7_75t_L g2288 ( 
.A(n_1925),
.B(n_1401),
.Y(n_2288)
);

INVx8_ASAP7_75t_L g2289 ( 
.A(n_1998),
.Y(n_2289)
);

NAND2xp5_ASAP7_75t_SL g2290 ( 
.A(n_2100),
.B(n_1427),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_2144),
.Y(n_2291)
);

INVx2_ASAP7_75t_L g2292 ( 
.A(n_2081),
.Y(n_2292)
);

NAND3xp33_ASAP7_75t_L g2293 ( 
.A(n_2110),
.B(n_1411),
.C(n_1410),
.Y(n_2293)
);

NAND2xp5_ASAP7_75t_SL g2294 ( 
.A(n_2096),
.B(n_1452),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_2147),
.Y(n_2295)
);

INVx1_ASAP7_75t_L g2296 ( 
.A(n_2148),
.Y(n_2296)
);

AOI22xp33_ASAP7_75t_L g2297 ( 
.A1(n_1917),
.A2(n_1499),
.B1(n_1428),
.B2(n_1429),
.Y(n_2297)
);

NOR2xp33_ASAP7_75t_L g2298 ( 
.A(n_1924),
.B(n_1422),
.Y(n_2298)
);

NAND2xp5_ASAP7_75t_L g2299 ( 
.A(n_2149),
.B(n_2152),
.Y(n_2299)
);

NAND2xp5_ASAP7_75t_SL g2300 ( 
.A(n_1911),
.B(n_1467),
.Y(n_2300)
);

INVx1_ASAP7_75t_L g2301 ( 
.A(n_2157),
.Y(n_2301)
);

NAND2xp5_ASAP7_75t_L g2302 ( 
.A(n_2016),
.B(n_1433),
.Y(n_2302)
);

NAND2xp5_ASAP7_75t_L g2303 ( 
.A(n_2037),
.B(n_1437),
.Y(n_2303)
);

HB1xp67_ASAP7_75t_L g2304 ( 
.A(n_1998),
.Y(n_2304)
);

NOR2xp33_ASAP7_75t_L g2305 ( 
.A(n_2025),
.B(n_1450),
.Y(n_2305)
);

O2A1O1Ixp5_ASAP7_75t_L g2306 ( 
.A1(n_1935),
.A2(n_1421),
.B(n_1423),
.C(n_1418),
.Y(n_2306)
);

NAND2xp5_ASAP7_75t_SL g2307 ( 
.A(n_1986),
.B(n_1476),
.Y(n_2307)
);

INVx1_ASAP7_75t_SL g2308 ( 
.A(n_1918),
.Y(n_2308)
);

INVx2_ASAP7_75t_L g2309 ( 
.A(n_2084),
.Y(n_2309)
);

NOR2xp33_ASAP7_75t_L g2310 ( 
.A(n_2052),
.B(n_1462),
.Y(n_2310)
);

AO221x1_ASAP7_75t_L g2311 ( 
.A1(n_2120),
.A2(n_1372),
.B1(n_1383),
.B2(n_1059),
.C(n_981),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_2028),
.Y(n_2312)
);

INVx2_ASAP7_75t_SL g2313 ( 
.A(n_2088),
.Y(n_2313)
);

INVx2_ASAP7_75t_L g2314 ( 
.A(n_2089),
.Y(n_2314)
);

INVxp67_ASAP7_75t_L g2315 ( 
.A(n_1940),
.Y(n_2315)
);

NOR2xp33_ASAP7_75t_L g2316 ( 
.A(n_2130),
.B(n_1464),
.Y(n_2316)
);

AND2x4_ASAP7_75t_L g2317 ( 
.A(n_1876),
.B(n_1026),
.Y(n_2317)
);

NAND2xp5_ASAP7_75t_SL g2318 ( 
.A(n_1952),
.B(n_1481),
.Y(n_2318)
);

BUFx6f_ASAP7_75t_SL g2319 ( 
.A(n_2113),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_2029),
.Y(n_2320)
);

NAND2xp5_ASAP7_75t_L g2321 ( 
.A(n_1917),
.B(n_1475),
.Y(n_2321)
);

HB1xp67_ASAP7_75t_L g2322 ( 
.A(n_1980),
.Y(n_2322)
);

AND2x2_ASAP7_75t_L g2323 ( 
.A(n_1989),
.B(n_1373),
.Y(n_2323)
);

BUFx2_ASAP7_75t_L g2324 ( 
.A(n_1989),
.Y(n_2324)
);

AND2x4_ASAP7_75t_L g2325 ( 
.A(n_1884),
.B(n_1883),
.Y(n_2325)
);

INVx2_ASAP7_75t_L g2326 ( 
.A(n_2111),
.Y(n_2326)
);

AND2x2_ASAP7_75t_L g2327 ( 
.A(n_1953),
.B(n_1390),
.Y(n_2327)
);

NAND2xp5_ASAP7_75t_L g2328 ( 
.A(n_2030),
.B(n_1483),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_2031),
.Y(n_2329)
);

INVx4_ASAP7_75t_L g2330 ( 
.A(n_1988),
.Y(n_2330)
);

INVx2_ASAP7_75t_L g2331 ( 
.A(n_2114),
.Y(n_2331)
);

NAND2xp5_ASAP7_75t_SL g2332 ( 
.A(n_1897),
.B(n_1494),
.Y(n_2332)
);

INVx3_ASAP7_75t_L g2333 ( 
.A(n_2032),
.Y(n_2333)
);

INVx2_ASAP7_75t_L g2334 ( 
.A(n_2117),
.Y(n_2334)
);

NAND2xp5_ASAP7_75t_L g2335 ( 
.A(n_2040),
.B(n_1488),
.Y(n_2335)
);

NOR2xp33_ASAP7_75t_L g2336 ( 
.A(n_2137),
.B(n_1491),
.Y(n_2336)
);

NAND2xp5_ASAP7_75t_L g2337 ( 
.A(n_2043),
.B(n_1497),
.Y(n_2337)
);

NAND2x1p5_ASAP7_75t_L g2338 ( 
.A(n_2093),
.B(n_2099),
.Y(n_2338)
);

INVx3_ASAP7_75t_L g2339 ( 
.A(n_2032),
.Y(n_2339)
);

NAND2xp5_ASAP7_75t_L g2340 ( 
.A(n_2045),
.B(n_1500),
.Y(n_2340)
);

NAND2xp5_ASAP7_75t_SL g2341 ( 
.A(n_1962),
.B(n_2083),
.Y(n_2341)
);

BUFx6f_ASAP7_75t_L g2342 ( 
.A(n_2033),
.Y(n_2342)
);

INVx2_ASAP7_75t_L g2343 ( 
.A(n_2033),
.Y(n_2343)
);

NAND2xp5_ASAP7_75t_L g2344 ( 
.A(n_2048),
.B(n_1914),
.Y(n_2344)
);

NAND2xp5_ASAP7_75t_L g2345 ( 
.A(n_2079),
.B(n_1527),
.Y(n_2345)
);

NAND2xp5_ASAP7_75t_L g2346 ( 
.A(n_2163),
.B(n_1895),
.Y(n_2346)
);

O2A1O1Ixp33_ASAP7_75t_L g2347 ( 
.A1(n_2086),
.A2(n_1440),
.B(n_1458),
.C(n_1438),
.Y(n_2347)
);

INVx1_ASAP7_75t_L g2348 ( 
.A(n_1995),
.Y(n_2348)
);

AND2x2_ASAP7_75t_L g2349 ( 
.A(n_1927),
.B(n_1431),
.Y(n_2349)
);

INVx2_ASAP7_75t_SL g2350 ( 
.A(n_2124),
.Y(n_2350)
);

INVx1_ASAP7_75t_L g2351 ( 
.A(n_2015),
.Y(n_2351)
);

OR2x2_ASAP7_75t_L g2352 ( 
.A(n_2116),
.B(n_959),
.Y(n_2352)
);

NAND2xp5_ASAP7_75t_SL g2353 ( 
.A(n_1884),
.B(n_961),
.Y(n_2353)
);

AND2x2_ASAP7_75t_L g2354 ( 
.A(n_1934),
.B(n_1515),
.Y(n_2354)
);

NAND2xp5_ASAP7_75t_SL g2355 ( 
.A(n_2061),
.B(n_966),
.Y(n_2355)
);

AND2x2_ASAP7_75t_SL g2356 ( 
.A(n_2129),
.B(n_1460),
.Y(n_2356)
);

NAND3xp33_ASAP7_75t_L g2357 ( 
.A(n_2049),
.B(n_968),
.C(n_967),
.Y(n_2357)
);

NAND2xp5_ASAP7_75t_L g2358 ( 
.A(n_2058),
.B(n_1505),
.Y(n_2358)
);

INVx2_ASAP7_75t_SL g2359 ( 
.A(n_2073),
.Y(n_2359)
);

INVx8_ASAP7_75t_L g2360 ( 
.A(n_1964),
.Y(n_2360)
);

NOR3xp33_ASAP7_75t_L g2361 ( 
.A(n_2103),
.B(n_974),
.C(n_971),
.Y(n_2361)
);

NAND2xp5_ASAP7_75t_SL g2362 ( 
.A(n_1912),
.B(n_979),
.Y(n_2362)
);

NOR2xp33_ASAP7_75t_L g2363 ( 
.A(n_1983),
.B(n_983),
.Y(n_2363)
);

INVx2_ASAP7_75t_L g2364 ( 
.A(n_2041),
.Y(n_2364)
);

NOR2xp33_ASAP7_75t_L g2365 ( 
.A(n_2055),
.B(n_984),
.Y(n_2365)
);

NOR2xp33_ASAP7_75t_L g2366 ( 
.A(n_2082),
.B(n_992),
.Y(n_2366)
);

AND2x2_ASAP7_75t_L g2367 ( 
.A(n_2092),
.B(n_2054),
.Y(n_2367)
);

NOR2xp33_ASAP7_75t_L g2368 ( 
.A(n_1978),
.B(n_993),
.Y(n_2368)
);

BUFx10_ASAP7_75t_L g2369 ( 
.A(n_1907),
.Y(n_2369)
);

INVx2_ASAP7_75t_SL g2370 ( 
.A(n_2113),
.Y(n_2370)
);

NAND2xp5_ASAP7_75t_L g2371 ( 
.A(n_2063),
.B(n_1519),
.Y(n_2371)
);

NAND2xp5_ASAP7_75t_L g2372 ( 
.A(n_2038),
.B(n_1485),
.Y(n_2372)
);

INVx2_ASAP7_75t_L g2373 ( 
.A(n_2041),
.Y(n_2373)
);

NAND2xp5_ASAP7_75t_SL g2374 ( 
.A(n_2102),
.B(n_994),
.Y(n_2374)
);

NAND2xp5_ASAP7_75t_SL g2375 ( 
.A(n_2118),
.B(n_1001),
.Y(n_2375)
);

NAND2xp5_ASAP7_75t_SL g2376 ( 
.A(n_1920),
.B(n_1003),
.Y(n_2376)
);

NAND2xp33_ASAP7_75t_L g2377 ( 
.A(n_1951),
.B(n_1214),
.Y(n_2377)
);

AND2x2_ASAP7_75t_L g2378 ( 
.A(n_2093),
.B(n_1020),
.Y(n_2378)
);

AOI22xp5_ASAP7_75t_L g2379 ( 
.A1(n_2074),
.A2(n_1008),
.B1(n_1016),
.B2(n_1011),
.Y(n_2379)
);

NAND2xp5_ASAP7_75t_L g2380 ( 
.A(n_1937),
.B(n_1518),
.Y(n_2380)
);

NAND2xp5_ASAP7_75t_SL g2381 ( 
.A(n_2085),
.B(n_1018),
.Y(n_2381)
);

NOR2xp33_ASAP7_75t_L g2382 ( 
.A(n_1904),
.B(n_2094),
.Y(n_2382)
);

AOI22xp5_ASAP7_75t_L g2383 ( 
.A1(n_2009),
.A2(n_1030),
.B1(n_1031),
.B2(n_1024),
.Y(n_2383)
);

NAND2xp5_ASAP7_75t_SL g2384 ( 
.A(n_1971),
.B(n_1032),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_2046),
.Y(n_2385)
);

NAND2x1_ASAP7_75t_L g2386 ( 
.A(n_1939),
.B(n_981),
.Y(n_2386)
);

INVxp67_ASAP7_75t_L g2387 ( 
.A(n_1891),
.Y(n_2387)
);

NAND2xp5_ASAP7_75t_L g2388 ( 
.A(n_1943),
.B(n_1514),
.Y(n_2388)
);

NAND3xp33_ASAP7_75t_L g2389 ( 
.A(n_2060),
.B(n_1055),
.C(n_1051),
.Y(n_2389)
);

NOR2xp33_ASAP7_75t_L g2390 ( 
.A(n_2087),
.B(n_1069),
.Y(n_2390)
);

NAND2xp5_ASAP7_75t_SL g2391 ( 
.A(n_2041),
.B(n_1074),
.Y(n_2391)
);

INVxp67_ASAP7_75t_L g2392 ( 
.A(n_2122),
.Y(n_2392)
);

O2A1O1Ixp5_ASAP7_75t_L g2393 ( 
.A1(n_1981),
.A2(n_1490),
.B(n_1517),
.C(n_1487),
.Y(n_2393)
);

AND2x2_ASAP7_75t_L g2394 ( 
.A(n_2091),
.B(n_1020),
.Y(n_2394)
);

NAND2xp5_ASAP7_75t_SL g2395 ( 
.A(n_2044),
.B(n_1098),
.Y(n_2395)
);

INVx1_ASAP7_75t_L g2396 ( 
.A(n_2050),
.Y(n_2396)
);

INVx1_ASAP7_75t_L g2397 ( 
.A(n_2051),
.Y(n_2397)
);

INVx2_ASAP7_75t_L g2398 ( 
.A(n_2044),
.Y(n_2398)
);

NAND3xp33_ASAP7_75t_SL g2399 ( 
.A(n_2123),
.B(n_1502),
.C(n_1498),
.Y(n_2399)
);

AND2x4_ASAP7_75t_L g2400 ( 
.A(n_1908),
.B(n_1027),
.Y(n_2400)
);

INVx2_ASAP7_75t_L g2401 ( 
.A(n_2044),
.Y(n_2401)
);

INVx2_ASAP7_75t_L g2402 ( 
.A(n_2057),
.Y(n_2402)
);

INVx2_ASAP7_75t_L g2403 ( 
.A(n_2057),
.Y(n_2403)
);

NAND2xp5_ASAP7_75t_SL g2404 ( 
.A(n_2057),
.B(n_1100),
.Y(n_2404)
);

INVx2_ASAP7_75t_SL g2405 ( 
.A(n_2011),
.Y(n_2405)
);

NAND2xp5_ASAP7_75t_L g2406 ( 
.A(n_2021),
.B(n_1102),
.Y(n_2406)
);

INVx2_ASAP7_75t_L g2407 ( 
.A(n_2026),
.Y(n_2407)
);

NAND2x1_ASAP7_75t_L g2408 ( 
.A(n_1946),
.B(n_981),
.Y(n_2408)
);

AND2x4_ASAP7_75t_L g2409 ( 
.A(n_1885),
.B(n_1044),
.Y(n_2409)
);

INVx2_ASAP7_75t_L g2410 ( 
.A(n_2042),
.Y(n_2410)
);

NAND2xp33_ASAP7_75t_L g2411 ( 
.A(n_2127),
.B(n_1214),
.Y(n_2411)
);

NAND2xp5_ASAP7_75t_SL g2412 ( 
.A(n_1913),
.B(n_1107),
.Y(n_2412)
);

INVx1_ASAP7_75t_L g2413 ( 
.A(n_2059),
.Y(n_2413)
);

BUFx3_ASAP7_75t_L g2414 ( 
.A(n_1969),
.Y(n_2414)
);

INVx1_ASAP7_75t_L g2415 ( 
.A(n_2119),
.Y(n_2415)
);

NAND2xp5_ASAP7_75t_L g2416 ( 
.A(n_2072),
.B(n_1117),
.Y(n_2416)
);

AND2x4_ASAP7_75t_L g2417 ( 
.A(n_1885),
.B(n_1910),
.Y(n_2417)
);

AND2x2_ASAP7_75t_L g2418 ( 
.A(n_2097),
.B(n_1062),
.Y(n_2418)
);

NAND2xp5_ASAP7_75t_L g2419 ( 
.A(n_2017),
.B(n_1118),
.Y(n_2419)
);

INVx2_ASAP7_75t_L g2420 ( 
.A(n_2047),
.Y(n_2420)
);

NAND2xp5_ASAP7_75t_SL g2421 ( 
.A(n_1916),
.B(n_1127),
.Y(n_2421)
);

NAND2xp5_ASAP7_75t_L g2422 ( 
.A(n_2065),
.B(n_1133),
.Y(n_2422)
);

OR2x6_ASAP7_75t_L g2423 ( 
.A(n_1910),
.B(n_1915),
.Y(n_2423)
);

NAND2xp5_ASAP7_75t_SL g2424 ( 
.A(n_1929),
.B(n_1155),
.Y(n_2424)
);

AOI22xp33_ASAP7_75t_L g2425 ( 
.A1(n_2077),
.A2(n_1372),
.B1(n_1383),
.B2(n_1059),
.Y(n_2425)
);

NAND2xp5_ASAP7_75t_L g2426 ( 
.A(n_2125),
.B(n_1162),
.Y(n_2426)
);

NAND2xp5_ASAP7_75t_SL g2427 ( 
.A(n_1942),
.B(n_1163),
.Y(n_2427)
);

BUFx3_ASAP7_75t_L g2428 ( 
.A(n_1969),
.Y(n_2428)
);

INVx1_ASAP7_75t_L g2429 ( 
.A(n_2121),
.Y(n_2429)
);

INVxp67_ASAP7_75t_L g2430 ( 
.A(n_2155),
.Y(n_2430)
);

BUFx6f_ASAP7_75t_L g2431 ( 
.A(n_2132),
.Y(n_2431)
);

NAND2xp5_ASAP7_75t_SL g2432 ( 
.A(n_1945),
.B(n_1169),
.Y(n_2432)
);

NAND2xp5_ASAP7_75t_L g2433 ( 
.A(n_2156),
.B(n_2159),
.Y(n_2433)
);

NAND2xp5_ASAP7_75t_L g2434 ( 
.A(n_2078),
.B(n_1172),
.Y(n_2434)
);

AND2x4_ASAP7_75t_L g2435 ( 
.A(n_1915),
.B(n_1046),
.Y(n_2435)
);

INVx2_ASAP7_75t_L g2436 ( 
.A(n_2056),
.Y(n_2436)
);

NAND2xp5_ASAP7_75t_L g2437 ( 
.A(n_2098),
.B(n_2107),
.Y(n_2437)
);

INVx1_ASAP7_75t_L g2438 ( 
.A(n_2064),
.Y(n_2438)
);

AOI22xp33_ASAP7_75t_L g2439 ( 
.A1(n_2066),
.A2(n_1372),
.B1(n_1383),
.B2(n_1059),
.Y(n_2439)
);

NOR2xp33_ASAP7_75t_L g2440 ( 
.A(n_1947),
.B(n_1197),
.Y(n_2440)
);

AND2x2_ASAP7_75t_L g2441 ( 
.A(n_1947),
.B(n_1062),
.Y(n_2441)
);

AOI22xp33_ASAP7_75t_L g2442 ( 
.A1(n_2070),
.A2(n_1405),
.B1(n_1456),
.B2(n_1403),
.Y(n_2442)
);

A2O1A1Ixp33_ASAP7_75t_L g2443 ( 
.A1(n_2076),
.A2(n_1050),
.B(n_1058),
.C(n_1056),
.Y(n_2443)
);

NAND2xp5_ASAP7_75t_L g2444 ( 
.A(n_1991),
.B(n_1204),
.Y(n_2444)
);

NAND2xp5_ASAP7_75t_L g2445 ( 
.A(n_1963),
.B(n_1205),
.Y(n_2445)
);

NAND2xp5_ASAP7_75t_L g2446 ( 
.A(n_1963),
.B(n_1213),
.Y(n_2446)
);

INVx2_ASAP7_75t_L g2447 ( 
.A(n_2141),
.Y(n_2447)
);

NAND2xp5_ASAP7_75t_SL g2448 ( 
.A(n_1965),
.B(n_1229),
.Y(n_2448)
);

INVx2_ASAP7_75t_L g2449 ( 
.A(n_2143),
.Y(n_2449)
);

INVxp67_ASAP7_75t_SL g2450 ( 
.A(n_2146),
.Y(n_2450)
);

NAND2xp5_ASAP7_75t_L g2451 ( 
.A(n_1954),
.B(n_1236),
.Y(n_2451)
);

NAND2xp5_ASAP7_75t_L g2452 ( 
.A(n_1957),
.B(n_1240),
.Y(n_2452)
);

NAND2xp5_ASAP7_75t_L g2453 ( 
.A(n_1961),
.B(n_1242),
.Y(n_2453)
);

AO221x1_ASAP7_75t_L g2454 ( 
.A1(n_2150),
.A2(n_1403),
.B1(n_1470),
.B2(n_1456),
.C(n_1405),
.Y(n_2454)
);

NAND2xp5_ASAP7_75t_SL g2455 ( 
.A(n_1966),
.B(n_1245),
.Y(n_2455)
);

NAND2xp5_ASAP7_75t_L g2456 ( 
.A(n_1967),
.B(n_1266),
.Y(n_2456)
);

NAND2xp33_ASAP7_75t_L g2457 ( 
.A(n_2153),
.B(n_1214),
.Y(n_2457)
);

NOR2xp33_ASAP7_75t_L g2458 ( 
.A(n_1992),
.B(n_1275),
.Y(n_2458)
);

AND3x2_ASAP7_75t_L g2459 ( 
.A(n_1973),
.B(n_1083),
.C(n_1078),
.Y(n_2459)
);

NOR2xp33_ASAP7_75t_L g2460 ( 
.A(n_2150),
.B(n_1278),
.Y(n_2460)
);

INVx1_ASAP7_75t_L g2461 ( 
.A(n_2018),
.Y(n_2461)
);

AND2x2_ASAP7_75t_L g2462 ( 
.A(n_2018),
.B(n_1147),
.Y(n_2462)
);

AND2x2_ASAP7_75t_L g2463 ( 
.A(n_1969),
.B(n_1147),
.Y(n_2463)
);

AOI22xp33_ASAP7_75t_L g2464 ( 
.A1(n_1975),
.A2(n_1405),
.B1(n_1456),
.B2(n_1403),
.Y(n_2464)
);

NAND2xp5_ASAP7_75t_SL g2465 ( 
.A(n_1974),
.B(n_1279),
.Y(n_2465)
);

INVx1_ASAP7_75t_L g2466 ( 
.A(n_1976),
.Y(n_2466)
);

NAND2xp5_ASAP7_75t_L g2467 ( 
.A(n_1977),
.B(n_1285),
.Y(n_2467)
);

NAND2xp5_ASAP7_75t_SL g2468 ( 
.A(n_1979),
.B(n_1293),
.Y(n_2468)
);

INVx2_ASAP7_75t_L g2469 ( 
.A(n_2162),
.Y(n_2469)
);

NAND2xp5_ASAP7_75t_L g2470 ( 
.A(n_2151),
.B(n_1294),
.Y(n_2470)
);

NAND2xp5_ASAP7_75t_L g2471 ( 
.A(n_2151),
.B(n_1314),
.Y(n_2471)
);

NAND2xp5_ASAP7_75t_L g2472 ( 
.A(n_1984),
.B(n_1319),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_1990),
.Y(n_2473)
);

AOI22xp5_ASAP7_75t_L g2474 ( 
.A1(n_2075),
.A2(n_1330),
.B1(n_1349),
.B2(n_1328),
.Y(n_2474)
);

NAND2xp5_ASAP7_75t_SL g2475 ( 
.A(n_2004),
.B(n_1354),
.Y(n_2475)
);

NAND2xp5_ASAP7_75t_L g2476 ( 
.A(n_2007),
.B(n_1356),
.Y(n_2476)
);

INVx1_ASAP7_75t_L g2477 ( 
.A(n_2020),
.Y(n_2477)
);

NAND2xp5_ASAP7_75t_L g2478 ( 
.A(n_2160),
.B(n_1364),
.Y(n_2478)
);

NAND2xp5_ASAP7_75t_L g2479 ( 
.A(n_2160),
.B(n_1369),
.Y(n_2479)
);

NAND2xp5_ASAP7_75t_SL g2480 ( 
.A(n_2160),
.B(n_1378),
.Y(n_2480)
);

NAND2xp5_ASAP7_75t_L g2481 ( 
.A(n_2164),
.B(n_1380),
.Y(n_2481)
);

NAND2xp5_ASAP7_75t_L g2482 ( 
.A(n_1909),
.B(n_1384),
.Y(n_2482)
);

NAND2xp5_ASAP7_75t_L g2483 ( 
.A(n_1909),
.B(n_1385),
.Y(n_2483)
);

NAND2xp5_ASAP7_75t_SL g2484 ( 
.A(n_1887),
.B(n_1389),
.Y(n_2484)
);

INVx2_ASAP7_75t_L g2485 ( 
.A(n_1896),
.Y(n_2485)
);

AOI22xp5_ASAP7_75t_L g2486 ( 
.A1(n_2019),
.A2(n_1397),
.B1(n_1400),
.B2(n_1395),
.Y(n_2486)
);

INVx8_ASAP7_75t_L g2487 ( 
.A(n_1997),
.Y(n_2487)
);

NOR2xp67_ASAP7_75t_L g2488 ( 
.A(n_1890),
.B(n_4),
.Y(n_2488)
);

NAND2xp5_ASAP7_75t_L g2489 ( 
.A(n_1909),
.B(n_1404),
.Y(n_2489)
);

INVx2_ASAP7_75t_SL g2490 ( 
.A(n_1894),
.Y(n_2490)
);

NAND2xp5_ASAP7_75t_L g2491 ( 
.A(n_1909),
.B(n_1406),
.Y(n_2491)
);

NAND2xp5_ASAP7_75t_L g2492 ( 
.A(n_1909),
.B(n_1408),
.Y(n_2492)
);

NOR2xp33_ASAP7_75t_L g2493 ( 
.A(n_2019),
.B(n_1409),
.Y(n_2493)
);

INVx2_ASAP7_75t_SL g2494 ( 
.A(n_1894),
.Y(n_2494)
);

INVx1_ASAP7_75t_L g2495 ( 
.A(n_1996),
.Y(n_2495)
);

NOR2xp33_ASAP7_75t_L g2496 ( 
.A(n_2019),
.B(n_1413),
.Y(n_2496)
);

NAND2xp5_ASAP7_75t_L g2497 ( 
.A(n_1909),
.B(n_1414),
.Y(n_2497)
);

AND2x2_ASAP7_75t_L g2498 ( 
.A(n_1887),
.B(n_1192),
.Y(n_2498)
);

NAND2xp5_ASAP7_75t_L g2499 ( 
.A(n_1909),
.B(n_1415),
.Y(n_2499)
);

BUFx2_ASAP7_75t_L g2500 ( 
.A(n_1894),
.Y(n_2500)
);

NAND2xp5_ASAP7_75t_L g2501 ( 
.A(n_1909),
.B(n_1417),
.Y(n_2501)
);

AOI22xp33_ASAP7_75t_L g2502 ( 
.A1(n_2039),
.A2(n_1405),
.B1(n_1456),
.B2(n_1403),
.Y(n_2502)
);

AOI221xp5_ASAP7_75t_L g2503 ( 
.A1(n_1879),
.A2(n_1084),
.B1(n_1116),
.B2(n_1113),
.C(n_1097),
.Y(n_2503)
);

NOR2xp33_ASAP7_75t_L g2504 ( 
.A(n_2019),
.B(n_1419),
.Y(n_2504)
);

OR2x2_ASAP7_75t_L g2505 ( 
.A(n_1887),
.B(n_1420),
.Y(n_2505)
);

INVx1_ASAP7_75t_L g2506 ( 
.A(n_1996),
.Y(n_2506)
);

NAND2xp5_ASAP7_75t_L g2507 ( 
.A(n_1909),
.B(n_1436),
.Y(n_2507)
);

AOI22xp5_ASAP7_75t_L g2508 ( 
.A1(n_2019),
.A2(n_1443),
.B1(n_1445),
.B2(n_1441),
.Y(n_2508)
);

INVx2_ASAP7_75t_L g2509 ( 
.A(n_1896),
.Y(n_2509)
);

NOR2xp33_ASAP7_75t_L g2510 ( 
.A(n_2019),
.B(n_1451),
.Y(n_2510)
);

INVxp67_ASAP7_75t_L g2511 ( 
.A(n_2138),
.Y(n_2511)
);

NAND2xp5_ASAP7_75t_L g2512 ( 
.A(n_1909),
.B(n_1446),
.Y(n_2512)
);

NAND2xp5_ASAP7_75t_SL g2513 ( 
.A(n_1887),
.B(n_1459),
.Y(n_2513)
);

INVx1_ASAP7_75t_L g2514 ( 
.A(n_1996),
.Y(n_2514)
);

NAND2xp5_ASAP7_75t_SL g2515 ( 
.A(n_1887),
.B(n_1465),
.Y(n_2515)
);

NAND2xp5_ASAP7_75t_L g2516 ( 
.A(n_1909),
.B(n_1469),
.Y(n_2516)
);

NAND2xp5_ASAP7_75t_L g2517 ( 
.A(n_1909),
.B(n_1471),
.Y(n_2517)
);

INVx1_ASAP7_75t_L g2518 ( 
.A(n_1996),
.Y(n_2518)
);

NAND2xp5_ASAP7_75t_L g2519 ( 
.A(n_1909),
.B(n_1472),
.Y(n_2519)
);

INVx1_ASAP7_75t_L g2520 ( 
.A(n_1996),
.Y(n_2520)
);

INVx2_ASAP7_75t_L g2521 ( 
.A(n_1896),
.Y(n_2521)
);

AOI22xp5_ASAP7_75t_L g2522 ( 
.A1(n_2019),
.A2(n_1492),
.B1(n_1493),
.B2(n_1482),
.Y(n_2522)
);

INVx2_ASAP7_75t_L g2523 ( 
.A(n_1896),
.Y(n_2523)
);

NAND2xp5_ASAP7_75t_SL g2524 ( 
.A(n_1887),
.B(n_1495),
.Y(n_2524)
);

NAND2xp5_ASAP7_75t_L g2525 ( 
.A(n_1909),
.B(n_1507),
.Y(n_2525)
);

HB1xp67_ASAP7_75t_L g2526 ( 
.A(n_1887),
.Y(n_2526)
);

HB1xp67_ASAP7_75t_L g2527 ( 
.A(n_1887),
.Y(n_2527)
);

NAND2xp5_ASAP7_75t_L g2528 ( 
.A(n_1909),
.B(n_1508),
.Y(n_2528)
);

INVx1_ASAP7_75t_L g2529 ( 
.A(n_1996),
.Y(n_2529)
);

INVx2_ASAP7_75t_L g2530 ( 
.A(n_1896),
.Y(n_2530)
);

INVx1_ASAP7_75t_L g2531 ( 
.A(n_1996),
.Y(n_2531)
);

NAND2xp5_ASAP7_75t_L g2532 ( 
.A(n_1909),
.B(n_1532),
.Y(n_2532)
);

INVx2_ASAP7_75t_L g2533 ( 
.A(n_1896),
.Y(n_2533)
);

NAND2xp5_ASAP7_75t_L g2534 ( 
.A(n_1909),
.B(n_1136),
.Y(n_2534)
);

INVx1_ASAP7_75t_L g2535 ( 
.A(n_1996),
.Y(n_2535)
);

NAND3xp33_ASAP7_75t_L g2536 ( 
.A(n_2255),
.B(n_1470),
.C(n_1288),
.Y(n_2536)
);

OAI21xp5_ASAP7_75t_L g2537 ( 
.A1(n_2182),
.A2(n_1150),
.B(n_1141),
.Y(n_2537)
);

NAND2xp5_ASAP7_75t_SL g2538 ( 
.A(n_2262),
.B(n_1192),
.Y(n_2538)
);

NAND2xp5_ASAP7_75t_L g2539 ( 
.A(n_2264),
.B(n_2197),
.Y(n_2539)
);

AOI21xp33_ASAP7_75t_L g2540 ( 
.A1(n_2221),
.A2(n_1157),
.B(n_1156),
.Y(n_2540)
);

NAND2xp5_ASAP7_75t_L g2541 ( 
.A(n_2229),
.B(n_1504),
.Y(n_2541)
);

NAND2xp5_ASAP7_75t_L g2542 ( 
.A(n_2205),
.B(n_1516),
.Y(n_2542)
);

BUFx2_ASAP7_75t_L g2543 ( 
.A(n_2526),
.Y(n_2543)
);

NAND2xp5_ASAP7_75t_L g2544 ( 
.A(n_2234),
.B(n_1520),
.Y(n_2544)
);

HB1xp67_ASAP7_75t_L g2545 ( 
.A(n_2527),
.Y(n_2545)
);

INVx2_ASAP7_75t_L g2546 ( 
.A(n_2254),
.Y(n_2546)
);

O2A1O1Ixp33_ASAP7_75t_L g2547 ( 
.A1(n_2248),
.A2(n_1183),
.B(n_1211),
.C(n_1180),
.Y(n_2547)
);

BUFx6f_ASAP7_75t_L g2548 ( 
.A(n_2233),
.Y(n_2548)
);

AOI22xp5_ASAP7_75t_L g2549 ( 
.A1(n_2213),
.A2(n_1338),
.B1(n_1480),
.B2(n_1289),
.Y(n_2549)
);

OAI21xp5_ASAP7_75t_L g2550 ( 
.A1(n_2461),
.A2(n_1468),
.B(n_1463),
.Y(n_2550)
);

AOI21xp5_ASAP7_75t_L g2551 ( 
.A1(n_2450),
.A2(n_1227),
.B(n_1217),
.Y(n_2551)
);

OAI22xp5_ASAP7_75t_L g2552 ( 
.A1(n_2299),
.A2(n_1470),
.B1(n_1231),
.B2(n_1235),
.Y(n_2552)
);

NOR2xp33_ASAP7_75t_L g2553 ( 
.A(n_2511),
.B(n_1289),
.Y(n_2553)
);

INVx5_ASAP7_75t_L g2554 ( 
.A(n_2281),
.Y(n_2554)
);

AOI21xp5_ASAP7_75t_L g2555 ( 
.A1(n_2447),
.A2(n_2469),
.B(n_2449),
.Y(n_2555)
);

NAND2xp5_ASAP7_75t_SL g2556 ( 
.A(n_2209),
.B(n_1338),
.Y(n_2556)
);

AOI21xp5_ASAP7_75t_L g2557 ( 
.A1(n_2437),
.A2(n_1244),
.B(n_1230),
.Y(n_2557)
);

INVx4_ASAP7_75t_L g2558 ( 
.A(n_2281),
.Y(n_2558)
);

INVx2_ASAP7_75t_L g2559 ( 
.A(n_2173),
.Y(n_2559)
);

OAI21xp33_ASAP7_75t_L g2560 ( 
.A1(n_2259),
.A2(n_1263),
.B(n_1247),
.Y(n_2560)
);

OAI21xp5_ASAP7_75t_L g2561 ( 
.A1(n_2252),
.A2(n_1297),
.B(n_1284),
.Y(n_2561)
);

OR2x6_ASAP7_75t_L g2562 ( 
.A(n_2487),
.B(n_1039),
.Y(n_2562)
);

AOI21xp5_ASAP7_75t_L g2563 ( 
.A1(n_2481),
.A2(n_1351),
.B(n_1307),
.Y(n_2563)
);

INVx1_ASAP7_75t_L g2564 ( 
.A(n_2218),
.Y(n_2564)
);

INVx1_ASAP7_75t_L g2565 ( 
.A(n_2224),
.Y(n_2565)
);

NOR2xp33_ASAP7_75t_L g2566 ( 
.A(n_2241),
.B(n_1480),
.Y(n_2566)
);

NOR2xp33_ASAP7_75t_L g2567 ( 
.A(n_2226),
.B(n_1444),
.Y(n_2567)
);

OAI21xp5_ASAP7_75t_L g2568 ( 
.A1(n_2348),
.A2(n_1392),
.B(n_1375),
.Y(n_2568)
);

NAND2xp5_ASAP7_75t_L g2569 ( 
.A(n_2225),
.B(n_1474),
.Y(n_2569)
);

INVx3_ASAP7_75t_L g2570 ( 
.A(n_2231),
.Y(n_2570)
);

AOI22xp5_ASAP7_75t_L g2571 ( 
.A1(n_2210),
.A2(n_1407),
.B1(n_1412),
.B2(n_1399),
.Y(n_2571)
);

NOR2xp33_ASAP7_75t_L g2572 ( 
.A(n_2228),
.B(n_1486),
.Y(n_2572)
);

NOR2xp33_ASAP7_75t_L g2573 ( 
.A(n_2349),
.B(n_1496),
.Y(n_2573)
);

AOI21xp5_ASAP7_75t_L g2574 ( 
.A1(n_2411),
.A2(n_1426),
.B(n_1425),
.Y(n_2574)
);

OAI22xp5_ASAP7_75t_L g2575 ( 
.A1(n_2344),
.A2(n_2387),
.B1(n_2392),
.B2(n_2309),
.Y(n_2575)
);

AND2x2_ASAP7_75t_L g2576 ( 
.A(n_2327),
.B(n_2493),
.Y(n_2576)
);

NOR2xp33_ASAP7_75t_L g2577 ( 
.A(n_2354),
.B(n_1534),
.Y(n_2577)
);

NAND2xp5_ASAP7_75t_L g2578 ( 
.A(n_2180),
.B(n_1430),
.Y(n_2578)
);

INVx2_ASAP7_75t_L g2579 ( 
.A(n_2186),
.Y(n_2579)
);

NAND2xp5_ASAP7_75t_L g2580 ( 
.A(n_2495),
.B(n_1449),
.Y(n_2580)
);

NAND2xp5_ASAP7_75t_SL g2581 ( 
.A(n_2256),
.B(n_1470),
.Y(n_2581)
);

AOI21x1_ASAP7_75t_L g2582 ( 
.A1(n_2167),
.A2(n_1052),
.B(n_1039),
.Y(n_2582)
);

AOI21xp5_ASAP7_75t_L g2583 ( 
.A1(n_2457),
.A2(n_1484),
.B(n_1478),
.Y(n_2583)
);

AOI21xp5_ASAP7_75t_L g2584 ( 
.A1(n_2261),
.A2(n_1501),
.B(n_1121),
.Y(n_2584)
);

AOI21xp5_ASAP7_75t_L g2585 ( 
.A1(n_2270),
.A2(n_1121),
.B(n_1052),
.Y(n_2585)
);

AOI21xp5_ASAP7_75t_L g2586 ( 
.A1(n_2385),
.A2(n_1174),
.B(n_1168),
.Y(n_2586)
);

NOR2xp67_ASAP7_75t_L g2587 ( 
.A(n_2330),
.B(n_4),
.Y(n_2587)
);

NAND2xp5_ASAP7_75t_L g2588 ( 
.A(n_2506),
.B(n_2514),
.Y(n_2588)
);

NAND2xp5_ASAP7_75t_L g2589 ( 
.A(n_2518),
.B(n_1168),
.Y(n_2589)
);

NOR2xp33_ASAP7_75t_L g2590 ( 
.A(n_2269),
.B(n_1174),
.Y(n_2590)
);

AO21x1_ASAP7_75t_L g2591 ( 
.A1(n_2200),
.A2(n_1298),
.B(n_1264),
.Y(n_2591)
);

NAND2xp5_ASAP7_75t_L g2592 ( 
.A(n_2520),
.B(n_1264),
.Y(n_2592)
);

NOR2xp33_ASAP7_75t_L g2593 ( 
.A(n_2285),
.B(n_1298),
.Y(n_2593)
);

AOI21xp33_ASAP7_75t_L g2594 ( 
.A1(n_2496),
.A2(n_1457),
.B(n_1342),
.Y(n_2594)
);

OAI21xp5_ASAP7_75t_L g2595 ( 
.A1(n_2306),
.A2(n_1457),
.B(n_1342),
.Y(n_2595)
);

NAND2xp5_ASAP7_75t_L g2596 ( 
.A(n_2529),
.B(n_1489),
.Y(n_2596)
);

AOI21xp5_ASAP7_75t_L g2597 ( 
.A1(n_2396),
.A2(n_1503),
.B(n_1489),
.Y(n_2597)
);

NOR2xp67_ASAP7_75t_L g2598 ( 
.A(n_2330),
.B(n_5),
.Y(n_2598)
);

INVx1_ASAP7_75t_L g2599 ( 
.A(n_2531),
.Y(n_2599)
);

INVx1_ASAP7_75t_L g2600 ( 
.A(n_2535),
.Y(n_2600)
);

NAND2xp5_ASAP7_75t_L g2601 ( 
.A(n_2347),
.B(n_1503),
.Y(n_2601)
);

INVx2_ASAP7_75t_L g2602 ( 
.A(n_2292),
.Y(n_2602)
);

NAND2xp5_ASAP7_75t_L g2603 ( 
.A(n_2188),
.B(n_1512),
.Y(n_2603)
);

INVx2_ASAP7_75t_L g2604 ( 
.A(n_2314),
.Y(n_2604)
);

AOI33xp33_ASAP7_75t_L g2605 ( 
.A1(n_2503),
.A2(n_1512),
.A3(n_7),
.B1(n_9),
.B2(n_5),
.B3(n_6),
.Y(n_2605)
);

AOI22xp5_ASAP7_75t_L g2606 ( 
.A1(n_2268),
.A2(n_1288),
.B1(n_1281),
.B2(n_8),
.Y(n_2606)
);

OAI21xp5_ASAP7_75t_L g2607 ( 
.A1(n_2393),
.A2(n_1288),
.B(n_1281),
.Y(n_2607)
);

AOI21xp5_ASAP7_75t_L g2608 ( 
.A1(n_2397),
.A2(n_1288),
.B(n_1281),
.Y(n_2608)
);

NOR2xp33_ASAP7_75t_L g2609 ( 
.A(n_2277),
.B(n_6),
.Y(n_2609)
);

O2A1O1Ixp5_ASAP7_75t_L g2610 ( 
.A1(n_2341),
.A2(n_1281),
.B(n_8),
.C(n_6),
.Y(n_2610)
);

NAND2xp5_ASAP7_75t_L g2611 ( 
.A(n_2189),
.B(n_7),
.Y(n_2611)
);

NAND2xp5_ASAP7_75t_L g2612 ( 
.A(n_2191),
.B(n_7),
.Y(n_2612)
);

INVx1_ASAP7_75t_L g2613 ( 
.A(n_2244),
.Y(n_2613)
);

AOI22xp5_ASAP7_75t_L g2614 ( 
.A1(n_2198),
.A2(n_12),
.B1(n_10),
.B2(n_11),
.Y(n_2614)
);

OAI22xp5_ASAP7_75t_L g2615 ( 
.A1(n_2326),
.A2(n_12),
.B1(n_10),
.B2(n_11),
.Y(n_2615)
);

NAND2xp5_ASAP7_75t_L g2616 ( 
.A(n_2196),
.B(n_10),
.Y(n_2616)
);

NAND2xp5_ASAP7_75t_L g2617 ( 
.A(n_2208),
.B(n_11),
.Y(n_2617)
);

NAND2xp5_ASAP7_75t_L g2618 ( 
.A(n_2230),
.B(n_2237),
.Y(n_2618)
);

AOI21xp5_ASAP7_75t_L g2619 ( 
.A1(n_2413),
.A2(n_2172),
.B(n_2168),
.Y(n_2619)
);

INVx1_ASAP7_75t_L g2620 ( 
.A(n_2250),
.Y(n_2620)
);

NAND2xp33_ASAP7_75t_L g2621 ( 
.A(n_2249),
.B(n_14),
.Y(n_2621)
);

NAND2xp5_ASAP7_75t_L g2622 ( 
.A(n_2280),
.B(n_13),
.Y(n_2622)
);

NAND2xp5_ASAP7_75t_L g2623 ( 
.A(n_2358),
.B(n_13),
.Y(n_2623)
);

NAND2xp5_ASAP7_75t_L g2624 ( 
.A(n_2371),
.B(n_13),
.Y(n_2624)
);

NOR2xp33_ASAP7_75t_L g2625 ( 
.A(n_2305),
.B(n_14),
.Y(n_2625)
);

BUFx12f_ASAP7_75t_L g2626 ( 
.A(n_2232),
.Y(n_2626)
);

NAND2xp5_ASAP7_75t_L g2627 ( 
.A(n_2345),
.B(n_15),
.Y(n_2627)
);

NAND2xp5_ASAP7_75t_SL g2628 ( 
.A(n_2308),
.B(n_16),
.Y(n_2628)
);

AOI21xp5_ASAP7_75t_L g2629 ( 
.A1(n_2177),
.A2(n_15),
.B(n_16),
.Y(n_2629)
);

NOR2xp33_ASAP7_75t_L g2630 ( 
.A(n_2324),
.B(n_17),
.Y(n_2630)
);

NAND2xp5_ASAP7_75t_L g2631 ( 
.A(n_2534),
.B(n_18),
.Y(n_2631)
);

AOI21xp5_ASAP7_75t_L g2632 ( 
.A1(n_2485),
.A2(n_20),
.B(n_21),
.Y(n_2632)
);

INVx1_ASAP7_75t_L g2633 ( 
.A(n_2263),
.Y(n_2633)
);

INVx2_ASAP7_75t_L g2634 ( 
.A(n_2331),
.Y(n_2634)
);

NAND2xp5_ASAP7_75t_SL g2635 ( 
.A(n_2249),
.B(n_21),
.Y(n_2635)
);

OAI21xp33_ASAP7_75t_L g2636 ( 
.A1(n_2310),
.A2(n_20),
.B(n_21),
.Y(n_2636)
);

AND2x2_ASAP7_75t_L g2637 ( 
.A(n_2504),
.B(n_20),
.Y(n_2637)
);

OAI21xp33_ASAP7_75t_L g2638 ( 
.A1(n_2276),
.A2(n_22),
.B(n_23),
.Y(n_2638)
);

AOI21xp5_ASAP7_75t_L g2639 ( 
.A1(n_2509),
.A2(n_22),
.B(n_23),
.Y(n_2639)
);

AOI21xp5_ASAP7_75t_L g2640 ( 
.A1(n_2521),
.A2(n_2530),
.B(n_2523),
.Y(n_2640)
);

INVx2_ASAP7_75t_L g2641 ( 
.A(n_2334),
.Y(n_2641)
);

NOR2xp33_ASAP7_75t_SL g2642 ( 
.A(n_2289),
.B(n_22),
.Y(n_2642)
);

AOI21xp5_ASAP7_75t_L g2643 ( 
.A1(n_2533),
.A2(n_23),
.B(n_24),
.Y(n_2643)
);

O2A1O1Ixp33_ASAP7_75t_L g2644 ( 
.A1(n_2443),
.A2(n_26),
.B(n_24),
.C(n_25),
.Y(n_2644)
);

NAND2xp5_ASAP7_75t_L g2645 ( 
.A(n_2204),
.B(n_24),
.Y(n_2645)
);

NOR2xp33_ASAP7_75t_L g2646 ( 
.A(n_2315),
.B(n_25),
.Y(n_2646)
);

AND2x2_ASAP7_75t_L g2647 ( 
.A(n_2510),
.B(n_2243),
.Y(n_2647)
);

NAND2xp5_ASAP7_75t_L g2648 ( 
.A(n_2302),
.B(n_2303),
.Y(n_2648)
);

NOR2xp33_ASAP7_75t_L g2649 ( 
.A(n_2169),
.B(n_25),
.Y(n_2649)
);

HB1xp67_ASAP7_75t_L g2650 ( 
.A(n_2500),
.Y(n_2650)
);

O2A1O1Ixp33_ASAP7_75t_L g2651 ( 
.A1(n_2251),
.A2(n_29),
.B(n_27),
.C(n_28),
.Y(n_2651)
);

NOR3xp33_ASAP7_75t_L g2652 ( 
.A(n_2399),
.B(n_29),
.C(n_28),
.Y(n_2652)
);

INVx1_ASAP7_75t_L g2653 ( 
.A(n_2279),
.Y(n_2653)
);

INVx1_ASAP7_75t_L g2654 ( 
.A(n_2291),
.Y(n_2654)
);

O2A1O1Ixp33_ASAP7_75t_L g2655 ( 
.A1(n_2346),
.A2(n_29),
.B(n_27),
.C(n_28),
.Y(n_2655)
);

AND2x2_ASAP7_75t_L g2656 ( 
.A(n_2194),
.B(n_27),
.Y(n_2656)
);

OAI21xp5_ASAP7_75t_L g2657 ( 
.A1(n_2351),
.A2(n_30),
.B(n_31),
.Y(n_2657)
);

NAND2xp5_ASAP7_75t_L g2658 ( 
.A(n_2242),
.B(n_30),
.Y(n_2658)
);

NAND2xp5_ASAP7_75t_L g2659 ( 
.A(n_2247),
.B(n_32),
.Y(n_2659)
);

NAND2xp5_ASAP7_75t_SL g2660 ( 
.A(n_2249),
.B(n_33),
.Y(n_2660)
);

BUFx12f_ASAP7_75t_L g2661 ( 
.A(n_2232),
.Y(n_2661)
);

INVx3_ASAP7_75t_L g2662 ( 
.A(n_2231),
.Y(n_2662)
);

BUFx4f_ASAP7_75t_L g2663 ( 
.A(n_2487),
.Y(n_2663)
);

NAND2xp5_ASAP7_75t_L g2664 ( 
.A(n_2171),
.B(n_32),
.Y(n_2664)
);

NAND2xp5_ASAP7_75t_L g2665 ( 
.A(n_2170),
.B(n_32),
.Y(n_2665)
);

INVx1_ASAP7_75t_L g2666 ( 
.A(n_2295),
.Y(n_2666)
);

BUFx2_ASAP7_75t_L g2667 ( 
.A(n_2260),
.Y(n_2667)
);

BUFx12f_ASAP7_75t_L g2668 ( 
.A(n_2369),
.Y(n_2668)
);

NAND2xp5_ASAP7_75t_SL g2669 ( 
.A(n_2249),
.B(n_34),
.Y(n_2669)
);

AOI21xp5_ASAP7_75t_L g2670 ( 
.A1(n_2377),
.A2(n_33),
.B(n_34),
.Y(n_2670)
);

AOI21xp5_ASAP7_75t_L g2671 ( 
.A1(n_2431),
.A2(n_33),
.B(n_34),
.Y(n_2671)
);

CKINVDCx5p33_ASAP7_75t_R g2672 ( 
.A(n_2360),
.Y(n_2672)
);

NOR2x1p5_ASAP7_75t_L g2673 ( 
.A(n_2207),
.B(n_35),
.Y(n_2673)
);

INVx3_ASAP7_75t_L g2674 ( 
.A(n_2249),
.Y(n_2674)
);

NAND2xp5_ASAP7_75t_L g2675 ( 
.A(n_2175),
.B(n_35),
.Y(n_2675)
);

NAND2xp5_ASAP7_75t_SL g2676 ( 
.A(n_2203),
.B(n_36),
.Y(n_2676)
);

OAI21xp5_ASAP7_75t_L g2677 ( 
.A1(n_2185),
.A2(n_2202),
.B(n_2195),
.Y(n_2677)
);

NAND2xp5_ASAP7_75t_L g2678 ( 
.A(n_2321),
.B(n_2367),
.Y(n_2678)
);

NAND2xp5_ASAP7_75t_L g2679 ( 
.A(n_2178),
.B(n_35),
.Y(n_2679)
);

AND2x2_ASAP7_75t_L g2680 ( 
.A(n_2498),
.B(n_36),
.Y(n_2680)
);

INVx2_ASAP7_75t_L g2681 ( 
.A(n_2211),
.Y(n_2681)
);

OAI21xp5_ASAP7_75t_L g2682 ( 
.A1(n_2220),
.A2(n_36),
.B(n_37),
.Y(n_2682)
);

AOI21xp5_ASAP7_75t_L g2683 ( 
.A1(n_2431),
.A2(n_37),
.B(n_38),
.Y(n_2683)
);

NAND2xp5_ASAP7_75t_L g2684 ( 
.A(n_2181),
.B(n_37),
.Y(n_2684)
);

AOI21xp5_ASAP7_75t_L g2685 ( 
.A1(n_2431),
.A2(n_38),
.B(n_39),
.Y(n_2685)
);

NAND2xp5_ASAP7_75t_L g2686 ( 
.A(n_2183),
.B(n_38),
.Y(n_2686)
);

INVx2_ASAP7_75t_SL g2687 ( 
.A(n_2289),
.Y(n_2687)
);

AOI22xp5_ASAP7_75t_L g2688 ( 
.A1(n_2215),
.A2(n_41),
.B1(n_39),
.B2(n_40),
.Y(n_2688)
);

NAND2xp5_ASAP7_75t_L g2689 ( 
.A(n_2192),
.B(n_39),
.Y(n_2689)
);

AOI21xp5_ASAP7_75t_L g2690 ( 
.A1(n_2267),
.A2(n_40),
.B(n_41),
.Y(n_2690)
);

AND2x2_ASAP7_75t_L g2691 ( 
.A(n_2253),
.B(n_40),
.Y(n_2691)
);

INVx1_ASAP7_75t_L g2692 ( 
.A(n_2296),
.Y(n_2692)
);

NAND2xp5_ASAP7_75t_L g2693 ( 
.A(n_2193),
.B(n_41),
.Y(n_2693)
);

INVx2_ASAP7_75t_L g2694 ( 
.A(n_2236),
.Y(n_2694)
);

NAND2xp5_ASAP7_75t_L g2695 ( 
.A(n_2297),
.B(n_42),
.Y(n_2695)
);

NAND2xp5_ASAP7_75t_L g2696 ( 
.A(n_2240),
.B(n_42),
.Y(n_2696)
);

NAND2xp5_ASAP7_75t_L g2697 ( 
.A(n_2246),
.B(n_42),
.Y(n_2697)
);

NOR3xp33_ASAP7_75t_L g2698 ( 
.A(n_2199),
.B(n_45),
.C(n_44),
.Y(n_2698)
);

OAI21xp5_ASAP7_75t_L g2699 ( 
.A1(n_2238),
.A2(n_43),
.B(n_44),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_2301),
.Y(n_2700)
);

NAND2xp5_ASAP7_75t_L g2701 ( 
.A(n_2312),
.B(n_43),
.Y(n_2701)
);

BUFx6f_ASAP7_75t_L g2702 ( 
.A(n_2233),
.Y(n_2702)
);

INVx1_ASAP7_75t_L g2703 ( 
.A(n_2320),
.Y(n_2703)
);

AOI21xp5_ASAP7_75t_L g2704 ( 
.A1(n_2275),
.A2(n_43),
.B(n_45),
.Y(n_2704)
);

AOI21xp5_ASAP7_75t_L g2705 ( 
.A1(n_2278),
.A2(n_45),
.B(n_46),
.Y(n_2705)
);

NAND2xp5_ASAP7_75t_L g2706 ( 
.A(n_2329),
.B(n_46),
.Y(n_2706)
);

AOI21xp5_ASAP7_75t_L g2707 ( 
.A1(n_2282),
.A2(n_46),
.B(n_47),
.Y(n_2707)
);

O2A1O1Ixp33_ASAP7_75t_L g2708 ( 
.A1(n_2212),
.A2(n_49),
.B(n_47),
.C(n_48),
.Y(n_2708)
);

OAI21xp5_ASAP7_75t_L g2709 ( 
.A1(n_2462),
.A2(n_48),
.B(n_49),
.Y(n_2709)
);

AOI21xp5_ASAP7_75t_L g2710 ( 
.A1(n_2283),
.A2(n_2328),
.B(n_2286),
.Y(n_2710)
);

INVx2_ASAP7_75t_L g2711 ( 
.A(n_2407),
.Y(n_2711)
);

NAND2xp5_ASAP7_75t_SL g2712 ( 
.A(n_2490),
.B(n_50),
.Y(n_2712)
);

AO21x1_ASAP7_75t_L g2713 ( 
.A1(n_2271),
.A2(n_2311),
.B(n_2307),
.Y(n_2713)
);

NAND2xp5_ASAP7_75t_SL g2714 ( 
.A(n_2494),
.B(n_50),
.Y(n_2714)
);

AOI21xp5_ASAP7_75t_L g2715 ( 
.A1(n_2335),
.A2(n_49),
.B(n_51),
.Y(n_2715)
);

BUFx3_ASAP7_75t_L g2716 ( 
.A(n_2360),
.Y(n_2716)
);

O2A1O1Ixp5_ASAP7_75t_L g2717 ( 
.A1(n_2391),
.A2(n_2395),
.B(n_2404),
.C(n_2284),
.Y(n_2717)
);

INVx3_ASAP7_75t_L g2718 ( 
.A(n_2417),
.Y(n_2718)
);

AND2x2_ASAP7_75t_L g2719 ( 
.A(n_2323),
.B(n_51),
.Y(n_2719)
);

INVx2_ASAP7_75t_SL g2720 ( 
.A(n_2201),
.Y(n_2720)
);

A2O1A1Ixp33_ASAP7_75t_L g2721 ( 
.A1(n_2488),
.A2(n_54),
.B(n_52),
.C(n_53),
.Y(n_2721)
);

INVx1_ASAP7_75t_L g2722 ( 
.A(n_2409),
.Y(n_2722)
);

OAI21xp5_ASAP7_75t_L g2723 ( 
.A1(n_2179),
.A2(n_52),
.B(n_53),
.Y(n_2723)
);

AOI21xp5_ASAP7_75t_L g2724 ( 
.A1(n_2337),
.A2(n_52),
.B(n_53),
.Y(n_2724)
);

OAI21xp33_ASAP7_75t_L g2725 ( 
.A1(n_2298),
.A2(n_54),
.B(n_55),
.Y(n_2725)
);

NAND2xp5_ASAP7_75t_L g2726 ( 
.A(n_2340),
.B(n_54),
.Y(n_2726)
);

NAND2xp5_ASAP7_75t_L g2727 ( 
.A(n_2217),
.B(n_55),
.Y(n_2727)
);

NOR2xp33_ASAP7_75t_L g2728 ( 
.A(n_2304),
.B(n_56),
.Y(n_2728)
);

AND2x6_ASAP7_75t_L g2729 ( 
.A(n_2233),
.B(n_2245),
.Y(n_2729)
);

NOR2xp33_ASAP7_75t_L g2730 ( 
.A(n_2505),
.B(n_57),
.Y(n_2730)
);

BUFx2_ASAP7_75t_L g2731 ( 
.A(n_2260),
.Y(n_2731)
);

NAND2xp5_ASAP7_75t_L g2732 ( 
.A(n_2223),
.B(n_57),
.Y(n_2732)
);

INVx1_ASAP7_75t_L g2733 ( 
.A(n_2409),
.Y(n_2733)
);

AO21x1_ASAP7_75t_L g2734 ( 
.A1(n_2300),
.A2(n_2466),
.B(n_2318),
.Y(n_2734)
);

NAND2xp5_ASAP7_75t_SL g2735 ( 
.A(n_2356),
.B(n_58),
.Y(n_2735)
);

OAI21xp5_ASAP7_75t_L g2736 ( 
.A1(n_2235),
.A2(n_57),
.B(n_58),
.Y(n_2736)
);

O2A1O1Ixp33_ASAP7_75t_L g2737 ( 
.A1(n_2482),
.A2(n_60),
.B(n_58),
.C(n_59),
.Y(n_2737)
);

O2A1O1Ixp33_ASAP7_75t_L g2738 ( 
.A1(n_2483),
.A2(n_61),
.B(n_59),
.C(n_60),
.Y(n_2738)
);

O2A1O1Ixp5_ASAP7_75t_L g2739 ( 
.A1(n_2274),
.A2(n_61),
.B(n_59),
.C(n_60),
.Y(n_2739)
);

OAI21xp5_ASAP7_75t_L g2740 ( 
.A1(n_2438),
.A2(n_61),
.B(n_62),
.Y(n_2740)
);

AOI21xp5_ASAP7_75t_L g2741 ( 
.A1(n_2381),
.A2(n_62),
.B(n_63),
.Y(n_2741)
);

NAND2xp5_ASAP7_75t_L g2742 ( 
.A(n_2214),
.B(n_62),
.Y(n_2742)
);

INVx2_ASAP7_75t_L g2743 ( 
.A(n_2410),
.Y(n_2743)
);

NAND2xp5_ASAP7_75t_L g2744 ( 
.A(n_2214),
.B(n_63),
.Y(n_2744)
);

AOI21xp5_ASAP7_75t_L g2745 ( 
.A1(n_2245),
.A2(n_63),
.B(n_64),
.Y(n_2745)
);

OAI22xp5_ASAP7_75t_L g2746 ( 
.A1(n_2245),
.A2(n_66),
.B1(n_64),
.B2(n_65),
.Y(n_2746)
);

OAI21xp5_ASAP7_75t_L g2747 ( 
.A1(n_2257),
.A2(n_66),
.B(n_67),
.Y(n_2747)
);

NAND2xp5_ASAP7_75t_L g2748 ( 
.A(n_2489),
.B(n_67),
.Y(n_2748)
);

NAND2xp5_ASAP7_75t_L g2749 ( 
.A(n_2491),
.B(n_2492),
.Y(n_2749)
);

NOR3xp33_ASAP7_75t_L g2750 ( 
.A(n_2357),
.B(n_69),
.C(n_68),
.Y(n_2750)
);

AOI21xp5_ASAP7_75t_L g2751 ( 
.A1(n_2258),
.A2(n_2384),
.B(n_2416),
.Y(n_2751)
);

OAI21xp5_ASAP7_75t_L g2752 ( 
.A1(n_2420),
.A2(n_70),
.B(n_71),
.Y(n_2752)
);

AND2x2_ASAP7_75t_L g2753 ( 
.A(n_2184),
.B(n_72),
.Y(n_2753)
);

NOR2xp33_ASAP7_75t_L g2754 ( 
.A(n_2497),
.B(n_72),
.Y(n_2754)
);

NAND2xp5_ASAP7_75t_SL g2755 ( 
.A(n_2313),
.B(n_74),
.Y(n_2755)
);

NAND2xp5_ASAP7_75t_L g2756 ( 
.A(n_2499),
.B(n_2501),
.Y(n_2756)
);

CKINVDCx8_ASAP7_75t_R g2757 ( 
.A(n_2239),
.Y(n_2757)
);

INVx1_ASAP7_75t_L g2758 ( 
.A(n_2435),
.Y(n_2758)
);

AOI33xp33_ASAP7_75t_L g2759 ( 
.A1(n_2418),
.A2(n_75),
.A3(n_77),
.B1(n_73),
.B2(n_74),
.B3(n_76),
.Y(n_2759)
);

OAI22xp33_ASAP7_75t_L g2760 ( 
.A1(n_2239),
.A2(n_75),
.B1(n_73),
.B2(n_74),
.Y(n_2760)
);

A2O1A1Ixp33_ASAP7_75t_L g2761 ( 
.A1(n_2316),
.A2(n_78),
.B(n_76),
.C(n_77),
.Y(n_2761)
);

OAI22xp5_ASAP7_75t_L g2762 ( 
.A1(n_2380),
.A2(n_79),
.B1(n_76),
.B2(n_78),
.Y(n_2762)
);

AOI21xp5_ASAP7_75t_L g2763 ( 
.A1(n_2375),
.A2(n_78),
.B(n_79),
.Y(n_2763)
);

NAND2xp5_ASAP7_75t_L g2764 ( 
.A(n_2507),
.B(n_80),
.Y(n_2764)
);

OAI321xp33_ASAP7_75t_L g2765 ( 
.A1(n_2502),
.A2(n_82),
.A3(n_84),
.B1(n_80),
.B2(n_81),
.C(n_83),
.Y(n_2765)
);

NAND2xp5_ASAP7_75t_L g2766 ( 
.A(n_2512),
.B(n_80),
.Y(n_2766)
);

NAND2xp5_ASAP7_75t_L g2767 ( 
.A(n_2516),
.B(n_81),
.Y(n_2767)
);

O2A1O1Ixp33_ASAP7_75t_L g2768 ( 
.A1(n_2517),
.A2(n_83),
.B(n_81),
.C(n_82),
.Y(n_2768)
);

INVx3_ASAP7_75t_L g2769 ( 
.A(n_2417),
.Y(n_2769)
);

A2O1A1Ixp33_ASAP7_75t_L g2770 ( 
.A1(n_2336),
.A2(n_85),
.B(n_82),
.C(n_83),
.Y(n_2770)
);

O2A1O1Ixp33_ASAP7_75t_L g2771 ( 
.A1(n_2519),
.A2(n_2525),
.B(n_2532),
.C(n_2528),
.Y(n_2771)
);

AOI21xp5_ASAP7_75t_L g2772 ( 
.A1(n_2355),
.A2(n_85),
.B(n_86),
.Y(n_2772)
);

AOI21xp5_ASAP7_75t_L g2773 ( 
.A1(n_2434),
.A2(n_87),
.B(n_88),
.Y(n_2773)
);

AOI21xp5_ASAP7_75t_L g2774 ( 
.A1(n_2343),
.A2(n_87),
.B(n_88),
.Y(n_2774)
);

HB1xp67_ASAP7_75t_L g2775 ( 
.A(n_2322),
.Y(n_2775)
);

NAND2xp5_ASAP7_75t_L g2776 ( 
.A(n_2388),
.B(n_88),
.Y(n_2776)
);

CKINVDCx6p67_ASAP7_75t_R g2777 ( 
.A(n_2369),
.Y(n_2777)
);

BUFx4f_ASAP7_75t_L g2778 ( 
.A(n_2287),
.Y(n_2778)
);

AOI21xp5_ASAP7_75t_L g2779 ( 
.A1(n_2364),
.A2(n_89),
.B(n_90),
.Y(n_2779)
);

NOR2xp33_ASAP7_75t_L g2780 ( 
.A(n_2484),
.B(n_89),
.Y(n_2780)
);

AOI21xp5_ASAP7_75t_L g2781 ( 
.A1(n_2373),
.A2(n_90),
.B(n_91),
.Y(n_2781)
);

OAI321xp33_ASAP7_75t_L g2782 ( 
.A1(n_2425),
.A2(n_92),
.A3(n_94),
.B1(n_90),
.B2(n_91),
.C(n_93),
.Y(n_2782)
);

AOI21xp5_ASAP7_75t_L g2783 ( 
.A1(n_2398),
.A2(n_91),
.B(n_92),
.Y(n_2783)
);

INVx1_ASAP7_75t_L g2784 ( 
.A(n_2435),
.Y(n_2784)
);

A2O1A1Ixp33_ASAP7_75t_L g2785 ( 
.A1(n_2190),
.A2(n_95),
.B(n_93),
.C(n_94),
.Y(n_2785)
);

OAI21xp5_ASAP7_75t_L g2786 ( 
.A1(n_2436),
.A2(n_93),
.B(n_94),
.Y(n_2786)
);

NAND2xp5_ASAP7_75t_L g2787 ( 
.A(n_2372),
.B(n_95),
.Y(n_2787)
);

AOI21xp5_ASAP7_75t_L g2788 ( 
.A1(n_2401),
.A2(n_95),
.B(n_96),
.Y(n_2788)
);

XOR2x2_ASAP7_75t_L g2789 ( 
.A(n_2265),
.B(n_96),
.Y(n_2789)
);

NAND2xp5_ASAP7_75t_L g2790 ( 
.A(n_2288),
.B(n_96),
.Y(n_2790)
);

AOI21xp5_ASAP7_75t_L g2791 ( 
.A1(n_2402),
.A2(n_97),
.B(n_98),
.Y(n_2791)
);

NOR3xp33_ASAP7_75t_L g2792 ( 
.A(n_2206),
.B(n_99),
.C(n_98),
.Y(n_2792)
);

INVx1_ASAP7_75t_SL g2793 ( 
.A(n_2187),
.Y(n_2793)
);

NOR3xp33_ASAP7_75t_L g2794 ( 
.A(n_2293),
.B(n_2216),
.C(n_2513),
.Y(n_2794)
);

A2O1A1Ixp33_ASAP7_75t_L g2795 ( 
.A1(n_2176),
.A2(n_100),
.B(n_97),
.C(n_99),
.Y(n_2795)
);

NAND2xp5_ASAP7_75t_L g2796 ( 
.A(n_2325),
.B(n_99),
.Y(n_2796)
);

AOI21xp5_ASAP7_75t_L g2797 ( 
.A1(n_2403),
.A2(n_100),
.B(n_101),
.Y(n_2797)
);

AOI21xp5_ASAP7_75t_L g2798 ( 
.A1(n_2376),
.A2(n_100),
.B(n_101),
.Y(n_2798)
);

AND2x2_ASAP7_75t_SL g2799 ( 
.A(n_2352),
.B(n_101),
.Y(n_2799)
);

AOI21xp5_ASAP7_75t_L g2800 ( 
.A1(n_2294),
.A2(n_102),
.B(n_103),
.Y(n_2800)
);

NAND2xp5_ASAP7_75t_SL g2801 ( 
.A(n_2486),
.B(n_103),
.Y(n_2801)
);

BUFx8_ASAP7_75t_L g2802 ( 
.A(n_2319),
.Y(n_2802)
);

NOR2xp33_ASAP7_75t_L g2803 ( 
.A(n_2515),
.B(n_102),
.Y(n_2803)
);

BUFx6f_ASAP7_75t_L g2804 ( 
.A(n_2273),
.Y(n_2804)
);

AOI21xp5_ASAP7_75t_L g2805 ( 
.A1(n_2451),
.A2(n_102),
.B(n_104),
.Y(n_2805)
);

NAND2xp5_ASAP7_75t_L g2806 ( 
.A(n_2325),
.B(n_105),
.Y(n_2806)
);

NOR2xp33_ASAP7_75t_R g2807 ( 
.A(n_2350),
.B(n_105),
.Y(n_2807)
);

NAND2xp5_ASAP7_75t_L g2808 ( 
.A(n_2508),
.B(n_106),
.Y(n_2808)
);

AOI21xp5_ASAP7_75t_L g2809 ( 
.A1(n_2452),
.A2(n_2456),
.B(n_2453),
.Y(n_2809)
);

NAND2xp5_ASAP7_75t_L g2810 ( 
.A(n_2522),
.B(n_106),
.Y(n_2810)
);

NOR2xp33_ASAP7_75t_L g2811 ( 
.A(n_2524),
.B(n_107),
.Y(n_2811)
);

OAI22xp5_ASAP7_75t_L g2812 ( 
.A1(n_2389),
.A2(n_109),
.B1(n_107),
.B2(n_108),
.Y(n_2812)
);

INVx1_ASAP7_75t_L g2813 ( 
.A(n_2317),
.Y(n_2813)
);

NAND2xp5_ASAP7_75t_L g2814 ( 
.A(n_2317),
.B(n_107),
.Y(n_2814)
);

AOI21xp5_ASAP7_75t_L g2815 ( 
.A1(n_2467),
.A2(n_109),
.B(n_110),
.Y(n_2815)
);

AOI21xp5_ASAP7_75t_L g2816 ( 
.A1(n_2444),
.A2(n_109),
.B(n_110),
.Y(n_2816)
);

NAND2xp5_ASAP7_75t_SL g2817 ( 
.A(n_2361),
.B(n_111),
.Y(n_2817)
);

OAI22xp5_ASAP7_75t_L g2818 ( 
.A1(n_2333),
.A2(n_112),
.B1(n_110),
.B2(n_111),
.Y(n_2818)
);

AOI21xp5_ASAP7_75t_L g2819 ( 
.A1(n_2222),
.A2(n_2362),
.B(n_2415),
.Y(n_2819)
);

NAND2xp5_ASAP7_75t_L g2820 ( 
.A(n_2394),
.B(n_111),
.Y(n_2820)
);

BUFx6f_ASAP7_75t_L g2821 ( 
.A(n_2273),
.Y(n_2821)
);

BUFx6f_ASAP7_75t_L g2822 ( 
.A(n_2273),
.Y(n_2822)
);

AOI21xp5_ASAP7_75t_L g2823 ( 
.A1(n_2429),
.A2(n_112),
.B(n_113),
.Y(n_2823)
);

INVx5_ASAP7_75t_L g2824 ( 
.A(n_2227),
.Y(n_2824)
);

NAND2xp5_ASAP7_75t_SL g2825 ( 
.A(n_2440),
.B(n_114),
.Y(n_2825)
);

AOI22xp5_ASAP7_75t_L g2826 ( 
.A1(n_2363),
.A2(n_115),
.B1(n_113),
.B2(n_114),
.Y(n_2826)
);

INVx1_ASAP7_75t_L g2827 ( 
.A(n_2400),
.Y(n_2827)
);

NOR2xp33_ASAP7_75t_L g2828 ( 
.A(n_2374),
.B(n_113),
.Y(n_2828)
);

NAND2xp5_ASAP7_75t_L g2829 ( 
.A(n_2366),
.B(n_114),
.Y(n_2829)
);

NOR2x1_ASAP7_75t_R g2830 ( 
.A(n_2414),
.B(n_115),
.Y(n_2830)
);

AND2x2_ASAP7_75t_L g2831 ( 
.A(n_2378),
.B(n_115),
.Y(n_2831)
);

INVx2_ASAP7_75t_L g2832 ( 
.A(n_2473),
.Y(n_2832)
);

BUFx12f_ASAP7_75t_L g2833 ( 
.A(n_2219),
.Y(n_2833)
);

NAND2xp5_ASAP7_75t_L g2834 ( 
.A(n_2383),
.B(n_116),
.Y(n_2834)
);

NAND2xp5_ASAP7_75t_SL g2835 ( 
.A(n_2359),
.B(n_117),
.Y(n_2835)
);

AOI21xp33_ASAP7_75t_L g2836 ( 
.A1(n_2365),
.A2(n_116),
.B(n_117),
.Y(n_2836)
);

INVx1_ASAP7_75t_L g2837 ( 
.A(n_2400),
.Y(n_2837)
);

INVx1_ASAP7_75t_L g2838 ( 
.A(n_2470),
.Y(n_2838)
);

AOI21xp5_ASAP7_75t_L g2839 ( 
.A1(n_2477),
.A2(n_116),
.B(n_117),
.Y(n_2839)
);

AOI21xp5_ASAP7_75t_L g2840 ( 
.A1(n_2353),
.A2(n_118),
.B(n_119),
.Y(n_2840)
);

NOR2x1p5_ASAP7_75t_L g2841 ( 
.A(n_2428),
.B(n_2266),
.Y(n_2841)
);

NAND2xp5_ASAP7_75t_L g2842 ( 
.A(n_2382),
.B(n_118),
.Y(n_2842)
);

HB1xp67_ASAP7_75t_L g2843 ( 
.A(n_2423),
.Y(n_2843)
);

AND2x2_ASAP7_75t_L g2844 ( 
.A(n_2441),
.B(n_118),
.Y(n_2844)
);

NAND2xp5_ASAP7_75t_SL g2845 ( 
.A(n_2390),
.B(n_120),
.Y(n_2845)
);

INVx1_ASAP7_75t_L g2846 ( 
.A(n_2471),
.Y(n_2846)
);

NOR2xp33_ASAP7_75t_L g2847 ( 
.A(n_2332),
.B(n_2272),
.Y(n_2847)
);

AOI21xp5_ASAP7_75t_L g2848 ( 
.A1(n_2419),
.A2(n_119),
.B(n_120),
.Y(n_2848)
);

AOI22xp5_ASAP7_75t_L g2849 ( 
.A1(n_2368),
.A2(n_122),
.B1(n_119),
.B2(n_121),
.Y(n_2849)
);

NAND2xp5_ASAP7_75t_L g2850 ( 
.A(n_2379),
.B(n_121),
.Y(n_2850)
);

NAND2xp5_ASAP7_75t_L g2851 ( 
.A(n_2227),
.B(n_121),
.Y(n_2851)
);

NOR2xp67_ASAP7_75t_L g2852 ( 
.A(n_2370),
.B(n_123),
.Y(n_2852)
);

INVx3_ASAP7_75t_L g2853 ( 
.A(n_2333),
.Y(n_2853)
);

NAND2xp5_ASAP7_75t_SL g2854 ( 
.A(n_2342),
.B(n_124),
.Y(n_2854)
);

NOR2xp67_ASAP7_75t_L g2855 ( 
.A(n_2478),
.B(n_123),
.Y(n_2855)
);

OAI22xp5_ASAP7_75t_L g2856 ( 
.A1(n_2339),
.A2(n_125),
.B1(n_123),
.B2(n_124),
.Y(n_2856)
);

OAI22xp5_ASAP7_75t_L g2857 ( 
.A1(n_2339),
.A2(n_127),
.B1(n_125),
.B2(n_126),
.Y(n_2857)
);

INVx1_ASAP7_75t_L g2858 ( 
.A(n_2445),
.Y(n_2858)
);

AO21x1_ASAP7_75t_L g2859 ( 
.A1(n_2454),
.A2(n_712),
.B(n_710),
.Y(n_2859)
);

AND2x2_ASAP7_75t_L g2860 ( 
.A(n_2463),
.B(n_125),
.Y(n_2860)
);

O2A1O1Ixp33_ASAP7_75t_L g2861 ( 
.A1(n_2406),
.A2(n_128),
.B(n_126),
.C(n_127),
.Y(n_2861)
);

NAND2x1p5_ASAP7_75t_L g2862 ( 
.A(n_2342),
.B(n_126),
.Y(n_2862)
);

AOI21xp5_ASAP7_75t_L g2863 ( 
.A1(n_2472),
.A2(n_127),
.B(n_128),
.Y(n_2863)
);

AOI21xp5_ASAP7_75t_L g2864 ( 
.A1(n_2476),
.A2(n_129),
.B(n_131),
.Y(n_2864)
);

OAI21xp5_ASAP7_75t_L g2865 ( 
.A1(n_2422),
.A2(n_129),
.B(n_131),
.Y(n_2865)
);

AOI21xp5_ASAP7_75t_L g2866 ( 
.A1(n_2446),
.A2(n_129),
.B(n_131),
.Y(n_2866)
);

NOR2xp33_ASAP7_75t_R g2867 ( 
.A(n_2319),
.B(n_132),
.Y(n_2867)
);

AOI21xp5_ASAP7_75t_L g2868 ( 
.A1(n_2342),
.A2(n_132),
.B(n_133),
.Y(n_2868)
);

INVx3_ASAP7_75t_L g2869 ( 
.A(n_2423),
.Y(n_2869)
);

OR2x6_ASAP7_75t_L g2870 ( 
.A(n_2338),
.B(n_132),
.Y(n_2870)
);

INVx1_ASAP7_75t_L g2871 ( 
.A(n_2459),
.Y(n_2871)
);

NAND2xp5_ASAP7_75t_L g2872 ( 
.A(n_2227),
.B(n_133),
.Y(n_2872)
);

NOR2xp33_ASAP7_75t_L g2873 ( 
.A(n_2458),
.B(n_133),
.Y(n_2873)
);

A2O1A1Ixp33_ASAP7_75t_L g2874 ( 
.A1(n_2460),
.A2(n_136),
.B(n_134),
.C(n_135),
.Y(n_2874)
);

A2O1A1Ixp33_ASAP7_75t_L g2875 ( 
.A1(n_2174),
.A2(n_136),
.B(n_134),
.C(n_135),
.Y(n_2875)
);

AOI21xp5_ASAP7_75t_L g2876 ( 
.A1(n_2412),
.A2(n_134),
.B(n_135),
.Y(n_2876)
);

AOI22xp5_ASAP7_75t_L g2877 ( 
.A1(n_2227),
.A2(n_139),
.B1(n_137),
.B2(n_138),
.Y(n_2877)
);

NAND2xp5_ASAP7_75t_SL g2878 ( 
.A(n_2474),
.B(n_138),
.Y(n_2878)
);

AOI21xp5_ASAP7_75t_L g2879 ( 
.A1(n_2421),
.A2(n_137),
.B(n_138),
.Y(n_2879)
);

NAND2xp5_ASAP7_75t_L g2880 ( 
.A(n_2290),
.B(n_137),
.Y(n_2880)
);

AND2x2_ASAP7_75t_L g2881 ( 
.A(n_2405),
.B(n_139),
.Y(n_2881)
);

INVx8_ASAP7_75t_L g2882 ( 
.A(n_2430),
.Y(n_2882)
);

INVx2_ASAP7_75t_L g2883 ( 
.A(n_2386),
.Y(n_2883)
);

CKINVDCx20_ASAP7_75t_R g2884 ( 
.A(n_2479),
.Y(n_2884)
);

BUFx6f_ASAP7_75t_L g2885 ( 
.A(n_2433),
.Y(n_2885)
);

CKINVDCx10_ASAP7_75t_R g2886 ( 
.A(n_2480),
.Y(n_2886)
);

INVx1_ASAP7_75t_L g2887 ( 
.A(n_2426),
.Y(n_2887)
);

AOI21xp5_ASAP7_75t_L g2888 ( 
.A1(n_2424),
.A2(n_139),
.B(n_140),
.Y(n_2888)
);

NAND2xp5_ASAP7_75t_L g2889 ( 
.A(n_2427),
.B(n_140),
.Y(n_2889)
);

INVxp67_ASAP7_75t_L g2890 ( 
.A(n_2432),
.Y(n_2890)
);

INVx1_ASAP7_75t_L g2891 ( 
.A(n_2448),
.Y(n_2891)
);

BUFx3_ASAP7_75t_L g2892 ( 
.A(n_2408),
.Y(n_2892)
);

NOR2xp33_ASAP7_75t_L g2893 ( 
.A(n_2455),
.B(n_140),
.Y(n_2893)
);

AOI21xp33_ASAP7_75t_L g2894 ( 
.A1(n_2465),
.A2(n_141),
.B(n_142),
.Y(n_2894)
);

INVx1_ASAP7_75t_L g2895 ( 
.A(n_2468),
.Y(n_2895)
);

A2O1A1Ixp33_ASAP7_75t_L g2896 ( 
.A1(n_2439),
.A2(n_143),
.B(n_141),
.C(n_142),
.Y(n_2896)
);

NAND2xp5_ASAP7_75t_L g2897 ( 
.A(n_2475),
.B(n_142),
.Y(n_2897)
);

INVx1_ASAP7_75t_L g2898 ( 
.A(n_2442),
.Y(n_2898)
);

NOR2x1p5_ASAP7_75t_L g2899 ( 
.A(n_2464),
.B(n_143),
.Y(n_2899)
);

NAND2xp5_ASAP7_75t_L g2900 ( 
.A(n_2264),
.B(n_143),
.Y(n_2900)
);

AND2x2_ASAP7_75t_L g2901 ( 
.A(n_2210),
.B(n_144),
.Y(n_2901)
);

A2O1A1Ixp33_ASAP7_75t_L g2902 ( 
.A1(n_2248),
.A2(n_146),
.B(n_144),
.C(n_145),
.Y(n_2902)
);

OAI21xp5_ASAP7_75t_L g2903 ( 
.A1(n_2182),
.A2(n_144),
.B(n_145),
.Y(n_2903)
);

NAND2xp5_ASAP7_75t_L g2904 ( 
.A(n_2264),
.B(n_145),
.Y(n_2904)
);

NAND2xp5_ASAP7_75t_L g2905 ( 
.A(n_2264),
.B(n_146),
.Y(n_2905)
);

NAND2xp5_ASAP7_75t_L g2906 ( 
.A(n_2264),
.B(n_147),
.Y(n_2906)
);

NAND2xp5_ASAP7_75t_L g2907 ( 
.A(n_2264),
.B(n_147),
.Y(n_2907)
);

AND2x2_ASAP7_75t_L g2908 ( 
.A(n_2210),
.B(n_147),
.Y(n_2908)
);

INVx3_ASAP7_75t_L g2909 ( 
.A(n_2231),
.Y(n_2909)
);

AOI21xp33_ASAP7_75t_L g2910 ( 
.A1(n_2221),
.A2(n_148),
.B(n_149),
.Y(n_2910)
);

NAND2xp5_ASAP7_75t_SL g2911 ( 
.A(n_2262),
.B(n_149),
.Y(n_2911)
);

INVx1_ASAP7_75t_L g2912 ( 
.A(n_2205),
.Y(n_2912)
);

NAND2xp5_ASAP7_75t_L g2913 ( 
.A(n_2264),
.B(n_148),
.Y(n_2913)
);

INVx1_ASAP7_75t_L g2914 ( 
.A(n_2205),
.Y(n_2914)
);

NAND2xp5_ASAP7_75t_L g2915 ( 
.A(n_2264),
.B(n_148),
.Y(n_2915)
);

AOI21xp5_ASAP7_75t_L g2916 ( 
.A1(n_2450),
.A2(n_149),
.B(n_150),
.Y(n_2916)
);

AOI21xp5_ASAP7_75t_L g2917 ( 
.A1(n_2450),
.A2(n_150),
.B(n_151),
.Y(n_2917)
);

NAND2xp5_ASAP7_75t_SL g2918 ( 
.A(n_2262),
.B(n_152),
.Y(n_2918)
);

AOI21xp5_ASAP7_75t_L g2919 ( 
.A1(n_2450),
.A2(n_151),
.B(n_152),
.Y(n_2919)
);

OAI321xp33_ASAP7_75t_L g2920 ( 
.A1(n_2341),
.A2(n_155),
.A3(n_157),
.B1(n_153),
.B2(n_154),
.C(n_156),
.Y(n_2920)
);

AOI21xp5_ASAP7_75t_L g2921 ( 
.A1(n_2450),
.A2(n_153),
.B(n_154),
.Y(n_2921)
);

AND2x4_ASAP7_75t_L g2922 ( 
.A(n_2231),
.B(n_153),
.Y(n_2922)
);

OR2x2_ASAP7_75t_L g2923 ( 
.A(n_2215),
.B(n_154),
.Y(n_2923)
);

BUFx4f_ASAP7_75t_L g2924 ( 
.A(n_2281),
.Y(n_2924)
);

A2O1A1Ixp33_ASAP7_75t_L g2925 ( 
.A1(n_2248),
.A2(n_157),
.B(n_155),
.C(n_156),
.Y(n_2925)
);

BUFx3_ASAP7_75t_L g2926 ( 
.A(n_2281),
.Y(n_2926)
);

A2O1A1Ixp33_ASAP7_75t_L g2927 ( 
.A1(n_2248),
.A2(n_159),
.B(n_157),
.C(n_158),
.Y(n_2927)
);

NAND2xp5_ASAP7_75t_L g2928 ( 
.A(n_2264),
.B(n_158),
.Y(n_2928)
);

AND2x4_ASAP7_75t_L g2929 ( 
.A(n_2231),
.B(n_160),
.Y(n_2929)
);

AOI21x1_ASAP7_75t_L g2930 ( 
.A1(n_2461),
.A2(n_160),
.B(n_161),
.Y(n_2930)
);

NAND2xp5_ASAP7_75t_L g2931 ( 
.A(n_2264),
.B(n_160),
.Y(n_2931)
);

BUFx3_ASAP7_75t_L g2932 ( 
.A(n_2281),
.Y(n_2932)
);

NAND2xp5_ASAP7_75t_L g2933 ( 
.A(n_2264),
.B(n_161),
.Y(n_2933)
);

NAND2xp5_ASAP7_75t_L g2934 ( 
.A(n_2264),
.B(n_162),
.Y(n_2934)
);

INVx1_ASAP7_75t_L g2935 ( 
.A(n_2205),
.Y(n_2935)
);

INVx2_ASAP7_75t_L g2936 ( 
.A(n_2254),
.Y(n_2936)
);

AOI21xp5_ASAP7_75t_L g2937 ( 
.A1(n_2450),
.A2(n_162),
.B(n_163),
.Y(n_2937)
);

NOR2x1_ASAP7_75t_L g2938 ( 
.A(n_2330),
.B(n_162),
.Y(n_2938)
);

BUFx3_ASAP7_75t_L g2939 ( 
.A(n_2281),
.Y(n_2939)
);

INVx1_ASAP7_75t_L g2940 ( 
.A(n_2205),
.Y(n_2940)
);

NAND2xp5_ASAP7_75t_L g2941 ( 
.A(n_2264),
.B(n_163),
.Y(n_2941)
);

AND2x2_ASAP7_75t_L g2942 ( 
.A(n_2210),
.B(n_163),
.Y(n_2942)
);

AO21x1_ASAP7_75t_L g2943 ( 
.A1(n_2461),
.A2(n_712),
.B(n_710),
.Y(n_2943)
);

NAND2xp5_ASAP7_75t_L g2944 ( 
.A(n_2264),
.B(n_164),
.Y(n_2944)
);

INVxp67_ASAP7_75t_L g2945 ( 
.A(n_2526),
.Y(n_2945)
);

AOI21xp5_ASAP7_75t_L g2946 ( 
.A1(n_2450),
.A2(n_164),
.B(n_165),
.Y(n_2946)
);

O2A1O1Ixp33_ASAP7_75t_L g2947 ( 
.A1(n_2248),
.A2(n_166),
.B(n_164),
.C(n_165),
.Y(n_2947)
);

AND2x2_ASAP7_75t_L g2948 ( 
.A(n_2210),
.B(n_166),
.Y(n_2948)
);

INVx1_ASAP7_75t_SL g2949 ( 
.A(n_2526),
.Y(n_2949)
);

NAND2xp5_ASAP7_75t_SL g2950 ( 
.A(n_2262),
.B(n_168),
.Y(n_2950)
);

AOI21xp5_ASAP7_75t_L g2951 ( 
.A1(n_2450),
.A2(n_167),
.B(n_168),
.Y(n_2951)
);

INVx1_ASAP7_75t_L g2952 ( 
.A(n_2205),
.Y(n_2952)
);

AOI21xp5_ASAP7_75t_L g2953 ( 
.A1(n_2450),
.A2(n_167),
.B(n_169),
.Y(n_2953)
);

BUFx6f_ASAP7_75t_L g2954 ( 
.A(n_2233),
.Y(n_2954)
);

INVx3_ASAP7_75t_L g2955 ( 
.A(n_2231),
.Y(n_2955)
);

A2O1A1Ixp33_ASAP7_75t_L g2956 ( 
.A1(n_2248),
.A2(n_170),
.B(n_167),
.C(n_169),
.Y(n_2956)
);

INVx1_ASAP7_75t_L g2957 ( 
.A(n_2205),
.Y(n_2957)
);

INVx1_ASAP7_75t_L g2958 ( 
.A(n_2205),
.Y(n_2958)
);

A2O1A1Ixp33_ASAP7_75t_L g2959 ( 
.A1(n_2248),
.A2(n_172),
.B(n_170),
.C(n_171),
.Y(n_2959)
);

NAND2xp5_ASAP7_75t_L g2960 ( 
.A(n_2264),
.B(n_170),
.Y(n_2960)
);

OAI21xp5_ASAP7_75t_L g2961 ( 
.A1(n_2182),
.A2(n_172),
.B(n_173),
.Y(n_2961)
);

AOI21xp5_ASAP7_75t_L g2962 ( 
.A1(n_2450),
.A2(n_172),
.B(n_173),
.Y(n_2962)
);

A2O1A1Ixp33_ASAP7_75t_L g2963 ( 
.A1(n_2248),
.A2(n_176),
.B(n_174),
.C(n_175),
.Y(n_2963)
);

NAND2xp5_ASAP7_75t_L g2964 ( 
.A(n_2264),
.B(n_174),
.Y(n_2964)
);

O2A1O1Ixp33_ASAP7_75t_L g2965 ( 
.A1(n_2248),
.A2(n_176),
.B(n_174),
.C(n_175),
.Y(n_2965)
);

AOI21xp5_ASAP7_75t_L g2966 ( 
.A1(n_2450),
.A2(n_175),
.B(n_177),
.Y(n_2966)
);

AOI21xp5_ASAP7_75t_L g2967 ( 
.A1(n_2450),
.A2(n_177),
.B(n_178),
.Y(n_2967)
);

BUFx3_ASAP7_75t_L g2968 ( 
.A(n_2281),
.Y(n_2968)
);

OAI21xp5_ASAP7_75t_L g2969 ( 
.A1(n_2182),
.A2(n_177),
.B(n_178),
.Y(n_2969)
);

HB1xp67_ASAP7_75t_L g2970 ( 
.A(n_2526),
.Y(n_2970)
);

NOR2xp33_ASAP7_75t_L g2971 ( 
.A(n_2229),
.B(n_178),
.Y(n_2971)
);

OAI21xp5_ASAP7_75t_L g2972 ( 
.A1(n_2182),
.A2(n_179),
.B(n_180),
.Y(n_2972)
);

AOI22xp5_ASAP7_75t_L g2973 ( 
.A1(n_2213),
.A2(n_181),
.B1(n_179),
.B2(n_180),
.Y(n_2973)
);

A2O1A1Ixp33_ASAP7_75t_L g2974 ( 
.A1(n_2248),
.A2(n_182),
.B(n_180),
.C(n_181),
.Y(n_2974)
);

O2A1O1Ixp33_ASAP7_75t_L g2975 ( 
.A1(n_2248),
.A2(n_184),
.B(n_182),
.C(n_183),
.Y(n_2975)
);

AOI22xp5_ASAP7_75t_L g2976 ( 
.A1(n_2213),
.A2(n_185),
.B1(n_183),
.B2(n_184),
.Y(n_2976)
);

NOR2xp33_ASAP7_75t_L g2977 ( 
.A(n_2229),
.B(n_184),
.Y(n_2977)
);

O2A1O1Ixp33_ASAP7_75t_L g2978 ( 
.A1(n_2248),
.A2(n_187),
.B(n_185),
.C(n_186),
.Y(n_2978)
);

INVx3_ASAP7_75t_L g2979 ( 
.A(n_2231),
.Y(n_2979)
);

NAND2xp5_ASAP7_75t_L g2980 ( 
.A(n_2264),
.B(n_185),
.Y(n_2980)
);

NAND2xp5_ASAP7_75t_L g2981 ( 
.A(n_2264),
.B(n_186),
.Y(n_2981)
);

INVx2_ASAP7_75t_L g2982 ( 
.A(n_2254),
.Y(n_2982)
);

NOR2xp33_ASAP7_75t_SL g2983 ( 
.A(n_2262),
.B(n_186),
.Y(n_2983)
);

NOR2xp33_ASAP7_75t_L g2984 ( 
.A(n_2229),
.B(n_187),
.Y(n_2984)
);

NAND2xp5_ASAP7_75t_L g2985 ( 
.A(n_2264),
.B(n_187),
.Y(n_2985)
);

OAI21xp5_ASAP7_75t_L g2986 ( 
.A1(n_2461),
.A2(n_188),
.B(n_189),
.Y(n_2986)
);

INVx1_ASAP7_75t_SL g2987 ( 
.A(n_2526),
.Y(n_2987)
);

INVx1_ASAP7_75t_L g2988 ( 
.A(n_2205),
.Y(n_2988)
);

INVx1_ASAP7_75t_L g2989 ( 
.A(n_2205),
.Y(n_2989)
);

OR2x2_ASAP7_75t_L g2990 ( 
.A(n_2215),
.B(n_188),
.Y(n_2990)
);

NOR2xp67_ASAP7_75t_L g2991 ( 
.A(n_2511),
.B(n_188),
.Y(n_2991)
);

AOI21xp5_ASAP7_75t_L g2992 ( 
.A1(n_2450),
.A2(n_189),
.B(n_190),
.Y(n_2992)
);

AOI21xp5_ASAP7_75t_L g2993 ( 
.A1(n_2450),
.A2(n_189),
.B(n_190),
.Y(n_2993)
);

NAND2xp5_ASAP7_75t_L g2994 ( 
.A(n_2264),
.B(n_190),
.Y(n_2994)
);

NAND3xp33_ASAP7_75t_SL g2995 ( 
.A(n_2213),
.B(n_191),
.C(n_192),
.Y(n_2995)
);

OAI21xp5_ASAP7_75t_L g2996 ( 
.A1(n_2182),
.A2(n_191),
.B(n_192),
.Y(n_2996)
);

NAND2xp5_ASAP7_75t_L g2997 ( 
.A(n_2264),
.B(n_193),
.Y(n_2997)
);

INVx1_ASAP7_75t_L g2998 ( 
.A(n_2205),
.Y(n_2998)
);

NAND2xp5_ASAP7_75t_L g2999 ( 
.A(n_2264),
.B(n_195),
.Y(n_2999)
);

BUFx3_ASAP7_75t_L g3000 ( 
.A(n_2281),
.Y(n_3000)
);

HB1xp67_ASAP7_75t_L g3001 ( 
.A(n_2526),
.Y(n_3001)
);

NAND2xp5_ASAP7_75t_L g3002 ( 
.A(n_2264),
.B(n_195),
.Y(n_3002)
);

A2O1A1Ixp33_ASAP7_75t_L g3003 ( 
.A1(n_2248),
.A2(n_198),
.B(n_196),
.C(n_197),
.Y(n_3003)
);

NAND2xp5_ASAP7_75t_L g3004 ( 
.A(n_2264),
.B(n_196),
.Y(n_3004)
);

HB1xp67_ASAP7_75t_L g3005 ( 
.A(n_2526),
.Y(n_3005)
);

NOR2xp33_ASAP7_75t_L g3006 ( 
.A(n_2229),
.B(n_198),
.Y(n_3006)
);

AOI21xp5_ASAP7_75t_L g3007 ( 
.A1(n_2450),
.A2(n_199),
.B(n_200),
.Y(n_3007)
);

OAI22xp5_ASAP7_75t_L g3008 ( 
.A1(n_2197),
.A2(n_201),
.B1(n_199),
.B2(n_200),
.Y(n_3008)
);

NAND2xp5_ASAP7_75t_L g3009 ( 
.A(n_2264),
.B(n_199),
.Y(n_3009)
);

OAI21xp5_ASAP7_75t_L g3010 ( 
.A1(n_2182),
.A2(n_201),
.B(n_202),
.Y(n_3010)
);

OAI21xp5_ASAP7_75t_L g3011 ( 
.A1(n_2182),
.A2(n_201),
.B(n_202),
.Y(n_3011)
);

OR2x2_ASAP7_75t_L g3012 ( 
.A(n_2215),
.B(n_203),
.Y(n_3012)
);

AOI21xp5_ASAP7_75t_L g3013 ( 
.A1(n_2450),
.A2(n_203),
.B(n_204),
.Y(n_3013)
);

AND2x4_ASAP7_75t_L g3014 ( 
.A(n_2231),
.B(n_203),
.Y(n_3014)
);

AOI22xp5_ASAP7_75t_L g3015 ( 
.A1(n_2213),
.A2(n_206),
.B1(n_204),
.B2(n_205),
.Y(n_3015)
);

BUFx6f_ASAP7_75t_L g3016 ( 
.A(n_2233),
.Y(n_3016)
);

CKINVDCx5p33_ASAP7_75t_R g3017 ( 
.A(n_2281),
.Y(n_3017)
);

AOI21x1_ASAP7_75t_L g3018 ( 
.A1(n_2461),
.A2(n_205),
.B(n_206),
.Y(n_3018)
);

INVx1_ASAP7_75t_L g3019 ( 
.A(n_2205),
.Y(n_3019)
);

NOR2xp33_ASAP7_75t_L g3020 ( 
.A(n_2229),
.B(n_206),
.Y(n_3020)
);

NAND2xp5_ASAP7_75t_L g3021 ( 
.A(n_2264),
.B(n_207),
.Y(n_3021)
);

O2A1O1Ixp33_ASAP7_75t_L g3022 ( 
.A1(n_2248),
.A2(n_209),
.B(n_207),
.C(n_208),
.Y(n_3022)
);

NOR2xp33_ASAP7_75t_L g3023 ( 
.A(n_2229),
.B(n_207),
.Y(n_3023)
);

O2A1O1Ixp33_ASAP7_75t_L g3024 ( 
.A1(n_2248),
.A2(n_210),
.B(n_208),
.C(n_209),
.Y(n_3024)
);

AOI21xp5_ASAP7_75t_L g3025 ( 
.A1(n_2450),
.A2(n_208),
.B(n_209),
.Y(n_3025)
);

AOI21xp5_ASAP7_75t_L g3026 ( 
.A1(n_2450),
.A2(n_210),
.B(n_211),
.Y(n_3026)
);

INVx4_ASAP7_75t_L g3027 ( 
.A(n_2281),
.Y(n_3027)
);

INVx2_ASAP7_75t_L g3028 ( 
.A(n_2254),
.Y(n_3028)
);

INVx1_ASAP7_75t_SL g3029 ( 
.A(n_2526),
.Y(n_3029)
);

AOI21xp5_ASAP7_75t_L g3030 ( 
.A1(n_2450),
.A2(n_211),
.B(n_212),
.Y(n_3030)
);

INVx1_ASAP7_75t_L g3031 ( 
.A(n_2205),
.Y(n_3031)
);

INVx2_ASAP7_75t_L g3032 ( 
.A(n_2254),
.Y(n_3032)
);

O2A1O1Ixp33_ASAP7_75t_L g3033 ( 
.A1(n_2248),
.A2(n_213),
.B(n_211),
.C(n_212),
.Y(n_3033)
);

INVx3_ASAP7_75t_L g3034 ( 
.A(n_2231),
.Y(n_3034)
);

O2A1O1Ixp33_ASAP7_75t_L g3035 ( 
.A1(n_2248),
.A2(n_214),
.B(n_212),
.C(n_213),
.Y(n_3035)
);

AOI21xp5_ASAP7_75t_L g3036 ( 
.A1(n_2450),
.A2(n_213),
.B(n_214),
.Y(n_3036)
);

NAND2xp5_ASAP7_75t_L g3037 ( 
.A(n_2264),
.B(n_215),
.Y(n_3037)
);

INVx1_ASAP7_75t_L g3038 ( 
.A(n_2205),
.Y(n_3038)
);

AOI21x1_ASAP7_75t_L g3039 ( 
.A1(n_2461),
.A2(n_215),
.B(n_216),
.Y(n_3039)
);

OAI22xp5_ASAP7_75t_L g3040 ( 
.A1(n_2197),
.A2(n_218),
.B1(n_215),
.B2(n_217),
.Y(n_3040)
);

AOI21xp5_ASAP7_75t_L g3041 ( 
.A1(n_2450),
.A2(n_218),
.B(n_219),
.Y(n_3041)
);

BUFx4f_ASAP7_75t_L g3042 ( 
.A(n_2281),
.Y(n_3042)
);

NAND2xp5_ASAP7_75t_L g3043 ( 
.A(n_2264),
.B(n_218),
.Y(n_3043)
);

AOI22xp5_ASAP7_75t_L g3044 ( 
.A1(n_2213),
.A2(n_221),
.B1(n_219),
.B2(n_220),
.Y(n_3044)
);

AOI21xp5_ASAP7_75t_L g3045 ( 
.A1(n_2450),
.A2(n_219),
.B(n_220),
.Y(n_3045)
);

AOI21xp5_ASAP7_75t_L g3046 ( 
.A1(n_2450),
.A2(n_220),
.B(n_221),
.Y(n_3046)
);

NAND2xp5_ASAP7_75t_L g3047 ( 
.A(n_2264),
.B(n_221),
.Y(n_3047)
);

AOI21xp5_ASAP7_75t_L g3048 ( 
.A1(n_2450),
.A2(n_222),
.B(n_223),
.Y(n_3048)
);

INVx2_ASAP7_75t_SL g3049 ( 
.A(n_2281),
.Y(n_3049)
);

INVx6_ASAP7_75t_L g3050 ( 
.A(n_2281),
.Y(n_3050)
);

OAI22xp5_ASAP7_75t_L g3051 ( 
.A1(n_2197),
.A2(n_224),
.B1(n_222),
.B2(n_223),
.Y(n_3051)
);

NAND2xp5_ASAP7_75t_L g3052 ( 
.A(n_2264),
.B(n_223),
.Y(n_3052)
);

AOI21xp5_ASAP7_75t_L g3053 ( 
.A1(n_2450),
.A2(n_224),
.B(n_225),
.Y(n_3053)
);

AOI21xp5_ASAP7_75t_L g3054 ( 
.A1(n_2450),
.A2(n_225),
.B(n_226),
.Y(n_3054)
);

NAND2xp5_ASAP7_75t_L g3055 ( 
.A(n_2264),
.B(n_226),
.Y(n_3055)
);

BUFx8_ASAP7_75t_SL g3056 ( 
.A(n_2239),
.Y(n_3056)
);

NAND2xp5_ASAP7_75t_SL g3057 ( 
.A(n_2262),
.B(n_228),
.Y(n_3057)
);

INVx2_ASAP7_75t_L g3058 ( 
.A(n_2254),
.Y(n_3058)
);

BUFx2_ASAP7_75t_L g3059 ( 
.A(n_2526),
.Y(n_3059)
);

NOR2xp33_ASAP7_75t_L g3060 ( 
.A(n_2229),
.B(n_227),
.Y(n_3060)
);

OAI21xp5_ASAP7_75t_L g3061 ( 
.A1(n_2182),
.A2(n_227),
.B(n_228),
.Y(n_3061)
);

INVx2_ASAP7_75t_L g3062 ( 
.A(n_2254),
.Y(n_3062)
);

O2A1O1Ixp33_ASAP7_75t_L g3063 ( 
.A1(n_2248),
.A2(n_230),
.B(n_227),
.C(n_229),
.Y(n_3063)
);

NAND2xp5_ASAP7_75t_L g3064 ( 
.A(n_2264),
.B(n_229),
.Y(n_3064)
);

AND2x4_ASAP7_75t_L g3065 ( 
.A(n_2231),
.B(n_231),
.Y(n_3065)
);

BUFx6f_ASAP7_75t_L g3066 ( 
.A(n_2233),
.Y(n_3066)
);

INVx1_ASAP7_75t_L g3067 ( 
.A(n_2205),
.Y(n_3067)
);

NOR2xp33_ASAP7_75t_L g3068 ( 
.A(n_2229),
.B(n_231),
.Y(n_3068)
);

NAND2xp5_ASAP7_75t_SL g3069 ( 
.A(n_2262),
.B(n_233),
.Y(n_3069)
);

INVx1_ASAP7_75t_L g3070 ( 
.A(n_2205),
.Y(n_3070)
);

NOR2x1_ASAP7_75t_L g3071 ( 
.A(n_2330),
.B(n_232),
.Y(n_3071)
);

AOI21xp5_ASAP7_75t_L g3072 ( 
.A1(n_2450),
.A2(n_232),
.B(n_233),
.Y(n_3072)
);

NAND2xp5_ASAP7_75t_L g3073 ( 
.A(n_2264),
.B(n_232),
.Y(n_3073)
);

AND2x2_ASAP7_75t_L g3074 ( 
.A(n_2210),
.B(n_234),
.Y(n_3074)
);

INVx1_ASAP7_75t_L g3075 ( 
.A(n_2205),
.Y(n_3075)
);

AOI21xp5_ASAP7_75t_L g3076 ( 
.A1(n_2450),
.A2(n_234),
.B(n_235),
.Y(n_3076)
);

OAI22xp5_ASAP7_75t_L g3077 ( 
.A1(n_2197),
.A2(n_237),
.B1(n_235),
.B2(n_236),
.Y(n_3077)
);

INVx2_ASAP7_75t_L g3078 ( 
.A(n_2254),
.Y(n_3078)
);

INVx3_ASAP7_75t_L g3079 ( 
.A(n_2231),
.Y(n_3079)
);

NAND2xp5_ASAP7_75t_L g3080 ( 
.A(n_2264),
.B(n_235),
.Y(n_3080)
);

AOI22xp5_ASAP7_75t_L g3081 ( 
.A1(n_2213),
.A2(n_238),
.B1(n_236),
.B2(n_237),
.Y(n_3081)
);

NAND2xp5_ASAP7_75t_L g3082 ( 
.A(n_2264),
.B(n_236),
.Y(n_3082)
);

NAND2xp5_ASAP7_75t_L g3083 ( 
.A(n_2264),
.B(n_237),
.Y(n_3083)
);

INVx2_ASAP7_75t_L g3084 ( 
.A(n_2254),
.Y(n_3084)
);

OAI21xp5_ASAP7_75t_L g3085 ( 
.A1(n_2182),
.A2(n_238),
.B(n_239),
.Y(n_3085)
);

AND2x2_ASAP7_75t_SL g3086 ( 
.A(n_2213),
.B(n_238),
.Y(n_3086)
);

CKINVDCx5p33_ASAP7_75t_R g3087 ( 
.A(n_2281),
.Y(n_3087)
);

O2A1O1Ixp5_ASAP7_75t_L g3088 ( 
.A1(n_2341),
.A2(n_242),
.B(n_240),
.C(n_241),
.Y(n_3088)
);

OAI21xp5_ASAP7_75t_L g3089 ( 
.A1(n_2182),
.A2(n_240),
.B(n_241),
.Y(n_3089)
);

NOR2xp33_ASAP7_75t_L g3090 ( 
.A(n_2229),
.B(n_240),
.Y(n_3090)
);

AOI21xp5_ASAP7_75t_L g3091 ( 
.A1(n_2450),
.A2(n_241),
.B(n_242),
.Y(n_3091)
);

AOI21xp5_ASAP7_75t_L g3092 ( 
.A1(n_2450),
.A2(n_243),
.B(n_244),
.Y(n_3092)
);

AOI21xp5_ASAP7_75t_L g3093 ( 
.A1(n_2450),
.A2(n_243),
.B(n_244),
.Y(n_3093)
);

AOI21xp5_ASAP7_75t_L g3094 ( 
.A1(n_2450),
.A2(n_243),
.B(n_244),
.Y(n_3094)
);

AOI21xp5_ASAP7_75t_L g3095 ( 
.A1(n_2450),
.A2(n_245),
.B(n_246),
.Y(n_3095)
);

INVx2_ASAP7_75t_L g3096 ( 
.A(n_2254),
.Y(n_3096)
);

O2A1O1Ixp33_ASAP7_75t_L g3097 ( 
.A1(n_2248),
.A2(n_247),
.B(n_245),
.C(n_246),
.Y(n_3097)
);

OAI22xp5_ASAP7_75t_L g3098 ( 
.A1(n_2197),
.A2(n_248),
.B1(n_245),
.B2(n_247),
.Y(n_3098)
);

AOI21xp5_ASAP7_75t_L g3099 ( 
.A1(n_2450),
.A2(n_248),
.B(n_249),
.Y(n_3099)
);

NAND2xp5_ASAP7_75t_L g3100 ( 
.A(n_2264),
.B(n_251),
.Y(n_3100)
);

AOI33xp33_ASAP7_75t_L g3101 ( 
.A1(n_2503),
.A2(n_253),
.A3(n_255),
.B1(n_251),
.B2(n_252),
.B3(n_254),
.Y(n_3101)
);

OAI22xp5_ASAP7_75t_L g3102 ( 
.A1(n_2197),
.A2(n_253),
.B1(n_251),
.B2(n_252),
.Y(n_3102)
);

NAND2xp5_ASAP7_75t_SL g3103 ( 
.A(n_2262),
.B(n_255),
.Y(n_3103)
);

AOI21xp5_ASAP7_75t_L g3104 ( 
.A1(n_2450),
.A2(n_254),
.B(n_255),
.Y(n_3104)
);

AOI21xp5_ASAP7_75t_L g3105 ( 
.A1(n_2450),
.A2(n_256),
.B(n_257),
.Y(n_3105)
);

NAND2xp5_ASAP7_75t_L g3106 ( 
.A(n_2264),
.B(n_256),
.Y(n_3106)
);

OAI21xp5_ASAP7_75t_L g3107 ( 
.A1(n_2461),
.A2(n_256),
.B(n_257),
.Y(n_3107)
);

AOI21xp5_ASAP7_75t_L g3108 ( 
.A1(n_2450),
.A2(n_257),
.B(n_258),
.Y(n_3108)
);

NOR2x1_ASAP7_75t_SL g3109 ( 
.A(n_2239),
.B(n_259),
.Y(n_3109)
);

AND2x2_ASAP7_75t_L g3110 ( 
.A(n_2210),
.B(n_258),
.Y(n_3110)
);

OAI21xp5_ASAP7_75t_L g3111 ( 
.A1(n_2461),
.A2(n_259),
.B(n_260),
.Y(n_3111)
);

CKINVDCx5p33_ASAP7_75t_R g3112 ( 
.A(n_2281),
.Y(n_3112)
);

AOI21xp5_ASAP7_75t_L g3113 ( 
.A1(n_2450),
.A2(n_260),
.B(n_261),
.Y(n_3113)
);

AOI21xp5_ASAP7_75t_L g3114 ( 
.A1(n_2450),
.A2(n_260),
.B(n_261),
.Y(n_3114)
);

OAI21xp5_ASAP7_75t_L g3115 ( 
.A1(n_2461),
.A2(n_261),
.B(n_262),
.Y(n_3115)
);

BUFx6f_ASAP7_75t_L g3116 ( 
.A(n_2233),
.Y(n_3116)
);

INVx1_ASAP7_75t_L g3117 ( 
.A(n_2205),
.Y(n_3117)
);

NAND2xp5_ASAP7_75t_L g3118 ( 
.A(n_2264),
.B(n_262),
.Y(n_3118)
);

INVxp67_ASAP7_75t_L g3119 ( 
.A(n_2526),
.Y(n_3119)
);

NAND2xp5_ASAP7_75t_L g3120 ( 
.A(n_2264),
.B(n_263),
.Y(n_3120)
);

OAI21xp5_ASAP7_75t_L g3121 ( 
.A1(n_2461),
.A2(n_263),
.B(n_264),
.Y(n_3121)
);

AO21x1_ASAP7_75t_L g3122 ( 
.A1(n_2461),
.A2(n_714),
.B(n_713),
.Y(n_3122)
);

AND2x4_ASAP7_75t_L g3123 ( 
.A(n_2231),
.B(n_264),
.Y(n_3123)
);

BUFx2_ASAP7_75t_L g3124 ( 
.A(n_2526),
.Y(n_3124)
);

NAND2xp5_ASAP7_75t_L g3125 ( 
.A(n_2264),
.B(n_264),
.Y(n_3125)
);

OAI21xp5_ASAP7_75t_L g3126 ( 
.A1(n_2461),
.A2(n_265),
.B(n_266),
.Y(n_3126)
);

AOI21xp5_ASAP7_75t_L g3127 ( 
.A1(n_2450),
.A2(n_265),
.B(n_266),
.Y(n_3127)
);

AOI21xp5_ASAP7_75t_L g3128 ( 
.A1(n_2450),
.A2(n_267),
.B(n_268),
.Y(n_3128)
);

AOI22xp33_ASAP7_75t_L g3129 ( 
.A1(n_2212),
.A2(n_269),
.B1(n_267),
.B2(n_268),
.Y(n_3129)
);

AND2x2_ASAP7_75t_L g3130 ( 
.A(n_2210),
.B(n_267),
.Y(n_3130)
);

AOI21xp5_ASAP7_75t_L g3131 ( 
.A1(n_2450),
.A2(n_268),
.B(n_269),
.Y(n_3131)
);

HB1xp67_ASAP7_75t_L g3132 ( 
.A(n_2526),
.Y(n_3132)
);

AND2x4_ASAP7_75t_L g3133 ( 
.A(n_2231),
.B(n_270),
.Y(n_3133)
);

NAND2xp5_ASAP7_75t_L g3134 ( 
.A(n_2264),
.B(n_270),
.Y(n_3134)
);

AOI21xp5_ASAP7_75t_L g3135 ( 
.A1(n_2450),
.A2(n_271),
.B(n_272),
.Y(n_3135)
);

NAND2xp5_ASAP7_75t_L g3136 ( 
.A(n_2264),
.B(n_271),
.Y(n_3136)
);

AOI21xp5_ASAP7_75t_L g3137 ( 
.A1(n_2450),
.A2(n_272),
.B(n_273),
.Y(n_3137)
);

AOI21xp5_ASAP7_75t_L g3138 ( 
.A1(n_2450),
.A2(n_272),
.B(n_273),
.Y(n_3138)
);

INVx2_ASAP7_75t_L g3139 ( 
.A(n_2254),
.Y(n_3139)
);

OAI21xp5_ASAP7_75t_L g3140 ( 
.A1(n_2182),
.A2(n_273),
.B(n_274),
.Y(n_3140)
);

NOR2xp33_ASAP7_75t_L g3141 ( 
.A(n_2229),
.B(n_274),
.Y(n_3141)
);

INVx1_ASAP7_75t_L g3142 ( 
.A(n_2205),
.Y(n_3142)
);

O2A1O1Ixp33_ASAP7_75t_L g3143 ( 
.A1(n_2248),
.A2(n_276),
.B(n_274),
.C(n_275),
.Y(n_3143)
);

INVx1_ASAP7_75t_L g3144 ( 
.A(n_2205),
.Y(n_3144)
);

AOI21xp5_ASAP7_75t_L g3145 ( 
.A1(n_2450),
.A2(n_275),
.B(n_276),
.Y(n_3145)
);

OAI21xp5_ASAP7_75t_L g3146 ( 
.A1(n_2182),
.A2(n_276),
.B(n_277),
.Y(n_3146)
);

NAND2xp5_ASAP7_75t_SL g3147 ( 
.A(n_2262),
.B(n_278),
.Y(n_3147)
);

NAND2xp5_ASAP7_75t_SL g3148 ( 
.A(n_2262),
.B(n_278),
.Y(n_3148)
);

AOI21xp5_ASAP7_75t_L g3149 ( 
.A1(n_2450),
.A2(n_277),
.B(n_278),
.Y(n_3149)
);

NAND2xp33_ASAP7_75t_SL g3150 ( 
.A(n_2231),
.B(n_277),
.Y(n_3150)
);

AOI21xp5_ASAP7_75t_L g3151 ( 
.A1(n_2450),
.A2(n_279),
.B(n_280),
.Y(n_3151)
);

AOI21xp5_ASAP7_75t_L g3152 ( 
.A1(n_2450),
.A2(n_279),
.B(n_280),
.Y(n_3152)
);

AOI21xp5_ASAP7_75t_L g3153 ( 
.A1(n_2450),
.A2(n_279),
.B(n_280),
.Y(n_3153)
);

NAND2xp5_ASAP7_75t_SL g3154 ( 
.A(n_2262),
.B(n_282),
.Y(n_3154)
);

INVx1_ASAP7_75t_L g3155 ( 
.A(n_2205),
.Y(n_3155)
);

OAI21x1_ASAP7_75t_L g3156 ( 
.A1(n_2447),
.A2(n_715),
.B(n_714),
.Y(n_3156)
);

AOI22xp5_ASAP7_75t_L g3157 ( 
.A1(n_2213),
.A2(n_283),
.B1(n_281),
.B2(n_282),
.Y(n_3157)
);

OAI21xp5_ASAP7_75t_L g3158 ( 
.A1(n_2182),
.A2(n_281),
.B(n_282),
.Y(n_3158)
);

AND2x2_ASAP7_75t_L g3159 ( 
.A(n_2210),
.B(n_281),
.Y(n_3159)
);

INVx1_ASAP7_75t_L g3160 ( 
.A(n_2564),
.Y(n_3160)
);

INVx2_ASAP7_75t_L g3161 ( 
.A(n_2546),
.Y(n_3161)
);

BUFx8_ASAP7_75t_L g3162 ( 
.A(n_2626),
.Y(n_3162)
);

NAND2xp5_ASAP7_75t_L g3163 ( 
.A(n_2678),
.B(n_283),
.Y(n_3163)
);

INVx2_ASAP7_75t_L g3164 ( 
.A(n_2936),
.Y(n_3164)
);

AOI21xp5_ASAP7_75t_L g3165 ( 
.A1(n_2710),
.A2(n_283),
.B(n_285),
.Y(n_3165)
);

INVx1_ASAP7_75t_L g3166 ( 
.A(n_2565),
.Y(n_3166)
);

INVx1_ASAP7_75t_L g3167 ( 
.A(n_2912),
.Y(n_3167)
);

BUFx8_ASAP7_75t_SL g3168 ( 
.A(n_2661),
.Y(n_3168)
);

NAND2xp5_ASAP7_75t_L g3169 ( 
.A(n_2575),
.B(n_285),
.Y(n_3169)
);

AOI21xp5_ASAP7_75t_L g3170 ( 
.A1(n_2809),
.A2(n_286),
.B(n_287),
.Y(n_3170)
);

BUFx3_ASAP7_75t_L g3171 ( 
.A(n_2663),
.Y(n_3171)
);

NAND2xp5_ASAP7_75t_SL g3172 ( 
.A(n_2983),
.B(n_2949),
.Y(n_3172)
);

OAI21xp33_ASAP7_75t_L g3173 ( 
.A1(n_2983),
.A2(n_286),
.B(n_287),
.Y(n_3173)
);

NAND3xp33_ASAP7_75t_L g3174 ( 
.A(n_2652),
.B(n_286),
.C(n_288),
.Y(n_3174)
);

BUFx6f_ASAP7_75t_L g3175 ( 
.A(n_2804),
.Y(n_3175)
);

OAI22xp5_ASAP7_75t_L g3176 ( 
.A1(n_2539),
.A2(n_291),
.B1(n_288),
.B2(n_290),
.Y(n_3176)
);

BUFx2_ASAP7_75t_L g3177 ( 
.A(n_2663),
.Y(n_3177)
);

BUFx6f_ASAP7_75t_L g3178 ( 
.A(n_2804),
.Y(n_3178)
);

NAND2xp5_ASAP7_75t_SL g3179 ( 
.A(n_2949),
.B(n_717),
.Y(n_3179)
);

INVx1_ASAP7_75t_L g3180 ( 
.A(n_2914),
.Y(n_3180)
);

OAI22xp5_ASAP7_75t_L g3181 ( 
.A1(n_3086),
.A2(n_291),
.B1(n_288),
.B2(n_290),
.Y(n_3181)
);

INVx2_ASAP7_75t_L g3182 ( 
.A(n_2982),
.Y(n_3182)
);

AOI21xp5_ASAP7_75t_L g3183 ( 
.A1(n_2621),
.A2(n_291),
.B(n_292),
.Y(n_3183)
);

AOI21xp5_ASAP7_75t_L g3184 ( 
.A1(n_2555),
.A2(n_293),
.B(n_294),
.Y(n_3184)
);

INVx2_ASAP7_75t_L g3185 ( 
.A(n_3028),
.Y(n_3185)
);

AOI21xp5_ASAP7_75t_L g3186 ( 
.A1(n_2619),
.A2(n_293),
.B(n_294),
.Y(n_3186)
);

NOR2xp33_ASAP7_75t_L g3187 ( 
.A(n_2576),
.B(n_295),
.Y(n_3187)
);

CKINVDCx16_ASAP7_75t_R g3188 ( 
.A(n_2558),
.Y(n_3188)
);

AOI21xp5_ASAP7_75t_L g3189 ( 
.A1(n_2751),
.A2(n_2640),
.B(n_2771),
.Y(n_3189)
);

AOI22xp5_ASAP7_75t_L g3190 ( 
.A1(n_2647),
.A2(n_297),
.B1(n_295),
.B2(n_296),
.Y(n_3190)
);

INVx2_ASAP7_75t_L g3191 ( 
.A(n_3032),
.Y(n_3191)
);

AND2x2_ASAP7_75t_SL g3192 ( 
.A(n_2924),
.B(n_3042),
.Y(n_3192)
);

NAND2xp5_ASAP7_75t_L g3193 ( 
.A(n_2618),
.B(n_296),
.Y(n_3193)
);

INVx2_ASAP7_75t_L g3194 ( 
.A(n_3058),
.Y(n_3194)
);

AOI21x1_ASAP7_75t_L g3195 ( 
.A1(n_2582),
.A2(n_297),
.B(n_298),
.Y(n_3195)
);

NOR2xp33_ASAP7_75t_L g3196 ( 
.A(n_2793),
.B(n_297),
.Y(n_3196)
);

AOI22xp33_ASAP7_75t_L g3197 ( 
.A1(n_2799),
.A2(n_2778),
.B1(n_2794),
.B2(n_2609),
.Y(n_3197)
);

OAI22xp5_ASAP7_75t_L g3198 ( 
.A1(n_2870),
.A2(n_300),
.B1(n_298),
.B2(n_299),
.Y(n_3198)
);

AOI22xp33_ASAP7_75t_L g3199 ( 
.A1(n_2778),
.A2(n_300),
.B1(n_298),
.B2(n_299),
.Y(n_3199)
);

NOR2xp33_ASAP7_75t_L g3200 ( 
.A(n_2793),
.B(n_300),
.Y(n_3200)
);

INVx2_ASAP7_75t_L g3201 ( 
.A(n_3062),
.Y(n_3201)
);

INVxp67_ASAP7_75t_L g3202 ( 
.A(n_2543),
.Y(n_3202)
);

NOR2xp33_ASAP7_75t_L g3203 ( 
.A(n_2566),
.B(n_2749),
.Y(n_3203)
);

INVx2_ASAP7_75t_L g3204 ( 
.A(n_3078),
.Y(n_3204)
);

BUFx2_ASAP7_75t_L g3205 ( 
.A(n_2924),
.Y(n_3205)
);

AOI21xp5_ASAP7_75t_L g3206 ( 
.A1(n_2900),
.A2(n_301),
.B(n_302),
.Y(n_3206)
);

OAI21xp33_ASAP7_75t_L g3207 ( 
.A1(n_2572),
.A2(n_301),
.B(n_302),
.Y(n_3207)
);

NOR2xp67_ASAP7_75t_L g3208 ( 
.A(n_2554),
.B(n_303),
.Y(n_3208)
);

INVx2_ASAP7_75t_L g3209 ( 
.A(n_3084),
.Y(n_3209)
);

O2A1O1Ixp33_ASAP7_75t_L g3210 ( 
.A1(n_2540),
.A2(n_305),
.B(n_303),
.C(n_304),
.Y(n_3210)
);

NOR2xp33_ASAP7_75t_L g3211 ( 
.A(n_2756),
.B(n_2757),
.Y(n_3211)
);

NAND2xp5_ASAP7_75t_L g3212 ( 
.A(n_2935),
.B(n_303),
.Y(n_3212)
);

AOI21x1_ASAP7_75t_L g3213 ( 
.A1(n_2713),
.A2(n_304),
.B(n_305),
.Y(n_3213)
);

OAI21x1_ASAP7_75t_L g3214 ( 
.A1(n_2674),
.A2(n_305),
.B(n_306),
.Y(n_3214)
);

AOI22xp33_ASAP7_75t_L g3215 ( 
.A1(n_2625),
.A2(n_308),
.B1(n_306),
.B2(n_307),
.Y(n_3215)
);

INVx1_ASAP7_75t_SL g3216 ( 
.A(n_2987),
.Y(n_3216)
);

BUFx2_ASAP7_75t_L g3217 ( 
.A(n_3042),
.Y(n_3217)
);

CKINVDCx6p67_ASAP7_75t_R g3218 ( 
.A(n_2554),
.Y(n_3218)
);

BUFx12f_ASAP7_75t_L g3219 ( 
.A(n_3017),
.Y(n_3219)
);

CKINVDCx5p33_ASAP7_75t_R g3220 ( 
.A(n_3087),
.Y(n_3220)
);

AOI21xp5_ASAP7_75t_L g3221 ( 
.A1(n_2904),
.A2(n_306),
.B(n_307),
.Y(n_3221)
);

AOI21xp5_ASAP7_75t_L g3222 ( 
.A1(n_2905),
.A2(n_307),
.B(n_308),
.Y(n_3222)
);

O2A1O1Ixp33_ASAP7_75t_L g3223 ( 
.A1(n_2547),
.A2(n_310),
.B(n_308),
.C(n_309),
.Y(n_3223)
);

NAND2xp5_ASAP7_75t_L g3224 ( 
.A(n_2940),
.B(n_309),
.Y(n_3224)
);

INVx2_ASAP7_75t_L g3225 ( 
.A(n_3096),
.Y(n_3225)
);

INVx2_ASAP7_75t_L g3226 ( 
.A(n_3139),
.Y(n_3226)
);

OAI22xp5_ASAP7_75t_L g3227 ( 
.A1(n_2870),
.A2(n_312),
.B1(n_309),
.B2(n_310),
.Y(n_3227)
);

AOI21xp5_ASAP7_75t_L g3228 ( 
.A1(n_2906),
.A2(n_310),
.B(n_312),
.Y(n_3228)
);

BUFx12f_ASAP7_75t_L g3229 ( 
.A(n_3112),
.Y(n_3229)
);

AOI21xp5_ASAP7_75t_L g3230 ( 
.A1(n_2907),
.A2(n_312),
.B(n_313),
.Y(n_3230)
);

NAND2xp5_ASAP7_75t_L g3231 ( 
.A(n_2952),
.B(n_314),
.Y(n_3231)
);

INVx2_ASAP7_75t_L g3232 ( 
.A(n_2559),
.Y(n_3232)
);

INVx2_ASAP7_75t_L g3233 ( 
.A(n_2579),
.Y(n_3233)
);

INVxp67_ASAP7_75t_L g3234 ( 
.A(n_3059),
.Y(n_3234)
);

A2O1A1Ixp33_ASAP7_75t_L g3235 ( 
.A1(n_2873),
.A2(n_317),
.B(n_314),
.C(n_316),
.Y(n_3235)
);

AOI21xp5_ASAP7_75t_L g3236 ( 
.A1(n_2913),
.A2(n_314),
.B(n_316),
.Y(n_3236)
);

BUFx6f_ASAP7_75t_L g3237 ( 
.A(n_2804),
.Y(n_3237)
);

O2A1O1Ixp33_ASAP7_75t_L g3238 ( 
.A1(n_2708),
.A2(n_2594),
.B(n_2785),
.C(n_2795),
.Y(n_3238)
);

INVx1_ASAP7_75t_L g3239 ( 
.A(n_2957),
.Y(n_3239)
);

AOI21xp5_ASAP7_75t_L g3240 ( 
.A1(n_2915),
.A2(n_316),
.B(n_317),
.Y(n_3240)
);

NOR2xp33_ASAP7_75t_L g3241 ( 
.A(n_2720),
.B(n_317),
.Y(n_3241)
);

NOR3xp33_ASAP7_75t_SL g3242 ( 
.A(n_2672),
.B(n_318),
.C(n_319),
.Y(n_3242)
);

BUFx12f_ASAP7_75t_L g3243 ( 
.A(n_2558),
.Y(n_3243)
);

OAI21xp33_ASAP7_75t_L g3244 ( 
.A1(n_2638),
.A2(n_318),
.B(n_319),
.Y(n_3244)
);

A2O1A1Ixp33_ASAP7_75t_L g3245 ( 
.A1(n_2636),
.A2(n_320),
.B(n_318),
.C(n_319),
.Y(n_3245)
);

O2A1O1Ixp33_ASAP7_75t_L g3246 ( 
.A1(n_2910),
.A2(n_322),
.B(n_320),
.C(n_321),
.Y(n_3246)
);

INVx3_ASAP7_75t_L g3247 ( 
.A(n_2554),
.Y(n_3247)
);

INVx1_ASAP7_75t_L g3248 ( 
.A(n_2958),
.Y(n_3248)
);

AOI21xp5_ASAP7_75t_L g3249 ( 
.A1(n_2928),
.A2(n_320),
.B(n_321),
.Y(n_3249)
);

NAND2xp5_ASAP7_75t_SL g3250 ( 
.A(n_2987),
.B(n_717),
.Y(n_3250)
);

BUFx6f_ASAP7_75t_L g3251 ( 
.A(n_2821),
.Y(n_3251)
);

AOI21xp5_ASAP7_75t_L g3252 ( 
.A1(n_2931),
.A2(n_321),
.B(n_323),
.Y(n_3252)
);

AOI21xp5_ASAP7_75t_L g3253 ( 
.A1(n_2933),
.A2(n_323),
.B(n_324),
.Y(n_3253)
);

OR2x6_ASAP7_75t_L g3254 ( 
.A(n_3027),
.B(n_323),
.Y(n_3254)
);

AOI21xp5_ASAP7_75t_L g3255 ( 
.A1(n_2934),
.A2(n_324),
.B(n_325),
.Y(n_3255)
);

OR2x2_ASAP7_75t_L g3256 ( 
.A(n_3029),
.B(n_3124),
.Y(n_3256)
);

INVx1_ASAP7_75t_L g3257 ( 
.A(n_2988),
.Y(n_3257)
);

A2O1A1Ixp33_ASAP7_75t_SL g3258 ( 
.A1(n_2754),
.A2(n_328),
.B(n_325),
.C(n_326),
.Y(n_3258)
);

O2A1O1Ixp33_ASAP7_75t_L g3259 ( 
.A1(n_2721),
.A2(n_328),
.B(n_325),
.C(n_326),
.Y(n_3259)
);

INVx3_ASAP7_75t_L g3260 ( 
.A(n_2554),
.Y(n_3260)
);

A2O1A1Ixp33_ASAP7_75t_L g3261 ( 
.A1(n_3150),
.A2(n_330),
.B(n_326),
.C(n_329),
.Y(n_3261)
);

NAND2xp5_ASAP7_75t_L g3262 ( 
.A(n_2989),
.B(n_329),
.Y(n_3262)
);

CKINVDCx5p33_ASAP7_75t_R g3263 ( 
.A(n_3056),
.Y(n_3263)
);

NOR2xp33_ASAP7_75t_SL g3264 ( 
.A(n_3027),
.B(n_329),
.Y(n_3264)
);

A2O1A1Ixp33_ASAP7_75t_L g3265 ( 
.A1(n_2725),
.A2(n_332),
.B(n_330),
.C(n_331),
.Y(n_3265)
);

AOI21xp5_ASAP7_75t_L g3266 ( 
.A1(n_2941),
.A2(n_330),
.B(n_331),
.Y(n_3266)
);

INVx3_ASAP7_75t_L g3267 ( 
.A(n_2824),
.Y(n_3267)
);

NOR2xp33_ASAP7_75t_L g3268 ( 
.A(n_3029),
.B(n_332),
.Y(n_3268)
);

INVx4_ASAP7_75t_L g3269 ( 
.A(n_3050),
.Y(n_3269)
);

AOI21xp5_ASAP7_75t_L g3270 ( 
.A1(n_2944),
.A2(n_332),
.B(n_333),
.Y(n_3270)
);

INVx2_ASAP7_75t_L g3271 ( 
.A(n_2602),
.Y(n_3271)
);

NOR2xp67_ASAP7_75t_SL g3272 ( 
.A(n_3050),
.B(n_333),
.Y(n_3272)
);

INVx2_ASAP7_75t_L g3273 ( 
.A(n_2604),
.Y(n_3273)
);

NAND2xp5_ASAP7_75t_L g3274 ( 
.A(n_2998),
.B(n_333),
.Y(n_3274)
);

BUFx6f_ASAP7_75t_L g3275 ( 
.A(n_2821),
.Y(n_3275)
);

NAND3xp33_ASAP7_75t_SL g3276 ( 
.A(n_2642),
.B(n_334),
.C(n_335),
.Y(n_3276)
);

AOI21xp5_ASAP7_75t_L g3277 ( 
.A1(n_2960),
.A2(n_334),
.B(n_335),
.Y(n_3277)
);

NAND2xp5_ASAP7_75t_SL g3278 ( 
.A(n_2642),
.B(n_718),
.Y(n_3278)
);

CKINVDCx20_ASAP7_75t_R g3279 ( 
.A(n_2926),
.Y(n_3279)
);

AND2x2_ASAP7_75t_L g3280 ( 
.A(n_2901),
.B(n_335),
.Y(n_3280)
);

INVx1_ASAP7_75t_L g3281 ( 
.A(n_3019),
.Y(n_3281)
);

AOI21xp5_ASAP7_75t_L g3282 ( 
.A1(n_2964),
.A2(n_336),
.B(n_337),
.Y(n_3282)
);

INVx1_ASAP7_75t_L g3283 ( 
.A(n_3031),
.Y(n_3283)
);

NAND2xp5_ASAP7_75t_L g3284 ( 
.A(n_3038),
.B(n_336),
.Y(n_3284)
);

A2O1A1Ixp33_ASAP7_75t_L g3285 ( 
.A1(n_2651),
.A2(n_338),
.B(n_336),
.C(n_337),
.Y(n_3285)
);

AOI21xp5_ASAP7_75t_L g3286 ( 
.A1(n_2980),
.A2(n_337),
.B(n_338),
.Y(n_3286)
);

INVx5_ASAP7_75t_L g3287 ( 
.A(n_2870),
.Y(n_3287)
);

OAI22xp5_ASAP7_75t_L g3288 ( 
.A1(n_2824),
.A2(n_340),
.B1(n_338),
.B2(n_339),
.Y(n_3288)
);

INVx4_ASAP7_75t_L g3289 ( 
.A(n_2932),
.Y(n_3289)
);

AND2x2_ASAP7_75t_L g3290 ( 
.A(n_2908),
.B(n_339),
.Y(n_3290)
);

INVx3_ASAP7_75t_L g3291 ( 
.A(n_2824),
.Y(n_3291)
);

NAND2xp5_ASAP7_75t_SL g3292 ( 
.A(n_2824),
.B(n_718),
.Y(n_3292)
);

AOI21xp5_ASAP7_75t_L g3293 ( 
.A1(n_2981),
.A2(n_339),
.B(n_341),
.Y(n_3293)
);

AOI22xp33_ASAP7_75t_L g3294 ( 
.A1(n_2719),
.A2(n_2858),
.B1(n_2730),
.B2(n_2971),
.Y(n_3294)
);

NAND2xp5_ASAP7_75t_L g3295 ( 
.A(n_3067),
.B(n_341),
.Y(n_3295)
);

AOI21xp5_ASAP7_75t_L g3296 ( 
.A1(n_2985),
.A2(n_341),
.B(n_342),
.Y(n_3296)
);

INVx4_ASAP7_75t_L g3297 ( 
.A(n_2939),
.Y(n_3297)
);

AOI21xp5_ASAP7_75t_L g3298 ( 
.A1(n_2994),
.A2(n_342),
.B(n_343),
.Y(n_3298)
);

NAND3xp33_ASAP7_75t_SL g3299 ( 
.A(n_2867),
.B(n_342),
.C(n_343),
.Y(n_3299)
);

NAND2xp5_ASAP7_75t_L g3300 ( 
.A(n_3070),
.B(n_343),
.Y(n_3300)
);

NAND2xp5_ASAP7_75t_L g3301 ( 
.A(n_3075),
.B(n_344),
.Y(n_3301)
);

NAND2xp5_ASAP7_75t_SL g3302 ( 
.A(n_2807),
.B(n_719),
.Y(n_3302)
);

NAND2xp5_ASAP7_75t_L g3303 ( 
.A(n_3117),
.B(n_344),
.Y(n_3303)
);

NAND2xp5_ASAP7_75t_SL g3304 ( 
.A(n_2852),
.B(n_2991),
.Y(n_3304)
);

OAI22xp5_ASAP7_75t_L g3305 ( 
.A1(n_2562),
.A2(n_346),
.B1(n_344),
.B2(n_345),
.Y(n_3305)
);

INVx2_ASAP7_75t_L g3306 ( 
.A(n_2634),
.Y(n_3306)
);

AOI33xp33_ASAP7_75t_L g3307 ( 
.A1(n_2571),
.A2(n_347),
.A3(n_349),
.B1(n_345),
.B2(n_346),
.B3(n_348),
.Y(n_3307)
);

NAND2xp5_ASAP7_75t_SL g3308 ( 
.A(n_2945),
.B(n_719),
.Y(n_3308)
);

BUFx6f_ASAP7_75t_L g3309 ( 
.A(n_2821),
.Y(n_3309)
);

AOI21xp5_ASAP7_75t_L g3310 ( 
.A1(n_2997),
.A2(n_345),
.B(n_347),
.Y(n_3310)
);

OAI21xp5_ASAP7_75t_L g3311 ( 
.A1(n_2563),
.A2(n_348),
.B(n_349),
.Y(n_3311)
);

OAI22xp5_ASAP7_75t_L g3312 ( 
.A1(n_2562),
.A2(n_352),
.B1(n_350),
.B2(n_351),
.Y(n_3312)
);

INVx2_ASAP7_75t_L g3313 ( 
.A(n_2641),
.Y(n_3313)
);

INVx2_ASAP7_75t_L g3314 ( 
.A(n_3142),
.Y(n_3314)
);

INVx1_ASAP7_75t_L g3315 ( 
.A(n_3144),
.Y(n_3315)
);

NAND2xp5_ASAP7_75t_SL g3316 ( 
.A(n_3119),
.B(n_720),
.Y(n_3316)
);

INVx5_ASAP7_75t_L g3317 ( 
.A(n_2562),
.Y(n_3317)
);

A2O1A1Ixp33_ASAP7_75t_L g3318 ( 
.A1(n_2747),
.A2(n_352),
.B(n_350),
.C(n_351),
.Y(n_3318)
);

NOR2xp33_ASAP7_75t_L g3319 ( 
.A(n_2650),
.B(n_350),
.Y(n_3319)
);

NAND2xp5_ASAP7_75t_L g3320 ( 
.A(n_3155),
.B(n_351),
.Y(n_3320)
);

INVx1_ASAP7_75t_L g3321 ( 
.A(n_2599),
.Y(n_3321)
);

NAND2xp5_ASAP7_75t_L g3322 ( 
.A(n_2561),
.B(n_352),
.Y(n_3322)
);

BUFx8_ASAP7_75t_L g3323 ( 
.A(n_2667),
.Y(n_3323)
);

NAND2xp5_ASAP7_75t_L g3324 ( 
.A(n_2600),
.B(n_353),
.Y(n_3324)
);

INVx1_ASAP7_75t_L g3325 ( 
.A(n_2613),
.Y(n_3325)
);

INVx1_ASAP7_75t_L g3326 ( 
.A(n_2620),
.Y(n_3326)
);

O2A1O1Ixp33_ASAP7_75t_L g3327 ( 
.A1(n_2836),
.A2(n_355),
.B(n_353),
.C(n_354),
.Y(n_3327)
);

A2O1A1Ixp33_ASAP7_75t_L g3328 ( 
.A1(n_2690),
.A2(n_356),
.B(n_354),
.C(n_355),
.Y(n_3328)
);

NAND3xp33_ASAP7_75t_SL g3329 ( 
.A(n_2792),
.B(n_354),
.C(n_356),
.Y(n_3329)
);

INVx2_ASAP7_75t_L g3330 ( 
.A(n_2633),
.Y(n_3330)
);

INVx1_ASAP7_75t_L g3331 ( 
.A(n_2653),
.Y(n_3331)
);

INVx1_ASAP7_75t_L g3332 ( 
.A(n_2654),
.Y(n_3332)
);

NAND2xp5_ASAP7_75t_SL g3333 ( 
.A(n_2922),
.B(n_720),
.Y(n_3333)
);

NOR3xp33_ASAP7_75t_SL g3334 ( 
.A(n_2995),
.B(n_2760),
.C(n_2735),
.Y(n_3334)
);

NAND2xp5_ASAP7_75t_SL g3335 ( 
.A(n_2922),
.B(n_721),
.Y(n_3335)
);

NAND2x1p5_ASAP7_75t_L g3336 ( 
.A(n_2968),
.B(n_356),
.Y(n_3336)
);

A2O1A1Ixp33_ASAP7_75t_L g3337 ( 
.A1(n_2704),
.A2(n_359),
.B(n_357),
.C(n_358),
.Y(n_3337)
);

AOI22xp5_ASAP7_75t_L g3338 ( 
.A1(n_2884),
.A2(n_359),
.B1(n_357),
.B2(n_358),
.Y(n_3338)
);

INVx1_ASAP7_75t_L g3339 ( 
.A(n_2666),
.Y(n_3339)
);

AOI21xp5_ASAP7_75t_L g3340 ( 
.A1(n_2999),
.A2(n_357),
.B(n_358),
.Y(n_3340)
);

INVx1_ASAP7_75t_L g3341 ( 
.A(n_2692),
.Y(n_3341)
);

NAND2xp5_ASAP7_75t_SL g3342 ( 
.A(n_2929),
.B(n_722),
.Y(n_3342)
);

INVx2_ASAP7_75t_L g3343 ( 
.A(n_2700),
.Y(n_3343)
);

BUFx2_ASAP7_75t_L g3344 ( 
.A(n_3000),
.Y(n_3344)
);

INVxp67_ASAP7_75t_L g3345 ( 
.A(n_2545),
.Y(n_3345)
);

NOR2xp33_ASAP7_75t_L g3346 ( 
.A(n_2775),
.B(n_359),
.Y(n_3346)
);

AOI21xp5_ASAP7_75t_L g3347 ( 
.A1(n_3002),
.A2(n_360),
.B(n_361),
.Y(n_3347)
);

BUFx2_ASAP7_75t_L g3348 ( 
.A(n_2970),
.Y(n_3348)
);

A2O1A1Ixp33_ASAP7_75t_SL g3349 ( 
.A1(n_2573),
.A2(n_362),
.B(n_360),
.C(n_361),
.Y(n_3349)
);

OAI21x1_ASAP7_75t_L g3350 ( 
.A1(n_2674),
.A2(n_360),
.B(n_361),
.Y(n_3350)
);

OAI22x1_ASAP7_75t_L g3351 ( 
.A1(n_2673),
.A2(n_364),
.B1(n_362),
.B2(n_363),
.Y(n_3351)
);

AOI21x1_ASAP7_75t_L g3352 ( 
.A1(n_2591),
.A2(n_2859),
.B(n_2930),
.Y(n_3352)
);

NOR2x1_ASAP7_75t_L g3353 ( 
.A(n_2716),
.B(n_362),
.Y(n_3353)
);

BUFx6f_ASAP7_75t_L g3354 ( 
.A(n_2822),
.Y(n_3354)
);

OR2x2_ASAP7_75t_L g3355 ( 
.A(n_3001),
.B(n_3005),
.Y(n_3355)
);

NAND2xp5_ASAP7_75t_L g3356 ( 
.A(n_2942),
.B(n_363),
.Y(n_3356)
);

NOR2xp33_ASAP7_75t_R g3357 ( 
.A(n_2802),
.B(n_2731),
.Y(n_3357)
);

NAND2xp5_ASAP7_75t_L g3358 ( 
.A(n_2948),
.B(n_364),
.Y(n_3358)
);

AOI22xp33_ASAP7_75t_L g3359 ( 
.A1(n_2977),
.A2(n_367),
.B1(n_364),
.B2(n_365),
.Y(n_3359)
);

A2O1A1Ixp33_ASAP7_75t_L g3360 ( 
.A1(n_2705),
.A2(n_368),
.B(n_365),
.C(n_367),
.Y(n_3360)
);

AOI21xp5_ASAP7_75t_L g3361 ( 
.A1(n_3004),
.A2(n_367),
.B(n_368),
.Y(n_3361)
);

OR2x6_ASAP7_75t_SL g3362 ( 
.A(n_2923),
.B(n_368),
.Y(n_3362)
);

INVx1_ASAP7_75t_L g3363 ( 
.A(n_2703),
.Y(n_3363)
);

NOR2xp33_ASAP7_75t_R g3364 ( 
.A(n_2802),
.B(n_369),
.Y(n_3364)
);

NOR2xp33_ASAP7_75t_L g3365 ( 
.A(n_3132),
.B(n_2538),
.Y(n_3365)
);

INVx3_ASAP7_75t_SL g3366 ( 
.A(n_2777),
.Y(n_3366)
);

O2A1O1Ixp33_ASAP7_75t_L g3367 ( 
.A1(n_2628),
.A2(n_371),
.B(n_369),
.C(n_370),
.Y(n_3367)
);

AO22x1_ASAP7_75t_L g3368 ( 
.A1(n_2929),
.A2(n_371),
.B1(n_369),
.B2(n_370),
.Y(n_3368)
);

CKINVDCx16_ASAP7_75t_R g3369 ( 
.A(n_2668),
.Y(n_3369)
);

AOI222xp33_ASAP7_75t_L g3370 ( 
.A1(n_2789),
.A2(n_373),
.B1(n_375),
.B2(n_371),
.C1(n_372),
.C2(n_374),
.Y(n_3370)
);

NAND2x2_ASAP7_75t_L g3371 ( 
.A(n_2841),
.B(n_372),
.Y(n_3371)
);

INVx1_ASAP7_75t_L g3372 ( 
.A(n_2701),
.Y(n_3372)
);

NAND2xp5_ASAP7_75t_L g3373 ( 
.A(n_3074),
.B(n_373),
.Y(n_3373)
);

AOI22xp5_ASAP7_75t_L g3374 ( 
.A1(n_2656),
.A2(n_376),
.B1(n_374),
.B2(n_375),
.Y(n_3374)
);

INVx1_ASAP7_75t_L g3375 ( 
.A(n_2706),
.Y(n_3375)
);

NAND2xp5_ASAP7_75t_SL g3376 ( 
.A(n_3014),
.B(n_722),
.Y(n_3376)
);

INVx4_ASAP7_75t_L g3377 ( 
.A(n_3049),
.Y(n_3377)
);

AOI21xp5_ASAP7_75t_L g3378 ( 
.A1(n_3009),
.A2(n_374),
.B(n_375),
.Y(n_3378)
);

OAI21xp33_ASAP7_75t_L g3379 ( 
.A1(n_2560),
.A2(n_376),
.B(n_377),
.Y(n_3379)
);

NOR2xp33_ASAP7_75t_R g3380 ( 
.A(n_2833),
.B(n_376),
.Y(n_3380)
);

OAI22xp5_ASAP7_75t_L g3381 ( 
.A1(n_2588),
.A2(n_379),
.B1(n_377),
.B2(n_378),
.Y(n_3381)
);

AOI22x1_ASAP7_75t_L g3382 ( 
.A1(n_2608),
.A2(n_2670),
.B1(n_2715),
.B2(n_2707),
.Y(n_3382)
);

AOI21xp5_ASAP7_75t_L g3383 ( 
.A1(n_3021),
.A2(n_378),
.B(n_379),
.Y(n_3383)
);

AOI21xp5_ASAP7_75t_L g3384 ( 
.A1(n_3037),
.A2(n_378),
.B(n_380),
.Y(n_3384)
);

NAND2xp5_ASAP7_75t_L g3385 ( 
.A(n_3110),
.B(n_380),
.Y(n_3385)
);

INVx2_ASAP7_75t_L g3386 ( 
.A(n_2681),
.Y(n_3386)
);

OAI21xp5_ASAP7_75t_L g3387 ( 
.A1(n_2557),
.A2(n_380),
.B(n_381),
.Y(n_3387)
);

INVxp67_ASAP7_75t_L g3388 ( 
.A(n_2830),
.Y(n_3388)
);

AOI21xp5_ASAP7_75t_L g3389 ( 
.A1(n_3043),
.A2(n_381),
.B(n_382),
.Y(n_3389)
);

INVxp67_ASAP7_75t_SL g3390 ( 
.A(n_2862),
.Y(n_3390)
);

INVx1_ASAP7_75t_SL g3391 ( 
.A(n_3014),
.Y(n_3391)
);

OAI22xp5_ASAP7_75t_L g3392 ( 
.A1(n_2877),
.A2(n_384),
.B1(n_382),
.B2(n_383),
.Y(n_3392)
);

INVx1_ASAP7_75t_L g3393 ( 
.A(n_2611),
.Y(n_3393)
);

NOR2xp33_ASAP7_75t_L g3394 ( 
.A(n_2887),
.B(n_383),
.Y(n_3394)
);

AOI21xp5_ASAP7_75t_L g3395 ( 
.A1(n_3047),
.A2(n_384),
.B(n_385),
.Y(n_3395)
);

AOI22xp5_ASAP7_75t_L g3396 ( 
.A1(n_2567),
.A2(n_387),
.B1(n_385),
.B2(n_386),
.Y(n_3396)
);

AND2x2_ASAP7_75t_L g3397 ( 
.A(n_3130),
.B(n_386),
.Y(n_3397)
);

INVx2_ASAP7_75t_SL g3398 ( 
.A(n_2882),
.Y(n_3398)
);

NAND2xp5_ASAP7_75t_SL g3399 ( 
.A(n_3065),
.B(n_723),
.Y(n_3399)
);

OAI22xp5_ASAP7_75t_L g3400 ( 
.A1(n_2614),
.A2(n_391),
.B1(n_389),
.B2(n_390),
.Y(n_3400)
);

BUFx3_ASAP7_75t_L g3401 ( 
.A(n_2882),
.Y(n_3401)
);

NAND2xp5_ASAP7_75t_L g3402 ( 
.A(n_3159),
.B(n_389),
.Y(n_3402)
);

NAND2xp5_ASAP7_75t_L g3403 ( 
.A(n_2568),
.B(n_389),
.Y(n_3403)
);

NAND2xp5_ASAP7_75t_SL g3404 ( 
.A(n_3065),
.B(n_723),
.Y(n_3404)
);

AOI221xp5_ASAP7_75t_L g3405 ( 
.A1(n_2577),
.A2(n_393),
.B1(n_390),
.B2(n_392),
.C(n_394),
.Y(n_3405)
);

OAI22x1_ASAP7_75t_L g3406 ( 
.A1(n_2973),
.A2(n_394),
.B1(n_392),
.B2(n_393),
.Y(n_3406)
);

OR2x2_ASAP7_75t_L g3407 ( 
.A(n_2990),
.B(n_394),
.Y(n_3407)
);

AOI21xp5_ASAP7_75t_L g3408 ( 
.A1(n_3052),
.A2(n_395),
.B(n_396),
.Y(n_3408)
);

NOR2xp33_ASAP7_75t_L g3409 ( 
.A(n_2549),
.B(n_395),
.Y(n_3409)
);

AOI21xp5_ASAP7_75t_L g3410 ( 
.A1(n_3055),
.A2(n_395),
.B(n_396),
.Y(n_3410)
);

NOR2xp33_ASAP7_75t_L g3411 ( 
.A(n_2553),
.B(n_396),
.Y(n_3411)
);

OAI21x1_ASAP7_75t_L g3412 ( 
.A1(n_3156),
.A2(n_397),
.B(n_398),
.Y(n_3412)
);

O2A1O1Ixp5_ASAP7_75t_L g3413 ( 
.A1(n_2607),
.A2(n_399),
.B(n_397),
.C(n_398),
.Y(n_3413)
);

NAND2xp5_ASAP7_75t_L g3414 ( 
.A(n_2648),
.B(n_397),
.Y(n_3414)
);

NAND2xp5_ASAP7_75t_L g3415 ( 
.A(n_2838),
.B(n_398),
.Y(n_3415)
);

A2O1A1Ixp33_ASAP7_75t_L g3416 ( 
.A1(n_2724),
.A2(n_401),
.B(n_399),
.C(n_400),
.Y(n_3416)
);

BUFx2_ASAP7_75t_L g3417 ( 
.A(n_3123),
.Y(n_3417)
);

BUFx4f_ASAP7_75t_L g3418 ( 
.A(n_3123),
.Y(n_3418)
);

CKINVDCx14_ASAP7_75t_R g3419 ( 
.A(n_3012),
.Y(n_3419)
);

INVx1_ASAP7_75t_SL g3420 ( 
.A(n_3133),
.Y(n_3420)
);

NAND2xp5_ASAP7_75t_L g3421 ( 
.A(n_2846),
.B(n_400),
.Y(n_3421)
);

INVx1_ASAP7_75t_L g3422 ( 
.A(n_2612),
.Y(n_3422)
);

BUFx6f_ASAP7_75t_L g3423 ( 
.A(n_2822),
.Y(n_3423)
);

NAND2xp5_ASAP7_75t_L g3424 ( 
.A(n_2691),
.B(n_400),
.Y(n_3424)
);

NAND2xp5_ASAP7_75t_SL g3425 ( 
.A(n_3133),
.B(n_724),
.Y(n_3425)
);

AOI21xp5_ASAP7_75t_L g3426 ( 
.A1(n_3064),
.A2(n_401),
.B(n_402),
.Y(n_3426)
);

A2O1A1Ixp33_ASAP7_75t_L g3427 ( 
.A1(n_2737),
.A2(n_404),
.B(n_402),
.C(n_403),
.Y(n_3427)
);

NAND2xp5_ASAP7_75t_L g3428 ( 
.A(n_2631),
.B(n_402),
.Y(n_3428)
);

INVx5_ASAP7_75t_L g3429 ( 
.A(n_2729),
.Y(n_3429)
);

NAND3xp33_ASAP7_75t_SL g3430 ( 
.A(n_2759),
.B(n_403),
.C(n_404),
.Y(n_3430)
);

BUFx6f_ASAP7_75t_L g3431 ( 
.A(n_2822),
.Y(n_3431)
);

A2O1A1Ixp33_ASAP7_75t_L g3432 ( 
.A1(n_2738),
.A2(n_407),
.B(n_405),
.C(n_406),
.Y(n_3432)
);

CKINVDCx16_ASAP7_75t_R g3433 ( 
.A(n_2687),
.Y(n_3433)
);

INVx3_ASAP7_75t_L g3434 ( 
.A(n_2570),
.Y(n_3434)
);

A2O1A1Ixp33_ASAP7_75t_L g3435 ( 
.A1(n_2768),
.A2(n_408),
.B(n_405),
.C(n_407),
.Y(n_3435)
);

AND2x2_ASAP7_75t_L g3436 ( 
.A(n_3109),
.B(n_407),
.Y(n_3436)
);

NAND2xp5_ASAP7_75t_SL g3437 ( 
.A(n_2570),
.B(n_724),
.Y(n_3437)
);

CKINVDCx6p67_ASAP7_75t_R g3438 ( 
.A(n_2886),
.Y(n_3438)
);

INVx2_ASAP7_75t_L g3439 ( 
.A(n_2694),
.Y(n_3439)
);

BUFx6f_ASAP7_75t_L g3440 ( 
.A(n_2548),
.Y(n_3440)
);

NOR2xp33_ASAP7_75t_L g3441 ( 
.A(n_2827),
.B(n_408),
.Y(n_3441)
);

NAND2xp5_ASAP7_75t_L g3442 ( 
.A(n_2605),
.B(n_409),
.Y(n_3442)
);

BUFx2_ASAP7_75t_L g3443 ( 
.A(n_2662),
.Y(n_3443)
);

NAND2xp5_ASAP7_75t_L g3444 ( 
.A(n_2984),
.B(n_3006),
.Y(n_3444)
);

O2A1O1Ixp33_ASAP7_75t_L g3445 ( 
.A1(n_2825),
.A2(n_411),
.B(n_409),
.C(n_410),
.Y(n_3445)
);

INVx1_ASAP7_75t_L g3446 ( 
.A(n_2616),
.Y(n_3446)
);

OAI22xp5_ASAP7_75t_L g3447 ( 
.A1(n_3008),
.A2(n_414),
.B1(n_412),
.B2(n_413),
.Y(n_3447)
);

INVx2_ASAP7_75t_L g3448 ( 
.A(n_2711),
.Y(n_3448)
);

INVx1_ASAP7_75t_L g3449 ( 
.A(n_3101),
.Y(n_3449)
);

OAI22xp5_ASAP7_75t_L g3450 ( 
.A1(n_3040),
.A2(n_416),
.B1(n_412),
.B2(n_415),
.Y(n_3450)
);

A2O1A1Ixp33_ASAP7_75t_L g3451 ( 
.A1(n_2773),
.A2(n_418),
.B(n_415),
.C(n_417),
.Y(n_3451)
);

A2O1A1Ixp33_ASAP7_75t_SL g3452 ( 
.A1(n_2649),
.A2(n_2780),
.B(n_2811),
.C(n_2803),
.Y(n_3452)
);

AOI21xp5_ASAP7_75t_L g3453 ( 
.A1(n_3073),
.A2(n_415),
.B(n_417),
.Y(n_3453)
);

AND2x2_ASAP7_75t_L g3454 ( 
.A(n_2680),
.B(n_417),
.Y(n_3454)
);

NOR2xp33_ASAP7_75t_R g3455 ( 
.A(n_2882),
.B(n_418),
.Y(n_3455)
);

BUFx3_ASAP7_75t_L g3456 ( 
.A(n_2869),
.Y(n_3456)
);

INVx1_ASAP7_75t_L g3457 ( 
.A(n_2742),
.Y(n_3457)
);

NAND2xp5_ASAP7_75t_L g3458 ( 
.A(n_3020),
.B(n_418),
.Y(n_3458)
);

NAND2xp5_ASAP7_75t_SL g3459 ( 
.A(n_2662),
.B(n_725),
.Y(n_3459)
);

OAI22xp5_ASAP7_75t_L g3460 ( 
.A1(n_3051),
.A2(n_421),
.B1(n_419),
.B2(n_420),
.Y(n_3460)
);

BUFx12f_ASAP7_75t_L g3461 ( 
.A(n_2881),
.Y(n_3461)
);

INVx1_ASAP7_75t_L g3462 ( 
.A(n_2744),
.Y(n_3462)
);

NAND3xp33_ASAP7_75t_SL g3463 ( 
.A(n_2976),
.B(n_419),
.C(n_420),
.Y(n_3463)
);

AOI21xp5_ASAP7_75t_L g3464 ( 
.A1(n_3080),
.A2(n_3083),
.B(n_3082),
.Y(n_3464)
);

O2A1O1Ixp33_ASAP7_75t_L g3465 ( 
.A1(n_2845),
.A2(n_423),
.B(n_421),
.C(n_422),
.Y(n_3465)
);

INVx1_ASAP7_75t_L g3466 ( 
.A(n_2814),
.Y(n_3466)
);

AOI21xp5_ASAP7_75t_L g3467 ( 
.A1(n_3100),
.A2(n_422),
.B(n_423),
.Y(n_3467)
);

AOI21xp5_ASAP7_75t_L g3468 ( 
.A1(n_3106),
.A2(n_3120),
.B(n_3118),
.Y(n_3468)
);

AOI21xp5_ASAP7_75t_L g3469 ( 
.A1(n_3125),
.A2(n_423),
.B(n_424),
.Y(n_3469)
);

OAI22xp5_ASAP7_75t_L g3470 ( 
.A1(n_3077),
.A2(n_426),
.B1(n_424),
.B2(n_425),
.Y(n_3470)
);

AOI21xp5_ASAP7_75t_L g3471 ( 
.A1(n_3134),
.A2(n_424),
.B(n_425),
.Y(n_3471)
);

BUFx6f_ASAP7_75t_L g3472 ( 
.A(n_2548),
.Y(n_3472)
);

INVx6_ASAP7_75t_L g3473 ( 
.A(n_2885),
.Y(n_3473)
);

INVx1_ASAP7_75t_L g3474 ( 
.A(n_2796),
.Y(n_3474)
);

NAND2xp5_ASAP7_75t_SL g3475 ( 
.A(n_2909),
.B(n_726),
.Y(n_3475)
);

INVx4_ASAP7_75t_L g3476 ( 
.A(n_2909),
.Y(n_3476)
);

OAI21xp5_ASAP7_75t_L g3477 ( 
.A1(n_2551),
.A2(n_425),
.B(n_426),
.Y(n_3477)
);

INVx1_ASAP7_75t_L g3478 ( 
.A(n_2806),
.Y(n_3478)
);

AOI221xp5_ASAP7_75t_L g3479 ( 
.A1(n_3023),
.A2(n_429),
.B1(n_427),
.B2(n_428),
.C(n_430),
.Y(n_3479)
);

AOI21xp5_ASAP7_75t_L g3480 ( 
.A1(n_3136),
.A2(n_427),
.B(n_428),
.Y(n_3480)
);

HB1xp67_ASAP7_75t_L g3481 ( 
.A(n_2718),
.Y(n_3481)
);

NAND2xp5_ASAP7_75t_L g3482 ( 
.A(n_3060),
.B(n_429),
.Y(n_3482)
);

A2O1A1Ixp33_ASAP7_75t_L g3483 ( 
.A1(n_2947),
.A2(n_2965),
.B(n_2978),
.C(n_2975),
.Y(n_3483)
);

AOI21xp5_ASAP7_75t_L g3484 ( 
.A1(n_2679),
.A2(n_429),
.B(n_430),
.Y(n_3484)
);

NAND2xp5_ASAP7_75t_L g3485 ( 
.A(n_3068),
.B(n_431),
.Y(n_3485)
);

INVx4_ASAP7_75t_L g3486 ( 
.A(n_2955),
.Y(n_3486)
);

OAI22xp5_ASAP7_75t_L g3487 ( 
.A1(n_3098),
.A2(n_433),
.B1(n_431),
.B2(n_432),
.Y(n_3487)
);

AOI21xp5_ASAP7_75t_L g3488 ( 
.A1(n_2684),
.A2(n_431),
.B(n_434),
.Y(n_3488)
);

A2O1A1Ixp33_ASAP7_75t_L g3489 ( 
.A1(n_3022),
.A2(n_436),
.B(n_434),
.C(n_435),
.Y(n_3489)
);

AOI21xp5_ASAP7_75t_L g3490 ( 
.A1(n_2686),
.A2(n_434),
.B(n_435),
.Y(n_3490)
);

INVx2_ASAP7_75t_L g3491 ( 
.A(n_2743),
.Y(n_3491)
);

A2O1A1Ixp33_ASAP7_75t_SL g3492 ( 
.A1(n_2903),
.A2(n_437),
.B(n_435),
.C(n_436),
.Y(n_3492)
);

INVx1_ASAP7_75t_L g3493 ( 
.A(n_2589),
.Y(n_3493)
);

OAI21xp5_ASAP7_75t_L g3494 ( 
.A1(n_2689),
.A2(n_436),
.B(n_437),
.Y(n_3494)
);

NAND2xp33_ASAP7_75t_SL g3495 ( 
.A(n_2899),
.B(n_2911),
.Y(n_3495)
);

NOR3xp33_ASAP7_75t_SL g3496 ( 
.A(n_2817),
.B(n_437),
.C(n_438),
.Y(n_3496)
);

NOR2xp33_ASAP7_75t_L g3497 ( 
.A(n_2837),
.B(n_438),
.Y(n_3497)
);

CKINVDCx20_ASAP7_75t_R g3498 ( 
.A(n_2843),
.Y(n_3498)
);

O2A1O1Ixp5_ASAP7_75t_L g3499 ( 
.A1(n_2734),
.A2(n_440),
.B(n_438),
.C(n_439),
.Y(n_3499)
);

AOI21xp5_ASAP7_75t_L g3500 ( 
.A1(n_2693),
.A2(n_439),
.B(n_440),
.Y(n_3500)
);

A2O1A1Ixp33_ASAP7_75t_L g3501 ( 
.A1(n_3024),
.A2(n_443),
.B(n_439),
.C(n_441),
.Y(n_3501)
);

CKINVDCx20_ASAP7_75t_R g3502 ( 
.A(n_3015),
.Y(n_3502)
);

NAND2x1p5_ASAP7_75t_L g3503 ( 
.A(n_2955),
.B(n_441),
.Y(n_3503)
);

OAI21xp33_ASAP7_75t_L g3504 ( 
.A1(n_3090),
.A2(n_443),
.B(n_444),
.Y(n_3504)
);

OAI21xp33_ASAP7_75t_L g3505 ( 
.A1(n_3141),
.A2(n_444),
.B(n_445),
.Y(n_3505)
);

O2A1O1Ixp33_ASAP7_75t_L g3506 ( 
.A1(n_2761),
.A2(n_447),
.B(n_445),
.C(n_446),
.Y(n_3506)
);

NOR2xp33_ASAP7_75t_R g3507 ( 
.A(n_2979),
.B(n_446),
.Y(n_3507)
);

OAI22xp5_ASAP7_75t_L g3508 ( 
.A1(n_3102),
.A2(n_448),
.B1(n_446),
.B2(n_447),
.Y(n_3508)
);

AOI21xp5_ASAP7_75t_L g3509 ( 
.A1(n_2617),
.A2(n_447),
.B(n_448),
.Y(n_3509)
);

AOI21xp5_ASAP7_75t_L g3510 ( 
.A1(n_2819),
.A2(n_448),
.B(n_449),
.Y(n_3510)
);

A2O1A1Ixp33_ASAP7_75t_SL g3511 ( 
.A1(n_2961),
.A2(n_451),
.B(n_449),
.C(n_450),
.Y(n_3511)
);

AOI21xp5_ASAP7_75t_L g3512 ( 
.A1(n_2726),
.A2(n_449),
.B(n_450),
.Y(n_3512)
);

INVx2_ASAP7_75t_L g3513 ( 
.A(n_2832),
.Y(n_3513)
);

A2O1A1Ixp33_ASAP7_75t_L g3514 ( 
.A1(n_3033),
.A2(n_452),
.B(n_450),
.C(n_451),
.Y(n_3514)
);

INVx1_ASAP7_75t_L g3515 ( 
.A(n_2592),
.Y(n_3515)
);

INVx4_ASAP7_75t_L g3516 ( 
.A(n_2979),
.Y(n_3516)
);

A2O1A1Ixp33_ASAP7_75t_L g3517 ( 
.A1(n_3035),
.A2(n_453),
.B(n_451),
.C(n_452),
.Y(n_3517)
);

NAND2xp5_ASAP7_75t_SL g3518 ( 
.A(n_3034),
.B(n_726),
.Y(n_3518)
);

OR2x2_ASAP7_75t_L g3519 ( 
.A(n_2541),
.B(n_453),
.Y(n_3519)
);

NAND2xp5_ASAP7_75t_L g3520 ( 
.A(n_2601),
.B(n_453),
.Y(n_3520)
);

AOI21xp33_ASAP7_75t_L g3521 ( 
.A1(n_2665),
.A2(n_454),
.B(n_456),
.Y(n_3521)
);

O2A1O1Ixp33_ASAP7_75t_L g3522 ( 
.A1(n_2770),
.A2(n_457),
.B(n_454),
.C(n_456),
.Y(n_3522)
);

AOI21xp5_ASAP7_75t_L g3523 ( 
.A1(n_2677),
.A2(n_456),
.B(n_457),
.Y(n_3523)
);

A2O1A1Ixp33_ASAP7_75t_SL g3524 ( 
.A1(n_2969),
.A2(n_459),
.B(n_457),
.C(n_458),
.Y(n_3524)
);

INVx3_ASAP7_75t_L g3525 ( 
.A(n_3034),
.Y(n_3525)
);

NAND2xp5_ASAP7_75t_L g3526 ( 
.A(n_2813),
.B(n_458),
.Y(n_3526)
);

OA22x2_ASAP7_75t_L g3527 ( 
.A1(n_2688),
.A2(n_461),
.B1(n_459),
.B2(n_460),
.Y(n_3527)
);

AND2x4_ASAP7_75t_L g3528 ( 
.A(n_3079),
.B(n_2718),
.Y(n_3528)
);

AOI21xp5_ASAP7_75t_L g3529 ( 
.A1(n_2727),
.A2(n_459),
.B(n_460),
.Y(n_3529)
);

INVx1_ASAP7_75t_L g3530 ( 
.A(n_2596),
.Y(n_3530)
);

AOI21xp5_ASAP7_75t_L g3531 ( 
.A1(n_2675),
.A2(n_2764),
.B(n_2748),
.Y(n_3531)
);

INVx2_ASAP7_75t_L g3532 ( 
.A(n_3018),
.Y(n_3532)
);

AOI21xp5_ASAP7_75t_L g3533 ( 
.A1(n_2766),
.A2(n_460),
.B(n_461),
.Y(n_3533)
);

A2O1A1Ixp33_ASAP7_75t_L g3534 ( 
.A1(n_3063),
.A2(n_463),
.B(n_461),
.C(n_462),
.Y(n_3534)
);

NOR2x1p5_ASAP7_75t_SL g3535 ( 
.A(n_3039),
.B(n_727),
.Y(n_3535)
);

NAND2xp5_ASAP7_75t_L g3536 ( 
.A(n_2753),
.B(n_2627),
.Y(n_3536)
);

INVx3_ASAP7_75t_L g3537 ( 
.A(n_3079),
.Y(n_3537)
);

O2A1O1Ixp33_ASAP7_75t_SL g3538 ( 
.A1(n_2635),
.A2(n_465),
.B(n_463),
.C(n_464),
.Y(n_3538)
);

INVx1_ASAP7_75t_L g3539 ( 
.A(n_2603),
.Y(n_3539)
);

O2A1O1Ixp5_ASAP7_75t_L g3540 ( 
.A1(n_2581),
.A2(n_465),
.B(n_463),
.C(n_464),
.Y(n_3540)
);

NOR3xp33_ASAP7_75t_L g3541 ( 
.A(n_2918),
.B(n_464),
.C(n_466),
.Y(n_3541)
);

OAI22xp5_ASAP7_75t_L g3542 ( 
.A1(n_2826),
.A2(n_468),
.B1(n_466),
.B2(n_467),
.Y(n_3542)
);

AND2x4_ASAP7_75t_L g3543 ( 
.A(n_2769),
.B(n_466),
.Y(n_3543)
);

NAND2xp5_ASAP7_75t_L g3544 ( 
.A(n_2722),
.B(n_467),
.Y(n_3544)
);

NAND2xp5_ASAP7_75t_SL g3545 ( 
.A(n_2587),
.B(n_728),
.Y(n_3545)
);

INVx1_ASAP7_75t_L g3546 ( 
.A(n_2762),
.Y(n_3546)
);

CKINVDCx5p33_ASAP7_75t_R g3547 ( 
.A(n_2630),
.Y(n_3547)
);

NOR2xp33_ASAP7_75t_SL g3548 ( 
.A(n_2709),
.B(n_467),
.Y(n_3548)
);

OAI22xp5_ASAP7_75t_L g3549 ( 
.A1(n_2849),
.A2(n_470),
.B1(n_468),
.B2(n_469),
.Y(n_3549)
);

AOI21xp5_ASAP7_75t_L g3550 ( 
.A1(n_2767),
.A2(n_468),
.B(n_470),
.Y(n_3550)
);

INVx1_ASAP7_75t_SL g3551 ( 
.A(n_2869),
.Y(n_3551)
);

INVx1_ASAP7_75t_L g3552 ( 
.A(n_2733),
.Y(n_3552)
);

NAND2xp5_ASAP7_75t_L g3553 ( 
.A(n_2758),
.B(n_470),
.Y(n_3553)
);

INVx3_ASAP7_75t_L g3554 ( 
.A(n_2729),
.Y(n_3554)
);

AOI21xp5_ASAP7_75t_L g3555 ( 
.A1(n_2645),
.A2(n_471),
.B(n_472),
.Y(n_3555)
);

BUFx4f_ASAP7_75t_L g3556 ( 
.A(n_2871),
.Y(n_3556)
);

BUFx6f_ASAP7_75t_L g3557 ( 
.A(n_2548),
.Y(n_3557)
);

BUFx6f_ASAP7_75t_SL g3558 ( 
.A(n_2784),
.Y(n_3558)
);

BUFx6f_ASAP7_75t_L g3559 ( 
.A(n_2702),
.Y(n_3559)
);

AOI21x1_ASAP7_75t_L g3560 ( 
.A1(n_2574),
.A2(n_471),
.B(n_472),
.Y(n_3560)
);

INVx2_ASAP7_75t_L g3561 ( 
.A(n_2885),
.Y(n_3561)
);

NAND2xp5_ASAP7_75t_L g3562 ( 
.A(n_2831),
.B(n_471),
.Y(n_3562)
);

INVx2_ASAP7_75t_L g3563 ( 
.A(n_2885),
.Y(n_3563)
);

NOR2xp33_ASAP7_75t_L g3564 ( 
.A(n_2890),
.B(n_473),
.Y(n_3564)
);

NAND2xp5_ASAP7_75t_L g3565 ( 
.A(n_2844),
.B(n_473),
.Y(n_3565)
);

NOR2x1p5_ASAP7_75t_L g3566 ( 
.A(n_2851),
.B(n_473),
.Y(n_3566)
);

OR2x2_ASAP7_75t_L g3567 ( 
.A(n_2646),
.B(n_474),
.Y(n_3567)
);

NOR2xp33_ASAP7_75t_L g3568 ( 
.A(n_2847),
.B(n_474),
.Y(n_3568)
);

OAI22xp33_ASAP7_75t_L g3569 ( 
.A1(n_3044),
.A2(n_476),
.B1(n_474),
.B2(n_475),
.Y(n_3569)
);

BUFx2_ASAP7_75t_L g3570 ( 
.A(n_2769),
.Y(n_3570)
);

INVx1_ASAP7_75t_L g3571 ( 
.A(n_2818),
.Y(n_3571)
);

NOR2xp33_ASAP7_75t_L g3572 ( 
.A(n_2556),
.B(n_475),
.Y(n_3572)
);

A2O1A1Ixp33_ASAP7_75t_L g3573 ( 
.A1(n_3097),
.A2(n_478),
.B(n_476),
.C(n_477),
.Y(n_3573)
);

NAND2xp5_ASAP7_75t_L g3574 ( 
.A(n_2860),
.B(n_476),
.Y(n_3574)
);

INVxp67_ASAP7_75t_L g3575 ( 
.A(n_2728),
.Y(n_3575)
);

A2O1A1Ixp33_ASAP7_75t_L g3576 ( 
.A1(n_3143),
.A2(n_479),
.B(n_477),
.C(n_478),
.Y(n_3576)
);

NAND2xp5_ASAP7_75t_L g3577 ( 
.A(n_2696),
.B(n_477),
.Y(n_3577)
);

INVx2_ASAP7_75t_L g3578 ( 
.A(n_2739),
.Y(n_3578)
);

OAI21xp5_ASAP7_75t_L g3579 ( 
.A1(n_2790),
.A2(n_478),
.B(n_479),
.Y(n_3579)
);

HB1xp67_ASAP7_75t_L g3580 ( 
.A(n_2872),
.Y(n_3580)
);

NAND2xp5_ASAP7_75t_SL g3581 ( 
.A(n_2598),
.B(n_728),
.Y(n_3581)
);

NOR2xp33_ASAP7_75t_R g3582 ( 
.A(n_2853),
.B(n_479),
.Y(n_3582)
);

NAND2xp5_ASAP7_75t_L g3583 ( 
.A(n_2697),
.B(n_480),
.Y(n_3583)
);

O2A1O1Ixp33_ASAP7_75t_L g3584 ( 
.A1(n_2874),
.A2(n_3148),
.B(n_3154),
.C(n_3147),
.Y(n_3584)
);

AOI21xp5_ASAP7_75t_L g3585 ( 
.A1(n_2537),
.A2(n_480),
.B(n_481),
.Y(n_3585)
);

INVx4_ASAP7_75t_L g3586 ( 
.A(n_2729),
.Y(n_3586)
);

NOR2xp33_ASAP7_75t_L g3587 ( 
.A(n_2820),
.B(n_480),
.Y(n_3587)
);

INVx2_ASAP7_75t_L g3588 ( 
.A(n_2610),
.Y(n_3588)
);

NAND2xp5_ASAP7_75t_L g3589 ( 
.A(n_2637),
.B(n_2542),
.Y(n_3589)
);

AOI21xp5_ASAP7_75t_L g3590 ( 
.A1(n_2898),
.A2(n_481),
.B(n_482),
.Y(n_3590)
);

HB1xp67_ASAP7_75t_L g3591 ( 
.A(n_2855),
.Y(n_3591)
);

INVx1_ASAP7_75t_L g3592 ( 
.A(n_2856),
.Y(n_3592)
);

INVx1_ASAP7_75t_L g3593 ( 
.A(n_2857),
.Y(n_3593)
);

AOI21xp5_ASAP7_75t_L g3594 ( 
.A1(n_2536),
.A2(n_481),
.B(n_482),
.Y(n_3594)
);

OAI22xp5_ASAP7_75t_L g3595 ( 
.A1(n_3081),
.A2(n_485),
.B1(n_483),
.B2(n_484),
.Y(n_3595)
);

O2A1O1Ixp33_ASAP7_75t_L g3596 ( 
.A1(n_2950),
.A2(n_486),
.B(n_484),
.C(n_485),
.Y(n_3596)
);

BUFx6f_ASAP7_75t_L g3597 ( 
.A(n_2702),
.Y(n_3597)
);

NOR2xp33_ASAP7_75t_L g3598 ( 
.A(n_2891),
.B(n_484),
.Y(n_3598)
);

NAND2xp5_ASAP7_75t_L g3599 ( 
.A(n_2544),
.B(n_485),
.Y(n_3599)
);

NAND2xp5_ASAP7_75t_SL g3600 ( 
.A(n_3057),
.B(n_729),
.Y(n_3600)
);

BUFx2_ASAP7_75t_L g3601 ( 
.A(n_2853),
.Y(n_3601)
);

OR2x6_ASAP7_75t_L g3602 ( 
.A(n_2938),
.B(n_487),
.Y(n_3602)
);

AOI21xp5_ASAP7_75t_L g3603 ( 
.A1(n_2536),
.A2(n_487),
.B(n_488),
.Y(n_3603)
);

AOI22xp5_ASAP7_75t_L g3604 ( 
.A1(n_3069),
.A2(n_489),
.B1(n_487),
.B2(n_488),
.Y(n_3604)
);

OAI21xp5_ASAP7_75t_L g3605 ( 
.A1(n_2695),
.A2(n_489),
.B(n_490),
.Y(n_3605)
);

INVx2_ASAP7_75t_L g3606 ( 
.A(n_3088),
.Y(n_3606)
);

INVxp67_ASAP7_75t_L g3607 ( 
.A(n_2828),
.Y(n_3607)
);

INVx2_ASAP7_75t_L g3608 ( 
.A(n_2623),
.Y(n_3608)
);

A2O1A1Ixp33_ASAP7_75t_L g3609 ( 
.A1(n_2865),
.A2(n_492),
.B(n_490),
.C(n_491),
.Y(n_3609)
);

OAI22xp5_ASAP7_75t_L g3610 ( 
.A1(n_3157),
.A2(n_492),
.B1(n_490),
.B2(n_491),
.Y(n_3610)
);

OR2x2_ASAP7_75t_L g3611 ( 
.A(n_2664),
.B(n_2829),
.Y(n_3611)
);

AOI21xp5_ASAP7_75t_L g3612 ( 
.A1(n_2624),
.A2(n_492),
.B(n_493),
.Y(n_3612)
);

INVxp67_ASAP7_75t_SL g3613 ( 
.A(n_2702),
.Y(n_3613)
);

INVx1_ASAP7_75t_L g3614 ( 
.A(n_2880),
.Y(n_3614)
);

INVx1_ASAP7_75t_L g3615 ( 
.A(n_2615),
.Y(n_3615)
);

INVx2_ASAP7_75t_L g3616 ( 
.A(n_2660),
.Y(n_3616)
);

NOR3xp33_ASAP7_75t_SL g3617 ( 
.A(n_2920),
.B(n_493),
.C(n_494),
.Y(n_3617)
);

AOI21xp5_ASAP7_75t_L g3618 ( 
.A1(n_2550),
.A2(n_494),
.B(n_495),
.Y(n_3618)
);

INVx1_ASAP7_75t_L g3619 ( 
.A(n_2889),
.Y(n_3619)
);

AOI21xp5_ASAP7_75t_L g3620 ( 
.A1(n_2550),
.A2(n_494),
.B(n_496),
.Y(n_3620)
);

OAI22xp5_ASAP7_75t_L g3621 ( 
.A1(n_2606),
.A2(n_499),
.B1(n_497),
.B2(n_498),
.Y(n_3621)
);

INVx5_ASAP7_75t_L g3622 ( 
.A(n_2729),
.Y(n_3622)
);

AOI21xp5_ASAP7_75t_L g3623 ( 
.A1(n_2585),
.A2(n_497),
.B(n_498),
.Y(n_3623)
);

O2A1O1Ixp33_ASAP7_75t_L g3624 ( 
.A1(n_3103),
.A2(n_500),
.B(n_497),
.C(n_499),
.Y(n_3624)
);

NAND2xp5_ASAP7_75t_L g3625 ( 
.A(n_2569),
.B(n_500),
.Y(n_3625)
);

AOI21xp5_ASAP7_75t_L g3626 ( 
.A1(n_2669),
.A2(n_500),
.B(n_501),
.Y(n_3626)
);

OR2x2_ASAP7_75t_L g3627 ( 
.A(n_2808),
.B(n_501),
.Y(n_3627)
);

NAND2xp5_ASAP7_75t_L g3628 ( 
.A(n_2578),
.B(n_501),
.Y(n_3628)
);

AOI21xp5_ASAP7_75t_L g3629 ( 
.A1(n_2776),
.A2(n_502),
.B(n_503),
.Y(n_3629)
);

INVx2_ASAP7_75t_L g3630 ( 
.A(n_2787),
.Y(n_3630)
);

O2A1O1Ixp33_ASAP7_75t_L g3631 ( 
.A1(n_2902),
.A2(n_504),
.B(n_502),
.C(n_503),
.Y(n_3631)
);

HB1xp67_ASAP7_75t_L g3632 ( 
.A(n_2746),
.Y(n_3632)
);

AO22x1_ASAP7_75t_L g3633 ( 
.A1(n_2709),
.A2(n_506),
.B1(n_504),
.B2(n_505),
.Y(n_3633)
);

NAND2xp5_ASAP7_75t_SL g3634 ( 
.A(n_2657),
.B(n_730),
.Y(n_3634)
);

OAI22x1_ASAP7_75t_L g3635 ( 
.A1(n_3071),
.A2(n_507),
.B1(n_505),
.B2(n_506),
.Y(n_3635)
);

O2A1O1Ixp33_ASAP7_75t_L g3636 ( 
.A1(n_2925),
.A2(n_507),
.B(n_505),
.C(n_506),
.Y(n_3636)
);

O2A1O1Ixp33_ASAP7_75t_L g3637 ( 
.A1(n_2927),
.A2(n_510),
.B(n_508),
.C(n_509),
.Y(n_3637)
);

NAND2xp5_ASAP7_75t_L g3638 ( 
.A(n_2580),
.B(n_508),
.Y(n_3638)
);

NOR2xp33_ASAP7_75t_L g3639 ( 
.A(n_2895),
.B(n_509),
.Y(n_3639)
);

NOR2xp67_ASAP7_75t_L g3640 ( 
.A(n_2920),
.B(n_510),
.Y(n_3640)
);

NOR3xp33_ASAP7_75t_SL g3641 ( 
.A(n_2755),
.B(n_510),
.C(n_511),
.Y(n_3641)
);

A2O1A1Ixp33_ASAP7_75t_SL g3642 ( 
.A1(n_2972),
.A2(n_513),
.B(n_511),
.C(n_512),
.Y(n_3642)
);

AOI21xp5_ASAP7_75t_L g3643 ( 
.A1(n_2583),
.A2(n_512),
.B(n_513),
.Y(n_3643)
);

HB1xp67_ASAP7_75t_L g3644 ( 
.A(n_2676),
.Y(n_3644)
);

AOI21xp5_ASAP7_75t_L g3645 ( 
.A1(n_2842),
.A2(n_514),
.B(n_515),
.Y(n_3645)
);

INVxp67_ASAP7_75t_SL g3646 ( 
.A(n_2954),
.Y(n_3646)
);

A2O1A1Ixp33_ASAP7_75t_L g3647 ( 
.A1(n_2655),
.A2(n_516),
.B(n_514),
.C(n_515),
.Y(n_3647)
);

BUFx2_ASAP7_75t_L g3648 ( 
.A(n_2996),
.Y(n_3648)
);

BUFx6f_ASAP7_75t_L g3649 ( 
.A(n_2954),
.Y(n_3649)
);

CKINVDCx14_ASAP7_75t_R g3650 ( 
.A(n_2590),
.Y(n_3650)
);

NAND2xp5_ASAP7_75t_L g3651 ( 
.A(n_2658),
.B(n_515),
.Y(n_3651)
);

BUFx2_ASAP7_75t_L g3652 ( 
.A(n_3010),
.Y(n_3652)
);

NAND2xp5_ASAP7_75t_L g3653 ( 
.A(n_2659),
.B(n_516),
.Y(n_3653)
);

BUFx2_ASAP7_75t_L g3654 ( 
.A(n_3011),
.Y(n_3654)
);

NOR2xp33_ASAP7_75t_L g3655 ( 
.A(n_2593),
.B(n_517),
.Y(n_3655)
);

CKINVDCx20_ASAP7_75t_R g3656 ( 
.A(n_2712),
.Y(n_3656)
);

BUFx3_ASAP7_75t_L g3657 ( 
.A(n_2892),
.Y(n_3657)
);

HB1xp67_ASAP7_75t_L g3658 ( 
.A(n_2714),
.Y(n_3658)
);

BUFx2_ASAP7_75t_SL g3659 ( 
.A(n_2835),
.Y(n_3659)
);

NAND2xp5_ASAP7_75t_L g3660 ( 
.A(n_2622),
.B(n_517),
.Y(n_3660)
);

INVx2_ASAP7_75t_L g3661 ( 
.A(n_2854),
.Y(n_3661)
);

INVx1_ASAP7_75t_L g3662 ( 
.A(n_2897),
.Y(n_3662)
);

BUFx2_ASAP7_75t_L g3663 ( 
.A(n_3061),
.Y(n_3663)
);

AND2x4_ASAP7_75t_L g3664 ( 
.A(n_2723),
.B(n_517),
.Y(n_3664)
);

NAND2xp5_ASAP7_75t_SL g3665 ( 
.A(n_2954),
.B(n_3016),
.Y(n_3665)
);

NAND2xp5_ASAP7_75t_SL g3666 ( 
.A(n_3016),
.B(n_730),
.Y(n_3666)
);

A2O1A1Ixp33_ASAP7_75t_L g3667 ( 
.A1(n_2816),
.A2(n_520),
.B(n_518),
.C(n_519),
.Y(n_3667)
);

NOR2xp33_ASAP7_75t_L g3668 ( 
.A(n_2878),
.B(n_518),
.Y(n_3668)
);

OR2x2_ASAP7_75t_L g3669 ( 
.A(n_2810),
.B(n_518),
.Y(n_3669)
);

O2A1O1Ixp33_ASAP7_75t_L g3670 ( 
.A1(n_2956),
.A2(n_521),
.B(n_519),
.C(n_520),
.Y(n_3670)
);

O2A1O1Ixp33_ASAP7_75t_L g3671 ( 
.A1(n_2959),
.A2(n_523),
.B(n_521),
.C(n_522),
.Y(n_3671)
);

A2O1A1Ixp33_ASAP7_75t_L g3672 ( 
.A1(n_2861),
.A2(n_2805),
.B(n_2815),
.C(n_2866),
.Y(n_3672)
);

NAND2xp5_ASAP7_75t_L g3673 ( 
.A(n_3129),
.B(n_521),
.Y(n_3673)
);

AOI21xp5_ASAP7_75t_L g3674 ( 
.A1(n_3016),
.A2(n_522),
.B(n_523),
.Y(n_3674)
);

NAND2xp5_ASAP7_75t_SL g3675 ( 
.A(n_3066),
.B(n_731),
.Y(n_3675)
);

NAND2xp5_ASAP7_75t_L g3676 ( 
.A(n_2732),
.B(n_522),
.Y(n_3676)
);

AND2x2_ASAP7_75t_L g3677 ( 
.A(n_2740),
.B(n_2698),
.Y(n_3677)
);

NOR2xp33_ASAP7_75t_L g3678 ( 
.A(n_2850),
.B(n_523),
.Y(n_3678)
);

A2O1A1Ixp33_ASAP7_75t_SL g3679 ( 
.A1(n_3085),
.A2(n_526),
.B(n_524),
.C(n_525),
.Y(n_3679)
);

O2A1O1Ixp33_ASAP7_75t_L g3680 ( 
.A1(n_2963),
.A2(n_526),
.B(n_524),
.C(n_525),
.Y(n_3680)
);

INVx2_ASAP7_75t_L g3681 ( 
.A(n_2834),
.Y(n_3681)
);

CKINVDCx8_ASAP7_75t_R g3682 ( 
.A(n_2893),
.Y(n_3682)
);

CKINVDCx5p33_ASAP7_75t_R g3683 ( 
.A(n_2812),
.Y(n_3683)
);

OAI22xp5_ASAP7_75t_L g3684 ( 
.A1(n_2723),
.A2(n_2736),
.B1(n_3003),
.B2(n_2974),
.Y(n_3684)
);

INVx1_ASAP7_75t_L g3685 ( 
.A(n_2595),
.Y(n_3685)
);

NOR2x1_ASAP7_75t_L g3686 ( 
.A(n_2752),
.B(n_524),
.Y(n_3686)
);

AOI21xp5_ASAP7_75t_L g3687 ( 
.A1(n_3066),
.A2(n_526),
.B(n_527),
.Y(n_3687)
);

BUFx6f_ASAP7_75t_L g3688 ( 
.A(n_3066),
.Y(n_3688)
);

A2O1A1Ixp33_ASAP7_75t_L g3689 ( 
.A1(n_2863),
.A2(n_529),
.B(n_527),
.C(n_528),
.Y(n_3689)
);

OAI21x1_ASAP7_75t_L g3690 ( 
.A1(n_3189),
.A2(n_2683),
.B(n_2671),
.Y(n_3690)
);

AO32x2_ASAP7_75t_L g3691 ( 
.A1(n_3181),
.A2(n_2552),
.A3(n_2943),
.B1(n_3122),
.B2(n_3107),
.Y(n_3691)
);

AOI21xp5_ASAP7_75t_L g3692 ( 
.A1(n_3464),
.A2(n_3116),
.B(n_3107),
.Y(n_3692)
);

INVx1_ASAP7_75t_L g3693 ( 
.A(n_3160),
.Y(n_3693)
);

AOI21xp5_ASAP7_75t_L g3694 ( 
.A1(n_3468),
.A2(n_3116),
.B(n_3111),
.Y(n_3694)
);

OAI21x1_ASAP7_75t_L g3695 ( 
.A1(n_3532),
.A2(n_2685),
.B(n_2745),
.Y(n_3695)
);

BUFx6f_ASAP7_75t_L g3696 ( 
.A(n_3243),
.Y(n_3696)
);

BUFx6f_ASAP7_75t_L g3697 ( 
.A(n_3192),
.Y(n_3697)
);

O2A1O1Ixp33_ASAP7_75t_L g3698 ( 
.A1(n_3452),
.A2(n_2801),
.B(n_2875),
.C(n_2644),
.Y(n_3698)
);

AOI21x1_ASAP7_75t_L g3699 ( 
.A1(n_3352),
.A2(n_3111),
.B(n_2986),
.Y(n_3699)
);

BUFx4f_ASAP7_75t_L g3700 ( 
.A(n_3366),
.Y(n_3700)
);

AOI21xp5_ASAP7_75t_L g3701 ( 
.A1(n_3531),
.A2(n_3116),
.B(n_3115),
.Y(n_3701)
);

AND2x2_ASAP7_75t_L g3702 ( 
.A(n_3370),
.B(n_2894),
.Y(n_3702)
);

CKINVDCx20_ASAP7_75t_R g3703 ( 
.A(n_3162),
.Y(n_3703)
);

NAND2xp5_ASAP7_75t_L g3704 ( 
.A(n_3203),
.B(n_2586),
.Y(n_3704)
);

AOI21xp5_ASAP7_75t_L g3705 ( 
.A1(n_3672),
.A2(n_3115),
.B(n_2986),
.Y(n_3705)
);

HB1xp67_ASAP7_75t_L g3706 ( 
.A(n_3256),
.Y(n_3706)
);

AOI22xp33_ASAP7_75t_L g3707 ( 
.A1(n_3419),
.A2(n_2750),
.B1(n_2736),
.B2(n_2699),
.Y(n_3707)
);

OAI22xp5_ASAP7_75t_L g3708 ( 
.A1(n_3287),
.A2(n_2682),
.B1(n_2786),
.B2(n_3121),
.Y(n_3708)
);

OA21x2_ASAP7_75t_L g3709 ( 
.A1(n_3412),
.A2(n_3126),
.B(n_3121),
.Y(n_3709)
);

AOI21xp5_ASAP7_75t_L g3710 ( 
.A1(n_3685),
.A2(n_3126),
.B(n_3158),
.Y(n_3710)
);

AOI21x1_ASAP7_75t_L g3711 ( 
.A1(n_3172),
.A2(n_2632),
.B(n_2629),
.Y(n_3711)
);

OA21x2_ASAP7_75t_L g3712 ( 
.A1(n_3648),
.A2(n_3140),
.B(n_3089),
.Y(n_3712)
);

OAI21xp5_ASAP7_75t_L g3713 ( 
.A1(n_3483),
.A2(n_2772),
.B(n_2741),
.Y(n_3713)
);

AND2x4_ASAP7_75t_L g3714 ( 
.A(n_3287),
.B(n_2840),
.Y(n_3714)
);

BUFx6f_ASAP7_75t_L g3715 ( 
.A(n_3218),
.Y(n_3715)
);

OA21x2_ASAP7_75t_L g3716 ( 
.A1(n_3652),
.A2(n_3146),
.B(n_2643),
.Y(n_3716)
);

AOI21xp5_ASAP7_75t_L g3717 ( 
.A1(n_3684),
.A2(n_2717),
.B(n_2597),
.Y(n_3717)
);

AND2x2_ASAP7_75t_L g3718 ( 
.A(n_3280),
.B(n_528),
.Y(n_3718)
);

OA21x2_ASAP7_75t_L g3719 ( 
.A1(n_3654),
.A2(n_2639),
.B(n_2916),
.Y(n_3719)
);

OAI21x1_ASAP7_75t_L g3720 ( 
.A1(n_3665),
.A2(n_2868),
.B(n_2883),
.Y(n_3720)
);

NAND2xp5_ASAP7_75t_SL g3721 ( 
.A(n_3287),
.B(n_2765),
.Y(n_3721)
);

AOI21xp5_ASAP7_75t_L g3722 ( 
.A1(n_3548),
.A2(n_2584),
.B(n_2917),
.Y(n_3722)
);

INVx2_ASAP7_75t_L g3723 ( 
.A(n_3232),
.Y(n_3723)
);

O2A1O1Ixp33_ASAP7_75t_L g3724 ( 
.A1(n_3444),
.A2(n_2896),
.B(n_2763),
.C(n_2800),
.Y(n_3724)
);

AOI21xp5_ASAP7_75t_L g3725 ( 
.A1(n_3588),
.A2(n_2921),
.B(n_2919),
.Y(n_3725)
);

OAI21x1_ASAP7_75t_L g3726 ( 
.A1(n_3382),
.A2(n_2779),
.B(n_2774),
.Y(n_3726)
);

OAI21xp33_ASAP7_75t_SL g3727 ( 
.A1(n_3640),
.A2(n_2946),
.B(n_2937),
.Y(n_3727)
);

AO31x2_ASAP7_75t_L g3728 ( 
.A1(n_3663),
.A2(n_2953),
.A3(n_2962),
.B(n_2951),
.Y(n_3728)
);

BUFx10_ASAP7_75t_L g3729 ( 
.A(n_3254),
.Y(n_3729)
);

AND2x2_ASAP7_75t_L g3730 ( 
.A(n_3290),
.B(n_529),
.Y(n_3730)
);

BUFx4f_ASAP7_75t_SL g3731 ( 
.A(n_3162),
.Y(n_3731)
);

AOI21xp5_ASAP7_75t_L g3732 ( 
.A1(n_3390),
.A2(n_2967),
.B(n_2966),
.Y(n_3732)
);

AOI21x1_ASAP7_75t_L g3733 ( 
.A1(n_3213),
.A2(n_2993),
.B(n_2992),
.Y(n_3733)
);

INVx1_ASAP7_75t_L g3734 ( 
.A(n_3166),
.Y(n_3734)
);

INVx2_ASAP7_75t_L g3735 ( 
.A(n_3233),
.Y(n_3735)
);

INVx1_ASAP7_75t_L g3736 ( 
.A(n_3167),
.Y(n_3736)
);

INVx2_ASAP7_75t_L g3737 ( 
.A(n_3513),
.Y(n_3737)
);

OAI21x1_ASAP7_75t_L g3738 ( 
.A1(n_3554),
.A2(n_2783),
.B(n_2781),
.Y(n_3738)
);

OAI21x1_ASAP7_75t_L g3739 ( 
.A1(n_3554),
.A2(n_2791),
.B(n_2788),
.Y(n_3739)
);

INVx1_ASAP7_75t_L g3740 ( 
.A(n_3180),
.Y(n_3740)
);

AOI221xp5_ASAP7_75t_L g3741 ( 
.A1(n_3187),
.A2(n_2848),
.B1(n_2864),
.B2(n_2765),
.C(n_2839),
.Y(n_3741)
);

BUFx2_ASAP7_75t_L g3742 ( 
.A(n_3418),
.Y(n_3742)
);

INVx1_ASAP7_75t_L g3743 ( 
.A(n_3239),
.Y(n_3743)
);

INVx2_ASAP7_75t_L g3744 ( 
.A(n_3314),
.Y(n_3744)
);

NAND2xp5_ASAP7_75t_L g3745 ( 
.A(n_3449),
.B(n_2798),
.Y(n_3745)
);

INVx3_ASAP7_75t_L g3746 ( 
.A(n_3188),
.Y(n_3746)
);

BUFx2_ASAP7_75t_L g3747 ( 
.A(n_3401),
.Y(n_3747)
);

AOI21xp5_ASAP7_75t_L g3748 ( 
.A1(n_3578),
.A2(n_3013),
.B(n_3007),
.Y(n_3748)
);

BUFx3_ASAP7_75t_L g3749 ( 
.A(n_3279),
.Y(n_3749)
);

AOI21xp5_ASAP7_75t_L g3750 ( 
.A1(n_3606),
.A2(n_3026),
.B(n_3025),
.Y(n_3750)
);

NAND2xp5_ASAP7_75t_L g3751 ( 
.A(n_3211),
.B(n_2876),
.Y(n_3751)
);

O2A1O1Ixp5_ASAP7_75t_L g3752 ( 
.A1(n_3634),
.A2(n_3036),
.B(n_3041),
.C(n_3030),
.Y(n_3752)
);

HB1xp67_ASAP7_75t_L g3753 ( 
.A(n_3348),
.Y(n_3753)
);

INVx1_ASAP7_75t_L g3754 ( 
.A(n_3248),
.Y(n_3754)
);

BUFx6f_ASAP7_75t_L g3755 ( 
.A(n_3171),
.Y(n_3755)
);

BUFx2_ASAP7_75t_L g3756 ( 
.A(n_3247),
.Y(n_3756)
);

AOI21xp5_ASAP7_75t_L g3757 ( 
.A1(n_3238),
.A2(n_3046),
.B(n_3045),
.Y(n_3757)
);

BUFx2_ASAP7_75t_L g3758 ( 
.A(n_3247),
.Y(n_3758)
);

OAI21xp33_ASAP7_75t_SL g3759 ( 
.A1(n_3686),
.A2(n_3053),
.B(n_3048),
.Y(n_3759)
);

OAI21x1_ASAP7_75t_L g3760 ( 
.A1(n_3195),
.A2(n_2797),
.B(n_3054),
.Y(n_3760)
);

AOI221x1_ASAP7_75t_L g3761 ( 
.A1(n_3173),
.A2(n_3076),
.B1(n_3092),
.B2(n_3091),
.C(n_3072),
.Y(n_3761)
);

NOR2xp33_ASAP7_75t_L g3762 ( 
.A(n_3682),
.B(n_2879),
.Y(n_3762)
);

OAI21x1_ASAP7_75t_L g3763 ( 
.A1(n_3267),
.A2(n_3094),
.B(n_3093),
.Y(n_3763)
);

INVx2_ASAP7_75t_L g3764 ( 
.A(n_3330),
.Y(n_3764)
);

AO32x2_ASAP7_75t_L g3765 ( 
.A1(n_3198),
.A2(n_2782),
.A3(n_3095),
.B1(n_3104),
.B2(n_3099),
.Y(n_3765)
);

CKINVDCx5p33_ASAP7_75t_R g3766 ( 
.A(n_3168),
.Y(n_3766)
);

AO31x2_ASAP7_75t_L g3767 ( 
.A1(n_3265),
.A2(n_3108),
.A3(n_3113),
.B(n_3105),
.Y(n_3767)
);

OAI21x1_ASAP7_75t_L g3768 ( 
.A1(n_3267),
.A2(n_3127),
.B(n_3114),
.Y(n_3768)
);

INVx1_ASAP7_75t_L g3769 ( 
.A(n_3257),
.Y(n_3769)
);

O2A1O1Ixp33_ASAP7_75t_L g3770 ( 
.A1(n_3349),
.A2(n_3258),
.B(n_3607),
.C(n_3299),
.Y(n_3770)
);

O2A1O1Ixp33_ASAP7_75t_L g3771 ( 
.A1(n_3489),
.A2(n_2888),
.B(n_2823),
.C(n_2782),
.Y(n_3771)
);

OAI21x1_ASAP7_75t_L g3772 ( 
.A1(n_3291),
.A2(n_3131),
.B(n_3128),
.Y(n_3772)
);

NOR2xp67_ASAP7_75t_L g3773 ( 
.A(n_3289),
.B(n_3135),
.Y(n_3773)
);

OAI22xp5_ASAP7_75t_L g3774 ( 
.A1(n_3362),
.A2(n_3138),
.B1(n_3145),
.B2(n_3137),
.Y(n_3774)
);

AND2x2_ASAP7_75t_L g3775 ( 
.A(n_3397),
.B(n_529),
.Y(n_3775)
);

CKINVDCx5p33_ASAP7_75t_R g3776 ( 
.A(n_3357),
.Y(n_3776)
);

OAI21xp5_ASAP7_75t_L g3777 ( 
.A1(n_3584),
.A2(n_3151),
.B(n_3149),
.Y(n_3777)
);

A2O1A1Ixp33_ASAP7_75t_L g3778 ( 
.A1(n_3495),
.A2(n_3153),
.B(n_3152),
.C(n_532),
.Y(n_3778)
);

AO31x2_ASAP7_75t_L g3779 ( 
.A1(n_3245),
.A2(n_533),
.A3(n_530),
.B(n_531),
.Y(n_3779)
);

BUFx6f_ASAP7_75t_L g3780 ( 
.A(n_3289),
.Y(n_3780)
);

AOI21xp5_ASAP7_75t_L g3781 ( 
.A1(n_3608),
.A2(n_530),
.B(n_533),
.Y(n_3781)
);

NOR2xp33_ASAP7_75t_L g3782 ( 
.A(n_3650),
.B(n_530),
.Y(n_3782)
);

NAND2x1_ASAP7_75t_L g3783 ( 
.A(n_3586),
.B(n_533),
.Y(n_3783)
);

AO31x2_ASAP7_75t_L g3784 ( 
.A1(n_3318),
.A2(n_536),
.A3(n_534),
.B(n_535),
.Y(n_3784)
);

NOR2xp33_ASAP7_75t_SL g3785 ( 
.A(n_3263),
.B(n_534),
.Y(n_3785)
);

NAND2xp5_ASAP7_75t_SL g3786 ( 
.A(n_3317),
.B(n_534),
.Y(n_3786)
);

NAND2xp5_ASAP7_75t_L g3787 ( 
.A(n_3294),
.B(n_3281),
.Y(n_3787)
);

NAND2xp5_ASAP7_75t_L g3788 ( 
.A(n_3283),
.B(n_535),
.Y(n_3788)
);

AOI221x1_ASAP7_75t_L g3789 ( 
.A1(n_3351),
.A2(n_537),
.B1(n_535),
.B2(n_536),
.C(n_538),
.Y(n_3789)
);

BUFx2_ASAP7_75t_L g3790 ( 
.A(n_3260),
.Y(n_3790)
);

OA21x2_ASAP7_75t_L g3791 ( 
.A1(n_3413),
.A2(n_538),
.B(n_539),
.Y(n_3791)
);

OAI22xp5_ASAP7_75t_L g3792 ( 
.A1(n_3317),
.A2(n_542),
.B1(n_540),
.B2(n_541),
.Y(n_3792)
);

OA21x2_ASAP7_75t_L g3793 ( 
.A1(n_3499),
.A2(n_540),
.B(n_541),
.Y(n_3793)
);

OAI21x1_ASAP7_75t_L g3794 ( 
.A1(n_3291),
.A2(n_544),
.B(n_543),
.Y(n_3794)
);

INVx1_ASAP7_75t_L g3795 ( 
.A(n_3315),
.Y(n_3795)
);

INVx1_ASAP7_75t_L g3796 ( 
.A(n_3321),
.Y(n_3796)
);

INVx1_ASAP7_75t_L g3797 ( 
.A(n_3325),
.Y(n_3797)
);

NAND2x1p5_ASAP7_75t_L g3798 ( 
.A(n_3317),
.B(n_540),
.Y(n_3798)
);

OAI21xp5_ASAP7_75t_L g3799 ( 
.A1(n_3165),
.A2(n_543),
.B(n_545),
.Y(n_3799)
);

INVx1_ASAP7_75t_L g3800 ( 
.A(n_3326),
.Y(n_3800)
);

INVxp67_ASAP7_75t_SL g3801 ( 
.A(n_3417),
.Y(n_3801)
);

BUFx6f_ASAP7_75t_L g3802 ( 
.A(n_3297),
.Y(n_3802)
);

OAI21x1_ASAP7_75t_L g3803 ( 
.A1(n_3214),
.A2(n_546),
.B(n_545),
.Y(n_3803)
);

OAI22x1_ASAP7_75t_L g3804 ( 
.A1(n_3336),
.A2(n_546),
.B1(n_543),
.B2(n_545),
.Y(n_3804)
);

NOR2x1_ASAP7_75t_R g3805 ( 
.A(n_3219),
.B(n_546),
.Y(n_3805)
);

AOI21xp5_ASAP7_75t_L g3806 ( 
.A1(n_3630),
.A2(n_547),
.B(n_548),
.Y(n_3806)
);

INVx1_ASAP7_75t_L g3807 ( 
.A(n_3331),
.Y(n_3807)
);

OAI21xp5_ASAP7_75t_L g3808 ( 
.A1(n_3170),
.A2(n_547),
.B(n_548),
.Y(n_3808)
);

NAND2xp5_ASAP7_75t_SL g3809 ( 
.A(n_3664),
.B(n_547),
.Y(n_3809)
);

NAND2xp5_ASAP7_75t_L g3810 ( 
.A(n_3332),
.B(n_548),
.Y(n_3810)
);

BUFx3_ASAP7_75t_L g3811 ( 
.A(n_3323),
.Y(n_3811)
);

AOI21xp5_ASAP7_75t_L g3812 ( 
.A1(n_3492),
.A2(n_549),
.B(n_550),
.Y(n_3812)
);

AOI21xp5_ASAP7_75t_L g3813 ( 
.A1(n_3511),
.A2(n_549),
.B(n_550),
.Y(n_3813)
);

AO21x1_ASAP7_75t_L g3814 ( 
.A1(n_3664),
.A2(n_550),
.B(n_551),
.Y(n_3814)
);

AOI21xp5_ASAP7_75t_L g3815 ( 
.A1(n_3524),
.A2(n_551),
.B(n_552),
.Y(n_3815)
);

INVx1_ASAP7_75t_L g3816 ( 
.A(n_3339),
.Y(n_3816)
);

AO31x2_ASAP7_75t_L g3817 ( 
.A1(n_3609),
.A2(n_553),
.A3(n_551),
.B(n_552),
.Y(n_3817)
);

AO31x2_ASAP7_75t_L g3818 ( 
.A1(n_3616),
.A2(n_554),
.A3(n_552),
.B(n_553),
.Y(n_3818)
);

AOI21xp33_ASAP7_75t_L g3819 ( 
.A1(n_3611),
.A2(n_553),
.B(n_554),
.Y(n_3819)
);

O2A1O1Ixp33_ASAP7_75t_L g3820 ( 
.A1(n_3501),
.A2(n_556),
.B(n_554),
.C(n_555),
.Y(n_3820)
);

NAND2xp33_ASAP7_75t_L g3821 ( 
.A(n_3507),
.B(n_555),
.Y(n_3821)
);

NOR2xp67_ASAP7_75t_SL g3822 ( 
.A(n_3429),
.B(n_555),
.Y(n_3822)
);

OAI21xp5_ASAP7_75t_L g3823 ( 
.A1(n_3334),
.A2(n_556),
.B(n_558),
.Y(n_3823)
);

BUFx12f_ASAP7_75t_L g3824 ( 
.A(n_3323),
.Y(n_3824)
);

NAND2xp5_ASAP7_75t_L g3825 ( 
.A(n_3341),
.B(n_556),
.Y(n_3825)
);

BUFx10_ASAP7_75t_L g3826 ( 
.A(n_3254),
.Y(n_3826)
);

INVx5_ASAP7_75t_L g3827 ( 
.A(n_3177),
.Y(n_3827)
);

O2A1O1Ixp33_ASAP7_75t_L g3828 ( 
.A1(n_3514),
.A2(n_560),
.B(n_558),
.C(n_559),
.Y(n_3828)
);

AOI21xp5_ASAP7_75t_L g3829 ( 
.A1(n_3642),
.A2(n_558),
.B(n_559),
.Y(n_3829)
);

INVx5_ASAP7_75t_L g3830 ( 
.A(n_3205),
.Y(n_3830)
);

AOI21xp5_ASAP7_75t_L g3831 ( 
.A1(n_3679),
.A2(n_559),
.B(n_560),
.Y(n_3831)
);

OAI21xp5_ASAP7_75t_L g3832 ( 
.A1(n_3540),
.A2(n_560),
.B(n_561),
.Y(n_3832)
);

AOI21xp5_ASAP7_75t_L g3833 ( 
.A1(n_3546),
.A2(n_561),
.B(n_562),
.Y(n_3833)
);

NOR2xp33_ASAP7_75t_L g3834 ( 
.A(n_3502),
.B(n_562),
.Y(n_3834)
);

NOR2xp33_ASAP7_75t_L g3835 ( 
.A(n_3656),
.B(n_563),
.Y(n_3835)
);

OAI21xp5_ASAP7_75t_L g3836 ( 
.A1(n_3183),
.A2(n_563),
.B(n_564),
.Y(n_3836)
);

INVx2_ASAP7_75t_L g3837 ( 
.A(n_3343),
.Y(n_3837)
);

A2O1A1Ixp33_ASAP7_75t_L g3838 ( 
.A1(n_3506),
.A2(n_3522),
.B(n_3636),
.C(n_3631),
.Y(n_3838)
);

OAI21x1_ASAP7_75t_L g3839 ( 
.A1(n_3350),
.A2(n_565),
.B(n_564),
.Y(n_3839)
);

NAND3xp33_ASAP7_75t_L g3840 ( 
.A(n_3242),
.B(n_3197),
.C(n_3264),
.Y(n_3840)
);

AOI22xp5_ASAP7_75t_L g3841 ( 
.A1(n_3683),
.A2(n_566),
.B1(n_563),
.B2(n_565),
.Y(n_3841)
);

OAI22xp5_ASAP7_75t_L g3842 ( 
.A1(n_3391),
.A2(n_3420),
.B1(n_3169),
.B2(n_3503),
.Y(n_3842)
);

OAI21x1_ASAP7_75t_L g3843 ( 
.A1(n_3613),
.A2(n_568),
.B(n_567),
.Y(n_3843)
);

CKINVDCx5p33_ASAP7_75t_R g3844 ( 
.A(n_3369),
.Y(n_3844)
);

HB1xp67_ASAP7_75t_L g3845 ( 
.A(n_3355),
.Y(n_3845)
);

NAND2xp5_ASAP7_75t_L g3846 ( 
.A(n_3363),
.B(n_566),
.Y(n_3846)
);

INVx1_ASAP7_75t_L g3847 ( 
.A(n_3552),
.Y(n_3847)
);

NAND2xp5_ASAP7_75t_L g3848 ( 
.A(n_3589),
.B(n_566),
.Y(n_3848)
);

A2O1A1Ixp33_ASAP7_75t_L g3849 ( 
.A1(n_3637),
.A2(n_569),
.B(n_567),
.C(n_568),
.Y(n_3849)
);

NAND2xp5_ASAP7_75t_L g3850 ( 
.A(n_3457),
.B(n_567),
.Y(n_3850)
);

AO31x2_ASAP7_75t_L g3851 ( 
.A1(n_3647),
.A2(n_571),
.A3(n_568),
.B(n_570),
.Y(n_3851)
);

O2A1O1Ixp33_ASAP7_75t_L g3852 ( 
.A1(n_3517),
.A2(n_3573),
.B(n_3576),
.C(n_3534),
.Y(n_3852)
);

INVx3_ASAP7_75t_L g3853 ( 
.A(n_3297),
.Y(n_3853)
);

INVx3_ASAP7_75t_L g3854 ( 
.A(n_3217),
.Y(n_3854)
);

CKINVDCx5p33_ASAP7_75t_R g3855 ( 
.A(n_3438),
.Y(n_3855)
);

NAND3xp33_ASAP7_75t_SL g3856 ( 
.A(n_3455),
.B(n_570),
.C(n_571),
.Y(n_3856)
);

OR2x6_ASAP7_75t_L g3857 ( 
.A(n_3229),
.B(n_3388),
.Y(n_3857)
);

OAI22xp5_ASAP7_75t_L g3858 ( 
.A1(n_3322),
.A2(n_574),
.B1(n_572),
.B2(n_573),
.Y(n_3858)
);

BUFx2_ASAP7_75t_L g3859 ( 
.A(n_3260),
.Y(n_3859)
);

NAND2xp5_ASAP7_75t_L g3860 ( 
.A(n_3462),
.B(n_572),
.Y(n_3860)
);

NAND2xp5_ASAP7_75t_L g3861 ( 
.A(n_3466),
.B(n_3372),
.Y(n_3861)
);

NAND2xp5_ASAP7_75t_L g3862 ( 
.A(n_3375),
.B(n_572),
.Y(n_3862)
);

AOI21xp5_ASAP7_75t_L g3863 ( 
.A1(n_3681),
.A2(n_573),
.B(n_574),
.Y(n_3863)
);

AOI22xp5_ASAP7_75t_L g3864 ( 
.A1(n_3575),
.A2(n_575),
.B1(n_573),
.B2(n_574),
.Y(n_3864)
);

AOI22xp5_ASAP7_75t_L g3865 ( 
.A1(n_3547),
.A2(n_578),
.B1(n_576),
.B2(n_577),
.Y(n_3865)
);

NOR2xp33_ASAP7_75t_L g3866 ( 
.A(n_3433),
.B(n_576),
.Y(n_3866)
);

OAI22xp33_ASAP7_75t_L g3867 ( 
.A1(n_3602),
.A2(n_578),
.B1(n_576),
.B2(n_577),
.Y(n_3867)
);

AO31x2_ASAP7_75t_L g3868 ( 
.A1(n_3615),
.A2(n_580),
.A3(n_577),
.B(n_579),
.Y(n_3868)
);

O2A1O1Ixp33_ASAP7_75t_L g3869 ( 
.A1(n_3285),
.A2(n_3427),
.B(n_3435),
.C(n_3432),
.Y(n_3869)
);

OAI21xp5_ASAP7_75t_L g3870 ( 
.A1(n_3677),
.A2(n_579),
.B(n_580),
.Y(n_3870)
);

A2O1A1Ixp33_ASAP7_75t_L g3871 ( 
.A1(n_3670),
.A2(n_582),
.B(n_579),
.C(n_581),
.Y(n_3871)
);

O2A1O1Ixp33_ASAP7_75t_L g3872 ( 
.A1(n_3223),
.A2(n_583),
.B(n_581),
.C(n_582),
.Y(n_3872)
);

OAI21xp5_ASAP7_75t_L g3873 ( 
.A1(n_3206),
.A2(n_581),
.B(n_583),
.Y(n_3873)
);

HB1xp67_ASAP7_75t_L g3874 ( 
.A(n_3216),
.Y(n_3874)
);

OAI21xp5_ASAP7_75t_L g3875 ( 
.A1(n_3221),
.A2(n_583),
.B(n_584),
.Y(n_3875)
);

BUFx2_ASAP7_75t_L g3876 ( 
.A(n_3398),
.Y(n_3876)
);

OAI21x1_ASAP7_75t_L g3877 ( 
.A1(n_3646),
.A2(n_584),
.B(n_585),
.Y(n_3877)
);

O2A1O1Ixp33_ASAP7_75t_L g3878 ( 
.A1(n_3329),
.A2(n_587),
.B(n_584),
.C(n_586),
.Y(n_3878)
);

OAI21x1_ASAP7_75t_L g3879 ( 
.A1(n_3561),
.A2(n_586),
.B(n_587),
.Y(n_3879)
);

INVx1_ASAP7_75t_L g3880 ( 
.A(n_3271),
.Y(n_3880)
);

AO31x2_ASAP7_75t_L g3881 ( 
.A1(n_3571),
.A2(n_590),
.A3(n_588),
.B(n_589),
.Y(n_3881)
);

AO31x2_ASAP7_75t_L g3882 ( 
.A1(n_3592),
.A2(n_590),
.A3(n_588),
.B(n_589),
.Y(n_3882)
);

OAI22xp5_ASAP7_75t_L g3883 ( 
.A1(n_3403),
.A2(n_592),
.B1(n_588),
.B2(n_591),
.Y(n_3883)
);

AOI21xp5_ASAP7_75t_L g3884 ( 
.A1(n_3393),
.A2(n_591),
.B(n_592),
.Y(n_3884)
);

AOI21xp5_ASAP7_75t_L g3885 ( 
.A1(n_3422),
.A2(n_591),
.B(n_592),
.Y(n_3885)
);

BUFx6f_ASAP7_75t_L g3886 ( 
.A(n_3344),
.Y(n_3886)
);

INVx2_ASAP7_75t_L g3887 ( 
.A(n_3273),
.Y(n_3887)
);

INVxp67_ASAP7_75t_SL g3888 ( 
.A(n_3202),
.Y(n_3888)
);

AO31x2_ASAP7_75t_L g3889 ( 
.A1(n_3593),
.A2(n_3523),
.A3(n_3563),
.B(n_3406),
.Y(n_3889)
);

OAI22xp5_ASAP7_75t_SL g3890 ( 
.A1(n_3602),
.A2(n_595),
.B1(n_593),
.B2(n_594),
.Y(n_3890)
);

AOI21xp5_ASAP7_75t_SL g3891 ( 
.A1(n_3586),
.A2(n_593),
.B(n_595),
.Y(n_3891)
);

INVx1_ASAP7_75t_L g3892 ( 
.A(n_3306),
.Y(n_3892)
);

BUFx10_ASAP7_75t_L g3893 ( 
.A(n_3220),
.Y(n_3893)
);

AOI22xp5_ASAP7_75t_L g3894 ( 
.A1(n_3409),
.A2(n_3411),
.B1(n_3655),
.B2(n_3568),
.Y(n_3894)
);

AND3x2_ASAP7_75t_L g3895 ( 
.A(n_3364),
.B(n_595),
.C(n_596),
.Y(n_3895)
);

INVx1_ASAP7_75t_SL g3896 ( 
.A(n_3498),
.Y(n_3896)
);

AOI221xp5_ASAP7_75t_SL g3897 ( 
.A1(n_3227),
.A2(n_598),
.B1(n_596),
.B2(n_597),
.C(n_599),
.Y(n_3897)
);

OAI22xp5_ASAP7_75t_L g3898 ( 
.A1(n_3566),
.A2(n_3261),
.B1(n_3374),
.B2(n_3536),
.Y(n_3898)
);

AOI21xp5_ASAP7_75t_SL g3899 ( 
.A1(n_3276),
.A2(n_597),
.B(n_598),
.Y(n_3899)
);

A2O1A1Ixp33_ASAP7_75t_L g3900 ( 
.A1(n_3671),
.A2(n_600),
.B(n_598),
.C(n_599),
.Y(n_3900)
);

AND2x6_ASAP7_75t_L g3901 ( 
.A(n_3543),
.B(n_599),
.Y(n_3901)
);

INVx1_ASAP7_75t_L g3902 ( 
.A(n_3313),
.Y(n_3902)
);

NOR2xp33_ASAP7_75t_L g3903 ( 
.A(n_3461),
.B(n_600),
.Y(n_3903)
);

OAI21x1_ASAP7_75t_L g3904 ( 
.A1(n_3560),
.A2(n_3661),
.B(n_3186),
.Y(n_3904)
);

NAND2x1_ASAP7_75t_L g3905 ( 
.A(n_3476),
.B(n_600),
.Y(n_3905)
);

AO31x2_ASAP7_75t_L g3906 ( 
.A1(n_3510),
.A2(n_603),
.A3(n_601),
.B(n_602),
.Y(n_3906)
);

AOI21xp5_ASAP7_75t_L g3907 ( 
.A1(n_3446),
.A2(n_601),
.B(n_602),
.Y(n_3907)
);

NOR2xp67_ASAP7_75t_L g3908 ( 
.A(n_3377),
.B(n_601),
.Y(n_3908)
);

AND2x2_ASAP7_75t_L g3909 ( 
.A(n_3454),
.B(n_602),
.Y(n_3909)
);

A2O1A1Ixp33_ASAP7_75t_L g3910 ( 
.A1(n_3680),
.A2(n_605),
.B(n_603),
.C(n_604),
.Y(n_3910)
);

BUFx3_ASAP7_75t_L g3911 ( 
.A(n_3269),
.Y(n_3911)
);

CKINVDCx11_ASAP7_75t_R g3912 ( 
.A(n_3371),
.Y(n_3912)
);

INVx2_ASAP7_75t_L g3913 ( 
.A(n_3161),
.Y(n_3913)
);

INVx2_ASAP7_75t_L g3914 ( 
.A(n_3164),
.Y(n_3914)
);

NAND2xp5_ASAP7_75t_L g3915 ( 
.A(n_3394),
.B(n_603),
.Y(n_3915)
);

INVx1_ASAP7_75t_L g3916 ( 
.A(n_3212),
.Y(n_3916)
);

INVxp67_ASAP7_75t_SL g3917 ( 
.A(n_3234),
.Y(n_3917)
);

A2O1A1Ixp33_ASAP7_75t_L g3918 ( 
.A1(n_3259),
.A2(n_606),
.B(n_604),
.C(n_605),
.Y(n_3918)
);

NOR2xp33_ASAP7_75t_SL g3919 ( 
.A(n_3269),
.B(n_3377),
.Y(n_3919)
);

INVx2_ASAP7_75t_L g3920 ( 
.A(n_3182),
.Y(n_3920)
);

AOI21xp5_ASAP7_75t_L g3921 ( 
.A1(n_3414),
.A2(n_604),
.B(n_605),
.Y(n_3921)
);

NAND2xp5_ASAP7_75t_L g3922 ( 
.A(n_3193),
.B(n_3474),
.Y(n_3922)
);

INVx1_ASAP7_75t_L g3923 ( 
.A(n_3224),
.Y(n_3923)
);

AOI21xp5_ASAP7_75t_L g3924 ( 
.A1(n_3520),
.A2(n_3304),
.B(n_3428),
.Y(n_3924)
);

INVx1_ASAP7_75t_L g3925 ( 
.A(n_3231),
.Y(n_3925)
);

NAND2xp5_ASAP7_75t_L g3926 ( 
.A(n_3478),
.B(n_3163),
.Y(n_3926)
);

AOI221x1_ASAP7_75t_L g3927 ( 
.A1(n_3244),
.A2(n_608),
.B1(n_606),
.B2(n_607),
.C(n_609),
.Y(n_3927)
);

INVx2_ASAP7_75t_L g3928 ( 
.A(n_3185),
.Y(n_3928)
);

OAI21x1_ASAP7_75t_L g3929 ( 
.A1(n_3434),
.A2(n_607),
.B(n_608),
.Y(n_3929)
);

INVx1_ASAP7_75t_L g3930 ( 
.A(n_3262),
.Y(n_3930)
);

INVx6_ASAP7_75t_L g3931 ( 
.A(n_3657),
.Y(n_3931)
);

OAI21x1_ASAP7_75t_L g3932 ( 
.A1(n_3434),
.A2(n_3537),
.B(n_3525),
.Y(n_3932)
);

AOI21xp5_ASAP7_75t_L g3933 ( 
.A1(n_3577),
.A2(n_609),
.B(n_610),
.Y(n_3933)
);

A2O1A1Ixp33_ASAP7_75t_L g3934 ( 
.A1(n_3207),
.A2(n_612),
.B(n_610),
.C(n_611),
.Y(n_3934)
);

NAND2xp5_ASAP7_75t_L g3935 ( 
.A(n_3519),
.B(n_3614),
.Y(n_3935)
);

AOI21xp5_ASAP7_75t_L g3936 ( 
.A1(n_3583),
.A2(n_610),
.B(n_611),
.Y(n_3936)
);

AOI22xp5_ASAP7_75t_L g3937 ( 
.A1(n_3564),
.A2(n_613),
.B1(n_611),
.B2(n_612),
.Y(n_3937)
);

NAND3xp33_ASAP7_75t_SL g3938 ( 
.A(n_3582),
.B(n_612),
.C(n_613),
.Y(n_3938)
);

OAI22xp5_ASAP7_75t_L g3939 ( 
.A1(n_3190),
.A2(n_615),
.B1(n_613),
.B2(n_614),
.Y(n_3939)
);

AO31x2_ASAP7_75t_L g3940 ( 
.A1(n_3689),
.A2(n_617),
.A3(n_614),
.B(n_616),
.Y(n_3940)
);

NOR2xp67_ASAP7_75t_L g3941 ( 
.A(n_3345),
.B(n_616),
.Y(n_3941)
);

A2O1A1Ixp33_ASAP7_75t_L g3942 ( 
.A1(n_3477),
.A2(n_618),
.B(n_616),
.C(n_617),
.Y(n_3942)
);

OR2x6_ASAP7_75t_L g3943 ( 
.A(n_3368),
.B(n_617),
.Y(n_3943)
);

NAND2xp5_ASAP7_75t_SL g3944 ( 
.A(n_3429),
.B(n_618),
.Y(n_3944)
);

AOI21xp5_ASAP7_75t_SL g3945 ( 
.A1(n_3278),
.A2(n_618),
.B(n_619),
.Y(n_3945)
);

NAND2xp5_ASAP7_75t_L g3946 ( 
.A(n_3424),
.B(n_619),
.Y(n_3946)
);

NAND2xp5_ASAP7_75t_L g3947 ( 
.A(n_3619),
.B(n_3662),
.Y(n_3947)
);

AOI22xp5_ASAP7_75t_L g3948 ( 
.A1(n_3572),
.A2(n_622),
.B1(n_620),
.B2(n_621),
.Y(n_3948)
);

AOI21xp5_ASAP7_75t_L g3949 ( 
.A1(n_3292),
.A2(n_620),
.B(n_621),
.Y(n_3949)
);

INVx2_ASAP7_75t_L g3950 ( 
.A(n_3191),
.Y(n_3950)
);

AOI21xp5_ASAP7_75t_L g3951 ( 
.A1(n_3633),
.A2(n_620),
.B(n_621),
.Y(n_3951)
);

INVx2_ASAP7_75t_L g3952 ( 
.A(n_3194),
.Y(n_3952)
);

BUFx10_ASAP7_75t_L g3953 ( 
.A(n_3558),
.Y(n_3953)
);

AOI21xp5_ASAP7_75t_L g3954 ( 
.A1(n_3651),
.A2(n_622),
.B(n_623),
.Y(n_3954)
);

OAI21x1_ASAP7_75t_L g3955 ( 
.A1(n_3525),
.A2(n_622),
.B(n_623),
.Y(n_3955)
);

AND2x2_ASAP7_75t_L g3956 ( 
.A(n_3196),
.B(n_623),
.Y(n_3956)
);

AOI21xp5_ASAP7_75t_L g3957 ( 
.A1(n_3653),
.A2(n_624),
.B(n_625),
.Y(n_3957)
);

OAI21xp5_ASAP7_75t_SL g3958 ( 
.A1(n_3338),
.A2(n_3302),
.B(n_3353),
.Y(n_3958)
);

AOI21xp5_ASAP7_75t_L g3959 ( 
.A1(n_3632),
.A2(n_624),
.B(n_625),
.Y(n_3959)
);

AOI21xp5_ASAP7_75t_L g3960 ( 
.A1(n_3538),
.A2(n_624),
.B(n_626),
.Y(n_3960)
);

INVx1_ASAP7_75t_L g3961 ( 
.A(n_3274),
.Y(n_3961)
);

BUFx2_ASAP7_75t_R g3962 ( 
.A(n_3659),
.Y(n_3962)
);

AOI21xp5_ASAP7_75t_L g3963 ( 
.A1(n_3493),
.A2(n_3530),
.B(n_3515),
.Y(n_3963)
);

OR2x2_ASAP7_75t_L g3964 ( 
.A(n_3407),
.B(n_626),
.Y(n_3964)
);

NAND2xp5_ASAP7_75t_SL g3965 ( 
.A(n_3429),
.B(n_626),
.Y(n_3965)
);

NAND2xp5_ASAP7_75t_L g3966 ( 
.A(n_3539),
.B(n_627),
.Y(n_3966)
);

INVx2_ASAP7_75t_SL g3967 ( 
.A(n_3556),
.Y(n_3967)
);

AOI21xp33_ASAP7_75t_SL g3968 ( 
.A1(n_3305),
.A2(n_627),
.B(n_628),
.Y(n_3968)
);

AOI21xp5_ASAP7_75t_L g3969 ( 
.A1(n_3660),
.A2(n_628),
.B(n_629),
.Y(n_3969)
);

AOI31xp67_ASAP7_75t_L g3970 ( 
.A1(n_3666),
.A2(n_3675),
.A3(n_3581),
.B(n_3545),
.Y(n_3970)
);

AND2x4_ASAP7_75t_L g3971 ( 
.A(n_3476),
.B(n_629),
.Y(n_3971)
);

OR2x2_ASAP7_75t_L g3972 ( 
.A(n_3356),
.B(n_629),
.Y(n_3972)
);

A2O1A1Ixp33_ASAP7_75t_L g3973 ( 
.A1(n_3387),
.A2(n_632),
.B(n_630),
.C(n_631),
.Y(n_3973)
);

NAND2xp5_ASAP7_75t_L g3974 ( 
.A(n_3307),
.B(n_630),
.Y(n_3974)
);

AOI21xp33_ASAP7_75t_L g3975 ( 
.A1(n_3591),
.A2(n_631),
.B(n_632),
.Y(n_3975)
);

AOI221x1_ASAP7_75t_L g3976 ( 
.A1(n_3504),
.A2(n_634),
.B1(n_631),
.B2(n_633),
.C(n_635),
.Y(n_3976)
);

AOI21xp5_ASAP7_75t_L g3977 ( 
.A1(n_3676),
.A2(n_633),
.B(n_634),
.Y(n_3977)
);

AOI22xp5_ASAP7_75t_L g3978 ( 
.A1(n_3333),
.A2(n_636),
.B1(n_633),
.B2(n_635),
.Y(n_3978)
);

AND2x4_ASAP7_75t_L g3979 ( 
.A(n_3486),
.B(n_635),
.Y(n_3979)
);

A2O1A1Ixp33_ASAP7_75t_L g3980 ( 
.A1(n_3311),
.A2(n_3618),
.B(n_3620),
.C(n_3585),
.Y(n_3980)
);

A2O1A1Ixp33_ASAP7_75t_L g3981 ( 
.A1(n_3465),
.A2(n_638),
.B(n_636),
.C(n_637),
.Y(n_3981)
);

NAND2xp5_ASAP7_75t_SL g3982 ( 
.A(n_3622),
.B(n_637),
.Y(n_3982)
);

INVx1_ASAP7_75t_L g3983 ( 
.A(n_3284),
.Y(n_3983)
);

BUFx2_ASAP7_75t_L g3984 ( 
.A(n_3486),
.Y(n_3984)
);

AO32x2_ASAP7_75t_L g3985 ( 
.A1(n_3312),
.A2(n_640),
.A3(n_638),
.B1(n_639),
.B2(n_641),
.Y(n_3985)
);

OAI21xp5_ASAP7_75t_L g3986 ( 
.A1(n_3222),
.A2(n_638),
.B(n_639),
.Y(n_3986)
);

AOI21x1_ASAP7_75t_L g3987 ( 
.A1(n_3580),
.A2(n_732),
.B(n_731),
.Y(n_3987)
);

BUFx6f_ASAP7_75t_L g3988 ( 
.A(n_3175),
.Y(n_3988)
);

INVx1_ASAP7_75t_L g3989 ( 
.A(n_3295),
.Y(n_3989)
);

INVx2_ASAP7_75t_SL g3990 ( 
.A(n_3456),
.Y(n_3990)
);

OAI21x1_ASAP7_75t_L g3991 ( 
.A1(n_3537),
.A2(n_639),
.B(n_640),
.Y(n_3991)
);

O2A1O1Ixp33_ASAP7_75t_L g3992 ( 
.A1(n_3235),
.A2(n_3482),
.B(n_3485),
.C(n_3458),
.Y(n_3992)
);

BUFx10_ASAP7_75t_L g3993 ( 
.A(n_3543),
.Y(n_3993)
);

AOI21xp33_ASAP7_75t_L g3994 ( 
.A1(n_3587),
.A2(n_641),
.B(n_642),
.Y(n_3994)
);

A2O1A1Ixp33_ASAP7_75t_L g3995 ( 
.A1(n_3445),
.A2(n_643),
.B(n_641),
.C(n_642),
.Y(n_3995)
);

A2O1A1Ixp33_ASAP7_75t_L g3996 ( 
.A1(n_3494),
.A2(n_644),
.B(n_642),
.C(n_643),
.Y(n_3996)
);

OAI21x1_ASAP7_75t_L g3997 ( 
.A1(n_3184),
.A2(n_644),
.B(n_645),
.Y(n_3997)
);

INVx5_ASAP7_75t_L g3998 ( 
.A(n_3622),
.Y(n_3998)
);

AOI21xp5_ASAP7_75t_L g3999 ( 
.A1(n_3175),
.A2(n_644),
.B(n_645),
.Y(n_3999)
);

OAI22xp5_ASAP7_75t_L g4000 ( 
.A1(n_3496),
.A2(n_648),
.B1(n_646),
.B2(n_647),
.Y(n_4000)
);

OAI22xp5_ASAP7_75t_L g4001 ( 
.A1(n_3396),
.A2(n_648),
.B1(n_646),
.B2(n_647),
.Y(n_4001)
);

OAI22xp33_ASAP7_75t_L g4002 ( 
.A1(n_3527),
.A2(n_648),
.B1(n_646),
.B2(n_647),
.Y(n_4002)
);

BUFx2_ASAP7_75t_L g4003 ( 
.A(n_3516),
.Y(n_4003)
);

INVx2_ASAP7_75t_L g4004 ( 
.A(n_3201),
.Y(n_4004)
);

AOI21xp5_ASAP7_75t_L g4005 ( 
.A1(n_3175),
.A2(n_649),
.B(n_650),
.Y(n_4005)
);

AOI221x1_ASAP7_75t_L g4006 ( 
.A1(n_3505),
.A2(n_651),
.B1(n_649),
.B2(n_650),
.C(n_652),
.Y(n_4006)
);

AOI21xp33_ASAP7_75t_L g4007 ( 
.A1(n_3644),
.A2(n_649),
.B(n_650),
.Y(n_4007)
);

NOR2xp33_ASAP7_75t_L g4008 ( 
.A(n_3365),
.B(n_651),
.Y(n_4008)
);

OR2x2_ASAP7_75t_L g4009 ( 
.A(n_3358),
.B(n_3373),
.Y(n_4009)
);

OAI21xp5_ASAP7_75t_L g4010 ( 
.A1(n_3228),
.A2(n_651),
.B(n_652),
.Y(n_4010)
);

NAND2xp5_ASAP7_75t_L g4011 ( 
.A(n_3678),
.B(n_652),
.Y(n_4011)
);

AO31x2_ASAP7_75t_L g4012 ( 
.A1(n_3328),
.A2(n_655),
.A3(n_653),
.B(n_654),
.Y(n_4012)
);

AOI221x1_ASAP7_75t_L g4013 ( 
.A1(n_3635),
.A2(n_655),
.B1(n_653),
.B2(n_654),
.C(n_656),
.Y(n_4013)
);

INVx2_ASAP7_75t_L g4014 ( 
.A(n_3204),
.Y(n_4014)
);

AOI21xp5_ASAP7_75t_L g4015 ( 
.A1(n_3178),
.A2(n_653),
.B(n_654),
.Y(n_4015)
);

BUFx2_ASAP7_75t_SL g4016 ( 
.A(n_3703),
.Y(n_4016)
);

CKINVDCx20_ASAP7_75t_R g4017 ( 
.A(n_3731),
.Y(n_4017)
);

INVx6_ASAP7_75t_L g4018 ( 
.A(n_3696),
.Y(n_4018)
);

AOI22xp33_ASAP7_75t_L g4019 ( 
.A1(n_3702),
.A2(n_3430),
.B1(n_3463),
.B2(n_3541),
.Y(n_4019)
);

INVx1_ASAP7_75t_L g4020 ( 
.A(n_3693),
.Y(n_4020)
);

CKINVDCx20_ASAP7_75t_R g4021 ( 
.A(n_3766),
.Y(n_4021)
);

AOI22xp33_ASAP7_75t_L g4022 ( 
.A1(n_3943),
.A2(n_3549),
.B1(n_3542),
.B2(n_3621),
.Y(n_4022)
);

BUFx6f_ASAP7_75t_L g4023 ( 
.A(n_3780),
.Y(n_4023)
);

CKINVDCx20_ASAP7_75t_R g4024 ( 
.A(n_3700),
.Y(n_4024)
);

BUFx2_ASAP7_75t_SL g4025 ( 
.A(n_3811),
.Y(n_4025)
);

AOI22xp5_ASAP7_75t_L g4026 ( 
.A1(n_3821),
.A2(n_3436),
.B1(n_3272),
.B2(n_3342),
.Y(n_4026)
);

INVx2_ASAP7_75t_L g4027 ( 
.A(n_3723),
.Y(n_4027)
);

BUFx3_ASAP7_75t_L g4028 ( 
.A(n_3780),
.Y(n_4028)
);

CKINVDCx5p33_ASAP7_75t_R g4029 ( 
.A(n_3824),
.Y(n_4029)
);

INVx1_ASAP7_75t_L g4030 ( 
.A(n_3734),
.Y(n_4030)
);

AOI22xp33_ASAP7_75t_L g4031 ( 
.A1(n_3943),
.A2(n_3447),
.B1(n_3460),
.B2(n_3450),
.Y(n_4031)
);

INVx1_ASAP7_75t_SL g4032 ( 
.A(n_3802),
.Y(n_4032)
);

INVx1_ASAP7_75t_L g4033 ( 
.A(n_3736),
.Y(n_4033)
);

AOI22xp33_ASAP7_75t_SL g4034 ( 
.A1(n_3901),
.A2(n_3380),
.B1(n_3443),
.B2(n_3658),
.Y(n_4034)
);

INVx8_ASAP7_75t_L g4035 ( 
.A(n_3696),
.Y(n_4035)
);

OAI22xp5_ASAP7_75t_L g4036 ( 
.A1(n_3707),
.A2(n_3617),
.B1(n_3641),
.B2(n_3199),
.Y(n_4036)
);

INVx2_ASAP7_75t_L g4037 ( 
.A(n_3735),
.Y(n_4037)
);

AOI22xp33_ASAP7_75t_SL g4038 ( 
.A1(n_3901),
.A2(n_3890),
.B1(n_3840),
.B2(n_3898),
.Y(n_4038)
);

INVx1_ASAP7_75t_L g4039 ( 
.A(n_3740),
.Y(n_4039)
);

OAI22xp33_ASAP7_75t_L g4040 ( 
.A1(n_3894),
.A2(n_3208),
.B1(n_3376),
.B2(n_3335),
.Y(n_4040)
);

AND2x2_ASAP7_75t_L g4041 ( 
.A(n_3718),
.B(n_3268),
.Y(n_4041)
);

AOI22xp33_ASAP7_75t_L g4042 ( 
.A1(n_3901),
.A2(n_3470),
.B1(n_3508),
.B2(n_3487),
.Y(n_4042)
);

INVx6_ASAP7_75t_L g4043 ( 
.A(n_3715),
.Y(n_4043)
);

INVx1_ASAP7_75t_SL g4044 ( 
.A(n_3802),
.Y(n_4044)
);

INVx6_ASAP7_75t_L g4045 ( 
.A(n_3715),
.Y(n_4045)
);

OAI22xp5_ASAP7_75t_L g4046 ( 
.A1(n_3721),
.A2(n_3404),
.B1(n_3425),
.B2(n_3399),
.Y(n_4046)
);

INVx1_ASAP7_75t_L g4047 ( 
.A(n_3743),
.Y(n_4047)
);

AOI22xp33_ASAP7_75t_L g4048 ( 
.A1(n_3938),
.A2(n_3174),
.B1(n_3400),
.B2(n_3392),
.Y(n_4048)
);

CKINVDCx5p33_ASAP7_75t_R g4049 ( 
.A(n_3776),
.Y(n_4049)
);

CKINVDCx20_ASAP7_75t_R g4050 ( 
.A(n_3844),
.Y(n_4050)
);

INVx6_ASAP7_75t_L g4051 ( 
.A(n_3893),
.Y(n_4051)
);

BUFx12f_ASAP7_75t_L g4052 ( 
.A(n_3855),
.Y(n_4052)
);

BUFx12f_ASAP7_75t_L g4053 ( 
.A(n_3953),
.Y(n_4053)
);

INVx2_ASAP7_75t_L g4054 ( 
.A(n_3737),
.Y(n_4054)
);

AOI22xp33_ASAP7_75t_L g4055 ( 
.A1(n_3856),
.A2(n_3668),
.B1(n_3610),
.B2(n_3595),
.Y(n_4055)
);

BUFx8_ASAP7_75t_L g4056 ( 
.A(n_3749),
.Y(n_4056)
);

INVx1_ASAP7_75t_L g4057 ( 
.A(n_3754),
.Y(n_4057)
);

AOI22xp5_ASAP7_75t_SL g4058 ( 
.A1(n_3746),
.A2(n_3319),
.B1(n_3346),
.B2(n_3200),
.Y(n_4058)
);

INVx2_ASAP7_75t_L g4059 ( 
.A(n_3887),
.Y(n_4059)
);

BUFx2_ASAP7_75t_L g4060 ( 
.A(n_3984),
.Y(n_4060)
);

BUFx8_ASAP7_75t_L g4061 ( 
.A(n_3755),
.Y(n_4061)
);

INVx1_ASAP7_75t_L g4062 ( 
.A(n_3769),
.Y(n_4062)
);

OAI22xp33_ASAP7_75t_L g4063 ( 
.A1(n_3785),
.A2(n_3604),
.B1(n_3516),
.B2(n_3288),
.Y(n_4063)
);

BUFx8_ASAP7_75t_SL g4064 ( 
.A(n_3857),
.Y(n_4064)
);

BUFx3_ASAP7_75t_L g4065 ( 
.A(n_3747),
.Y(n_4065)
);

OAI22xp5_ASAP7_75t_L g4066 ( 
.A1(n_3908),
.A2(n_3215),
.B1(n_3359),
.B2(n_3567),
.Y(n_4066)
);

INVx1_ASAP7_75t_L g4067 ( 
.A(n_3795),
.Y(n_4067)
);

AOI22xp33_ASAP7_75t_L g4068 ( 
.A1(n_3870),
.A2(n_3405),
.B1(n_3569),
.B2(n_3479),
.Y(n_4068)
);

BUFx6f_ASAP7_75t_L g4069 ( 
.A(n_3886),
.Y(n_4069)
);

BUFx6f_ASAP7_75t_L g4070 ( 
.A(n_3886),
.Y(n_4070)
);

INVx1_ASAP7_75t_L g4071 ( 
.A(n_3796),
.Y(n_4071)
);

AOI22xp33_ASAP7_75t_L g4072 ( 
.A1(n_3809),
.A2(n_3176),
.B1(n_3379),
.B2(n_3381),
.Y(n_4072)
);

INVx2_ASAP7_75t_L g4073 ( 
.A(n_3913),
.Y(n_4073)
);

BUFx3_ASAP7_75t_L g4074 ( 
.A(n_3853),
.Y(n_4074)
);

BUFx12f_ASAP7_75t_L g4075 ( 
.A(n_3857),
.Y(n_4075)
);

NAND2xp5_ASAP7_75t_L g4076 ( 
.A(n_3845),
.B(n_3787),
.Y(n_4076)
);

BUFx2_ASAP7_75t_L g4077 ( 
.A(n_4003),
.Y(n_4077)
);

CKINVDCx6p67_ASAP7_75t_R g4078 ( 
.A(n_3729),
.Y(n_4078)
);

BUFx10_ASAP7_75t_L g4079 ( 
.A(n_3755),
.Y(n_4079)
);

INVx2_ASAP7_75t_L g4080 ( 
.A(n_3914),
.Y(n_4080)
);

INVx6_ASAP7_75t_L g4081 ( 
.A(n_3827),
.Y(n_4081)
);

INVxp67_ASAP7_75t_SL g4082 ( 
.A(n_3753),
.Y(n_4082)
);

INVx2_ASAP7_75t_L g4083 ( 
.A(n_3920),
.Y(n_4083)
);

AOI22xp33_ASAP7_75t_L g4084 ( 
.A1(n_3762),
.A2(n_3579),
.B1(n_3673),
.B2(n_3442),
.Y(n_4084)
);

AOI22xp33_ASAP7_75t_SL g4085 ( 
.A1(n_3826),
.A2(n_3622),
.B1(n_3601),
.B2(n_3551),
.Y(n_4085)
);

INVx1_ASAP7_75t_L g4086 ( 
.A(n_3797),
.Y(n_4086)
);

CKINVDCx11_ASAP7_75t_R g4087 ( 
.A(n_3896),
.Y(n_4087)
);

BUFx3_ASAP7_75t_L g4088 ( 
.A(n_3931),
.Y(n_4088)
);

AOI22xp33_ASAP7_75t_L g4089 ( 
.A1(n_3774),
.A2(n_3521),
.B1(n_3600),
.B2(n_3179),
.Y(n_4089)
);

AOI22xp33_ASAP7_75t_L g4090 ( 
.A1(n_3912),
.A2(n_3250),
.B1(n_3639),
.B2(n_3598),
.Y(n_4090)
);

NAND2xp5_ASAP7_75t_L g4091 ( 
.A(n_3706),
.B(n_3441),
.Y(n_4091)
);

BUFx12f_ASAP7_75t_L g4092 ( 
.A(n_3742),
.Y(n_4092)
);

INVx3_ASAP7_75t_L g4093 ( 
.A(n_3911),
.Y(n_4093)
);

OAI22xp5_ASAP7_75t_L g4094 ( 
.A1(n_3962),
.A2(n_3605),
.B1(n_3667),
.B2(n_3360),
.Y(n_4094)
);

CKINVDCx20_ASAP7_75t_R g4095 ( 
.A(n_3931),
.Y(n_4095)
);

AOI22xp33_ASAP7_75t_SL g4096 ( 
.A1(n_3842),
.A2(n_3570),
.B1(n_3473),
.B2(n_3481),
.Y(n_4096)
);

BUFx2_ASAP7_75t_L g4097 ( 
.A(n_3756),
.Y(n_4097)
);

AND2x2_ASAP7_75t_L g4098 ( 
.A(n_3730),
.B(n_3209),
.Y(n_4098)
);

INVx1_ASAP7_75t_L g4099 ( 
.A(n_3800),
.Y(n_4099)
);

INVx1_ASAP7_75t_SL g4100 ( 
.A(n_3876),
.Y(n_4100)
);

INVx8_ASAP7_75t_L g4101 ( 
.A(n_3827),
.Y(n_4101)
);

AOI22xp33_ASAP7_75t_L g4102 ( 
.A1(n_3708),
.A2(n_3308),
.B1(n_3316),
.B2(n_3241),
.Y(n_4102)
);

CKINVDCx6p67_ASAP7_75t_R g4103 ( 
.A(n_3830),
.Y(n_4103)
);

OAI22x1_ASAP7_75t_L g4104 ( 
.A1(n_3782),
.A2(n_3459),
.B1(n_3475),
.B2(n_3437),
.Y(n_4104)
);

BUFx10_ASAP7_75t_L g4105 ( 
.A(n_3895),
.Y(n_4105)
);

BUFx3_ASAP7_75t_L g4106 ( 
.A(n_3830),
.Y(n_4106)
);

INVx2_ASAP7_75t_L g4107 ( 
.A(n_3928),
.Y(n_4107)
);

INVx6_ASAP7_75t_L g4108 ( 
.A(n_3993),
.Y(n_4108)
);

AOI22xp33_ASAP7_75t_SL g4109 ( 
.A1(n_3919),
.A2(n_3473),
.B1(n_3528),
.B2(n_3402),
.Y(n_4109)
);

BUFx12f_ASAP7_75t_L g4110 ( 
.A(n_3967),
.Y(n_4110)
);

INVx3_ASAP7_75t_L g4111 ( 
.A(n_3697),
.Y(n_4111)
);

INVx6_ASAP7_75t_L g4112 ( 
.A(n_3697),
.Y(n_4112)
);

INVx1_ASAP7_75t_L g4113 ( 
.A(n_3807),
.Y(n_4113)
);

AOI22xp33_ASAP7_75t_L g4114 ( 
.A1(n_3939),
.A2(n_3645),
.B1(n_3497),
.B2(n_3488),
.Y(n_4114)
);

CKINVDCx20_ASAP7_75t_R g4115 ( 
.A(n_3866),
.Y(n_4115)
);

BUFx2_ASAP7_75t_SL g4116 ( 
.A(n_3998),
.Y(n_4116)
);

INVx1_ASAP7_75t_L g4117 ( 
.A(n_3816),
.Y(n_4117)
);

OAI22xp5_ASAP7_75t_L g4118 ( 
.A1(n_3941),
.A2(n_3416),
.B1(n_3451),
.B2(n_3337),
.Y(n_4118)
);

NAND2xp5_ASAP7_75t_L g4119 ( 
.A(n_3861),
.B(n_3300),
.Y(n_4119)
);

BUFx12f_ASAP7_75t_L g4120 ( 
.A(n_3798),
.Y(n_4120)
);

CKINVDCx11_ASAP7_75t_R g4121 ( 
.A(n_3971),
.Y(n_4121)
);

AOI22xp33_ASAP7_75t_L g4122 ( 
.A1(n_4001),
.A2(n_3490),
.B1(n_3500),
.B2(n_3484),
.Y(n_4122)
);

INVx6_ASAP7_75t_L g4123 ( 
.A(n_3998),
.Y(n_4123)
);

OR2x2_ASAP7_75t_L g4124 ( 
.A(n_3964),
.B(n_3385),
.Y(n_4124)
);

INVx1_ASAP7_75t_L g4125 ( 
.A(n_3847),
.Y(n_4125)
);

AOI22xp33_ASAP7_75t_L g4126 ( 
.A1(n_3704),
.A2(n_4008),
.B1(n_3751),
.B2(n_3814),
.Y(n_4126)
);

AOI21xp5_ASAP7_75t_L g4127 ( 
.A1(n_3705),
.A2(n_3237),
.B(n_3178),
.Y(n_4127)
);

INVx1_ASAP7_75t_SL g4128 ( 
.A(n_3990),
.Y(n_4128)
);

OAI21xp5_ASAP7_75t_SL g4129 ( 
.A1(n_3958),
.A2(n_3367),
.B(n_3210),
.Y(n_4129)
);

AOI22xp33_ASAP7_75t_L g4130 ( 
.A1(n_3867),
.A2(n_3509),
.B1(n_3612),
.B2(n_3529),
.Y(n_4130)
);

INVx3_ASAP7_75t_L g4131 ( 
.A(n_3854),
.Y(n_4131)
);

AND2x2_ASAP7_75t_L g4132 ( 
.A(n_3775),
.B(n_3225),
.Y(n_4132)
);

BUFx10_ASAP7_75t_L g4133 ( 
.A(n_3903),
.Y(n_4133)
);

OAI21xp5_ASAP7_75t_SL g4134 ( 
.A1(n_3789),
.A2(n_3624),
.B(n_3596),
.Y(n_4134)
);

BUFx10_ASAP7_75t_L g4135 ( 
.A(n_3979),
.Y(n_4135)
);

NAND2x1p5_ASAP7_75t_L g4136 ( 
.A(n_3822),
.B(n_3528),
.Y(n_4136)
);

CKINVDCx11_ASAP7_75t_R g4137 ( 
.A(n_3805),
.Y(n_4137)
);

OAI21xp5_ASAP7_75t_L g4138 ( 
.A1(n_3770),
.A2(n_3590),
.B(n_3246),
.Y(n_4138)
);

OAI22xp33_ASAP7_75t_L g4139 ( 
.A1(n_3841),
.A2(n_3574),
.B1(n_3669),
.B2(n_3627),
.Y(n_4139)
);

AOI22xp33_ASAP7_75t_L g4140 ( 
.A1(n_3994),
.A2(n_3512),
.B1(n_3550),
.B2(n_3533),
.Y(n_4140)
);

AOI22xp33_ASAP7_75t_SL g4141 ( 
.A1(n_3801),
.A2(n_3565),
.B1(n_3562),
.B2(n_3599),
.Y(n_4141)
);

AOI22xp33_ASAP7_75t_L g4142 ( 
.A1(n_3834),
.A2(n_3629),
.B1(n_3555),
.B2(n_3518),
.Y(n_4142)
);

OR2x2_ASAP7_75t_L g4143 ( 
.A(n_3874),
.B(n_3226),
.Y(n_4143)
);

INVx2_ASAP7_75t_L g4144 ( 
.A(n_3950),
.Y(n_4144)
);

INVx1_ASAP7_75t_L g4145 ( 
.A(n_3744),
.Y(n_4145)
);

HB1xp67_ASAP7_75t_L g4146 ( 
.A(n_3758),
.Y(n_4146)
);

AOI22xp33_ASAP7_75t_L g4147 ( 
.A1(n_3956),
.A2(n_3230),
.B1(n_3240),
.B2(n_3236),
.Y(n_4147)
);

INVx1_ASAP7_75t_L g4148 ( 
.A(n_3764),
.Y(n_4148)
);

AOI22xp33_ASAP7_75t_SL g4149 ( 
.A1(n_3790),
.A2(n_3628),
.B1(n_3638),
.B2(n_3625),
.Y(n_4149)
);

BUFx6f_ASAP7_75t_L g4150 ( 
.A(n_3988),
.Y(n_4150)
);

OAI22xp33_ASAP7_75t_L g4151 ( 
.A1(n_3804),
.A2(n_3421),
.B1(n_3415),
.B2(n_3303),
.Y(n_4151)
);

INVx1_ASAP7_75t_SL g4152 ( 
.A(n_3909),
.Y(n_4152)
);

INVx2_ASAP7_75t_L g4153 ( 
.A(n_3952),
.Y(n_4153)
);

AOI22xp33_ASAP7_75t_L g4154 ( 
.A1(n_3974),
.A2(n_3252),
.B1(n_3253),
.B2(n_3249),
.Y(n_4154)
);

INVx1_ASAP7_75t_L g4155 ( 
.A(n_3837),
.Y(n_4155)
);

CKINVDCx6p67_ASAP7_75t_R g4156 ( 
.A(n_3859),
.Y(n_4156)
);

OAI21xp5_ASAP7_75t_SL g4157 ( 
.A1(n_3823),
.A2(n_3327),
.B(n_3643),
.Y(n_4157)
);

INVx1_ASAP7_75t_SL g4158 ( 
.A(n_3988),
.Y(n_4158)
);

INVx2_ASAP7_75t_L g4159 ( 
.A(n_4004),
.Y(n_4159)
);

INVx2_ASAP7_75t_L g4160 ( 
.A(n_4014),
.Y(n_4160)
);

AOI22xp5_ASAP7_75t_L g4161 ( 
.A1(n_4002),
.A2(n_3320),
.B1(n_3324),
.B2(n_3301),
.Y(n_4161)
);

BUFx3_ASAP7_75t_L g4162 ( 
.A(n_3880),
.Y(n_4162)
);

AOI22xp5_ASAP7_75t_L g4163 ( 
.A1(n_3835),
.A2(n_3544),
.B1(n_3553),
.B2(n_3526),
.Y(n_4163)
);

INVx2_ASAP7_75t_SL g4164 ( 
.A(n_3905),
.Y(n_4164)
);

AOI22xp33_ASAP7_75t_L g4165 ( 
.A1(n_3873),
.A2(n_3266),
.B1(n_3270),
.B2(n_3255),
.Y(n_4165)
);

INVx3_ASAP7_75t_L g4166 ( 
.A(n_3783),
.Y(n_4166)
);

AOI22xp33_ASAP7_75t_SL g4167 ( 
.A1(n_3888),
.A2(n_3237),
.B1(n_3251),
.B2(n_3178),
.Y(n_4167)
);

AOI22xp33_ASAP7_75t_SL g4168 ( 
.A1(n_3917),
.A2(n_3836),
.B1(n_3712),
.B2(n_3714),
.Y(n_4168)
);

AOI22xp33_ASAP7_75t_L g4169 ( 
.A1(n_3875),
.A2(n_3282),
.B1(n_3286),
.B2(n_3277),
.Y(n_4169)
);

INVx1_ASAP7_75t_L g4170 ( 
.A(n_3892),
.Y(n_4170)
);

INVx1_ASAP7_75t_L g4171 ( 
.A(n_3902),
.Y(n_4171)
);

INVx6_ASAP7_75t_L g4172 ( 
.A(n_4009),
.Y(n_4172)
);

AOI22xp33_ASAP7_75t_L g4173 ( 
.A1(n_3986),
.A2(n_3296),
.B1(n_3298),
.B2(n_3293),
.Y(n_4173)
);

BUFx8_ASAP7_75t_L g4174 ( 
.A(n_3985),
.Y(n_4174)
);

NAND2xp5_ASAP7_75t_L g4175 ( 
.A(n_3935),
.B(n_3386),
.Y(n_4175)
);

NAND2xp5_ASAP7_75t_L g4176 ( 
.A(n_3947),
.B(n_3439),
.Y(n_4176)
);

INVxp67_ASAP7_75t_SL g4177 ( 
.A(n_3932),
.Y(n_4177)
);

INVx1_ASAP7_75t_L g4178 ( 
.A(n_3881),
.Y(n_4178)
);

INVx1_ASAP7_75t_SL g4179 ( 
.A(n_3972),
.Y(n_4179)
);

INVx5_ASAP7_75t_L g4180 ( 
.A(n_3891),
.Y(n_4180)
);

BUFx6f_ASAP7_75t_L g4181 ( 
.A(n_3794),
.Y(n_4181)
);

AOI22xp33_ASAP7_75t_SL g4182 ( 
.A1(n_4010),
.A2(n_3251),
.B1(n_3275),
.B2(n_3237),
.Y(n_4182)
);

NAND2x1p5_ASAP7_75t_L g4183 ( 
.A(n_3944),
.B(n_3251),
.Y(n_4183)
);

AOI22xp33_ASAP7_75t_L g4184 ( 
.A1(n_3741),
.A2(n_3340),
.B1(n_3347),
.B2(n_3310),
.Y(n_4184)
);

BUFx10_ASAP7_75t_L g4185 ( 
.A(n_3916),
.Y(n_4185)
);

INVx1_ASAP7_75t_SL g4186 ( 
.A(n_3966),
.Y(n_4186)
);

AOI22xp33_ASAP7_75t_L g4187 ( 
.A1(n_3792),
.A2(n_4011),
.B1(n_3808),
.B2(n_3799),
.Y(n_4187)
);

AOI22xp33_ASAP7_75t_L g4188 ( 
.A1(n_3819),
.A2(n_3378),
.B1(n_3383),
.B2(n_3361),
.Y(n_4188)
);

CKINVDCx6p67_ASAP7_75t_R g4189 ( 
.A(n_3786),
.Y(n_4189)
);

BUFx6f_ASAP7_75t_L g4190 ( 
.A(n_3929),
.Y(n_4190)
);

BUFx6f_ASAP7_75t_L g4191 ( 
.A(n_3955),
.Y(n_4191)
);

INVx1_ASAP7_75t_L g4192 ( 
.A(n_3881),
.Y(n_4192)
);

AOI22xp33_ASAP7_75t_L g4193 ( 
.A1(n_3858),
.A2(n_3389),
.B1(n_3395),
.B2(n_3384),
.Y(n_4193)
);

CKINVDCx20_ASAP7_75t_R g4194 ( 
.A(n_3865),
.Y(n_4194)
);

BUFx3_ASAP7_75t_L g4195 ( 
.A(n_3991),
.Y(n_4195)
);

NAND2xp5_ASAP7_75t_L g4196 ( 
.A(n_3923),
.B(n_3448),
.Y(n_4196)
);

INVx2_ASAP7_75t_L g4197 ( 
.A(n_3803),
.Y(n_4197)
);

OAI22xp33_ASAP7_75t_L g4198 ( 
.A1(n_3978),
.A2(n_3626),
.B1(n_3603),
.B2(n_3594),
.Y(n_4198)
);

AOI22xp33_ASAP7_75t_L g4199 ( 
.A1(n_3925),
.A2(n_3410),
.B1(n_3426),
.B2(n_3408),
.Y(n_4199)
);

INVx2_ASAP7_75t_L g4200 ( 
.A(n_3839),
.Y(n_4200)
);

BUFx2_ASAP7_75t_L g4201 ( 
.A(n_3843),
.Y(n_4201)
);

INVx1_ASAP7_75t_L g4202 ( 
.A(n_3882),
.Y(n_4202)
);

AND2x2_ASAP7_75t_L g4203 ( 
.A(n_3848),
.B(n_3491),
.Y(n_4203)
);

AND2x2_ASAP7_75t_L g4204 ( 
.A(n_3930),
.B(n_655),
.Y(n_4204)
);

CKINVDCx20_ASAP7_75t_R g4205 ( 
.A(n_4000),
.Y(n_4205)
);

INVx1_ASAP7_75t_L g4206 ( 
.A(n_3882),
.Y(n_4206)
);

AOI22xp33_ASAP7_75t_L g4207 ( 
.A1(n_3961),
.A2(n_3467),
.B1(n_3469),
.B2(n_3453),
.Y(n_4207)
);

AOI22xp5_ASAP7_75t_L g4208 ( 
.A1(n_3983),
.A2(n_3480),
.B1(n_3471),
.B2(n_3623),
.Y(n_4208)
);

AOI22xp33_ASAP7_75t_L g4209 ( 
.A1(n_3989),
.A2(n_3687),
.B1(n_3674),
.B2(n_3309),
.Y(n_4209)
);

NAND2xp5_ASAP7_75t_L g4210 ( 
.A(n_3922),
.B(n_3926),
.Y(n_4210)
);

CKINVDCx5p33_ASAP7_75t_R g4211 ( 
.A(n_3864),
.Y(n_4211)
);

INVx2_ASAP7_75t_L g4212 ( 
.A(n_3818),
.Y(n_4212)
);

INVx6_ASAP7_75t_L g4213 ( 
.A(n_3773),
.Y(n_4213)
);

BUFx4f_ASAP7_75t_SL g4214 ( 
.A(n_3965),
.Y(n_4214)
);

BUFx6f_ASAP7_75t_L g4215 ( 
.A(n_3877),
.Y(n_4215)
);

CKINVDCx5p33_ASAP7_75t_R g4216 ( 
.A(n_3948),
.Y(n_4216)
);

INVx1_ASAP7_75t_L g4217 ( 
.A(n_3868),
.Y(n_4217)
);

INVx1_ASAP7_75t_L g4218 ( 
.A(n_3868),
.Y(n_4218)
);

INVx1_ASAP7_75t_L g4219 ( 
.A(n_3788),
.Y(n_4219)
);

AOI22xp33_ASAP7_75t_L g4220 ( 
.A1(n_3883),
.A2(n_3309),
.B1(n_3354),
.B2(n_3275),
.Y(n_4220)
);

BUFx6f_ASAP7_75t_L g4221 ( 
.A(n_3720),
.Y(n_4221)
);

NAND2xp5_ASAP7_75t_L g4222 ( 
.A(n_3963),
.B(n_3535),
.Y(n_4222)
);

INVx6_ASAP7_75t_L g4223 ( 
.A(n_3945),
.Y(n_4223)
);

INVx1_ASAP7_75t_L g4224 ( 
.A(n_3810),
.Y(n_4224)
);

BUFx3_ASAP7_75t_L g4225 ( 
.A(n_4061),
.Y(n_4225)
);

BUFx3_ASAP7_75t_L g4226 ( 
.A(n_4017),
.Y(n_4226)
);

INVxp67_ASAP7_75t_R g4227 ( 
.A(n_4064),
.Y(n_4227)
);

INVx1_ASAP7_75t_L g4228 ( 
.A(n_4020),
.Y(n_4228)
);

INVx2_ASAP7_75t_L g4229 ( 
.A(n_4027),
.Y(n_4229)
);

BUFx2_ASAP7_75t_L g4230 ( 
.A(n_4060),
.Y(n_4230)
);

AND2x4_ASAP7_75t_L g4231 ( 
.A(n_4097),
.B(n_3889),
.Y(n_4231)
);

BUFx2_ASAP7_75t_L g4232 ( 
.A(n_4077),
.Y(n_4232)
);

HB1xp67_ASAP7_75t_L g4233 ( 
.A(n_4162),
.Y(n_4233)
);

AND2x2_ASAP7_75t_L g4234 ( 
.A(n_4152),
.B(n_3889),
.Y(n_4234)
);

INVx1_ASAP7_75t_L g4235 ( 
.A(n_4178),
.Y(n_4235)
);

BUFx2_ASAP7_75t_L g4236 ( 
.A(n_4156),
.Y(n_4236)
);

INVx1_ASAP7_75t_L g4237 ( 
.A(n_4192),
.Y(n_4237)
);

INVx1_ASAP7_75t_L g4238 ( 
.A(n_4202),
.Y(n_4238)
);

INVx2_ASAP7_75t_L g4239 ( 
.A(n_4037),
.Y(n_4239)
);

INVx1_ASAP7_75t_L g4240 ( 
.A(n_4030),
.Y(n_4240)
);

AO21x2_ASAP7_75t_L g4241 ( 
.A1(n_4222),
.A2(n_3987),
.B(n_3717),
.Y(n_4241)
);

INVx1_ASAP7_75t_L g4242 ( 
.A(n_4033),
.Y(n_4242)
);

OAI21xp5_ASAP7_75t_L g4243 ( 
.A1(n_4038),
.A2(n_3924),
.B(n_3951),
.Y(n_4243)
);

NAND2x1p5_ASAP7_75t_L g4244 ( 
.A(n_4106),
.B(n_3982),
.Y(n_4244)
);

INVx1_ASAP7_75t_L g4245 ( 
.A(n_4039),
.Y(n_4245)
);

AOI22xp33_ASAP7_75t_L g4246 ( 
.A1(n_4205),
.A2(n_3713),
.B1(n_3777),
.B2(n_3915),
.Y(n_4246)
);

OAI21x1_ASAP7_75t_L g4247 ( 
.A1(n_4127),
.A2(n_3726),
.B(n_3694),
.Y(n_4247)
);

INVx1_ASAP7_75t_L g4248 ( 
.A(n_4047),
.Y(n_4248)
);

BUFx2_ASAP7_75t_L g4249 ( 
.A(n_4065),
.Y(n_4249)
);

INVx2_ASAP7_75t_L g4250 ( 
.A(n_4054),
.Y(n_4250)
);

NAND2xp5_ASAP7_75t_L g4251 ( 
.A(n_4076),
.B(n_3825),
.Y(n_4251)
);

INVx2_ASAP7_75t_L g4252 ( 
.A(n_4059),
.Y(n_4252)
);

INVx2_ASAP7_75t_L g4253 ( 
.A(n_4073),
.Y(n_4253)
);

NAND2xp5_ASAP7_75t_L g4254 ( 
.A(n_4145),
.B(n_3846),
.Y(n_4254)
);

INVx3_ASAP7_75t_L g4255 ( 
.A(n_4185),
.Y(n_4255)
);

INVx2_ASAP7_75t_SL g4256 ( 
.A(n_4023),
.Y(n_4256)
);

AND2x4_ASAP7_75t_L g4257 ( 
.A(n_4146),
.B(n_4028),
.Y(n_4257)
);

NAND2xp5_ASAP7_75t_L g4258 ( 
.A(n_4148),
.B(n_3862),
.Y(n_4258)
);

INVxp67_ASAP7_75t_L g4259 ( 
.A(n_4074),
.Y(n_4259)
);

INVx2_ASAP7_75t_L g4260 ( 
.A(n_4080),
.Y(n_4260)
);

INVx2_ASAP7_75t_L g4261 ( 
.A(n_4083),
.Y(n_4261)
);

INVx1_ASAP7_75t_L g4262 ( 
.A(n_4057),
.Y(n_4262)
);

INVx1_ASAP7_75t_L g4263 ( 
.A(n_4062),
.Y(n_4263)
);

INVx1_ASAP7_75t_L g4264 ( 
.A(n_4206),
.Y(n_4264)
);

NAND2xp5_ASAP7_75t_L g4265 ( 
.A(n_4155),
.B(n_3850),
.Y(n_4265)
);

OR2x2_ASAP7_75t_L g4266 ( 
.A(n_4082),
.B(n_3860),
.Y(n_4266)
);

INVx1_ASAP7_75t_L g4267 ( 
.A(n_4067),
.Y(n_4267)
);

INVx2_ASAP7_75t_L g4268 ( 
.A(n_4107),
.Y(n_4268)
);

INVx1_ASAP7_75t_L g4269 ( 
.A(n_4217),
.Y(n_4269)
);

INVx1_ASAP7_75t_SL g4270 ( 
.A(n_4032),
.Y(n_4270)
);

INVx2_ASAP7_75t_SL g4271 ( 
.A(n_4023),
.Y(n_4271)
);

AND2x2_ASAP7_75t_L g4272 ( 
.A(n_4098),
.B(n_3818),
.Y(n_4272)
);

INVx2_ASAP7_75t_L g4273 ( 
.A(n_4144),
.Y(n_4273)
);

AO21x2_ASAP7_75t_L g4274 ( 
.A1(n_4218),
.A2(n_3813),
.B(n_3812),
.Y(n_4274)
);

INVx1_ASAP7_75t_L g4275 ( 
.A(n_4071),
.Y(n_4275)
);

INVx1_ASAP7_75t_L g4276 ( 
.A(n_4086),
.Y(n_4276)
);

INVx1_ASAP7_75t_L g4277 ( 
.A(n_4099),
.Y(n_4277)
);

OR2x2_ASAP7_75t_L g4278 ( 
.A(n_4143),
.B(n_3946),
.Y(n_4278)
);

BUFx2_ASAP7_75t_L g4279 ( 
.A(n_4069),
.Y(n_4279)
);

INVx1_ASAP7_75t_L g4280 ( 
.A(n_4113),
.Y(n_4280)
);

BUFx2_ASAP7_75t_SL g4281 ( 
.A(n_4093),
.Y(n_4281)
);

INVx1_ASAP7_75t_L g4282 ( 
.A(n_4117),
.Y(n_4282)
);

INVx1_ASAP7_75t_L g4283 ( 
.A(n_4125),
.Y(n_4283)
);

AND2x4_ASAP7_75t_L g4284 ( 
.A(n_4069),
.B(n_4013),
.Y(n_4284)
);

INVx3_ASAP7_75t_L g4285 ( 
.A(n_4081),
.Y(n_4285)
);

AND2x2_ASAP7_75t_L g4286 ( 
.A(n_4132),
.B(n_3985),
.Y(n_4286)
);

HB1xp67_ASAP7_75t_SL g4287 ( 
.A(n_4025),
.Y(n_4287)
);

O2A1O1Ixp33_ASAP7_75t_L g4288 ( 
.A1(n_4151),
.A2(n_3992),
.B(n_3975),
.C(n_3996),
.Y(n_4288)
);

INVx3_ASAP7_75t_L g4289 ( 
.A(n_4081),
.Y(n_4289)
);

INVx2_ASAP7_75t_L g4290 ( 
.A(n_4153),
.Y(n_4290)
);

INVx1_ASAP7_75t_L g4291 ( 
.A(n_4170),
.Y(n_4291)
);

INVx2_ASAP7_75t_L g4292 ( 
.A(n_4159),
.Y(n_4292)
);

BUFx3_ASAP7_75t_L g4293 ( 
.A(n_4035),
.Y(n_4293)
);

INVx3_ASAP7_75t_L g4294 ( 
.A(n_4123),
.Y(n_4294)
);

INVx1_ASAP7_75t_L g4295 ( 
.A(n_4171),
.Y(n_4295)
);

BUFx3_ASAP7_75t_L g4296 ( 
.A(n_4035),
.Y(n_4296)
);

INVx2_ASAP7_75t_L g4297 ( 
.A(n_4160),
.Y(n_4297)
);

INVx2_ASAP7_75t_L g4298 ( 
.A(n_4176),
.Y(n_4298)
);

INVx1_ASAP7_75t_L g4299 ( 
.A(n_4196),
.Y(n_4299)
);

BUFx6f_ASAP7_75t_L g4300 ( 
.A(n_4101),
.Y(n_4300)
);

INVx2_ASAP7_75t_L g4301 ( 
.A(n_4172),
.Y(n_4301)
);

INVx1_ASAP7_75t_L g4302 ( 
.A(n_4212),
.Y(n_4302)
);

INVx1_ASAP7_75t_L g4303 ( 
.A(n_4172),
.Y(n_4303)
);

INVx2_ASAP7_75t_L g4304 ( 
.A(n_4203),
.Y(n_4304)
);

INVx1_ASAP7_75t_L g4305 ( 
.A(n_4210),
.Y(n_4305)
);

CKINVDCx5p33_ASAP7_75t_R g4306 ( 
.A(n_4029),
.Y(n_4306)
);

CKINVDCx20_ASAP7_75t_R g4307 ( 
.A(n_4021),
.Y(n_4307)
);

INVx2_ASAP7_75t_L g4308 ( 
.A(n_4175),
.Y(n_4308)
);

INVx2_ASAP7_75t_L g4309 ( 
.A(n_4150),
.Y(n_4309)
);

INVx1_ASAP7_75t_L g4310 ( 
.A(n_4219),
.Y(n_4310)
);

INVx2_ASAP7_75t_SL g4311 ( 
.A(n_4079),
.Y(n_4311)
);

INVxp67_ASAP7_75t_L g4312 ( 
.A(n_4116),
.Y(n_4312)
);

AOI21x1_ASAP7_75t_L g4313 ( 
.A1(n_4201),
.A2(n_3699),
.B(n_3692),
.Y(n_4313)
);

HB1xp67_ASAP7_75t_L g4314 ( 
.A(n_4100),
.Y(n_4314)
);

INVx1_ASAP7_75t_L g4315 ( 
.A(n_4224),
.Y(n_4315)
);

OA21x2_ASAP7_75t_L g4316 ( 
.A1(n_4197),
.A2(n_3927),
.B(n_3976),
.Y(n_4316)
);

INVx1_ASAP7_75t_SL g4317 ( 
.A(n_4044),
.Y(n_4317)
);

AND2x2_ASAP7_75t_L g4318 ( 
.A(n_4041),
.B(n_3779),
.Y(n_4318)
);

INVx1_ASAP7_75t_L g4319 ( 
.A(n_4204),
.Y(n_4319)
);

INVx2_ASAP7_75t_L g4320 ( 
.A(n_4150),
.Y(n_4320)
);

INVx3_ASAP7_75t_L g4321 ( 
.A(n_4123),
.Y(n_4321)
);

AND2x2_ASAP7_75t_L g4322 ( 
.A(n_4179),
.B(n_4070),
.Y(n_4322)
);

INVx3_ASAP7_75t_L g4323 ( 
.A(n_4213),
.Y(n_4323)
);

AO21x2_ASAP7_75t_L g4324 ( 
.A1(n_4040),
.A2(n_3829),
.B(n_3815),
.Y(n_4324)
);

AND2x2_ASAP7_75t_L g4325 ( 
.A(n_4070),
.B(n_3779),
.Y(n_4325)
);

INVx1_ASAP7_75t_L g4326 ( 
.A(n_4131),
.Y(n_4326)
);

OAI21x1_ASAP7_75t_L g4327 ( 
.A1(n_4200),
.A2(n_3701),
.B(n_3690),
.Y(n_4327)
);

HB1xp67_ASAP7_75t_L g4328 ( 
.A(n_4128),
.Y(n_4328)
);

BUFx2_ASAP7_75t_L g4329 ( 
.A(n_4101),
.Y(n_4329)
);

INVx1_ASAP7_75t_L g4330 ( 
.A(n_4091),
.Y(n_4330)
);

AO31x2_ASAP7_75t_L g4331 ( 
.A1(n_4118),
.A2(n_4006),
.A3(n_3710),
.B(n_3980),
.Y(n_4331)
);

AND2x4_ASAP7_75t_L g4332 ( 
.A(n_4164),
.B(n_3940),
.Y(n_4332)
);

OA21x2_ASAP7_75t_L g4333 ( 
.A1(n_4177),
.A2(n_3904),
.B(n_3695),
.Y(n_4333)
);

AND2x4_ASAP7_75t_L g4334 ( 
.A(n_4180),
.B(n_3940),
.Y(n_4334)
);

INVx2_ASAP7_75t_SL g4335 ( 
.A(n_4043),
.Y(n_4335)
);

BUFx8_ASAP7_75t_L g4336 ( 
.A(n_4075),
.Y(n_4336)
);

INVx1_ASAP7_75t_L g4337 ( 
.A(n_4186),
.Y(n_4337)
);

INVx1_ASAP7_75t_L g4338 ( 
.A(n_4124),
.Y(n_4338)
);

INVx1_ASAP7_75t_L g4339 ( 
.A(n_4174),
.Y(n_4339)
);

INVx1_ASAP7_75t_L g4340 ( 
.A(n_4119),
.Y(n_4340)
);

INVx2_ASAP7_75t_L g4341 ( 
.A(n_4158),
.Y(n_4341)
);

INVx1_ASAP7_75t_L g4342 ( 
.A(n_4103),
.Y(n_4342)
);

INVx2_ASAP7_75t_L g4343 ( 
.A(n_4213),
.Y(n_4343)
);

AOI22xp33_ASAP7_75t_L g4344 ( 
.A1(n_4036),
.A2(n_3959),
.B1(n_4007),
.B2(n_3832),
.Y(n_4344)
);

AOI22xp33_ASAP7_75t_L g4345 ( 
.A1(n_4194),
.A2(n_3732),
.B1(n_4005),
.B2(n_3999),
.Y(n_4345)
);

INVx1_ASAP7_75t_L g4346 ( 
.A(n_4135),
.Y(n_4346)
);

HB1xp67_ASAP7_75t_L g4347 ( 
.A(n_4166),
.Y(n_4347)
);

BUFx2_ASAP7_75t_L g4348 ( 
.A(n_4120),
.Y(n_4348)
);

INVx2_ASAP7_75t_L g4349 ( 
.A(n_4181),
.Y(n_4349)
);

INVx2_ASAP7_75t_L g4350 ( 
.A(n_4181),
.Y(n_4350)
);

INVx1_ASAP7_75t_L g4351 ( 
.A(n_4195),
.Y(n_4351)
);

CKINVDCx5p33_ASAP7_75t_R g4352 ( 
.A(n_4016),
.Y(n_4352)
);

INVx1_ASAP7_75t_L g4353 ( 
.A(n_4190),
.Y(n_4353)
);

BUFx3_ASAP7_75t_L g4354 ( 
.A(n_4095),
.Y(n_4354)
);

NAND4xp25_ASAP7_75t_L g4355 ( 
.A(n_4019),
.B(n_3897),
.C(n_3937),
.D(n_3872),
.Y(n_4355)
);

INVx1_ASAP7_75t_L g4356 ( 
.A(n_4111),
.Y(n_4356)
);

AO21x2_ASAP7_75t_L g4357 ( 
.A1(n_4138),
.A2(n_3831),
.B(n_3934),
.Y(n_4357)
);

INVx1_ASAP7_75t_L g4358 ( 
.A(n_4112),
.Y(n_4358)
);

AO21x1_ASAP7_75t_SL g4359 ( 
.A1(n_4220),
.A2(n_3727),
.B(n_3745),
.Y(n_4359)
);

INVx1_ASAP7_75t_L g4360 ( 
.A(n_4112),
.Y(n_4360)
);

INVxp67_ASAP7_75t_L g4361 ( 
.A(n_4088),
.Y(n_4361)
);

OAI21x1_ASAP7_75t_L g4362 ( 
.A1(n_4183),
.A2(n_3711),
.B(n_3760),
.Y(n_4362)
);

INVx2_ASAP7_75t_L g4363 ( 
.A(n_4215),
.Y(n_4363)
);

INVx2_ASAP7_75t_L g4364 ( 
.A(n_4215),
.Y(n_4364)
);

CKINVDCx20_ASAP7_75t_R g4365 ( 
.A(n_4024),
.Y(n_4365)
);

INVx1_ASAP7_75t_L g4366 ( 
.A(n_4190),
.Y(n_4366)
);

INVx2_ASAP7_75t_L g4367 ( 
.A(n_4191),
.Y(n_4367)
);

A2O1A1Ixp33_ASAP7_75t_L g4368 ( 
.A1(n_4255),
.A2(n_4034),
.B(n_4058),
.C(n_4026),
.Y(n_4368)
);

BUFx3_ASAP7_75t_L g4369 ( 
.A(n_4293),
.Y(n_4369)
);

AOI21xp5_ASAP7_75t_L g4370 ( 
.A1(n_4288),
.A2(n_4182),
.B(n_4167),
.Y(n_4370)
);

NAND2xp5_ASAP7_75t_L g4371 ( 
.A(n_4318),
.B(n_4126),
.Y(n_4371)
);

AND2x2_ASAP7_75t_L g4372 ( 
.A(n_4233),
.B(n_4096),
.Y(n_4372)
);

AND2x2_ASAP7_75t_L g4373 ( 
.A(n_4304),
.B(n_4168),
.Y(n_4373)
);

NAND2xp5_ASAP7_75t_L g4374 ( 
.A(n_4286),
.B(n_4141),
.Y(n_4374)
);

OR2x2_ASAP7_75t_L g4375 ( 
.A(n_4230),
.B(n_4078),
.Y(n_4375)
);

AND2x4_ASAP7_75t_L g4376 ( 
.A(n_4257),
.B(n_4180),
.Y(n_4376)
);

OAI21xp5_ASAP7_75t_L g4377 ( 
.A1(n_4243),
.A2(n_4129),
.B(n_4149),
.Y(n_4377)
);

AND2x2_ASAP7_75t_L g4378 ( 
.A(n_4232),
.B(n_4301),
.Y(n_4378)
);

NAND2xp5_ASAP7_75t_L g4379 ( 
.A(n_4330),
.B(n_4084),
.Y(n_4379)
);

AOI22xp5_ASAP7_75t_L g4380 ( 
.A1(n_4246),
.A2(n_4211),
.B1(n_4216),
.B2(n_4094),
.Y(n_4380)
);

INVx2_ASAP7_75t_L g4381 ( 
.A(n_4229),
.Y(n_4381)
);

CKINVDCx20_ASAP7_75t_R g4382 ( 
.A(n_4307),
.Y(n_4382)
);

OR2x6_ASAP7_75t_L g4383 ( 
.A(n_4281),
.B(n_4051),
.Y(n_4383)
);

OR2x2_ASAP7_75t_L g4384 ( 
.A(n_4308),
.B(n_4012),
.Y(n_4384)
);

AND2x4_ASAP7_75t_L g4385 ( 
.A(n_4257),
.B(n_4050),
.Y(n_4385)
);

OAI22xp5_ASAP7_75t_SL g4386 ( 
.A1(n_4339),
.A2(n_4051),
.B1(n_4115),
.B2(n_4053),
.Y(n_4386)
);

NOR2x1_ASAP7_75t_SL g4387 ( 
.A(n_4281),
.B(n_4092),
.Y(n_4387)
);

INVx3_ASAP7_75t_L g4388 ( 
.A(n_4300),
.Y(n_4388)
);

NAND2xp5_ASAP7_75t_L g4389 ( 
.A(n_4340),
.B(n_4187),
.Y(n_4389)
);

NAND2xp5_ASAP7_75t_L g4390 ( 
.A(n_4298),
.B(n_4139),
.Y(n_4390)
);

BUFx2_ASAP7_75t_L g4391 ( 
.A(n_4249),
.Y(n_4391)
);

AND2x2_ASAP7_75t_L g4392 ( 
.A(n_4303),
.B(n_4121),
.Y(n_4392)
);

AND2x2_ASAP7_75t_L g4393 ( 
.A(n_4322),
.B(n_4338),
.Y(n_4393)
);

AOI21xp5_ASAP7_75t_L g4394 ( 
.A1(n_4347),
.A2(n_4241),
.B(n_4063),
.Y(n_4394)
);

OAI31xp33_ASAP7_75t_SL g4395 ( 
.A1(n_4270),
.A2(n_4109),
.A3(n_4046),
.B(n_4085),
.Y(n_4395)
);

OA21x2_ASAP7_75t_L g4396 ( 
.A1(n_4231),
.A2(n_4157),
.B(n_4089),
.Y(n_4396)
);

NOR2xp33_ASAP7_75t_L g4397 ( 
.A(n_4312),
.B(n_4018),
.Y(n_4397)
);

OA21x2_ASAP7_75t_L g4398 ( 
.A1(n_4231),
.A2(n_4134),
.B(n_4090),
.Y(n_4398)
);

OR2x2_ASAP7_75t_L g4399 ( 
.A(n_4234),
.B(n_4337),
.Y(n_4399)
);

INVx3_ASAP7_75t_L g4400 ( 
.A(n_4300),
.Y(n_4400)
);

OAI22xp5_ASAP7_75t_L g4401 ( 
.A1(n_4287),
.A2(n_4189),
.B1(n_4214),
.B2(n_4022),
.Y(n_4401)
);

AO32x1_ASAP7_75t_L g4402 ( 
.A1(n_4343),
.A2(n_4066),
.A3(n_4105),
.B1(n_4087),
.B2(n_4223),
.Y(n_4402)
);

OR2x2_ASAP7_75t_L g4403 ( 
.A(n_4305),
.B(n_4228),
.Y(n_4403)
);

AND2x2_ASAP7_75t_L g4404 ( 
.A(n_4341),
.B(n_4043),
.Y(n_4404)
);

INVx2_ASAP7_75t_L g4405 ( 
.A(n_4239),
.Y(n_4405)
);

AND2x2_ASAP7_75t_L g4406 ( 
.A(n_4272),
.B(n_4045),
.Y(n_4406)
);

BUFx3_ASAP7_75t_L g4407 ( 
.A(n_4296),
.Y(n_4407)
);

AND2x2_ASAP7_75t_L g4408 ( 
.A(n_4314),
.B(n_4045),
.Y(n_4408)
);

INVx3_ASAP7_75t_L g4409 ( 
.A(n_4300),
.Y(n_4409)
);

INVx3_ASAP7_75t_L g4410 ( 
.A(n_4329),
.Y(n_4410)
);

OR2x6_ASAP7_75t_L g4411 ( 
.A(n_4236),
.B(n_4223),
.Y(n_4411)
);

OAI21xp5_ASAP7_75t_L g4412 ( 
.A1(n_4284),
.A2(n_3973),
.B(n_3942),
.Y(n_4412)
);

OAI21xp5_ASAP7_75t_L g4413 ( 
.A1(n_4284),
.A2(n_3899),
.B(n_3878),
.Y(n_4413)
);

O2A1O1Ixp33_ASAP7_75t_L g4414 ( 
.A1(n_4355),
.A2(n_3968),
.B(n_3995),
.C(n_3981),
.Y(n_4414)
);

INVx4_ASAP7_75t_L g4415 ( 
.A(n_4225),
.Y(n_4415)
);

NOR2x1_ASAP7_75t_SL g4416 ( 
.A(n_4359),
.B(n_4110),
.Y(n_4416)
);

OR2x2_ASAP7_75t_L g4417 ( 
.A(n_4240),
.B(n_4012),
.Y(n_4417)
);

INVx1_ASAP7_75t_L g4418 ( 
.A(n_4242),
.Y(n_4418)
);

AND2x4_ASAP7_75t_L g4419 ( 
.A(n_4255),
.B(n_4191),
.Y(n_4419)
);

AND2x4_ASAP7_75t_L g4420 ( 
.A(n_4279),
.B(n_4049),
.Y(n_4420)
);

AO32x2_ASAP7_75t_L g4421 ( 
.A1(n_4335),
.A2(n_4133),
.A3(n_3691),
.B1(n_4056),
.B2(n_4137),
.Y(n_4421)
);

OAI21x1_ASAP7_75t_SL g4422 ( 
.A1(n_4311),
.A2(n_4031),
.B(n_3960),
.Y(n_4422)
);

INVx4_ASAP7_75t_L g4423 ( 
.A(n_4348),
.Y(n_4423)
);

OAI21x1_ASAP7_75t_SL g4424 ( 
.A1(n_4227),
.A2(n_4042),
.B(n_4102),
.Y(n_4424)
);

INVx1_ASAP7_75t_L g4425 ( 
.A(n_4245),
.Y(n_4425)
);

AND2x2_ASAP7_75t_L g4426 ( 
.A(n_4328),
.B(n_4108),
.Y(n_4426)
);

NOR2xp33_ASAP7_75t_SL g4427 ( 
.A(n_4336),
.B(n_4052),
.Y(n_4427)
);

INVx2_ASAP7_75t_L g4428 ( 
.A(n_4250),
.Y(n_4428)
);

NOR2xp33_ASAP7_75t_L g4429 ( 
.A(n_4342),
.B(n_4018),
.Y(n_4429)
);

HB1xp67_ASAP7_75t_L g4430 ( 
.A(n_4317),
.Y(n_4430)
);

INVx3_ASAP7_75t_L g4431 ( 
.A(n_4336),
.Y(n_4431)
);

NAND2x1_ASAP7_75t_L g4432 ( 
.A(n_4334),
.B(n_4108),
.Y(n_4432)
);

OR2x2_ASAP7_75t_L g4433 ( 
.A(n_4248),
.B(n_3906),
.Y(n_4433)
);

NAND2xp5_ASAP7_75t_L g4434 ( 
.A(n_4299),
.B(n_3784),
.Y(n_4434)
);

OAI22xp5_ASAP7_75t_L g4435 ( 
.A1(n_4244),
.A2(n_4072),
.B1(n_4136),
.B2(n_4068),
.Y(n_4435)
);

OR2x2_ASAP7_75t_L g4436 ( 
.A(n_4262),
.B(n_3906),
.Y(n_4436)
);

OAI22xp5_ASAP7_75t_L g4437 ( 
.A1(n_4259),
.A2(n_4048),
.B1(n_4055),
.B2(n_4142),
.Y(n_4437)
);

INVx2_ASAP7_75t_L g4438 ( 
.A(n_4252),
.Y(n_4438)
);

OR2x2_ASAP7_75t_L g4439 ( 
.A(n_4263),
.B(n_3784),
.Y(n_4439)
);

OAI22xp5_ASAP7_75t_SL g4440 ( 
.A1(n_4352),
.A2(n_4104),
.B1(n_4169),
.B2(n_4165),
.Y(n_4440)
);

INVx2_ASAP7_75t_L g4441 ( 
.A(n_4253),
.Y(n_4441)
);

INVx3_ASAP7_75t_L g4442 ( 
.A(n_4354),
.Y(n_4442)
);

BUFx4f_ASAP7_75t_SL g4443 ( 
.A(n_4365),
.Y(n_4443)
);

AND2x2_ASAP7_75t_L g4444 ( 
.A(n_4326),
.B(n_4221),
.Y(n_4444)
);

OR2x6_ASAP7_75t_L g4445 ( 
.A(n_4285),
.B(n_3970),
.Y(n_4445)
);

INVxp67_ASAP7_75t_L g4446 ( 
.A(n_4310),
.Y(n_4446)
);

NAND2xp5_ASAP7_75t_L g4447 ( 
.A(n_4315),
.B(n_3817),
.Y(n_4447)
);

INVx2_ASAP7_75t_L g4448 ( 
.A(n_4260),
.Y(n_4448)
);

INVx1_ASAP7_75t_L g4449 ( 
.A(n_4267),
.Y(n_4449)
);

OAI21x1_ASAP7_75t_L g4450 ( 
.A1(n_4313),
.A2(n_3879),
.B(n_3733),
.Y(n_4450)
);

NAND2xp5_ASAP7_75t_L g4451 ( 
.A(n_4251),
.B(n_3817),
.Y(n_4451)
);

OAI211xp5_ASAP7_75t_L g4452 ( 
.A1(n_4344),
.A2(n_4163),
.B(n_4184),
.C(n_4173),
.Y(n_4452)
);

AOI221xp5_ASAP7_75t_L g4453 ( 
.A1(n_4319),
.A2(n_3936),
.B1(n_3933),
.B2(n_3977),
.C(n_3921),
.Y(n_4453)
);

A2O1A1Ixp33_ASAP7_75t_L g4454 ( 
.A1(n_4294),
.A2(n_3828),
.B(n_3820),
.C(n_3852),
.Y(n_4454)
);

OR2x6_ASAP7_75t_L g4455 ( 
.A(n_4285),
.B(n_4289),
.Y(n_4455)
);

INVx1_ASAP7_75t_L g4456 ( 
.A(n_4403),
.Y(n_4456)
);

CKINVDCx20_ASAP7_75t_R g4457 ( 
.A(n_4382),
.Y(n_4457)
);

OR2x2_ASAP7_75t_L g4458 ( 
.A(n_4399),
.B(n_4275),
.Y(n_4458)
);

NAND2x1_ASAP7_75t_L g4459 ( 
.A(n_4383),
.B(n_4334),
.Y(n_4459)
);

AND2x2_ASAP7_75t_L g4460 ( 
.A(n_4406),
.B(n_4325),
.Y(n_4460)
);

INVx1_ASAP7_75t_L g4461 ( 
.A(n_4403),
.Y(n_4461)
);

AOI22xp5_ASAP7_75t_L g4462 ( 
.A1(n_4437),
.A2(n_4345),
.B1(n_4332),
.B2(n_4208),
.Y(n_4462)
);

AND2x4_ASAP7_75t_L g4463 ( 
.A(n_4419),
.B(n_4444),
.Y(n_4463)
);

AND2x2_ASAP7_75t_L g4464 ( 
.A(n_4378),
.B(n_4276),
.Y(n_4464)
);

AND2x2_ASAP7_75t_L g4465 ( 
.A(n_4393),
.B(n_4277),
.Y(n_4465)
);

NAND2xp5_ASAP7_75t_L g4466 ( 
.A(n_4451),
.B(n_4280),
.Y(n_4466)
);

AOI22xp33_ASAP7_75t_L g4467 ( 
.A1(n_4440),
.A2(n_4332),
.B1(n_4324),
.B2(n_4357),
.Y(n_4467)
);

INVx2_ASAP7_75t_L g4468 ( 
.A(n_4391),
.Y(n_4468)
);

OR2x2_ASAP7_75t_L g4469 ( 
.A(n_4399),
.B(n_4282),
.Y(n_4469)
);

AND2x2_ASAP7_75t_L g4470 ( 
.A(n_4430),
.B(n_4283),
.Y(n_4470)
);

NAND2xp5_ASAP7_75t_L g4471 ( 
.A(n_4371),
.B(n_4291),
.Y(n_4471)
);

AND2x2_ASAP7_75t_L g4472 ( 
.A(n_4408),
.B(n_4346),
.Y(n_4472)
);

AND2x2_ASAP7_75t_L g4473 ( 
.A(n_4372),
.B(n_4426),
.Y(n_4473)
);

BUFx2_ASAP7_75t_L g4474 ( 
.A(n_4383),
.Y(n_4474)
);

INVx1_ASAP7_75t_L g4475 ( 
.A(n_4418),
.Y(n_4475)
);

AND2x2_ASAP7_75t_L g4476 ( 
.A(n_4404),
.B(n_4295),
.Y(n_4476)
);

HB1xp67_ASAP7_75t_L g4477 ( 
.A(n_4381),
.Y(n_4477)
);

INVx1_ASAP7_75t_L g4478 ( 
.A(n_4425),
.Y(n_4478)
);

INVx2_ASAP7_75t_L g4479 ( 
.A(n_4405),
.Y(n_4479)
);

HB1xp67_ASAP7_75t_L g4480 ( 
.A(n_4428),
.Y(n_4480)
);

OR2x2_ASAP7_75t_L g4481 ( 
.A(n_4438),
.B(n_4278),
.Y(n_4481)
);

AND2x2_ASAP7_75t_L g4482 ( 
.A(n_4373),
.B(n_4446),
.Y(n_4482)
);

INVx1_ASAP7_75t_L g4483 ( 
.A(n_4449),
.Y(n_4483)
);

NAND2xp5_ASAP7_75t_L g4484 ( 
.A(n_4434),
.B(n_4235),
.Y(n_4484)
);

INVx2_ASAP7_75t_L g4485 ( 
.A(n_4441),
.Y(n_4485)
);

BUFx2_ASAP7_75t_L g4486 ( 
.A(n_4423),
.Y(n_4486)
);

HB1xp67_ASAP7_75t_L g4487 ( 
.A(n_4448),
.Y(n_4487)
);

OAI222xp33_ASAP7_75t_L g4488 ( 
.A1(n_4411),
.A2(n_4266),
.B1(n_4361),
.B2(n_4289),
.C1(n_4356),
.C2(n_4323),
.Y(n_4488)
);

HB1xp67_ASAP7_75t_L g4489 ( 
.A(n_4410),
.Y(n_4489)
);

AND2x2_ASAP7_75t_L g4490 ( 
.A(n_4392),
.B(n_4323),
.Y(n_4490)
);

NAND2xp5_ASAP7_75t_L g4491 ( 
.A(n_4433),
.B(n_4235),
.Y(n_4491)
);

NAND2xp5_ASAP7_75t_L g4492 ( 
.A(n_4436),
.B(n_4237),
.Y(n_4492)
);

OR2x2_ASAP7_75t_L g4493 ( 
.A(n_4384),
.B(n_4261),
.Y(n_4493)
);

AND2x2_ASAP7_75t_L g4494 ( 
.A(n_4385),
.B(n_4351),
.Y(n_4494)
);

INVx5_ASAP7_75t_SL g4495 ( 
.A(n_4411),
.Y(n_4495)
);

INVxp67_ASAP7_75t_SL g4496 ( 
.A(n_4416),
.Y(n_4496)
);

OR2x2_ASAP7_75t_L g4497 ( 
.A(n_4374),
.B(n_4268),
.Y(n_4497)
);

OR2x2_ASAP7_75t_L g4498 ( 
.A(n_4379),
.B(n_4273),
.Y(n_4498)
);

INVx1_ASAP7_75t_L g4499 ( 
.A(n_4389),
.Y(n_4499)
);

AND2x2_ASAP7_75t_L g4500 ( 
.A(n_4442),
.B(n_4366),
.Y(n_4500)
);

AND2x2_ASAP7_75t_L g4501 ( 
.A(n_4396),
.B(n_4349),
.Y(n_4501)
);

AND2x2_ASAP7_75t_L g4502 ( 
.A(n_4398),
.B(n_4350),
.Y(n_4502)
);

AOI22xp33_ASAP7_75t_L g4503 ( 
.A1(n_4377),
.A2(n_4147),
.B1(n_4154),
.B2(n_4358),
.Y(n_4503)
);

AOI22xp33_ASAP7_75t_L g4504 ( 
.A1(n_4424),
.A2(n_4360),
.B1(n_4294),
.B2(n_4321),
.Y(n_4504)
);

INVx2_ASAP7_75t_L g4505 ( 
.A(n_4439),
.Y(n_4505)
);

INVx2_ASAP7_75t_SL g4506 ( 
.A(n_4369),
.Y(n_4506)
);

INVx1_ASAP7_75t_L g4507 ( 
.A(n_4390),
.Y(n_4507)
);

INVx1_ASAP7_75t_L g4508 ( 
.A(n_4417),
.Y(n_4508)
);

INVx1_ASAP7_75t_L g4509 ( 
.A(n_4447),
.Y(n_4509)
);

BUFx2_ASAP7_75t_L g4510 ( 
.A(n_4415),
.Y(n_4510)
);

INVx2_ASAP7_75t_L g4511 ( 
.A(n_4376),
.Y(n_4511)
);

OR2x2_ASAP7_75t_L g4512 ( 
.A(n_4375),
.B(n_4290),
.Y(n_4512)
);

INVx1_ASAP7_75t_L g4513 ( 
.A(n_4455),
.Y(n_4513)
);

NAND2xp5_ASAP7_75t_L g4514 ( 
.A(n_4394),
.B(n_4237),
.Y(n_4514)
);

INVx1_ASAP7_75t_L g4515 ( 
.A(n_4455),
.Y(n_4515)
);

INVx1_ASAP7_75t_L g4516 ( 
.A(n_4387),
.Y(n_4516)
);

NOR2xp33_ASAP7_75t_L g4517 ( 
.A(n_4431),
.B(n_4226),
.Y(n_4517)
);

AND2x2_ASAP7_75t_L g4518 ( 
.A(n_4420),
.B(n_4397),
.Y(n_4518)
);

AOI221xp5_ASAP7_75t_L g4519 ( 
.A1(n_4368),
.A2(n_4265),
.B1(n_4258),
.B2(n_4254),
.C(n_3957),
.Y(n_4519)
);

INVx2_ASAP7_75t_L g4520 ( 
.A(n_4432),
.Y(n_4520)
);

HB1xp67_ASAP7_75t_L g4521 ( 
.A(n_4407),
.Y(n_4521)
);

INVx2_ASAP7_75t_SL g4522 ( 
.A(n_4388),
.Y(n_4522)
);

HB1xp67_ASAP7_75t_L g4523 ( 
.A(n_4400),
.Y(n_4523)
);

INVx1_ASAP7_75t_L g4524 ( 
.A(n_4421),
.Y(n_4524)
);

OR2x2_ASAP7_75t_L g4525 ( 
.A(n_4409),
.B(n_4292),
.Y(n_4525)
);

INVx1_ASAP7_75t_L g4526 ( 
.A(n_4421),
.Y(n_4526)
);

INVx2_ASAP7_75t_L g4527 ( 
.A(n_4445),
.Y(n_4527)
);

AO21x2_ASAP7_75t_L g4528 ( 
.A1(n_4524),
.A2(n_4422),
.B(n_4370),
.Y(n_4528)
);

AO21x2_ASAP7_75t_L g4529 ( 
.A1(n_4526),
.A2(n_4413),
.B(n_4452),
.Y(n_4529)
);

NAND2xp5_ASAP7_75t_L g4530 ( 
.A(n_4509),
.B(n_4297),
.Y(n_4530)
);

INVx2_ASAP7_75t_SL g4531 ( 
.A(n_4510),
.Y(n_4531)
);

INVx1_ASAP7_75t_L g4532 ( 
.A(n_4498),
.Y(n_4532)
);

INVx2_ASAP7_75t_L g4533 ( 
.A(n_4477),
.Y(n_4533)
);

INVx1_ASAP7_75t_L g4534 ( 
.A(n_4458),
.Y(n_4534)
);

AND5x1_ASAP7_75t_L g4535 ( 
.A(n_4519),
.B(n_4427),
.C(n_4395),
.D(n_4462),
.E(n_4517),
.Y(n_4535)
);

AND2x4_ASAP7_75t_L g4536 ( 
.A(n_4496),
.B(n_4445),
.Y(n_4536)
);

INVx2_ASAP7_75t_L g4537 ( 
.A(n_4480),
.Y(n_4537)
);

NOR2xp33_ASAP7_75t_L g4538 ( 
.A(n_4486),
.B(n_4521),
.Y(n_4538)
);

OR2x2_ASAP7_75t_L g4539 ( 
.A(n_4481),
.B(n_4238),
.Y(n_4539)
);

AND2x2_ASAP7_75t_L g4540 ( 
.A(n_4473),
.B(n_4429),
.Y(n_4540)
);

AND2x2_ASAP7_75t_L g4541 ( 
.A(n_4513),
.B(n_4353),
.Y(n_4541)
);

INVx2_ASAP7_75t_L g4542 ( 
.A(n_4487),
.Y(n_4542)
);

AOI22xp33_ASAP7_75t_L g4543 ( 
.A1(n_4519),
.A2(n_4380),
.B1(n_4435),
.B2(n_4401),
.Y(n_4543)
);

INVx2_ASAP7_75t_L g4544 ( 
.A(n_4493),
.Y(n_4544)
);

INVx2_ASAP7_75t_SL g4545 ( 
.A(n_4506),
.Y(n_4545)
);

INVx1_ASAP7_75t_SL g4546 ( 
.A(n_4474),
.Y(n_4546)
);

INVx1_ASAP7_75t_L g4547 ( 
.A(n_4469),
.Y(n_4547)
);

HB1xp67_ASAP7_75t_L g4548 ( 
.A(n_4489),
.Y(n_4548)
);

INVx1_ASAP7_75t_SL g4549 ( 
.A(n_4523),
.Y(n_4549)
);

AND2x2_ASAP7_75t_L g4550 ( 
.A(n_4515),
.B(n_4353),
.Y(n_4550)
);

INVxp67_ASAP7_75t_SL g4551 ( 
.A(n_4496),
.Y(n_4551)
);

AOI22xp5_ASAP7_75t_L g4552 ( 
.A1(n_4462),
.A2(n_4386),
.B1(n_4412),
.B2(n_4321),
.Y(n_4552)
);

AND2x2_ASAP7_75t_L g4553 ( 
.A(n_4460),
.B(n_4363),
.Y(n_4553)
);

INVx2_ASAP7_75t_L g4554 ( 
.A(n_4479),
.Y(n_4554)
);

NAND2x1_ASAP7_75t_L g4555 ( 
.A(n_4516),
.B(n_4364),
.Y(n_4555)
);

OR2x2_ASAP7_75t_L g4556 ( 
.A(n_4497),
.B(n_4238),
.Y(n_4556)
);

AND2x2_ASAP7_75t_L g4557 ( 
.A(n_4494),
.B(n_4367),
.Y(n_4557)
);

INVx1_ASAP7_75t_L g4558 ( 
.A(n_4475),
.Y(n_4558)
);

NAND2xp5_ASAP7_75t_L g4559 ( 
.A(n_4499),
.B(n_4264),
.Y(n_4559)
);

INVx2_ASAP7_75t_L g4560 ( 
.A(n_4485),
.Y(n_4560)
);

OR2x2_ASAP7_75t_L g4561 ( 
.A(n_4471),
.B(n_4505),
.Y(n_4561)
);

HB1xp67_ASAP7_75t_L g4562 ( 
.A(n_4470),
.Y(n_4562)
);

BUFx3_ASAP7_75t_L g4563 ( 
.A(n_4457),
.Y(n_4563)
);

INVx3_ASAP7_75t_L g4564 ( 
.A(n_4459),
.Y(n_4564)
);

AND2x2_ASAP7_75t_L g4565 ( 
.A(n_4482),
.B(n_4309),
.Y(n_4565)
);

INVx1_ASAP7_75t_L g4566 ( 
.A(n_4478),
.Y(n_4566)
);

AND2x2_ASAP7_75t_L g4567 ( 
.A(n_4463),
.B(n_4320),
.Y(n_4567)
);

INVx2_ASAP7_75t_L g4568 ( 
.A(n_4525),
.Y(n_4568)
);

INVx1_ASAP7_75t_L g4569 ( 
.A(n_4483),
.Y(n_4569)
);

NAND4xp25_ASAP7_75t_SL g4570 ( 
.A(n_4504),
.B(n_4414),
.C(n_4443),
.D(n_4402),
.Y(n_4570)
);

HB1xp67_ASAP7_75t_L g4571 ( 
.A(n_4508),
.Y(n_4571)
);

AOI22xp33_ASAP7_75t_L g4572 ( 
.A1(n_4507),
.A2(n_4453),
.B1(n_4271),
.B2(n_4256),
.Y(n_4572)
);

AO21x2_ASAP7_75t_L g4573 ( 
.A1(n_4514),
.A2(n_4450),
.B(n_4313),
.Y(n_4573)
);

AOI22xp33_ASAP7_75t_L g4574 ( 
.A1(n_4503),
.A2(n_4269),
.B1(n_4264),
.B2(n_4199),
.Y(n_4574)
);

INVx1_ASAP7_75t_L g4575 ( 
.A(n_4456),
.Y(n_4575)
);

INVx1_ASAP7_75t_L g4576 ( 
.A(n_4461),
.Y(n_4576)
);

BUFx3_ASAP7_75t_L g4577 ( 
.A(n_4490),
.Y(n_4577)
);

AND2x2_ASAP7_75t_L g4578 ( 
.A(n_4463),
.B(n_4269),
.Y(n_4578)
);

AND2x2_ASAP7_75t_L g4579 ( 
.A(n_4511),
.B(n_4476),
.Y(n_4579)
);

AOI22xp33_ASAP7_75t_L g4580 ( 
.A1(n_4467),
.A2(n_4207),
.B1(n_4114),
.B2(n_4274),
.Y(n_4580)
);

INVx2_ASAP7_75t_L g4581 ( 
.A(n_4512),
.Y(n_4581)
);

OAI31xp33_ASAP7_75t_L g4582 ( 
.A1(n_4488),
.A2(n_4454),
.A3(n_4402),
.B(n_3918),
.Y(n_4582)
);

NAND2xp5_ASAP7_75t_L g4583 ( 
.A(n_4466),
.B(n_4491),
.Y(n_4583)
);

NAND2xp5_ASAP7_75t_L g4584 ( 
.A(n_4466),
.B(n_4331),
.Y(n_4584)
);

INVx2_ASAP7_75t_L g4585 ( 
.A(n_4468),
.Y(n_4585)
);

AND2x2_ASAP7_75t_L g4586 ( 
.A(n_4464),
.B(n_4500),
.Y(n_4586)
);

INVx1_ASAP7_75t_L g4587 ( 
.A(n_4491),
.Y(n_4587)
);

INVx1_ASAP7_75t_L g4588 ( 
.A(n_4492),
.Y(n_4588)
);

INVx2_ASAP7_75t_SL g4589 ( 
.A(n_4518),
.Y(n_4589)
);

INVx2_ASAP7_75t_L g4590 ( 
.A(n_4548),
.Y(n_4590)
);

INVx2_ASAP7_75t_L g4591 ( 
.A(n_4548),
.Y(n_4591)
);

NAND2xp5_ASAP7_75t_L g4592 ( 
.A(n_4584),
.B(n_4587),
.Y(n_4592)
);

AND2x2_ASAP7_75t_L g4593 ( 
.A(n_4551),
.B(n_4527),
.Y(n_4593)
);

INVx1_ASAP7_75t_L g4594 ( 
.A(n_4551),
.Y(n_4594)
);

INVx2_ASAP7_75t_L g4595 ( 
.A(n_4533),
.Y(n_4595)
);

INVx1_ASAP7_75t_L g4596 ( 
.A(n_4559),
.Y(n_4596)
);

INVx1_ASAP7_75t_L g4597 ( 
.A(n_4559),
.Y(n_4597)
);

INVx2_ASAP7_75t_L g4598 ( 
.A(n_4537),
.Y(n_4598)
);

HB1xp67_ASAP7_75t_L g4599 ( 
.A(n_4549),
.Y(n_4599)
);

NOR2xp33_ASAP7_75t_L g4600 ( 
.A(n_4546),
.B(n_4488),
.Y(n_4600)
);

INVx1_ASAP7_75t_L g4601 ( 
.A(n_4556),
.Y(n_4601)
);

OR2x2_ASAP7_75t_L g4602 ( 
.A(n_4583),
.B(n_4471),
.Y(n_4602)
);

INVx1_ASAP7_75t_L g4603 ( 
.A(n_4571),
.Y(n_4603)
);

HB1xp67_ASAP7_75t_L g4604 ( 
.A(n_4549),
.Y(n_4604)
);

AND2x2_ASAP7_75t_L g4605 ( 
.A(n_4546),
.B(n_4501),
.Y(n_4605)
);

INVx1_ASAP7_75t_L g4606 ( 
.A(n_4571),
.Y(n_4606)
);

AND2x2_ASAP7_75t_L g4607 ( 
.A(n_4562),
.B(n_4502),
.Y(n_4607)
);

INVx1_ASAP7_75t_L g4608 ( 
.A(n_4561),
.Y(n_4608)
);

OR2x2_ASAP7_75t_L g4609 ( 
.A(n_4583),
.B(n_4492),
.Y(n_4609)
);

INVx1_ASAP7_75t_L g4610 ( 
.A(n_4530),
.Y(n_4610)
);

INVx1_ASAP7_75t_L g4611 ( 
.A(n_4530),
.Y(n_4611)
);

INVx2_ASAP7_75t_L g4612 ( 
.A(n_4542),
.Y(n_4612)
);

BUFx3_ASAP7_75t_L g4613 ( 
.A(n_4563),
.Y(n_4613)
);

INVx1_ASAP7_75t_L g4614 ( 
.A(n_4588),
.Y(n_4614)
);

INVx1_ASAP7_75t_L g4615 ( 
.A(n_4532),
.Y(n_4615)
);

AND2x2_ASAP7_75t_L g4616 ( 
.A(n_4562),
.B(n_4472),
.Y(n_4616)
);

NAND2xp5_ASAP7_75t_L g4617 ( 
.A(n_4584),
.B(n_4484),
.Y(n_4617)
);

INVx1_ASAP7_75t_SL g4618 ( 
.A(n_4531),
.Y(n_4618)
);

OR2x2_ASAP7_75t_L g4619 ( 
.A(n_4539),
.B(n_4484),
.Y(n_4619)
);

INVx1_ASAP7_75t_L g4620 ( 
.A(n_4558),
.Y(n_4620)
);

AND2x4_ASAP7_75t_L g4621 ( 
.A(n_4536),
.B(n_4520),
.Y(n_4621)
);

INVx1_ASAP7_75t_L g4622 ( 
.A(n_4566),
.Y(n_4622)
);

AND2x2_ASAP7_75t_L g4623 ( 
.A(n_4578),
.B(n_4465),
.Y(n_4623)
);

OR2x2_ASAP7_75t_L g4624 ( 
.A(n_4544),
.B(n_4514),
.Y(n_4624)
);

NAND2xp5_ASAP7_75t_L g4625 ( 
.A(n_4529),
.B(n_4331),
.Y(n_4625)
);

INVx2_ASAP7_75t_SL g4626 ( 
.A(n_4613),
.Y(n_4626)
);

NAND2xp5_ASAP7_75t_L g4627 ( 
.A(n_4596),
.B(n_4529),
.Y(n_4627)
);

AND2x2_ASAP7_75t_L g4628 ( 
.A(n_4605),
.B(n_4536),
.Y(n_4628)
);

INVx1_ASAP7_75t_L g4629 ( 
.A(n_4599),
.Y(n_4629)
);

INVx2_ASAP7_75t_L g4630 ( 
.A(n_4599),
.Y(n_4630)
);

HB1xp67_ASAP7_75t_L g4631 ( 
.A(n_4604),
.Y(n_4631)
);

NAND2xp5_ASAP7_75t_L g4632 ( 
.A(n_4597),
.B(n_4528),
.Y(n_4632)
);

AND2x4_ASAP7_75t_SL g4633 ( 
.A(n_4616),
.B(n_4538),
.Y(n_4633)
);

AND2x2_ASAP7_75t_L g4634 ( 
.A(n_4607),
.B(n_4564),
.Y(n_4634)
);

OR2x2_ASAP7_75t_L g4635 ( 
.A(n_4602),
.B(n_4534),
.Y(n_4635)
);

OR2x2_ASAP7_75t_L g4636 ( 
.A(n_4609),
.B(n_4547),
.Y(n_4636)
);

INVx2_ASAP7_75t_L g4637 ( 
.A(n_4604),
.Y(n_4637)
);

OR2x2_ASAP7_75t_L g4638 ( 
.A(n_4617),
.B(n_4568),
.Y(n_4638)
);

INVx1_ASAP7_75t_L g4639 ( 
.A(n_4610),
.Y(n_4639)
);

INVx2_ASAP7_75t_L g4640 ( 
.A(n_4594),
.Y(n_4640)
);

INVx1_ASAP7_75t_L g4641 ( 
.A(n_4611),
.Y(n_4641)
);

HB1xp67_ASAP7_75t_L g4642 ( 
.A(n_4590),
.Y(n_4642)
);

INVx1_ASAP7_75t_L g4643 ( 
.A(n_4619),
.Y(n_4643)
);

INVx1_ASAP7_75t_L g4644 ( 
.A(n_4608),
.Y(n_4644)
);

NAND2xp5_ASAP7_75t_L g4645 ( 
.A(n_4614),
.B(n_4528),
.Y(n_4645)
);

NAND2xp5_ASAP7_75t_L g4646 ( 
.A(n_4617),
.B(n_4569),
.Y(n_4646)
);

INVx2_ASAP7_75t_L g4647 ( 
.A(n_4591),
.Y(n_4647)
);

AND2x2_ASAP7_75t_L g4648 ( 
.A(n_4621),
.B(n_4564),
.Y(n_4648)
);

INVx1_ASAP7_75t_L g4649 ( 
.A(n_4601),
.Y(n_4649)
);

INVx1_ASAP7_75t_L g4650 ( 
.A(n_4620),
.Y(n_4650)
);

AND2x2_ASAP7_75t_L g4651 ( 
.A(n_4621),
.B(n_4567),
.Y(n_4651)
);

INVx2_ASAP7_75t_L g4652 ( 
.A(n_4593),
.Y(n_4652)
);

INVx1_ASAP7_75t_L g4653 ( 
.A(n_4622),
.Y(n_4653)
);

NAND2xp5_ASAP7_75t_SL g4654 ( 
.A(n_4600),
.B(n_4618),
.Y(n_4654)
);

NAND4xp75_ASAP7_75t_L g4655 ( 
.A(n_4600),
.B(n_4582),
.C(n_4552),
.D(n_4625),
.Y(n_4655)
);

NAND2xp5_ASAP7_75t_L g4656 ( 
.A(n_4592),
.B(n_4575),
.Y(n_4656)
);

INVxp67_ASAP7_75t_L g4657 ( 
.A(n_4618),
.Y(n_4657)
);

O2A1O1Ixp33_ASAP7_75t_L g4658 ( 
.A1(n_4625),
.A2(n_4543),
.B(n_4582),
.C(n_4603),
.Y(n_4658)
);

AND2x2_ASAP7_75t_L g4659 ( 
.A(n_4623),
.B(n_4540),
.Y(n_4659)
);

INVx1_ASAP7_75t_L g4660 ( 
.A(n_4615),
.Y(n_4660)
);

AND2x2_ASAP7_75t_L g4661 ( 
.A(n_4624),
.B(n_4545),
.Y(n_4661)
);

OAI22xp33_ASAP7_75t_L g4662 ( 
.A1(n_4606),
.A2(n_4555),
.B1(n_4577),
.B2(n_4589),
.Y(n_4662)
);

INVx1_ASAP7_75t_L g4663 ( 
.A(n_4595),
.Y(n_4663)
);

AND2x4_ASAP7_75t_SL g4664 ( 
.A(n_4612),
.B(n_4557),
.Y(n_4664)
);

NAND2xp5_ASAP7_75t_L g4665 ( 
.A(n_4592),
.B(n_4574),
.Y(n_4665)
);

INVx1_ASAP7_75t_SL g4666 ( 
.A(n_4598),
.Y(n_4666)
);

NOR2xp33_ASAP7_75t_SL g4667 ( 
.A(n_4618),
.B(n_4570),
.Y(n_4667)
);

OAI22xp5_ASAP7_75t_SL g4668 ( 
.A1(n_4613),
.A2(n_4543),
.B1(n_4306),
.B2(n_4572),
.Y(n_4668)
);

INVx2_ASAP7_75t_L g4669 ( 
.A(n_4599),
.Y(n_4669)
);

INVx2_ASAP7_75t_L g4670 ( 
.A(n_4599),
.Y(n_4670)
);

INVx1_ASAP7_75t_L g4671 ( 
.A(n_4599),
.Y(n_4671)
);

AND2x2_ASAP7_75t_L g4672 ( 
.A(n_4605),
.B(n_4541),
.Y(n_4672)
);

OAI21xp33_ASAP7_75t_SL g4673 ( 
.A1(n_4654),
.A2(n_4570),
.B(n_4586),
.Y(n_4673)
);

AND2x2_ASAP7_75t_L g4674 ( 
.A(n_4628),
.B(n_4550),
.Y(n_4674)
);

INVx1_ASAP7_75t_L g4675 ( 
.A(n_4631),
.Y(n_4675)
);

INVx1_ASAP7_75t_L g4676 ( 
.A(n_4629),
.Y(n_4676)
);

NOR2xp33_ASAP7_75t_L g4677 ( 
.A(n_4626),
.B(n_4576),
.Y(n_4677)
);

NAND2xp5_ASAP7_75t_L g4678 ( 
.A(n_4657),
.B(n_4665),
.Y(n_4678)
);

NOR2x1_ASAP7_75t_L g4679 ( 
.A(n_4655),
.B(n_4573),
.Y(n_4679)
);

INVx1_ASAP7_75t_L g4680 ( 
.A(n_4671),
.Y(n_4680)
);

INVx1_ASAP7_75t_L g4681 ( 
.A(n_4630),
.Y(n_4681)
);

NAND2xp5_ASAP7_75t_L g4682 ( 
.A(n_4643),
.B(n_4580),
.Y(n_4682)
);

OR2x2_ASAP7_75t_L g4683 ( 
.A(n_4638),
.B(n_4581),
.Y(n_4683)
);

AND2x2_ASAP7_75t_L g4684 ( 
.A(n_4633),
.B(n_4648),
.Y(n_4684)
);

INVx1_ASAP7_75t_L g4685 ( 
.A(n_4637),
.Y(n_4685)
);

OR2x2_ASAP7_75t_L g4686 ( 
.A(n_4646),
.B(n_4585),
.Y(n_4686)
);

NAND2xp5_ASAP7_75t_L g4687 ( 
.A(n_4658),
.B(n_4580),
.Y(n_4687)
);

NAND2xp5_ASAP7_75t_L g4688 ( 
.A(n_4644),
.B(n_4572),
.Y(n_4688)
);

NAND2xp5_ASAP7_75t_L g4689 ( 
.A(n_4669),
.B(n_4574),
.Y(n_4689)
);

INVx1_ASAP7_75t_L g4690 ( 
.A(n_4670),
.Y(n_4690)
);

INVx1_ASAP7_75t_L g4691 ( 
.A(n_4635),
.Y(n_4691)
);

NAND2xp5_ASAP7_75t_SL g4692 ( 
.A(n_4667),
.B(n_4495),
.Y(n_4692)
);

INVx2_ASAP7_75t_SL g4693 ( 
.A(n_4664),
.Y(n_4693)
);

NAND2xp5_ASAP7_75t_L g4694 ( 
.A(n_4649),
.B(n_4579),
.Y(n_4694)
);

AND2x4_ASAP7_75t_L g4695 ( 
.A(n_4661),
.B(n_4535),
.Y(n_4695)
);

INVx1_ASAP7_75t_L g4696 ( 
.A(n_4636),
.Y(n_4696)
);

NOR2xp33_ASAP7_75t_L g4697 ( 
.A(n_4667),
.B(n_4565),
.Y(n_4697)
);

INVxp67_ASAP7_75t_SL g4698 ( 
.A(n_4645),
.Y(n_4698)
);

NAND2xp5_ASAP7_75t_L g4699 ( 
.A(n_4660),
.B(n_4573),
.Y(n_4699)
);

OR2x2_ASAP7_75t_L g4700 ( 
.A(n_4646),
.B(n_4554),
.Y(n_4700)
);

INVx1_ASAP7_75t_L g4701 ( 
.A(n_4650),
.Y(n_4701)
);

INVx2_ASAP7_75t_L g4702 ( 
.A(n_4652),
.Y(n_4702)
);

OR2x2_ASAP7_75t_L g4703 ( 
.A(n_4656),
.B(n_4560),
.Y(n_4703)
);

AND2x2_ASAP7_75t_L g4704 ( 
.A(n_4634),
.B(n_4651),
.Y(n_4704)
);

INVx1_ASAP7_75t_SL g4705 ( 
.A(n_4666),
.Y(n_4705)
);

NAND2xp5_ASAP7_75t_L g4706 ( 
.A(n_4666),
.B(n_4553),
.Y(n_4706)
);

INVx1_ASAP7_75t_L g4707 ( 
.A(n_4653),
.Y(n_4707)
);

NAND2xp33_ASAP7_75t_SL g4708 ( 
.A(n_4668),
.B(n_4522),
.Y(n_4708)
);

INVx1_ASAP7_75t_L g4709 ( 
.A(n_4639),
.Y(n_4709)
);

AND2x4_ASAP7_75t_L g4710 ( 
.A(n_4659),
.B(n_4647),
.Y(n_4710)
);

INVx1_ASAP7_75t_L g4711 ( 
.A(n_4641),
.Y(n_4711)
);

NOR2xp33_ASAP7_75t_L g4712 ( 
.A(n_4668),
.B(n_4495),
.Y(n_4712)
);

NAND2xp5_ASAP7_75t_L g4713 ( 
.A(n_4656),
.B(n_4495),
.Y(n_4713)
);

INVx1_ASAP7_75t_L g4714 ( 
.A(n_4642),
.Y(n_4714)
);

NAND2xp5_ASAP7_75t_L g4715 ( 
.A(n_4663),
.B(n_4331),
.Y(n_4715)
);

HB1xp67_ASAP7_75t_L g4716 ( 
.A(n_4640),
.Y(n_4716)
);

INVx1_ASAP7_75t_L g4717 ( 
.A(n_4632),
.Y(n_4717)
);

OR2x2_ASAP7_75t_L g4718 ( 
.A(n_4627),
.B(n_4316),
.Y(n_4718)
);

INVx1_ASAP7_75t_L g4719 ( 
.A(n_4632),
.Y(n_4719)
);

AND2x2_ASAP7_75t_L g4720 ( 
.A(n_4672),
.B(n_4316),
.Y(n_4720)
);

INVx1_ASAP7_75t_L g4721 ( 
.A(n_4645),
.Y(n_4721)
);

NAND2xp5_ASAP7_75t_L g4722 ( 
.A(n_4627),
.B(n_3851),
.Y(n_4722)
);

AND2x2_ASAP7_75t_L g4723 ( 
.A(n_4684),
.B(n_4662),
.Y(n_4723)
);

INVx1_ASAP7_75t_L g4724 ( 
.A(n_4714),
.Y(n_4724)
);

AOI321xp33_ASAP7_75t_L g4725 ( 
.A1(n_4687),
.A2(n_3869),
.A3(n_3969),
.B1(n_3954),
.B2(n_4015),
.C(n_3833),
.Y(n_4725)
);

INVx2_ASAP7_75t_L g4726 ( 
.A(n_4710),
.Y(n_4726)
);

INVx1_ASAP7_75t_SL g4727 ( 
.A(n_4705),
.Y(n_4727)
);

INVx1_ASAP7_75t_SL g4728 ( 
.A(n_4675),
.Y(n_4728)
);

INVxp67_ASAP7_75t_L g4729 ( 
.A(n_4678),
.Y(n_4729)
);

OAI22xp5_ASAP7_75t_L g4730 ( 
.A1(n_4692),
.A2(n_4209),
.B1(n_4130),
.B2(n_4188),
.Y(n_4730)
);

XNOR2xp5_ASAP7_75t_L g4731 ( 
.A(n_4693),
.B(n_656),
.Y(n_4731)
);

AOI22xp5_ASAP7_75t_L g4732 ( 
.A1(n_4673),
.A2(n_3759),
.B1(n_4161),
.B2(n_4140),
.Y(n_4732)
);

AOI32xp33_ASAP7_75t_L g4733 ( 
.A1(n_4679),
.A2(n_4198),
.A3(n_4122),
.B1(n_4193),
.B2(n_3997),
.Y(n_4733)
);

OAI22xp5_ASAP7_75t_L g4734 ( 
.A1(n_4712),
.A2(n_3838),
.B1(n_3871),
.B2(n_3849),
.Y(n_4734)
);

NAND2xp5_ASAP7_75t_SL g4735 ( 
.A(n_4708),
.B(n_3275),
.Y(n_4735)
);

OAI32xp33_ASAP7_75t_L g4736 ( 
.A1(n_4682),
.A2(n_4302),
.A3(n_3851),
.B1(n_3910),
.B2(n_3900),
.Y(n_4736)
);

INVxp67_ASAP7_75t_L g4737 ( 
.A(n_4677),
.Y(n_4737)
);

OAI22xp5_ASAP7_75t_L g4738 ( 
.A1(n_4697),
.A2(n_4302),
.B1(n_3778),
.B2(n_3757),
.Y(n_4738)
);

OAI22xp5_ASAP7_75t_L g4739 ( 
.A1(n_4695),
.A2(n_3716),
.B1(n_3722),
.B2(n_3719),
.Y(n_4739)
);

OAI221xp5_ASAP7_75t_L g4740 ( 
.A1(n_4689),
.A2(n_3698),
.B1(n_3885),
.B2(n_3907),
.C(n_3884),
.Y(n_4740)
);

INVx1_ASAP7_75t_L g4741 ( 
.A(n_4691),
.Y(n_4741)
);

INVx1_ASAP7_75t_L g4742 ( 
.A(n_4696),
.Y(n_4742)
);

NAND2xp5_ASAP7_75t_L g4743 ( 
.A(n_4676),
.B(n_3863),
.Y(n_4743)
);

AND2x2_ASAP7_75t_L g4744 ( 
.A(n_4704),
.B(n_3793),
.Y(n_4744)
);

NAND2xp5_ASAP7_75t_L g4745 ( 
.A(n_4680),
.B(n_3781),
.Y(n_4745)
);

NAND2xp5_ASAP7_75t_L g4746 ( 
.A(n_4688),
.B(n_3806),
.Y(n_4746)
);

AOI221xp5_ASAP7_75t_L g4747 ( 
.A1(n_4717),
.A2(n_3949),
.B1(n_3771),
.B2(n_3724),
.C(n_3752),
.Y(n_4747)
);

AOI22xp33_ASAP7_75t_SL g4748 ( 
.A1(n_4695),
.A2(n_4698),
.B1(n_4719),
.B2(n_4721),
.Y(n_4748)
);

A2O1A1Ixp33_ASAP7_75t_L g4749 ( 
.A1(n_4713),
.A2(n_3748),
.B(n_3750),
.C(n_3725),
.Y(n_4749)
);

OR2x2_ASAP7_75t_L g4750 ( 
.A(n_4681),
.B(n_4685),
.Y(n_4750)
);

INVx1_ASAP7_75t_L g4751 ( 
.A(n_4750),
.Y(n_4751)
);

NAND2xp5_ASAP7_75t_SL g4752 ( 
.A(n_4727),
.B(n_4690),
.Y(n_4752)
);

INVx1_ASAP7_75t_L g4753 ( 
.A(n_4731),
.Y(n_4753)
);

INVxp33_ASAP7_75t_L g4754 ( 
.A(n_4748),
.Y(n_4754)
);

INVx1_ASAP7_75t_L g4755 ( 
.A(n_4724),
.Y(n_4755)
);

AOI322xp5_ASAP7_75t_L g4756 ( 
.A1(n_4729),
.A2(n_4710),
.A3(n_4716),
.B1(n_4702),
.B2(n_4720),
.C1(n_4711),
.C2(n_4709),
.Y(n_4756)
);

OAI21xp5_ASAP7_75t_L g4757 ( 
.A1(n_4737),
.A2(n_4722),
.B(n_4707),
.Y(n_4757)
);

AND2x4_ASAP7_75t_L g4758 ( 
.A(n_4726),
.B(n_4674),
.Y(n_4758)
);

NAND2xp5_ASAP7_75t_L g4759 ( 
.A(n_4733),
.B(n_4701),
.Y(n_4759)
);

AND2x2_ASAP7_75t_SL g4760 ( 
.A(n_4723),
.B(n_4741),
.Y(n_4760)
);

NAND2x1_ASAP7_75t_L g4761 ( 
.A(n_4742),
.B(n_4706),
.Y(n_4761)
);

OAI22xp5_ASAP7_75t_L g4762 ( 
.A1(n_4728),
.A2(n_4694),
.B1(n_4686),
.B2(n_4683),
.Y(n_4762)
);

NAND2xp5_ASAP7_75t_L g4763 ( 
.A(n_4732),
.B(n_4703),
.Y(n_4763)
);

NOR2xp33_ASAP7_75t_SL g4764 ( 
.A(n_4730),
.B(n_4700),
.Y(n_4764)
);

NAND2xp5_ASAP7_75t_L g4765 ( 
.A(n_4746),
.B(n_4715),
.Y(n_4765)
);

AOI21xp33_ASAP7_75t_L g4766 ( 
.A1(n_4738),
.A2(n_4699),
.B(n_4718),
.Y(n_4766)
);

NAND2xp5_ASAP7_75t_L g4767 ( 
.A(n_4743),
.B(n_656),
.Y(n_4767)
);

AOI21xp33_ASAP7_75t_L g4768 ( 
.A1(n_4745),
.A2(n_4735),
.B(n_4739),
.Y(n_4768)
);

AOI21xp5_ASAP7_75t_L g4769 ( 
.A1(n_4734),
.A2(n_4362),
.B(n_3761),
.Y(n_4769)
);

NAND2xp5_ASAP7_75t_L g4770 ( 
.A(n_4744),
.B(n_657),
.Y(n_4770)
);

OAI211xp5_ASAP7_75t_L g4771 ( 
.A1(n_4725),
.A2(n_3791),
.B(n_660),
.C(n_658),
.Y(n_4771)
);

INVx1_ASAP7_75t_L g4772 ( 
.A(n_4725),
.Y(n_4772)
);

AOI322xp5_ASAP7_75t_L g4773 ( 
.A1(n_4747),
.A2(n_3691),
.A3(n_3765),
.B1(n_4221),
.B2(n_3728),
.C1(n_3767),
.C2(n_661),
.Y(n_4773)
);

AND2x2_ASAP7_75t_L g4774 ( 
.A(n_4749),
.B(n_659),
.Y(n_4774)
);

OA22x2_ASAP7_75t_L g4775 ( 
.A1(n_4736),
.A2(n_4247),
.B1(n_3768),
.B2(n_3772),
.Y(n_4775)
);

INVx1_ASAP7_75t_L g4776 ( 
.A(n_4740),
.Y(n_4776)
);

INVx1_ASAP7_75t_SL g4777 ( 
.A(n_4727),
.Y(n_4777)
);

OR2x2_ASAP7_75t_L g4778 ( 
.A(n_4727),
.B(n_659),
.Y(n_4778)
);

AOI22xp5_ASAP7_75t_L g4779 ( 
.A1(n_4727),
.A2(n_3709),
.B1(n_4333),
.B2(n_3763),
.Y(n_4779)
);

AND2x4_ASAP7_75t_L g4780 ( 
.A(n_4727),
.B(n_659),
.Y(n_4780)
);

INVxp67_ASAP7_75t_L g4781 ( 
.A(n_4731),
.Y(n_4781)
);

INVx1_ASAP7_75t_L g4782 ( 
.A(n_4750),
.Y(n_4782)
);

AND2x2_ASAP7_75t_L g4783 ( 
.A(n_4723),
.B(n_660),
.Y(n_4783)
);

INVx1_ASAP7_75t_L g4784 ( 
.A(n_4750),
.Y(n_4784)
);

NAND2xp5_ASAP7_75t_L g4785 ( 
.A(n_4727),
.B(n_660),
.Y(n_4785)
);

OAI21xp33_ASAP7_75t_SL g4786 ( 
.A1(n_4723),
.A2(n_4327),
.B(n_3739),
.Y(n_4786)
);

NAND2xp5_ASAP7_75t_L g4787 ( 
.A(n_4777),
.B(n_661),
.Y(n_4787)
);

INVx1_ASAP7_75t_L g4788 ( 
.A(n_4780),
.Y(n_4788)
);

NOR3xp33_ASAP7_75t_SL g4789 ( 
.A(n_4772),
.B(n_661),
.C(n_662),
.Y(n_4789)
);

INVx1_ASAP7_75t_SL g4790 ( 
.A(n_4780),
.Y(n_4790)
);

INVx1_ASAP7_75t_SL g4791 ( 
.A(n_4778),
.Y(n_4791)
);

AOI221xp5_ASAP7_75t_L g4792 ( 
.A1(n_4754),
.A2(n_664),
.B1(n_662),
.B2(n_663),
.C(n_665),
.Y(n_4792)
);

AOI22xp5_ASAP7_75t_L g4793 ( 
.A1(n_4764),
.A2(n_4333),
.B1(n_3738),
.B2(n_3354),
.Y(n_4793)
);

INVx1_ASAP7_75t_L g4794 ( 
.A(n_4785),
.Y(n_4794)
);

INVx3_ASAP7_75t_L g4795 ( 
.A(n_4758),
.Y(n_4795)
);

AOI22xp5_ASAP7_75t_L g4796 ( 
.A1(n_4783),
.A2(n_3354),
.B1(n_3423),
.B2(n_3309),
.Y(n_4796)
);

CKINVDCx5p33_ASAP7_75t_R g4797 ( 
.A(n_4781),
.Y(n_4797)
);

NOR2xp33_ASAP7_75t_L g4798 ( 
.A(n_4753),
.B(n_663),
.Y(n_4798)
);

INVxp67_ASAP7_75t_SL g4799 ( 
.A(n_4767),
.Y(n_4799)
);

INVx1_ASAP7_75t_L g4800 ( 
.A(n_4751),
.Y(n_4800)
);

NAND2xp5_ASAP7_75t_L g4801 ( 
.A(n_4756),
.B(n_666),
.Y(n_4801)
);

AND2x2_ASAP7_75t_L g4802 ( 
.A(n_4758),
.B(n_666),
.Y(n_4802)
);

NAND2xp5_ASAP7_75t_L g4803 ( 
.A(n_4776),
.B(n_666),
.Y(n_4803)
);

INVx2_ASAP7_75t_L g4804 ( 
.A(n_4752),
.Y(n_4804)
);

OR2x2_ASAP7_75t_L g4805 ( 
.A(n_4782),
.B(n_4784),
.Y(n_4805)
);

AOI21xp5_ASAP7_75t_L g4806 ( 
.A1(n_4760),
.A2(n_667),
.B(n_668),
.Y(n_4806)
);

INVx1_ASAP7_75t_L g4807 ( 
.A(n_4770),
.Y(n_4807)
);

INVx2_ASAP7_75t_L g4808 ( 
.A(n_4775),
.Y(n_4808)
);

AO21x2_ASAP7_75t_L g4809 ( 
.A1(n_4759),
.A2(n_668),
.B(n_669),
.Y(n_4809)
);

AND2x4_ASAP7_75t_L g4810 ( 
.A(n_4755),
.B(n_669),
.Y(n_4810)
);

AOI211xp5_ASAP7_75t_SL g4811 ( 
.A1(n_4771),
.A2(n_671),
.B(n_669),
.C(n_670),
.Y(n_4811)
);

OAI32xp33_ASAP7_75t_L g4812 ( 
.A1(n_4763),
.A2(n_672),
.A3(n_670),
.B1(n_671),
.B2(n_673),
.Y(n_4812)
);

OAI21xp5_ASAP7_75t_L g4813 ( 
.A1(n_4768),
.A2(n_671),
.B(n_672),
.Y(n_4813)
);

INVx1_ASAP7_75t_L g4814 ( 
.A(n_4762),
.Y(n_4814)
);

NAND2xp5_ASAP7_75t_L g4815 ( 
.A(n_4774),
.B(n_672),
.Y(n_4815)
);

INVx1_ASAP7_75t_L g4816 ( 
.A(n_4765),
.Y(n_4816)
);

NOR2xp33_ASAP7_75t_L g4817 ( 
.A(n_4761),
.B(n_673),
.Y(n_4817)
);

INVx1_ASAP7_75t_SL g4818 ( 
.A(n_4766),
.Y(n_4818)
);

OAI221xp5_ASAP7_75t_SL g4819 ( 
.A1(n_4786),
.A2(n_675),
.B1(n_673),
.B2(n_674),
.C(n_676),
.Y(n_4819)
);

INVx1_ASAP7_75t_L g4820 ( 
.A(n_4757),
.Y(n_4820)
);

NAND2xp5_ASAP7_75t_L g4821 ( 
.A(n_4769),
.B(n_674),
.Y(n_4821)
);

NAND2xp5_ASAP7_75t_L g4822 ( 
.A(n_4795),
.B(n_4779),
.Y(n_4822)
);

NAND4xp25_ASAP7_75t_L g4823 ( 
.A(n_4814),
.B(n_4773),
.C(n_676),
.D(n_674),
.Y(n_4823)
);

NOR2xp33_ASAP7_75t_L g4824 ( 
.A(n_4790),
.B(n_675),
.Y(n_4824)
);

AOI22xp33_ASAP7_75t_SL g4825 ( 
.A1(n_4818),
.A2(n_3431),
.B1(n_3423),
.B2(n_3440),
.Y(n_4825)
);

NOR2xp33_ASAP7_75t_L g4826 ( 
.A(n_4801),
.B(n_675),
.Y(n_4826)
);

NOR2xp33_ASAP7_75t_L g4827 ( 
.A(n_4797),
.B(n_676),
.Y(n_4827)
);

OAI221xp5_ASAP7_75t_L g4828 ( 
.A1(n_4811),
.A2(n_679),
.B1(n_677),
.B2(n_678),
.C(n_680),
.Y(n_4828)
);

INVxp67_ASAP7_75t_L g4829 ( 
.A(n_4817),
.Y(n_4829)
);

NOR3xp33_ASAP7_75t_L g4830 ( 
.A(n_4792),
.B(n_677),
.C(n_678),
.Y(n_4830)
);

NOR2xp33_ASAP7_75t_SL g4831 ( 
.A(n_4802),
.B(n_3423),
.Y(n_4831)
);

NOR2x1_ASAP7_75t_L g4832 ( 
.A(n_4787),
.B(n_677),
.Y(n_4832)
);

NAND3xp33_ASAP7_75t_L g4833 ( 
.A(n_4798),
.B(n_678),
.C(n_679),
.Y(n_4833)
);

NOR2x1p5_ASAP7_75t_L g4834 ( 
.A(n_4804),
.B(n_679),
.Y(n_4834)
);

NAND2xp5_ASAP7_75t_L g4835 ( 
.A(n_4789),
.B(n_680),
.Y(n_4835)
);

INVxp67_ASAP7_75t_L g4836 ( 
.A(n_4815),
.Y(n_4836)
);

OAI21xp5_ASAP7_75t_L g4837 ( 
.A1(n_4806),
.A2(n_680),
.B(n_681),
.Y(n_4837)
);

NAND3xp33_ASAP7_75t_SL g4838 ( 
.A(n_4813),
.B(n_681),
.C(n_682),
.Y(n_4838)
);

NOR2xp33_ASAP7_75t_L g4839 ( 
.A(n_4788),
.B(n_682),
.Y(n_4839)
);

NAND2xp5_ASAP7_75t_L g4840 ( 
.A(n_4810),
.B(n_683),
.Y(n_4840)
);

OAI21xp5_ASAP7_75t_L g4841 ( 
.A1(n_4803),
.A2(n_683),
.B(n_684),
.Y(n_4841)
);

NAND2xp5_ASAP7_75t_L g4842 ( 
.A(n_4810),
.B(n_683),
.Y(n_4842)
);

INVx1_ASAP7_75t_L g4843 ( 
.A(n_4805),
.Y(n_4843)
);

NOR2xp33_ASAP7_75t_SL g4844 ( 
.A(n_4791),
.B(n_4800),
.Y(n_4844)
);

NAND2xp5_ASAP7_75t_L g4845 ( 
.A(n_4809),
.B(n_684),
.Y(n_4845)
);

NOR2x1_ASAP7_75t_L g4846 ( 
.A(n_4821),
.B(n_685),
.Y(n_4846)
);

AOI221xp5_ASAP7_75t_L g4847 ( 
.A1(n_4819),
.A2(n_687),
.B1(n_685),
.B2(n_686),
.C(n_688),
.Y(n_4847)
);

INVx1_ASAP7_75t_L g4848 ( 
.A(n_4812),
.Y(n_4848)
);

NOR2xp33_ASAP7_75t_L g4849 ( 
.A(n_4820),
.B(n_685),
.Y(n_4849)
);

NAND4xp75_ASAP7_75t_L g4850 ( 
.A(n_4816),
.B(n_688),
.C(n_686),
.D(n_687),
.Y(n_4850)
);

INVx2_ASAP7_75t_L g4851 ( 
.A(n_4808),
.Y(n_4851)
);

NOR2xp33_ASAP7_75t_L g4852 ( 
.A(n_4807),
.B(n_687),
.Y(n_4852)
);

AOI21xp5_ASAP7_75t_L g4853 ( 
.A1(n_4799),
.A2(n_688),
.B(n_689),
.Y(n_4853)
);

OAI21xp33_ASAP7_75t_L g4854 ( 
.A1(n_4794),
.A2(n_689),
.B(n_690),
.Y(n_4854)
);

NOR3xp33_ASAP7_75t_L g4855 ( 
.A(n_4793),
.B(n_689),
.C(n_690),
.Y(n_4855)
);

XNOR2xp5_ASAP7_75t_L g4856 ( 
.A(n_4796),
.B(n_691),
.Y(n_4856)
);

HB1xp67_ASAP7_75t_L g4857 ( 
.A(n_4797),
.Y(n_4857)
);

INVx1_ASAP7_75t_L g4858 ( 
.A(n_4802),
.Y(n_4858)
);

INVx1_ASAP7_75t_L g4859 ( 
.A(n_4802),
.Y(n_4859)
);

OAI22xp5_ASAP7_75t_L g4860 ( 
.A1(n_4857),
.A2(n_3431),
.B1(n_3472),
.B2(n_3440),
.Y(n_4860)
);

AOI211xp5_ASAP7_75t_L g4861 ( 
.A1(n_4828),
.A2(n_694),
.B(n_692),
.C(n_693),
.Y(n_4861)
);

AOI22x1_ASAP7_75t_SL g4862 ( 
.A1(n_4848),
.A2(n_694),
.B1(n_692),
.B2(n_693),
.Y(n_4862)
);

NOR3xp33_ASAP7_75t_L g4863 ( 
.A(n_4827),
.B(n_693),
.C(n_695),
.Y(n_4863)
);

O2A1O1Ixp33_ASAP7_75t_L g4864 ( 
.A1(n_4845),
.A2(n_697),
.B(n_695),
.C(n_696),
.Y(n_4864)
);

AOI211xp5_ASAP7_75t_SL g4865 ( 
.A1(n_4849),
.A2(n_697),
.B(n_695),
.C(n_696),
.Y(n_4865)
);

AOI221xp5_ASAP7_75t_L g4866 ( 
.A1(n_4823),
.A2(n_700),
.B1(n_698),
.B2(n_699),
.C(n_701),
.Y(n_4866)
);

NAND4xp25_ASAP7_75t_SL g4867 ( 
.A(n_4843),
.B(n_700),
.C(n_698),
.D(n_699),
.Y(n_4867)
);

AOI221xp5_ASAP7_75t_L g4868 ( 
.A1(n_4851),
.A2(n_700),
.B1(n_698),
.B2(n_699),
.C(n_701),
.Y(n_4868)
);

AOI21xp5_ASAP7_75t_L g4869 ( 
.A1(n_4835),
.A2(n_4853),
.B(n_4838),
.Y(n_4869)
);

AOI221xp5_ASAP7_75t_L g4870 ( 
.A1(n_4829),
.A2(n_703),
.B1(n_701),
.B2(n_702),
.C(n_704),
.Y(n_4870)
);

OAI22xp33_ASAP7_75t_L g4871 ( 
.A1(n_4844),
.A2(n_3431),
.B1(n_3472),
.B2(n_3440),
.Y(n_4871)
);

AND4x1_ASAP7_75t_L g4872 ( 
.A(n_4824),
.B(n_704),
.C(n_702),
.D(n_703),
.Y(n_4872)
);

OAI211xp5_ASAP7_75t_SL g4873 ( 
.A1(n_4836),
.A2(n_706),
.B(n_703),
.C(n_705),
.Y(n_4873)
);

INVx1_ASAP7_75t_L g4874 ( 
.A(n_4840),
.Y(n_4874)
);

NAND3xp33_ASAP7_75t_L g4875 ( 
.A(n_4826),
.B(n_705),
.C(n_706),
.Y(n_4875)
);

AOI211xp5_ASAP7_75t_L g4876 ( 
.A1(n_4837),
.A2(n_707),
.B(n_705),
.C(n_706),
.Y(n_4876)
);

AOI22xp5_ASAP7_75t_L g4877 ( 
.A1(n_4830),
.A2(n_3472),
.B1(n_3559),
.B2(n_3557),
.Y(n_4877)
);

NAND2xp5_ASAP7_75t_L g4878 ( 
.A(n_4847),
.B(n_707),
.Y(n_4878)
);

NAND2xp5_ASAP7_75t_L g4879 ( 
.A(n_4839),
.B(n_707),
.Y(n_4879)
);

NAND3xp33_ASAP7_75t_L g4880 ( 
.A(n_4852),
.B(n_733),
.C(n_734),
.Y(n_4880)
);

NAND2xp5_ASAP7_75t_SL g4881 ( 
.A(n_4854),
.B(n_3557),
.Y(n_4881)
);

AOI22xp33_ASAP7_75t_L g4882 ( 
.A1(n_4855),
.A2(n_3559),
.B1(n_3597),
.B2(n_3557),
.Y(n_4882)
);

NAND2xp5_ASAP7_75t_L g4883 ( 
.A(n_4850),
.B(n_734),
.Y(n_4883)
);

AOI22xp5_ASAP7_75t_L g4884 ( 
.A1(n_4866),
.A2(n_4831),
.B1(n_4859),
.B2(n_4858),
.Y(n_4884)
);

INVx1_ASAP7_75t_L g4885 ( 
.A(n_4862),
.Y(n_4885)
);

INVx1_ASAP7_75t_L g4886 ( 
.A(n_4883),
.Y(n_4886)
);

OR3x1_ASAP7_75t_L g4887 ( 
.A(n_4873),
.B(n_4834),
.C(n_4846),
.Y(n_4887)
);

OAI221xp5_ASAP7_75t_L g4888 ( 
.A1(n_4861),
.A2(n_4868),
.B1(n_4876),
.B2(n_4863),
.C(n_4870),
.Y(n_4888)
);

HB1xp67_ASAP7_75t_L g4889 ( 
.A(n_4872),
.Y(n_4889)
);

OAI21xp5_ASAP7_75t_L g4890 ( 
.A1(n_4869),
.A2(n_4832),
.B(n_4822),
.Y(n_4890)
);

AND2x2_ASAP7_75t_L g4891 ( 
.A(n_4865),
.B(n_4841),
.Y(n_4891)
);

XNOR2xp5_ASAP7_75t_L g4892 ( 
.A(n_4875),
.B(n_4856),
.Y(n_4892)
);

AOI211xp5_ASAP7_75t_L g4893 ( 
.A1(n_4864),
.A2(n_4833),
.B(n_4842),
.C(n_4825),
.Y(n_4893)
);

AOI211xp5_ASAP7_75t_SL g4894 ( 
.A1(n_4878),
.A2(n_737),
.B(n_735),
.C(n_736),
.Y(n_4894)
);

NAND4xp75_ASAP7_75t_L g4895 ( 
.A(n_4874),
.B(n_737),
.C(n_735),
.D(n_736),
.Y(n_4895)
);

INVx1_ASAP7_75t_L g4896 ( 
.A(n_4879),
.Y(n_4896)
);

AOI211xp5_ASAP7_75t_L g4897 ( 
.A1(n_4867),
.A2(n_741),
.B(n_738),
.C(n_739),
.Y(n_4897)
);

AOI221xp5_ASAP7_75t_L g4898 ( 
.A1(n_4871),
.A2(n_3649),
.B1(n_3688),
.B2(n_3597),
.C(n_3559),
.Y(n_4898)
);

HB1xp67_ASAP7_75t_L g4899 ( 
.A(n_4881),
.Y(n_4899)
);

NOR2xp33_ASAP7_75t_L g4900 ( 
.A(n_4880),
.B(n_738),
.Y(n_4900)
);

NAND4xp25_ASAP7_75t_L g4901 ( 
.A(n_4877),
.B(n_744),
.C(n_739),
.D(n_743),
.Y(n_4901)
);

AOI222xp33_ASAP7_75t_L g4902 ( 
.A1(n_4860),
.A2(n_745),
.B1(n_747),
.B2(n_743),
.C1(n_744),
.C2(n_746),
.Y(n_4902)
);

OAI221xp5_ASAP7_75t_L g4903 ( 
.A1(n_4882),
.A2(n_749),
.B1(n_745),
.B2(n_747),
.C(n_750),
.Y(n_4903)
);

OAI21xp33_ASAP7_75t_L g4904 ( 
.A1(n_4866),
.A2(n_750),
.B(n_751),
.Y(n_4904)
);

AOI211xp5_ASAP7_75t_L g4905 ( 
.A1(n_4866),
.A2(n_753),
.B(n_751),
.C(n_752),
.Y(n_4905)
);

AOI221xp5_ASAP7_75t_L g4906 ( 
.A1(n_4866),
.A2(n_3688),
.B1(n_3649),
.B2(n_3597),
.C(n_754),
.Y(n_4906)
);

NAND2xp5_ASAP7_75t_L g4907 ( 
.A(n_4865),
.B(n_752),
.Y(n_4907)
);

INVx2_ASAP7_75t_L g4908 ( 
.A(n_4895),
.Y(n_4908)
);

OR2x2_ASAP7_75t_L g4909 ( 
.A(n_4907),
.B(n_753),
.Y(n_4909)
);

NAND2x1p5_ASAP7_75t_L g4910 ( 
.A(n_4885),
.B(n_3649),
.Y(n_4910)
);

AND2x4_ASAP7_75t_L g4911 ( 
.A(n_4899),
.B(n_754),
.Y(n_4911)
);

AND2x4_ASAP7_75t_L g4912 ( 
.A(n_4890),
.B(n_755),
.Y(n_4912)
);

NAND2xp5_ASAP7_75t_L g4913 ( 
.A(n_4897),
.B(n_755),
.Y(n_4913)
);

OAI22xp5_ASAP7_75t_L g4914 ( 
.A1(n_4887),
.A2(n_3688),
.B1(n_758),
.B2(n_756),
.Y(n_4914)
);

INVx1_ASAP7_75t_L g4915 ( 
.A(n_4889),
.Y(n_4915)
);

NOR2x1p5_ASAP7_75t_L g4916 ( 
.A(n_4901),
.B(n_757),
.Y(n_4916)
);

NAND2x1p5_ASAP7_75t_L g4917 ( 
.A(n_4886),
.B(n_757),
.Y(n_4917)
);

INVx1_ASAP7_75t_L g4918 ( 
.A(n_4891),
.Y(n_4918)
);

NOR2x1_ASAP7_75t_L g4919 ( 
.A(n_4896),
.B(n_4888),
.Y(n_4919)
);

NOR2x1_ASAP7_75t_L g4920 ( 
.A(n_4892),
.B(n_758),
.Y(n_4920)
);

BUFx2_ASAP7_75t_L g4921 ( 
.A(n_4884),
.Y(n_4921)
);

NOR2x1_ASAP7_75t_L g4922 ( 
.A(n_4900),
.B(n_759),
.Y(n_4922)
);

AND2x2_ASAP7_75t_L g4923 ( 
.A(n_4894),
.B(n_759),
.Y(n_4923)
);

AOI22xp5_ASAP7_75t_L g4924 ( 
.A1(n_4918),
.A2(n_4904),
.B1(n_4906),
.B2(n_4893),
.Y(n_4924)
);

NOR3xp33_ASAP7_75t_L g4925 ( 
.A(n_4915),
.B(n_4903),
.C(n_4905),
.Y(n_4925)
);

NOR3xp33_ASAP7_75t_L g4926 ( 
.A(n_4921),
.B(n_4902),
.C(n_4898),
.Y(n_4926)
);

OR2x2_ASAP7_75t_L g4927 ( 
.A(n_4914),
.B(n_760),
.Y(n_4927)
);

NOR2x1_ASAP7_75t_L g4928 ( 
.A(n_4920),
.B(n_760),
.Y(n_4928)
);

INVx4_ASAP7_75t_L g4929 ( 
.A(n_4911),
.Y(n_4929)
);

OR2x2_ASAP7_75t_L g4930 ( 
.A(n_4913),
.B(n_761),
.Y(n_4930)
);

AOI21xp5_ASAP7_75t_L g4931 ( 
.A1(n_4923),
.A2(n_761),
.B(n_763),
.Y(n_4931)
);

A2O1A1Ixp33_ASAP7_75t_L g4932 ( 
.A1(n_4919),
.A2(n_766),
.B(n_764),
.C(n_765),
.Y(n_4932)
);

AOI22xp5_ASAP7_75t_L g4933 ( 
.A1(n_4916),
.A2(n_4908),
.B1(n_4912),
.B2(n_4922),
.Y(n_4933)
);

OR2x6_ASAP7_75t_L g4934 ( 
.A(n_4910),
.B(n_765),
.Y(n_4934)
);

NAND2xp33_ASAP7_75t_SL g4935 ( 
.A(n_4909),
.B(n_766),
.Y(n_4935)
);

O2A1O1Ixp33_ASAP7_75t_L g4936 ( 
.A1(n_4917),
.A2(n_769),
.B(n_767),
.C(n_768),
.Y(n_4936)
);

OAI22xp5_ASAP7_75t_L g4937 ( 
.A1(n_4924),
.A2(n_772),
.B1(n_768),
.B2(n_771),
.Y(n_4937)
);

AOI221xp5_ASAP7_75t_L g4938 ( 
.A1(n_4926),
.A2(n_776),
.B1(n_773),
.B2(n_775),
.C(n_777),
.Y(n_4938)
);

AOI22xp5_ASAP7_75t_L g4939 ( 
.A1(n_4925),
.A2(n_778),
.B1(n_775),
.B2(n_777),
.Y(n_4939)
);

XNOR2xp5_ASAP7_75t_L g4940 ( 
.A(n_4933),
.B(n_4931),
.Y(n_4940)
);

INVx2_ASAP7_75t_L g4941 ( 
.A(n_4929),
.Y(n_4941)
);

NAND2xp5_ASAP7_75t_L g4942 ( 
.A(n_4932),
.B(n_779),
.Y(n_4942)
);

INVx1_ASAP7_75t_L g4943 ( 
.A(n_4927),
.Y(n_4943)
);

OAI22x1_ASAP7_75t_L g4944 ( 
.A1(n_4939),
.A2(n_4928),
.B1(n_4930),
.B2(n_4935),
.Y(n_4944)
);

OAI22xp5_ASAP7_75t_L g4945 ( 
.A1(n_4941),
.A2(n_4934),
.B1(n_4936),
.B2(n_782),
.Y(n_4945)
);

INVx1_ASAP7_75t_L g4946 ( 
.A(n_4942),
.Y(n_4946)
);

AOI22xp5_ASAP7_75t_L g4947 ( 
.A1(n_4943),
.A2(n_4938),
.B1(n_4937),
.B2(n_4940),
.Y(n_4947)
);

AOI22xp5_ASAP7_75t_L g4948 ( 
.A1(n_4941),
.A2(n_4934),
.B1(n_782),
.B2(n_779),
.Y(n_4948)
);

INVx1_ASAP7_75t_L g4949 ( 
.A(n_4941),
.Y(n_4949)
);

NAND2xp5_ASAP7_75t_L g4950 ( 
.A(n_4949),
.B(n_780),
.Y(n_4950)
);

XNOR2xp5_ASAP7_75t_L g4951 ( 
.A(n_4947),
.B(n_780),
.Y(n_4951)
);

OAI21x1_ASAP7_75t_SL g4952 ( 
.A1(n_4945),
.A2(n_783),
.B(n_785),
.Y(n_4952)
);

NAND4xp75_ASAP7_75t_L g4953 ( 
.A(n_4950),
.B(n_4946),
.C(n_4948),
.D(n_4944),
.Y(n_4953)
);

OAI22xp5_ASAP7_75t_L g4954 ( 
.A1(n_4951),
.A2(n_786),
.B1(n_783),
.B2(n_785),
.Y(n_4954)
);

NAND2xp5_ASAP7_75t_SL g4955 ( 
.A(n_4954),
.B(n_4952),
.Y(n_4955)
);

AOI221xp5_ASAP7_75t_L g4956 ( 
.A1(n_4953),
.A2(n_788),
.B1(n_786),
.B2(n_787),
.C(n_789),
.Y(n_4956)
);

AOI22xp33_ASAP7_75t_L g4957 ( 
.A1(n_4954),
.A2(n_791),
.B1(n_787),
.B2(n_790),
.Y(n_4957)
);

HB1xp67_ASAP7_75t_L g4958 ( 
.A(n_4956),
.Y(n_4958)
);

OAI22xp5_ASAP7_75t_L g4959 ( 
.A1(n_4955),
.A2(n_4957),
.B1(n_792),
.B2(n_790),
.Y(n_4959)
);

AOI21xp5_ASAP7_75t_L g4960 ( 
.A1(n_4955),
.A2(n_791),
.B(n_792),
.Y(n_4960)
);

NAND2xp5_ASAP7_75t_L g4961 ( 
.A(n_4960),
.B(n_793),
.Y(n_4961)
);

O2A1O1Ixp33_ASAP7_75t_L g4962 ( 
.A1(n_4958),
.A2(n_798),
.B(n_796),
.C(n_797),
.Y(n_4962)
);

OAI222xp33_ASAP7_75t_L g4963 ( 
.A1(n_4962),
.A2(n_4959),
.B1(n_798),
.B2(n_800),
.C1(n_796),
.C2(n_797),
.Y(n_4963)
);

AOI22xp5_ASAP7_75t_L g4964 ( 
.A1(n_4961),
.A2(n_3728),
.B1(n_801),
.B2(n_799),
.Y(n_4964)
);

AOI221xp5_ASAP7_75t_L g4965 ( 
.A1(n_4963),
.A2(n_801),
.B1(n_799),
.B2(n_800),
.C(n_802),
.Y(n_4965)
);

AOI211xp5_ASAP7_75t_L g4966 ( 
.A1(n_4965),
.A2(n_4964),
.B(n_803),
.C(n_802),
.Y(n_4966)
);


endmodule