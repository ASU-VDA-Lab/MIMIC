module fake_jpeg_13783_n_645 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_645);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_645;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_19;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_18),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_16),
.B(n_12),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_15),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_17),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_17),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

CKINVDCx14_ASAP7_75t_R g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx4f_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

INVx8_ASAP7_75t_SL g44 ( 
.A(n_15),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_8),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_7),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_6),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_2),
.B(n_3),
.Y(n_58)
);

BUFx16f_ASAP7_75t_L g59 ( 
.A(n_9),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_8),
.Y(n_60)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_57),
.Y(n_61)
);

INVx5_ASAP7_75t_L g217 ( 
.A(n_61),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_62),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_63),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_64),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g181 ( 
.A(n_65),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_22),
.B(n_15),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_66),
.B(n_73),
.Y(n_210)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_67),
.Y(n_149)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_68),
.Y(n_179)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g176 ( 
.A(n_69),
.Y(n_176)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_70),
.Y(n_173)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_71),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_22),
.B(n_14),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_72),
.B(n_103),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_28),
.B(n_0),
.Y(n_73)
);

INVx13_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

INVx4_ASAP7_75t_SL g138 ( 
.A(n_74),
.Y(n_138)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_75),
.Y(n_198)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g207 ( 
.A(n_76),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_58),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_77),
.B(n_78),
.Y(n_136)
);

AND2x2_ASAP7_75t_SL g78 ( 
.A(n_35),
.B(n_0),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_79),
.Y(n_204)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_23),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g130 ( 
.A(n_80),
.Y(n_130)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_20),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g175 ( 
.A(n_81),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_28),
.B(n_1),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_82),
.B(n_83),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_32),
.B(n_4),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_30),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_84),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_58),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_85),
.B(n_90),
.Y(n_147)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_30),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_86),
.Y(n_167)
);

BUFx10_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g146 ( 
.A(n_87),
.Y(n_146)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_39),
.Y(n_88)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_88),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_42),
.Y(n_89)
);

INVx5_ASAP7_75t_L g197 ( 
.A(n_89),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_51),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_30),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_91),
.Y(n_168)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_30),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_92),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_33),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_93),
.Y(n_188)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_21),
.Y(n_94)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_94),
.Y(n_135)
);

BUFx4f_ASAP7_75t_SL g95 ( 
.A(n_59),
.Y(n_95)
);

BUFx4f_ASAP7_75t_SL g150 ( 
.A(n_95),
.Y(n_150)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_59),
.Y(n_96)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_96),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_42),
.Y(n_97)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_97),
.Y(n_156)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_59),
.Y(n_98)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_98),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_33),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_99),
.Y(n_203)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_43),
.Y(n_100)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_100),
.Y(n_202)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_35),
.Y(n_101)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_101),
.Y(n_166)
);

NOR2xp67_ASAP7_75t_L g102 ( 
.A(n_20),
.B(n_4),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_102),
.B(n_115),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_32),
.B(n_5),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_35),
.Y(n_104)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_104),
.Y(n_185)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_59),
.Y(n_105)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_105),
.Y(n_172)
);

INVx2_ASAP7_75t_SL g106 ( 
.A(n_21),
.Y(n_106)
);

NAND2x1_ASAP7_75t_SL g184 ( 
.A(n_106),
.B(n_26),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_33),
.Y(n_107)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_107),
.Y(n_134)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_35),
.Y(n_108)
);

INVx2_ASAP7_75t_SL g196 ( 
.A(n_108),
.Y(n_196)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_35),
.Y(n_109)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_109),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_33),
.Y(n_110)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_110),
.Y(n_163)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_39),
.Y(n_111)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_111),
.Y(n_139)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_35),
.Y(n_112)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_112),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_48),
.Y(n_113)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_113),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_21),
.Y(n_114)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_114),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_36),
.B(n_5),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_36),
.B(n_5),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_116),
.B(n_27),
.Y(n_170)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_39),
.Y(n_117)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_117),
.Y(n_143)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_43),
.Y(n_118)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_118),
.Y(n_206)
);

BUFx12f_ASAP7_75t_L g119 ( 
.A(n_48),
.Y(n_119)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_119),
.Y(n_205)
);

INVx11_ASAP7_75t_L g120 ( 
.A(n_29),
.Y(n_120)
);

INVx11_ASAP7_75t_L g212 ( 
.A(n_120),
.Y(n_212)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_48),
.Y(n_121)
);

INVx6_ASAP7_75t_L g214 ( 
.A(n_121),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_48),
.Y(n_122)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_122),
.Y(n_140)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_54),
.Y(n_123)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_123),
.Y(n_211)
);

INVx11_ASAP7_75t_L g124 ( 
.A(n_29),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_124),
.Y(n_144)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_54),
.Y(n_125)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_125),
.Y(n_148)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_46),
.Y(n_126)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_126),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_39),
.Y(n_127)
);

INVx8_ASAP7_75t_L g161 ( 
.A(n_127),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_39),
.Y(n_128)
);

INVx8_ASAP7_75t_L g190 ( 
.A(n_128),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_54),
.Y(n_129)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_129),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_61),
.A2(n_20),
.B1(n_53),
.B2(n_56),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_141),
.A2(n_50),
.B1(n_56),
.B2(n_52),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_78),
.A2(n_38),
.B1(n_53),
.B2(n_49),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_145),
.B(n_160),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_124),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_152),
.B(n_155),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_87),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_87),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_159),
.B(n_164),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_106),
.A2(n_38),
.B1(n_53),
.B2(n_49),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_74),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_170),
.B(n_171),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_95),
.B(n_27),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_68),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_174),
.B(n_177),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_127),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_101),
.Y(n_178)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_178),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_128),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_180),
.B(n_192),
.Y(n_223)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_129),
.Y(n_183)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_183),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g290 ( 
.A(n_184),
.Y(n_290)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_125),
.Y(n_186)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_186),
.Y(n_286)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_94),
.Y(n_187)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_187),
.Y(n_289)
);

OR2x2_ASAP7_75t_L g192 ( 
.A(n_114),
.B(n_60),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_80),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_193),
.B(n_216),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_121),
.B(n_55),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_195),
.B(n_213),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_79),
.B(n_55),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_199),
.B(n_201),
.Y(n_222)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_86),
.Y(n_200)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_200),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_79),
.B(n_31),
.Y(n_201)
);

AOI21xp33_ASAP7_75t_L g208 ( 
.A1(n_68),
.A2(n_34),
.B(n_31),
.Y(n_208)
);

OR2x2_ASAP7_75t_L g224 ( 
.A(n_208),
.B(n_153),
.Y(n_224)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_104),
.Y(n_209)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_209),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_92),
.B(n_34),
.Y(n_213)
);

OR2x2_ASAP7_75t_L g216 ( 
.A(n_97),
.B(n_46),
.Y(n_216)
);

INVx6_ASAP7_75t_SL g218 ( 
.A(n_138),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_218),
.Y(n_315)
);

INVx5_ASAP7_75t_L g220 ( 
.A(n_181),
.Y(n_220)
);

INVx3_ASAP7_75t_L g305 ( 
.A(n_220),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_224),
.A2(n_225),
.B(n_25),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_147),
.A2(n_216),
.B(n_192),
.Y(n_225)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_138),
.Y(n_226)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_226),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_228),
.Y(n_335)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_205),
.Y(n_229)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_229),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_210),
.B(n_47),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_230),
.B(n_237),
.Y(n_299)
);

CKINVDCx9p33_ASAP7_75t_R g231 ( 
.A(n_150),
.Y(n_231)
);

BUFx12f_ASAP7_75t_L g326 ( 
.A(n_231),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_188),
.Y(n_233)
);

INVx6_ASAP7_75t_L g310 ( 
.A(n_233),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_142),
.B(n_47),
.Y(n_237)
);

BUFx12_ASAP7_75t_L g238 ( 
.A(n_150),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g294 ( 
.A(n_238),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_136),
.A2(n_122),
.B1(n_113),
.B2(n_110),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_239),
.A2(n_258),
.B1(n_277),
.B2(n_63),
.Y(n_336)
);

INVx13_ASAP7_75t_L g240 ( 
.A(n_175),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_240),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_184),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_241),
.B(n_246),
.Y(n_300)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_214),
.Y(n_242)
);

INVx3_ASAP7_75t_L g342 ( 
.A(n_242),
.Y(n_342)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_214),
.Y(n_243)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_243),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_157),
.B(n_60),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_244),
.B(n_245),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_202),
.B(n_45),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_206),
.Y(n_246)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_205),
.Y(n_247)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_247),
.Y(n_317)
);

BUFx8_ASAP7_75t_L g248 ( 
.A(n_212),
.Y(n_248)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_248),
.Y(n_325)
);

INVx5_ASAP7_75t_L g249 ( 
.A(n_181),
.Y(n_249)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_249),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_215),
.B(n_149),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_250),
.B(n_257),
.Y(n_351)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_135),
.Y(n_251)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_251),
.Y(n_303)
);

INVx5_ASAP7_75t_L g253 ( 
.A(n_181),
.Y(n_253)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_253),
.Y(n_330)
);

INVx5_ASAP7_75t_L g254 ( 
.A(n_156),
.Y(n_254)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_254),
.Y(n_345)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_182),
.Y(n_255)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_255),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_188),
.Y(n_256)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_256),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_173),
.B(n_89),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_141),
.A2(n_93),
.B1(n_107),
.B2(n_99),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_198),
.B(n_37),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_259),
.B(n_261),
.Y(n_352)
);

INVx5_ASAP7_75t_L g260 ( 
.A(n_156),
.Y(n_260)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_260),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_175),
.B(n_144),
.Y(n_261)
);

INVx8_ASAP7_75t_L g262 ( 
.A(n_182),
.Y(n_262)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_262),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_203),
.Y(n_263)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_263),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_130),
.A2(n_65),
.B1(n_89),
.B2(n_56),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_SL g319 ( 
.A1(n_264),
.A2(n_274),
.B1(n_276),
.B2(n_292),
.Y(n_319)
);

INVx5_ASAP7_75t_L g266 ( 
.A(n_197),
.Y(n_266)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_266),
.Y(n_338)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_131),
.Y(n_268)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_268),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_133),
.B(n_26),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_269),
.B(n_271),
.Y(n_302)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_154),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_270),
.B(n_278),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_158),
.B(n_119),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_139),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_272),
.B(n_273),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_143),
.B(n_172),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_203),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_194),
.B(n_119),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_275),
.B(n_280),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_132),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_162),
.A2(n_91),
.B1(n_84),
.B2(n_64),
.Y(n_277)
);

BUFx8_ASAP7_75t_L g278 ( 
.A(n_212),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_161),
.Y(n_280)
);

INVx5_ASAP7_75t_L g281 ( 
.A(n_185),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_281),
.B(n_282),
.Y(n_348)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_148),
.Y(n_282)
);

INVx4_ASAP7_75t_L g283 ( 
.A(n_185),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_283),
.B(n_285),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_194),
.B(n_24),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_284),
.B(n_287),
.Y(n_349)
);

INVx4_ASAP7_75t_L g285 ( 
.A(n_204),
.Y(n_285)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_217),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_196),
.B(n_191),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_288),
.B(n_291),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_196),
.B(n_24),
.Y(n_291)
);

INVx5_ASAP7_75t_L g292 ( 
.A(n_204),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_211),
.B(n_24),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_293),
.B(n_226),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_295),
.B(n_339),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_224),
.A2(n_134),
.B1(n_169),
.B2(n_163),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_297),
.A2(n_301),
.B1(n_308),
.B2(n_316),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_227),
.A2(n_290),
.B1(n_234),
.B2(n_223),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_222),
.B(n_235),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_307),
.B(n_322),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_228),
.A2(n_134),
.B1(n_169),
.B2(n_163),
.Y(n_308)
);

MAJx2_ASAP7_75t_L g309 ( 
.A(n_235),
.B(n_211),
.C(n_179),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_309),
.B(n_329),
.C(n_346),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_312),
.B(n_337),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_232),
.A2(n_151),
.B1(n_168),
.B2(n_165),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_219),
.B(n_166),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_267),
.A2(n_151),
.B1(n_168),
.B2(n_165),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_324),
.A2(n_336),
.B1(n_341),
.B2(n_347),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_SL g329 ( 
.A(n_236),
.B(n_179),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_SL g331 ( 
.A1(n_242),
.A2(n_130),
.B1(n_217),
.B2(n_146),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_331),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_240),
.A2(n_50),
.B(n_26),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g362 ( 
.A1(n_332),
.A2(n_300),
.B(n_313),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_265),
.B(n_167),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_334),
.B(n_343),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_231),
.Y(n_337)
);

AO22x2_ASAP7_75t_L g339 ( 
.A1(n_243),
.A2(n_146),
.B1(n_191),
.B2(n_189),
.Y(n_339)
);

AOI22xp33_ASAP7_75t_L g341 ( 
.A1(n_255),
.A2(n_140),
.B1(n_132),
.B2(n_137),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_264),
.A2(n_62),
.B1(n_167),
.B2(n_137),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_SL g346 ( 
.A(n_221),
.B(n_176),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_279),
.A2(n_140),
.B1(n_190),
.B2(n_161),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_238),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_350),
.B(n_229),
.Y(n_361)
);

INVx6_ASAP7_75t_L g355 ( 
.A(n_310),
.Y(n_355)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_355),
.Y(n_417)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_296),
.Y(n_356)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_356),
.Y(n_401)
);

INVx13_ASAP7_75t_L g358 ( 
.A(n_315),
.Y(n_358)
);

CKINVDCx14_ASAP7_75t_R g405 ( 
.A(n_358),
.Y(n_405)
);

INVx3_ASAP7_75t_SL g359 ( 
.A(n_310),
.Y(n_359)
);

INVxp33_ASAP7_75t_L g402 ( 
.A(n_359),
.Y(n_402)
);

INVx3_ASAP7_75t_L g360 ( 
.A(n_342),
.Y(n_360)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_360),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_361),
.B(n_376),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g431 ( 
.A(n_362),
.B(n_374),
.Y(n_431)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_334),
.Y(n_363)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_363),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_L g364 ( 
.A1(n_335),
.A2(n_268),
.B(n_270),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_L g406 ( 
.A1(n_364),
.A2(n_332),
.B(n_311),
.Y(n_406)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_296),
.Y(n_365)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_365),
.Y(n_426)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_344),
.Y(n_366)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_366),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_335),
.A2(n_262),
.B1(n_256),
.B2(n_274),
.Y(n_369)
);

AOI22xp33_ASAP7_75t_L g425 ( 
.A1(n_369),
.A2(n_375),
.B1(n_396),
.B2(n_397),
.Y(n_425)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_344),
.Y(n_370)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_370),
.Y(n_420)
);

AOI21xp5_ASAP7_75t_L g371 ( 
.A1(n_295),
.A2(n_349),
.B(n_319),
.Y(n_371)
);

AOI21xp5_ASAP7_75t_L g409 ( 
.A1(n_371),
.A2(n_311),
.B(n_320),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_348),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_373),
.B(n_377),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g374 ( 
.A(n_318),
.B(n_287),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_336),
.A2(n_276),
.B1(n_263),
.B2(n_233),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_351),
.B(n_266),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_333),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_326),
.Y(n_379)
);

CKINVDCx16_ASAP7_75t_R g437 ( 
.A(n_379),
.Y(n_437)
);

CKINVDCx12_ASAP7_75t_R g381 ( 
.A(n_294),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_381),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_307),
.B(n_286),
.C(n_252),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_382),
.B(n_393),
.C(n_368),
.Y(n_404)
);

OAI22xp33_ASAP7_75t_SL g383 ( 
.A1(n_309),
.A2(n_283),
.B1(n_247),
.B2(n_289),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_383),
.A2(n_399),
.B1(n_325),
.B2(n_314),
.Y(n_415)
);

INVx13_ASAP7_75t_L g384 ( 
.A(n_326),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_384),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_333),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_385),
.B(n_386),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_333),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_302),
.B(n_254),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_387),
.B(n_390),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_322),
.B(n_260),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_388),
.B(n_392),
.Y(n_428)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_304),
.Y(n_389)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_389),
.Y(n_422)
);

AND2x6_ASAP7_75t_L g390 ( 
.A(n_312),
.B(n_238),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_304),
.Y(n_391)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_391),
.Y(n_435)
);

INVx3_ASAP7_75t_L g392 ( 
.A(n_342),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_329),
.B(n_346),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_353),
.B(n_281),
.Y(n_394)
);

BUFx24_ASAP7_75t_SL g408 ( 
.A(n_394),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_298),
.Y(n_396)
);

CKINVDCx16_ASAP7_75t_R g397 ( 
.A(n_311),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_352),
.B(n_45),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_398),
.B(n_317),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_321),
.A2(n_190),
.B1(n_45),
.B2(n_52),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_380),
.A2(n_323),
.B1(n_343),
.B2(n_347),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_403),
.A2(n_410),
.B1(n_418),
.B2(n_424),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_404),
.B(n_407),
.C(n_416),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_406),
.B(n_354),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_368),
.B(n_299),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_L g473 ( 
.A1(n_409),
.A2(n_392),
.B(n_360),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_372),
.A2(n_320),
.B1(n_327),
.B2(n_298),
.Y(n_410)
);

OAI32xp33_ASAP7_75t_L g413 ( 
.A1(n_367),
.A2(n_339),
.A3(n_303),
.B1(n_306),
.B2(n_338),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_413),
.B(n_415),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_393),
.B(n_338),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_380),
.A2(n_327),
.B1(n_339),
.B2(n_306),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_367),
.B(n_382),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_419),
.B(n_433),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_L g424 ( 
.A1(n_372),
.A2(n_357),
.B1(n_362),
.B2(n_363),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_371),
.A2(n_339),
.B1(n_317),
.B2(n_345),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_427),
.A2(n_434),
.B1(n_378),
.B2(n_375),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_432),
.B(n_436),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_387),
.B(n_314),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_354),
.A2(n_345),
.B1(n_325),
.B2(n_340),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_398),
.B(n_340),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_417),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_440),
.B(n_448),
.Y(n_475)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_426),
.Y(n_441)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_441),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_412),
.B(n_373),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_SL g497 ( 
.A(n_443),
.B(n_449),
.Y(n_497)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_438),
.Y(n_445)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_445),
.Y(n_492)
);

OAI32xp33_ASAP7_75t_L g446 ( 
.A1(n_400),
.A2(n_354),
.A3(n_390),
.B1(n_366),
.B2(n_365),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_446),
.B(n_460),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_400),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_421),
.B(n_374),
.Y(n_449)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_450),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_SL g480 ( 
.A1(n_451),
.A2(n_454),
.B(n_465),
.Y(n_480)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_420),
.Y(n_452)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_452),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_406),
.B(n_364),
.Y(n_453)
);

INVxp67_ASAP7_75t_L g482 ( 
.A(n_453),
.Y(n_482)
);

AND2x6_ASAP7_75t_L g454 ( 
.A(n_430),
.B(n_379),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_405),
.B(n_374),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_455),
.B(n_464),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_411),
.B(n_377),
.Y(n_456)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_456),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_430),
.A2(n_395),
.B1(n_385),
.B2(n_386),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_457),
.A2(n_471),
.B1(n_472),
.B2(n_431),
.Y(n_478)
);

INVx13_ASAP7_75t_L g458 ( 
.A(n_437),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_458),
.Y(n_476)
);

INVx1_ASAP7_75t_SL g460 ( 
.A(n_431),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_422),
.Y(n_461)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_461),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_403),
.A2(n_369),
.B1(n_395),
.B2(n_359),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_462),
.A2(n_420),
.B1(n_401),
.B2(n_414),
.Y(n_477)
);

O2A1O1Ixp33_ASAP7_75t_L g463 ( 
.A1(n_431),
.A2(n_358),
.B(n_391),
.C(n_389),
.Y(n_463)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_463),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_408),
.B(n_428),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_427),
.B(n_356),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_417),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_466),
.B(n_468),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_423),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_467),
.B(n_326),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_432),
.B(n_396),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_422),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_469),
.B(n_474),
.Y(n_508)
);

INVx13_ASAP7_75t_L g470 ( 
.A(n_429),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_470),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_425),
.A2(n_415),
.B1(n_409),
.B2(n_423),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_404),
.A2(n_359),
.B1(n_355),
.B2(n_396),
.Y(n_472)
);

OAI21xp5_ASAP7_75t_SL g501 ( 
.A1(n_473),
.A2(n_305),
.B(n_249),
.Y(n_501)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_435),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g527 ( 
.A1(n_477),
.A2(n_465),
.B1(n_463),
.B2(n_461),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_SL g519 ( 
.A1(n_478),
.A2(n_487),
.B1(n_447),
.B2(n_460),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_471),
.A2(n_434),
.B1(n_418),
.B2(n_402),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_L g509 ( 
.A1(n_479),
.A2(n_481),
.B1(n_447),
.B2(n_462),
.Y(n_509)
);

AOI22x1_ASAP7_75t_L g481 ( 
.A1(n_444),
.A2(n_413),
.B1(n_401),
.B2(n_414),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_442),
.B(n_416),
.C(n_419),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_483),
.B(n_489),
.C(n_500),
.Y(n_512)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_442),
.B(n_439),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g517 ( 
.A(n_486),
.B(n_491),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_457),
.A2(n_402),
.B1(n_435),
.B2(n_433),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_439),
.B(n_407),
.C(n_436),
.Y(n_489)
);

OAI32xp33_ASAP7_75t_L g490 ( 
.A1(n_444),
.A2(n_330),
.A3(n_328),
.B1(n_189),
.B2(n_285),
.Y(n_490)
);

INVxp67_ASAP7_75t_L g521 ( 
.A(n_490),
.Y(n_521)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_446),
.B(n_294),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_SL g494 ( 
.A(n_451),
.B(n_384),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_SL g520 ( 
.A(n_494),
.B(n_507),
.Y(n_520)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_499),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_472),
.B(n_330),
.C(n_328),
.Y(n_500)
);

AOI21xp5_ASAP7_75t_L g516 ( 
.A1(n_501),
.A2(n_503),
.B(n_453),
.Y(n_516)
);

OAI21xp5_ASAP7_75t_SL g503 ( 
.A1(n_473),
.A2(n_305),
.B(n_253),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_456),
.B(n_292),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_505),
.B(n_278),
.Y(n_536)
);

XNOR2xp5_ASAP7_75t_SL g507 ( 
.A(n_451),
.B(n_220),
.Y(n_507)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_509),
.Y(n_544)
);

CKINVDCx16_ASAP7_75t_R g510 ( 
.A(n_508),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_510),
.B(n_513),
.Y(n_550)
);

CKINVDCx16_ASAP7_75t_R g513 ( 
.A(n_508),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_502),
.Y(n_514)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_514),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_502),
.B(n_468),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_515),
.B(n_518),
.Y(n_555)
);

AOI21xp5_ASAP7_75t_L g543 ( 
.A1(n_516),
.A2(n_529),
.B(n_503),
.Y(n_543)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_504),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g540 ( 
.A(n_519),
.B(n_522),
.Y(n_540)
);

XNOR2xp5_ASAP7_75t_L g522 ( 
.A(n_486),
.B(n_459),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g523 ( 
.A(n_489),
.B(n_483),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g549 ( 
.A(n_523),
.B(n_538),
.Y(n_549)
);

BUFx2_ASAP7_75t_L g524 ( 
.A(n_493),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_524),
.B(n_533),
.Y(n_553)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_504),
.Y(n_525)
);

INVx2_ASAP7_75t_SL g563 ( 
.A(n_525),
.Y(n_563)
);

OAI22xp5_ASAP7_75t_L g526 ( 
.A1(n_493),
.A2(n_450),
.B1(n_454),
.B2(n_469),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_L g541 ( 
.A1(n_526),
.A2(n_527),
.B1(n_528),
.B2(n_530),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_SL g528 ( 
.A1(n_478),
.A2(n_465),
.B1(n_474),
.B2(n_453),
.Y(n_528)
);

OAI21xp5_ASAP7_75t_L g529 ( 
.A1(n_482),
.A2(n_458),
.B(n_445),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_L g530 ( 
.A1(n_497),
.A2(n_441),
.B1(n_466),
.B2(n_470),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_L g531 ( 
.A1(n_491),
.A2(n_440),
.B1(n_19),
.B2(n_25),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_L g545 ( 
.A1(n_531),
.A2(n_535),
.B1(n_536),
.B2(n_537),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_482),
.B(n_507),
.C(n_487),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_532),
.B(n_500),
.C(n_481),
.Y(n_539)
);

HB1xp67_ASAP7_75t_L g533 ( 
.A(n_498),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_SL g534 ( 
.A1(n_485),
.A2(n_278),
.B1(n_248),
.B2(n_207),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_SL g542 ( 
.A1(n_534),
.A2(n_479),
.B1(n_476),
.B2(n_506),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_484),
.B(n_52),
.Y(n_535)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_488),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_L g538 ( 
.A(n_485),
.B(n_248),
.Y(n_538)
);

MAJx2_ASAP7_75t_L g583 ( 
.A(n_539),
.B(n_558),
.C(n_561),
.Y(n_583)
);

INVxp67_ASAP7_75t_L g578 ( 
.A(n_542),
.Y(n_578)
);

OAI21xp5_ASAP7_75t_L g581 ( 
.A1(n_543),
.A2(n_7),
.B(n_9),
.Y(n_581)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_512),
.B(n_480),
.C(n_494),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g577 ( 
.A(n_546),
.B(n_548),
.C(n_551),
.Y(n_577)
);

XNOR2xp5_ASAP7_75t_SL g547 ( 
.A(n_517),
.B(n_480),
.Y(n_547)
);

XOR2xp5_ASAP7_75t_L g565 ( 
.A(n_547),
.B(n_562),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_512),
.B(n_477),
.C(n_481),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_523),
.B(n_522),
.C(n_517),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_L g552 ( 
.A1(n_521),
.A2(n_506),
.B1(n_475),
.B2(n_496),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_552),
.B(n_6),
.Y(n_570)
);

OAI22xp5_ASAP7_75t_SL g556 ( 
.A1(n_521),
.A2(n_495),
.B1(n_496),
.B2(n_492),
.Y(n_556)
);

AOI322xp5_ASAP7_75t_L g564 ( 
.A1(n_556),
.A2(n_511),
.A3(n_527),
.B1(n_531),
.B2(n_524),
.C1(n_515),
.C2(n_534),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_532),
.B(n_495),
.C(n_501),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_557),
.B(n_559),
.Y(n_566)
);

XNOR2xp5_ASAP7_75t_L g558 ( 
.A(n_519),
.B(n_538),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g559 ( 
.A(n_529),
.B(n_492),
.C(n_488),
.Y(n_559)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_528),
.B(n_490),
.C(n_50),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_560),
.B(n_559),
.Y(n_575)
);

XNOR2xp5_ASAP7_75t_L g561 ( 
.A(n_520),
.B(n_40),
.Y(n_561)
);

XNOR2xp5_ASAP7_75t_L g562 ( 
.A(n_520),
.B(n_40),
.Y(n_562)
);

AOI22xp5_ASAP7_75t_L g588 ( 
.A1(n_564),
.A2(n_573),
.B1(n_579),
.B2(n_539),
.Y(n_588)
);

CKINVDCx20_ASAP7_75t_R g567 ( 
.A(n_555),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_567),
.B(n_572),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_553),
.B(n_516),
.Y(n_568)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_568),
.Y(n_586)
);

AOI21xp5_ASAP7_75t_L g569 ( 
.A1(n_544),
.A2(n_40),
.B(n_37),
.Y(n_569)
);

OAI21xp5_ASAP7_75t_SL g592 ( 
.A1(n_569),
.A2(n_576),
.B(n_584),
.Y(n_592)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_570),
.Y(n_589)
);

OAI221xp5_ASAP7_75t_L g571 ( 
.A1(n_550),
.A2(n_37),
.B1(n_25),
.B2(n_19),
.C(n_9),
.Y(n_571)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_571),
.Y(n_597)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_563),
.Y(n_572)
);

OAI22xp5_ASAP7_75t_SL g573 ( 
.A1(n_560),
.A2(n_19),
.B1(n_7),
.B2(n_8),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_563),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_574),
.B(n_575),
.Y(n_595)
);

CKINVDCx20_ASAP7_75t_R g576 ( 
.A(n_545),
.Y(n_576)
);

CKINVDCx14_ASAP7_75t_R g579 ( 
.A(n_541),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_554),
.B(n_6),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_SL g602 ( 
.A(n_580),
.B(n_582),
.Y(n_602)
);

XOR2xp5_ASAP7_75t_L g591 ( 
.A(n_581),
.B(n_562),
.Y(n_591)
);

CKINVDCx16_ASAP7_75t_R g582 ( 
.A(n_557),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_548),
.B(n_9),
.Y(n_584)
);

MAJIxp5_ASAP7_75t_L g587 ( 
.A(n_582),
.B(n_551),
.C(n_540),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_587),
.B(n_590),
.Y(n_603)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_588),
.Y(n_605)
);

MAJIxp5_ASAP7_75t_L g590 ( 
.A(n_566),
.B(n_540),
.C(n_546),
.Y(n_590)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_591),
.Y(n_610)
);

XOR2xp5_ASAP7_75t_L g593 ( 
.A(n_577),
.B(n_549),
.Y(n_593)
);

XNOR2xp5_ASAP7_75t_L g612 ( 
.A(n_593),
.B(n_565),
.Y(n_612)
);

OAI22xp5_ASAP7_75t_SL g594 ( 
.A1(n_578),
.A2(n_547),
.B1(n_558),
.B2(n_549),
.Y(n_594)
);

AOI22xp5_ASAP7_75t_L g606 ( 
.A1(n_594),
.A2(n_599),
.B1(n_573),
.B2(n_581),
.Y(n_606)
);

MAJIxp5_ASAP7_75t_L g596 ( 
.A(n_577),
.B(n_561),
.C(n_11),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_596),
.B(n_600),
.Y(n_607)
);

INVx6_ASAP7_75t_L g598 ( 
.A(n_576),
.Y(n_598)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_598),
.Y(n_613)
);

OAI22xp5_ASAP7_75t_SL g599 ( 
.A1(n_578),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_599)
);

MAJIxp5_ASAP7_75t_L g600 ( 
.A(n_583),
.B(n_10),
.C(n_13),
.Y(n_600)
);

MAJIxp5_ASAP7_75t_L g601 ( 
.A(n_583),
.B(n_10),
.C(n_13),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_601),
.B(n_13),
.Y(n_615)
);

OAI22xp5_ASAP7_75t_SL g604 ( 
.A1(n_588),
.A2(n_568),
.B1(n_570),
.B2(n_567),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_604),
.B(n_608),
.Y(n_622)
);

XOR2xp5_ASAP7_75t_L g623 ( 
.A(n_606),
.B(n_616),
.Y(n_623)
);

OAI22xp5_ASAP7_75t_L g608 ( 
.A1(n_597),
.A2(n_574),
.B1(n_572),
.B2(n_584),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_602),
.B(n_569),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_609),
.B(n_614),
.Y(n_624)
);

HB1xp67_ASAP7_75t_L g611 ( 
.A(n_595),
.Y(n_611)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_611),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_612),
.B(n_615),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_587),
.B(n_580),
.Y(n_614)
);

XOR2xp5_ASAP7_75t_L g616 ( 
.A(n_594),
.B(n_565),
.Y(n_616)
);

OAI21xp5_ASAP7_75t_L g617 ( 
.A1(n_605),
.A2(n_586),
.B(n_585),
.Y(n_617)
);

AOI32xp33_ASAP7_75t_L g629 ( 
.A1(n_617),
.A2(n_627),
.A3(n_607),
.B1(n_592),
.B2(n_589),
.Y(n_629)
);

CKINVDCx20_ASAP7_75t_R g618 ( 
.A(n_604),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_618),
.B(n_621),
.Y(n_634)
);

MAJIxp5_ASAP7_75t_L g620 ( 
.A(n_603),
.B(n_593),
.C(n_590),
.Y(n_620)
);

OR2x2_ASAP7_75t_L g633 ( 
.A(n_620),
.B(n_600),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_613),
.B(n_596),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_SL g626 ( 
.A(n_612),
.B(n_598),
.Y(n_626)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_626),
.Y(n_628)
);

OAI21xp5_ASAP7_75t_L g627 ( 
.A1(n_610),
.A2(n_592),
.B(n_601),
.Y(n_627)
);

OAI21x1_ASAP7_75t_L g637 ( 
.A1(n_629),
.A2(n_633),
.B(n_622),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_620),
.B(n_606),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_SL g635 ( 
.A(n_630),
.B(n_625),
.Y(n_635)
);

XOR2xp5_ASAP7_75t_L g631 ( 
.A(n_623),
.B(n_616),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_631),
.B(n_632),
.Y(n_638)
);

INVxp67_ASAP7_75t_SL g632 ( 
.A(n_617),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_635),
.B(n_636),
.Y(n_639)
);

MAJIxp5_ASAP7_75t_L g636 ( 
.A(n_628),
.B(n_624),
.C(n_623),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_637),
.B(n_634),
.Y(n_640)
);

AO221x1_ASAP7_75t_L g641 ( 
.A1(n_640),
.A2(n_634),
.B1(n_627),
.B2(n_638),
.C(n_619),
.Y(n_641)
);

MAJIxp5_ASAP7_75t_L g642 ( 
.A(n_641),
.B(n_639),
.C(n_599),
.Y(n_642)
);

MAJIxp5_ASAP7_75t_L g643 ( 
.A(n_642),
.B(n_591),
.C(n_571),
.Y(n_643)
);

XOR2xp5_ASAP7_75t_L g644 ( 
.A(n_643),
.B(n_14),
.Y(n_644)
);

BUFx24_ASAP7_75t_SL g645 ( 
.A(n_644),
.Y(n_645)
);


endmodule