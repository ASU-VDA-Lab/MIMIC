module fake_ariane_124_n_794 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_794);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_794;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_698;
wire n_695;
wire n_160;
wire n_180;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_176;
wire n_691;
wire n_404;
wire n_172;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_373;
wire n_299;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_771;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_245;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_760;
wire n_591;
wire n_690;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_244;
wire n_679;
wire n_643;
wire n_226;
wire n_781;
wire n_261;
wire n_220;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_286;
wire n_443;
wire n_586;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_524;
wire n_391;
wire n_349;
wire n_634;
wire n_466;
wire n_756;
wire n_346;
wire n_214;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_670;
wire n_607;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_162;
wire n_765;
wire n_264;
wire n_737;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_790;
wire n_363;
wire n_720;
wire n_354;
wire n_725;
wire n_419;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_338;
wire n_285;
wire n_473;
wire n_186;
wire n_202;
wire n_193;
wire n_761;
wire n_733;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_779;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_672;
wire n_487;
wire n_740;
wire n_167;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_259;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_578;
wire n_701;
wire n_625;
wire n_405;
wire n_557;
wire n_169;
wire n_173;
wire n_242;
wire n_645;
wire n_309;
wire n_320;
wire n_331;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_166;
wire n_253;
wire n_561;
wire n_770;
wire n_218;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_732;
wire n_369;
wire n_240;
wire n_224;
wire n_787;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_256;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_694;
wire n_689;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_248;
wire n_277;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_168;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_163;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_579;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_237;
wire n_780;
wire n_175;
wire n_711;
wire n_453;
wire n_734;
wire n_491;
wire n_181;
wire n_723;
wire n_616;
wire n_617;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_741;
wire n_747;
wire n_772;
wire n_371;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_178;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_249;
wire n_534;
wire n_212;
wire n_444;
wire n_355;
wire n_609;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_716;
wire n_742;
wire n_182;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_769;
wire n_577;
wire n_407;
wire n_774;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_280;
wire n_215;
wire n_252;
wire n_629;
wire n_664;
wire n_161;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_763;
wire n_655;
wire n_540;
wire n_216;
wire n_544;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_389;
wire n_657;
wire n_513;
wire n_288;
wire n_179;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_304;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_669;
wire n_785;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_793;
wire n_174;
wire n_275;
wire n_704;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_496;
wire n_739;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_792;
wire n_428;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_773;
wire n_165;
wire n_317;
wire n_243;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_749;
wire n_289;
wire n_542;
wire n_548;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_164;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_425;
wire n_431;
wire n_508;
wire n_624;
wire n_791;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_191;
wire n_382;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_558;
wire n_592;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_531;
wire n_783;
wire n_675;

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_128),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_52),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_125),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_69),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_75),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_6),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_101),
.Y(n_166)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_51),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_48),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_107),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_44),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_155),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_54),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_27),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_33),
.Y(n_174)
);

BUFx10_ASAP7_75t_L g175 ( 
.A(n_123),
.Y(n_175)
);

BUFx5_ASAP7_75t_L g176 ( 
.A(n_24),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_93),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_89),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_159),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_83),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_108),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_6),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_156),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_150),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_34),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_104),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_21),
.Y(n_187)
);

BUFx2_ASAP7_75t_L g188 ( 
.A(n_13),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_145),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_56),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_7),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_73),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_39),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_9),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_28),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_29),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_86),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_88),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_42),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_113),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_109),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_20),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_60),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_57),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_5),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_18),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_53),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_22),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_153),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_147),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_70),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_23),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_72),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_50),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_146),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_118),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_162),
.B(n_163),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_182),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_176),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_175),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_188),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_160),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_191),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g224 ( 
.A(n_198),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_194),
.Y(n_225)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_205),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_176),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_175),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_171),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_178),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_164),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_170),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_186),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_200),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_193),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_187),
.Y(n_236)
);

BUFx2_ASAP7_75t_L g237 ( 
.A(n_165),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_161),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_204),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_166),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_211),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_168),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_176),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_169),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_214),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_208),
.B(n_0),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_172),
.Y(n_247)
);

INVxp67_ASAP7_75t_SL g248 ( 
.A(n_213),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_176),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_173),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_187),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_174),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_177),
.Y(n_253)
);

NOR2xp67_ASAP7_75t_L g254 ( 
.A(n_187),
.B(n_0),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_179),
.Y(n_255)
);

INVxp33_ASAP7_75t_L g256 ( 
.A(n_187),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_180),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_181),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_183),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_184),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_185),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_223),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_225),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_231),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_236),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_251),
.B(n_224),
.Y(n_266)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_219),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_236),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_224),
.B(n_167),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_232),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_233),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_218),
.Y(n_272)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_219),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_236),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_236),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_227),
.Y(n_276)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_227),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_246),
.B(n_216),
.Y(n_278)
);

BUFx2_ASAP7_75t_L g279 ( 
.A(n_237),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_243),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_234),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_243),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_239),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_222),
.A2(n_210),
.B1(n_212),
.B2(n_215),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_241),
.B(n_189),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_249),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_247),
.B(n_190),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_249),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_245),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_256),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g291 ( 
.A(n_226),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_221),
.A2(n_209),
.B1(n_207),
.B2(n_206),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_257),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_256),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_248),
.B(n_192),
.Y(n_295)
);

NAND2x1_ASAP7_75t_L g296 ( 
.A(n_254),
.B(n_176),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_217),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_258),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_240),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_259),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_261),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_228),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_238),
.Y(n_303)
);

BUFx2_ASAP7_75t_L g304 ( 
.A(n_240),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_242),
.Y(n_305)
);

INVx1_ASAP7_75t_SL g306 ( 
.A(n_229),
.Y(n_306)
);

INVx3_ASAP7_75t_L g307 ( 
.A(n_244),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_250),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_252),
.B(n_195),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_253),
.B(n_196),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_262),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_267),
.Y(n_312)
);

NAND2xp33_ASAP7_75t_L g313 ( 
.A(n_305),
.B(n_253),
.Y(n_313)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_289),
.Y(n_314)
);

AND2x4_ASAP7_75t_L g315 ( 
.A(n_266),
.B(n_255),
.Y(n_315)
);

INVx4_ASAP7_75t_L g316 ( 
.A(n_289),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_263),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_289),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_276),
.B(n_220),
.Y(n_319)
);

AO22x2_ASAP7_75t_L g320 ( 
.A1(n_297),
.A2(n_222),
.B1(n_220),
.B2(n_235),
.Y(n_320)
);

AND2x6_ASAP7_75t_L g321 ( 
.A(n_266),
.B(n_176),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_289),
.Y(n_322)
);

AND2x6_ASAP7_75t_L g323 ( 
.A(n_307),
.B(n_17),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_289),
.Y(n_324)
);

INVx3_ASAP7_75t_L g325 ( 
.A(n_267),
.Y(n_325)
);

CKINVDCx11_ASAP7_75t_R g326 ( 
.A(n_299),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_264),
.Y(n_327)
);

INVx3_ASAP7_75t_L g328 ( 
.A(n_267),
.Y(n_328)
);

BUFx3_ASAP7_75t_L g329 ( 
.A(n_273),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_282),
.Y(n_330)
);

INVx3_ASAP7_75t_L g331 ( 
.A(n_273),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_301),
.B(n_293),
.Y(n_332)
);

INVx4_ASAP7_75t_L g333 ( 
.A(n_307),
.Y(n_333)
);

BUFx3_ASAP7_75t_L g334 ( 
.A(n_279),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_279),
.B(n_255),
.Y(n_335)
);

INVx3_ASAP7_75t_L g336 ( 
.A(n_273),
.Y(n_336)
);

INVx3_ASAP7_75t_L g337 ( 
.A(n_277),
.Y(n_337)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_277),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_301),
.B(n_260),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_293),
.B(n_260),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_270),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g342 ( 
.A(n_290),
.Y(n_342)
);

OR2x6_ASAP7_75t_L g343 ( 
.A(n_304),
.B(n_284),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_277),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_271),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_281),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_282),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_298),
.B(n_197),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_286),
.Y(n_349)
);

INVx3_ASAP7_75t_L g350 ( 
.A(n_286),
.Y(n_350)
);

BUFx10_ASAP7_75t_L g351 ( 
.A(n_308),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_306),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_283),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_276),
.B(n_199),
.Y(n_354)
);

INVx5_ASAP7_75t_L g355 ( 
.A(n_265),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_269),
.B(n_230),
.Y(n_356)
);

INVx3_ASAP7_75t_L g357 ( 
.A(n_288),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_269),
.B(n_291),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_304),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_288),
.Y(n_360)
);

AND2x4_ASAP7_75t_L g361 ( 
.A(n_294),
.B(n_1),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_274),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_305),
.B(n_201),
.Y(n_363)
);

INVx3_ASAP7_75t_L g364 ( 
.A(n_296),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_307),
.B(n_202),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_280),
.Y(n_366)
);

INVx1_ASAP7_75t_SL g367 ( 
.A(n_295),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_280),
.B(n_203),
.Y(n_368)
);

BUFx3_ASAP7_75t_L g369 ( 
.A(n_296),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_272),
.Y(n_370)
);

OR2x2_ASAP7_75t_L g371 ( 
.A(n_308),
.B(n_1),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_300),
.Y(n_372)
);

AND2x4_ASAP7_75t_L g373 ( 
.A(n_285),
.B(n_2),
.Y(n_373)
);

INVx2_ASAP7_75t_SL g374 ( 
.A(n_295),
.Y(n_374)
);

AND2x6_ASAP7_75t_L g375 ( 
.A(n_285),
.B(n_19),
.Y(n_375)
);

AND2x4_ASAP7_75t_L g376 ( 
.A(n_302),
.B(n_2),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_367),
.A2(n_278),
.B1(n_303),
.B2(n_310),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_366),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_334),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_329),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_349),
.Y(n_381)
);

NAND2xp33_ASAP7_75t_L g382 ( 
.A(n_323),
.B(n_309),
.Y(n_382)
);

OAI221xp5_ASAP7_75t_L g383 ( 
.A1(n_367),
.A2(n_292),
.B1(n_278),
.B2(n_287),
.C(n_275),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_333),
.A2(n_274),
.B1(n_275),
.B2(n_5),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_311),
.Y(n_385)
);

OAI22xp33_ASAP7_75t_SL g386 ( 
.A1(n_343),
.A2(n_3),
.B1(n_4),
.B2(n_7),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_317),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_327),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_341),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_332),
.B(n_265),
.Y(n_390)
);

AO22x2_ASAP7_75t_L g391 ( 
.A1(n_335),
.A2(n_3),
.B1(n_4),
.B2(n_8),
.Y(n_391)
);

AO22x2_ASAP7_75t_L g392 ( 
.A1(n_315),
.A2(n_356),
.B1(n_320),
.B2(n_373),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_329),
.Y(n_393)
);

AO22x2_ASAP7_75t_L g394 ( 
.A1(n_315),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_345),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_339),
.Y(n_396)
);

OAI221xp5_ASAP7_75t_L g397 ( 
.A1(n_374),
.A2(n_268),
.B1(n_265),
.B2(n_12),
.C(n_13),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_346),
.Y(n_398)
);

NAND2x1p5_ASAP7_75t_L g399 ( 
.A(n_358),
.B(n_265),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_353),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_325),
.Y(n_401)
);

AO22x2_ASAP7_75t_L g402 ( 
.A1(n_320),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_325),
.Y(n_403)
);

AO22x2_ASAP7_75t_L g404 ( 
.A1(n_320),
.A2(n_11),
.B1(n_14),
.B2(n_15),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_339),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_330),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_330),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_352),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_328),
.Y(n_409)
);

AOI22xp33_ASAP7_75t_L g410 ( 
.A1(n_321),
.A2(n_265),
.B1(n_268),
.B2(n_16),
.Y(n_410)
);

OAI22xp33_ASAP7_75t_SL g411 ( 
.A1(n_343),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_411)
);

NOR2xp67_ASAP7_75t_L g412 ( 
.A(n_370),
.B(n_25),
.Y(n_412)
);

BUFx3_ASAP7_75t_L g413 ( 
.A(n_326),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_328),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_331),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_326),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_331),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_336),
.Y(n_418)
);

AO22x2_ASAP7_75t_L g419 ( 
.A1(n_373),
.A2(n_26),
.B1(n_30),
.B2(n_31),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_332),
.B(n_268),
.Y(n_420)
);

OR2x6_ASAP7_75t_L g421 ( 
.A(n_343),
.B(n_376),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_336),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_330),
.Y(n_423)
);

AO22x2_ASAP7_75t_L g424 ( 
.A1(n_371),
.A2(n_32),
.B1(n_35),
.B2(n_36),
.Y(n_424)
);

NAND2x1p5_ASAP7_75t_L g425 ( 
.A(n_342),
.B(n_268),
.Y(n_425)
);

INVx3_ASAP7_75t_L g426 ( 
.A(n_369),
.Y(n_426)
);

NOR2xp67_ASAP7_75t_L g427 ( 
.A(n_340),
.B(n_37),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_340),
.B(n_268),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_330),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_347),
.Y(n_430)
);

AO22x2_ASAP7_75t_L g431 ( 
.A1(n_376),
.A2(n_38),
.B1(n_40),
.B2(n_41),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_347),
.Y(n_432)
);

CKINVDCx16_ASAP7_75t_R g433 ( 
.A(n_351),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_333),
.B(n_158),
.Y(n_434)
);

NAND2x1p5_ASAP7_75t_L g435 ( 
.A(n_361),
.B(n_43),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_R g436 ( 
.A(n_359),
.B(n_45),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_337),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_351),
.B(n_46),
.Y(n_438)
);

OAI221xp5_ASAP7_75t_L g439 ( 
.A1(n_372),
.A2(n_47),
.B1(n_49),
.B2(n_55),
.C(n_58),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_360),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_350),
.Y(n_441)
);

AO22x2_ASAP7_75t_L g442 ( 
.A1(n_361),
.A2(n_59),
.B1(n_61),
.B2(n_62),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_319),
.B(n_63),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_348),
.B(n_157),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_347),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_396),
.B(n_319),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_405),
.B(n_321),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_408),
.B(n_426),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_426),
.B(n_348),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_377),
.B(n_365),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_433),
.B(n_412),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_379),
.B(n_365),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_443),
.B(n_436),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_427),
.B(n_363),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_438),
.B(n_363),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_435),
.B(n_364),
.Y(n_456)
);

NAND2xp33_ASAP7_75t_SL g457 ( 
.A(n_444),
.B(n_354),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_385),
.B(n_321),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_380),
.B(n_364),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_393),
.B(n_369),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_428),
.B(n_354),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_387),
.B(n_321),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_399),
.B(n_368),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_388),
.B(n_368),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_389),
.B(n_337),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_395),
.B(n_398),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_400),
.B(n_338),
.Y(n_467)
);

AND2x4_ASAP7_75t_L g468 ( 
.A(n_421),
.B(n_321),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_386),
.B(n_338),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_411),
.B(n_318),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_410),
.B(n_318),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_378),
.B(n_318),
.Y(n_472)
);

AND2x4_ASAP7_75t_L g473 ( 
.A(n_421),
.B(n_375),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_378),
.B(n_318),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_401),
.B(n_313),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_434),
.B(n_441),
.Y(n_476)
);

NAND2xp33_ASAP7_75t_SL g477 ( 
.A(n_416),
.B(n_313),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_441),
.B(n_316),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_403),
.B(n_409),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_414),
.B(n_415),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_417),
.B(n_316),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_418),
.B(n_375),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_422),
.B(n_314),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_437),
.B(n_314),
.Y(n_484)
);

NAND2xp33_ASAP7_75t_SL g485 ( 
.A(n_384),
.B(n_312),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_425),
.B(n_344),
.Y(n_486)
);

NAND2xp33_ASAP7_75t_SL g487 ( 
.A(n_431),
.B(n_419),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_445),
.B(n_347),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_406),
.B(n_322),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_392),
.B(n_350),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_383),
.B(n_375),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_407),
.B(n_324),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_423),
.B(n_357),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_392),
.B(n_357),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_381),
.B(n_375),
.Y(n_495)
);

NAND2xp33_ASAP7_75t_SL g496 ( 
.A(n_431),
.B(n_419),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_429),
.B(n_355),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_430),
.B(n_355),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_432),
.B(n_355),
.Y(n_499)
);

AOI21xp5_ASAP7_75t_L g500 ( 
.A1(n_457),
.A2(n_382),
.B(n_390),
.Y(n_500)
);

AOI21xp5_ASAP7_75t_L g501 ( 
.A1(n_476),
.A2(n_420),
.B(n_442),
.Y(n_501)
);

AOI21x1_ASAP7_75t_L g502 ( 
.A1(n_454),
.A2(n_440),
.B(n_381),
.Y(n_502)
);

OAI21x1_ASAP7_75t_L g503 ( 
.A1(n_495),
.A2(n_440),
.B(n_362),
.Y(n_503)
);

BUFx2_ASAP7_75t_L g504 ( 
.A(n_477),
.Y(n_504)
);

AOI21x1_ASAP7_75t_SL g505 ( 
.A1(n_475),
.A2(n_424),
.B(n_323),
.Y(n_505)
);

NOR2xp67_ASAP7_75t_SL g506 ( 
.A(n_453),
.B(n_413),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_L g507 ( 
.A1(n_450),
.A2(n_442),
.B1(n_424),
.B2(n_391),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_466),
.Y(n_508)
);

INVx5_ASAP7_75t_L g509 ( 
.A(n_468),
.Y(n_509)
);

BUFx12f_ASAP7_75t_L g510 ( 
.A(n_468),
.Y(n_510)
);

AOI21xp5_ASAP7_75t_L g511 ( 
.A1(n_461),
.A2(n_439),
.B(n_397),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_490),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_446),
.B(n_391),
.Y(n_513)
);

OA21x2_ASAP7_75t_L g514 ( 
.A1(n_491),
.A2(n_482),
.B(n_471),
.Y(n_514)
);

BUFx6f_ASAP7_75t_SL g515 ( 
.A(n_473),
.Y(n_515)
);

INVxp67_ASAP7_75t_L g516 ( 
.A(n_452),
.Y(n_516)
);

AOI21xp5_ASAP7_75t_L g517 ( 
.A1(n_447),
.A2(n_355),
.B(n_323),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_473),
.B(n_394),
.Y(n_518)
);

OAI21xp5_ASAP7_75t_L g519 ( 
.A1(n_464),
.A2(n_323),
.B(n_375),
.Y(n_519)
);

OA22x2_ASAP7_75t_L g520 ( 
.A1(n_455),
.A2(n_404),
.B1(n_402),
.B2(n_394),
.Y(n_520)
);

OAI21xp5_ASAP7_75t_L g521 ( 
.A1(n_458),
.A2(n_462),
.B(n_469),
.Y(n_521)
);

AOI21xp5_ASAP7_75t_L g522 ( 
.A1(n_449),
.A2(n_323),
.B(n_404),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_494),
.Y(n_523)
);

AOI21xp33_ASAP7_75t_L g524 ( 
.A1(n_470),
.A2(n_402),
.B(n_65),
.Y(n_524)
);

OAI21x1_ASAP7_75t_L g525 ( 
.A1(n_472),
.A2(n_64),
.B(n_66),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_465),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_R g527 ( 
.A(n_487),
.B(n_67),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_496),
.B(n_68),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_448),
.B(n_71),
.Y(n_529)
);

AOI21xp5_ASAP7_75t_SL g530 ( 
.A1(n_456),
.A2(n_74),
.B(n_76),
.Y(n_530)
);

OAI21x1_ASAP7_75t_L g531 ( 
.A1(n_474),
.A2(n_77),
.B(n_78),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_451),
.B(n_79),
.Y(n_532)
);

OAI21x1_ASAP7_75t_L g533 ( 
.A1(n_488),
.A2(n_80),
.B(n_81),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_459),
.Y(n_534)
);

OA21x2_ASAP7_75t_L g535 ( 
.A1(n_463),
.A2(n_82),
.B(n_84),
.Y(n_535)
);

AOI21xp5_ASAP7_75t_L g536 ( 
.A1(n_478),
.A2(n_85),
.B(n_87),
.Y(n_536)
);

OAI21x1_ASAP7_75t_L g537 ( 
.A1(n_486),
.A2(n_90),
.B(n_91),
.Y(n_537)
);

AOI211x1_ASAP7_75t_L g538 ( 
.A1(n_467),
.A2(n_479),
.B(n_480),
.C(n_483),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_460),
.B(n_92),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_493),
.B(n_94),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_485),
.B(n_484),
.Y(n_541)
);

NOR2xp67_ASAP7_75t_L g542 ( 
.A(n_497),
.B(n_95),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_489),
.B(n_96),
.Y(n_543)
);

OAI21xp5_ASAP7_75t_L g544 ( 
.A1(n_511),
.A2(n_481),
.B(n_492),
.Y(n_544)
);

OAI21xp5_ASAP7_75t_L g545 ( 
.A1(n_501),
.A2(n_498),
.B(n_499),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_502),
.Y(n_546)
);

NAND3xp33_ASAP7_75t_SL g547 ( 
.A(n_507),
.B(n_97),
.C(n_98),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_503),
.Y(n_548)
);

OAI21x1_ASAP7_75t_L g549 ( 
.A1(n_500),
.A2(n_99),
.B(n_100),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_L g550 ( 
.A1(n_507),
.A2(n_102),
.B1(n_103),
.B2(n_105),
.Y(n_550)
);

OA21x2_ASAP7_75t_L g551 ( 
.A1(n_521),
.A2(n_106),
.B(n_110),
.Y(n_551)
);

INVx2_ASAP7_75t_SL g552 ( 
.A(n_509),
.Y(n_552)
);

OAI21x1_ASAP7_75t_L g553 ( 
.A1(n_517),
.A2(n_531),
.B(n_525),
.Y(n_553)
);

OR2x6_ASAP7_75t_L g554 ( 
.A(n_510),
.B(n_111),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_508),
.Y(n_555)
);

AOI21x1_ASAP7_75t_L g556 ( 
.A1(n_522),
.A2(n_112),
.B(n_114),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_512),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_523),
.Y(n_558)
);

BUFx3_ASAP7_75t_L g559 ( 
.A(n_509),
.Y(n_559)
);

A2O1A1Ixp33_ASAP7_75t_L g560 ( 
.A1(n_524),
.A2(n_115),
.B(n_116),
.C(n_117),
.Y(n_560)
);

NAND2x1p5_ASAP7_75t_L g561 ( 
.A(n_509),
.B(n_119),
.Y(n_561)
);

AND2x4_ASAP7_75t_L g562 ( 
.A(n_504),
.B(n_120),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_514),
.Y(n_563)
);

BUFx3_ASAP7_75t_L g564 ( 
.A(n_526),
.Y(n_564)
);

OAI21xp5_ASAP7_75t_L g565 ( 
.A1(n_521),
.A2(n_121),
.B(n_122),
.Y(n_565)
);

OAI21x1_ASAP7_75t_L g566 ( 
.A1(n_533),
.A2(n_124),
.B(n_126),
.Y(n_566)
);

AOI21xp5_ASAP7_75t_L g567 ( 
.A1(n_519),
.A2(n_127),
.B(n_129),
.Y(n_567)
);

AOI22xp33_ASAP7_75t_L g568 ( 
.A1(n_520),
.A2(n_130),
.B1(n_131),
.B2(n_132),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_534),
.Y(n_569)
);

BUFx6f_ASAP7_75t_L g570 ( 
.A(n_528),
.Y(n_570)
);

AO21x1_ASAP7_75t_L g571 ( 
.A1(n_524),
.A2(n_133),
.B(n_134),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g572 ( 
.A(n_528),
.Y(n_572)
);

OAI21x1_ASAP7_75t_L g573 ( 
.A1(n_537),
.A2(n_135),
.B(n_136),
.Y(n_573)
);

OAI21x1_ASAP7_75t_L g574 ( 
.A1(n_505),
.A2(n_137),
.B(n_138),
.Y(n_574)
);

INVx3_ASAP7_75t_L g575 ( 
.A(n_515),
.Y(n_575)
);

O2A1O1Ixp33_ASAP7_75t_L g576 ( 
.A1(n_541),
.A2(n_139),
.B(n_140),
.C(n_141),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_516),
.Y(n_577)
);

BUFx3_ASAP7_75t_L g578 ( 
.A(n_532),
.Y(n_578)
);

AOI21xp5_ASAP7_75t_L g579 ( 
.A1(n_519),
.A2(n_142),
.B(n_143),
.Y(n_579)
);

OAI22xp5_ASAP7_75t_L g580 ( 
.A1(n_513),
.A2(n_144),
.B1(n_148),
.B2(n_149),
.Y(n_580)
);

OR2x6_ASAP7_75t_L g581 ( 
.A(n_538),
.B(n_151),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_518),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_535),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_535),
.Y(n_584)
);

AO21x2_ASAP7_75t_L g585 ( 
.A1(n_583),
.A2(n_527),
.B(n_539),
.Y(n_585)
);

AOI22xp33_ASAP7_75t_L g586 ( 
.A1(n_568),
.A2(n_515),
.B1(n_506),
.B2(n_529),
.Y(n_586)
);

HB1xp67_ASAP7_75t_L g587 ( 
.A(n_564),
.Y(n_587)
);

OAI21x1_ASAP7_75t_L g588 ( 
.A1(n_553),
.A2(n_536),
.B(n_543),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_546),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_546),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_563),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_563),
.Y(n_592)
);

BUFx3_ASAP7_75t_L g593 ( 
.A(n_559),
.Y(n_593)
);

HB1xp67_ASAP7_75t_L g594 ( 
.A(n_564),
.Y(n_594)
);

BUFx3_ASAP7_75t_L g595 ( 
.A(n_559),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_577),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_569),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_569),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_555),
.Y(n_599)
);

HB1xp67_ASAP7_75t_L g600 ( 
.A(n_582),
.Y(n_600)
);

INVx3_ASAP7_75t_L g601 ( 
.A(n_574),
.Y(n_601)
);

OAI21x1_ASAP7_75t_L g602 ( 
.A1(n_553),
.A2(n_540),
.B(n_530),
.Y(n_602)
);

OAI21x1_ASAP7_75t_L g603 ( 
.A1(n_556),
.A2(n_542),
.B(n_152),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_548),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_548),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_570),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_583),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_570),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_570),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_584),
.Y(n_610)
);

OR2x6_ASAP7_75t_L g611 ( 
.A(n_570),
.B(n_154),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_578),
.B(n_562),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_572),
.Y(n_613)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_557),
.B(n_558),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_572),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_572),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_572),
.Y(n_617)
);

OR2x2_ASAP7_75t_L g618 ( 
.A(n_578),
.B(n_581),
.Y(n_618)
);

OAI21x1_ASAP7_75t_L g619 ( 
.A1(n_549),
.A2(n_574),
.B(n_566),
.Y(n_619)
);

BUFx6f_ASAP7_75t_L g620 ( 
.A(n_551),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_551),
.Y(n_621)
);

OA21x2_ASAP7_75t_L g622 ( 
.A1(n_545),
.A2(n_565),
.B(n_544),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_562),
.B(n_575),
.Y(n_623)
);

INVx3_ASAP7_75t_L g624 ( 
.A(n_551),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_581),
.Y(n_625)
);

AND2x2_ASAP7_75t_L g626 ( 
.A(n_562),
.B(n_581),
.Y(n_626)
);

BUFx2_ASAP7_75t_L g627 ( 
.A(n_549),
.Y(n_627)
);

AO21x2_ASAP7_75t_L g628 ( 
.A1(n_547),
.A2(n_560),
.B(n_571),
.Y(n_628)
);

INVx2_ASAP7_75t_SL g629 ( 
.A(n_575),
.Y(n_629)
);

BUFx3_ASAP7_75t_L g630 ( 
.A(n_552),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_573),
.Y(n_631)
);

NAND3xp33_ASAP7_75t_L g632 ( 
.A(n_568),
.B(n_560),
.C(n_550),
.Y(n_632)
);

OR2x6_ASAP7_75t_L g633 ( 
.A(n_561),
.B(n_552),
.Y(n_633)
);

XNOR2xp5_ASAP7_75t_L g634 ( 
.A(n_596),
.B(n_554),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_614),
.B(n_554),
.Y(n_635)
);

BUFx3_ASAP7_75t_L g636 ( 
.A(n_593),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_599),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_599),
.Y(n_638)
);

OR2x6_ASAP7_75t_L g639 ( 
.A(n_618),
.B(n_554),
.Y(n_639)
);

BUFx3_ASAP7_75t_L g640 ( 
.A(n_593),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_626),
.B(n_561),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_629),
.B(n_576),
.Y(n_642)
);

BUFx10_ASAP7_75t_L g643 ( 
.A(n_629),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_614),
.B(n_580),
.Y(n_644)
);

BUFx3_ASAP7_75t_L g645 ( 
.A(n_593),
.Y(n_645)
);

NAND2xp33_ASAP7_75t_R g646 ( 
.A(n_626),
.B(n_567),
.Y(n_646)
);

NAND2xp33_ASAP7_75t_R g647 ( 
.A(n_612),
.B(n_579),
.Y(n_647)
);

NAND2xp33_ASAP7_75t_R g648 ( 
.A(n_623),
.B(n_618),
.Y(n_648)
);

NAND2xp33_ASAP7_75t_R g649 ( 
.A(n_611),
.B(n_633),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_600),
.Y(n_650)
);

BUFx3_ASAP7_75t_L g651 ( 
.A(n_595),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_597),
.Y(n_652)
);

AND2x4_ASAP7_75t_L g653 ( 
.A(n_587),
.B(n_573),
.Y(n_653)
);

CKINVDCx16_ASAP7_75t_R g654 ( 
.A(n_595),
.Y(n_654)
);

NAND2xp33_ASAP7_75t_R g655 ( 
.A(n_611),
.B(n_566),
.Y(n_655)
);

AND2x4_ASAP7_75t_L g656 ( 
.A(n_594),
.B(n_595),
.Y(n_656)
);

AND2x4_ASAP7_75t_L g657 ( 
.A(n_630),
.B(n_625),
.Y(n_657)
);

AND2x4_ASAP7_75t_L g658 ( 
.A(n_630),
.B(n_625),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_586),
.B(n_630),
.Y(n_659)
);

OR2x4_ASAP7_75t_L g660 ( 
.A(n_606),
.B(n_608),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_597),
.Y(n_661)
);

NAND2xp33_ASAP7_75t_SL g662 ( 
.A(n_628),
.B(n_627),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_598),
.Y(n_663)
);

NAND2xp33_ASAP7_75t_R g664 ( 
.A(n_611),
.B(n_633),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_R g665 ( 
.A(n_606),
.B(n_609),
.Y(n_665)
);

NAND2xp33_ASAP7_75t_R g666 ( 
.A(n_611),
.B(n_633),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_R g667 ( 
.A(n_608),
.B(n_609),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_632),
.B(n_613),
.Y(n_668)
);

INVxp67_ASAP7_75t_L g669 ( 
.A(n_613),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_R g670 ( 
.A(n_616),
.B(n_617),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_589),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_616),
.B(n_617),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_589),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_638),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_650),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_671),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_657),
.B(n_617),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_654),
.B(n_622),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_656),
.B(n_615),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_657),
.B(n_622),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_637),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_656),
.B(n_622),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_665),
.B(n_620),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_671),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_668),
.B(n_628),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_673),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_673),
.Y(n_687)
);

AOI22xp33_ASAP7_75t_L g688 ( 
.A1(n_644),
.A2(n_628),
.B1(n_585),
.B2(n_622),
.Y(n_688)
);

INVx2_ASAP7_75t_SL g689 ( 
.A(n_660),
.Y(n_689)
);

OR2x2_ASAP7_75t_L g690 ( 
.A(n_672),
.B(n_615),
.Y(n_690)
);

OAI222xp33_ASAP7_75t_L g691 ( 
.A1(n_639),
.A2(n_659),
.B1(n_635),
.B2(n_641),
.C1(n_611),
.C2(n_634),
.Y(n_691)
);

OR2x2_ASAP7_75t_L g692 ( 
.A(n_669),
.B(n_590),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_636),
.B(n_590),
.Y(n_693)
);

BUFx3_ASAP7_75t_L g694 ( 
.A(n_640),
.Y(n_694)
);

OAI22xp5_ASAP7_75t_L g695 ( 
.A1(n_639),
.A2(n_633),
.B1(n_627),
.B2(n_620),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_652),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_645),
.B(n_598),
.Y(n_697)
);

OR2x2_ASAP7_75t_L g698 ( 
.A(n_658),
.B(n_605),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_658),
.B(n_624),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_663),
.Y(n_700)
);

AND2x4_ASAP7_75t_L g701 ( 
.A(n_651),
.B(n_633),
.Y(n_701)
);

AND2x4_ASAP7_75t_L g702 ( 
.A(n_653),
.B(n_604),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_661),
.Y(n_703)
);

OAI221xp5_ASAP7_75t_SL g704 ( 
.A1(n_642),
.A2(n_624),
.B1(n_621),
.B2(n_631),
.C(n_601),
.Y(n_704)
);

AND2x2_ASAP7_75t_L g705 ( 
.A(n_679),
.B(n_643),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_676),
.Y(n_706)
);

AND3x2_ASAP7_75t_L g707 ( 
.A(n_685),
.B(n_653),
.C(n_621),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_694),
.B(n_699),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_676),
.Y(n_709)
);

BUFx2_ASAP7_75t_L g710 ( 
.A(n_694),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_686),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_685),
.B(n_662),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_686),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_684),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_689),
.B(n_643),
.Y(n_715)
);

AOI221xp5_ASAP7_75t_L g716 ( 
.A1(n_704),
.A2(n_620),
.B1(n_624),
.B2(n_667),
.C(n_670),
.Y(n_716)
);

AOI211xp5_ASAP7_75t_L g717 ( 
.A1(n_689),
.A2(n_691),
.B(n_678),
.C(n_695),
.Y(n_717)
);

AND2x4_ASAP7_75t_L g718 ( 
.A(n_680),
.B(n_605),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_687),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_675),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_674),
.Y(n_721)
);

AO21x2_ASAP7_75t_L g722 ( 
.A1(n_682),
.A2(n_631),
.B(n_605),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_681),
.Y(n_723)
);

INVxp67_ASAP7_75t_L g724 ( 
.A(n_712),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_708),
.B(n_680),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_710),
.B(n_699),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_718),
.Y(n_727)
);

NAND2x1p5_ASAP7_75t_L g728 ( 
.A(n_715),
.B(n_683),
.Y(n_728)
);

AND2x2_ASAP7_75t_L g729 ( 
.A(n_705),
.B(n_677),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_718),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_720),
.B(n_688),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_712),
.B(n_688),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_721),
.Y(n_733)
);

AND2x2_ASAP7_75t_L g734 ( 
.A(n_715),
.B(n_677),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_723),
.B(n_701),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_714),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_706),
.Y(n_737)
);

A2O1A1Ixp33_ASAP7_75t_L g738 ( 
.A1(n_732),
.A2(n_716),
.B(n_717),
.C(n_683),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_724),
.B(n_732),
.Y(n_739)
);

AOI22xp5_ASAP7_75t_L g740 ( 
.A1(n_731),
.A2(n_716),
.B1(n_648),
.B2(n_655),
.Y(n_740)
);

AO221x2_ASAP7_75t_L g741 ( 
.A1(n_736),
.A2(n_719),
.B1(n_713),
.B2(n_711),
.C(n_709),
.Y(n_741)
);

INVxp67_ASAP7_75t_L g742 ( 
.A(n_731),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_724),
.Y(n_743)
);

AND2x2_ASAP7_75t_L g744 ( 
.A(n_743),
.B(n_726),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_741),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_738),
.B(n_728),
.Y(n_746)
);

INVx3_ASAP7_75t_L g747 ( 
.A(n_739),
.Y(n_747)
);

OAI22xp5_ASAP7_75t_L g748 ( 
.A1(n_740),
.A2(n_728),
.B1(n_734),
.B2(n_725),
.Y(n_748)
);

NAND2xp33_ASAP7_75t_L g749 ( 
.A(n_744),
.B(n_735),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_747),
.Y(n_750)
);

NOR2xp67_ASAP7_75t_SL g751 ( 
.A(n_746),
.B(n_730),
.Y(n_751)
);

AOI22xp5_ASAP7_75t_L g752 ( 
.A1(n_745),
.A2(n_742),
.B1(n_646),
.B2(n_647),
.Y(n_752)
);

HB1xp67_ASAP7_75t_L g753 ( 
.A(n_750),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_749),
.B(n_747),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_753),
.Y(n_755)
);

NOR2x1_ASAP7_75t_L g756 ( 
.A(n_754),
.B(n_748),
.Y(n_756)
);

INVx2_ASAP7_75t_SL g757 ( 
.A(n_754),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_755),
.B(n_752),
.Y(n_758)
);

NAND4xp25_ASAP7_75t_L g759 ( 
.A(n_756),
.B(n_751),
.C(n_666),
.D(n_649),
.Y(n_759)
);

NOR5xp2_ASAP7_75t_L g760 ( 
.A(n_757),
.B(n_696),
.C(n_700),
.D(n_707),
.E(n_703),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_755),
.B(n_729),
.Y(n_761)
);

INVx2_ASAP7_75t_SL g762 ( 
.A(n_757),
.Y(n_762)
);

AOI222xp33_ASAP7_75t_L g763 ( 
.A1(n_758),
.A2(n_761),
.B1(n_762),
.B2(n_759),
.C1(n_760),
.C2(n_620),
.Y(n_763)
);

AOI32xp33_ASAP7_75t_L g764 ( 
.A1(n_758),
.A2(n_624),
.A3(n_727),
.B1(n_619),
.B2(n_701),
.Y(n_764)
);

AOI211xp5_ASAP7_75t_L g765 ( 
.A1(n_758),
.A2(n_620),
.B(n_693),
.C(n_701),
.Y(n_765)
);

AOI221xp5_ASAP7_75t_L g766 ( 
.A1(n_758),
.A2(n_620),
.B1(n_737),
.B2(n_733),
.C(n_722),
.Y(n_766)
);

AOI211xp5_ASAP7_75t_SL g767 ( 
.A1(n_758),
.A2(n_601),
.B(n_697),
.C(n_692),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_763),
.B(n_702),
.Y(n_768)
);

NOR2x1p5_ASAP7_75t_L g769 ( 
.A(n_764),
.B(n_601),
.Y(n_769)
);

AND2x4_ASAP7_75t_L g770 ( 
.A(n_767),
.B(n_707),
.Y(n_770)
);

NAND4xp75_ASAP7_75t_L g771 ( 
.A(n_766),
.B(n_664),
.C(n_631),
.D(n_674),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_768),
.B(n_765),
.Y(n_772)
);

NAND2xp33_ASAP7_75t_R g773 ( 
.A(n_770),
.B(n_603),
.Y(n_773)
);

XNOR2xp5_ASAP7_75t_L g774 ( 
.A(n_769),
.B(n_722),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_771),
.B(n_702),
.Y(n_775)
);

NAND2xp33_ASAP7_75t_SL g776 ( 
.A(n_769),
.B(n_601),
.Y(n_776)
);

AOI22xp5_ASAP7_75t_L g777 ( 
.A1(n_773),
.A2(n_585),
.B1(n_702),
.B2(n_603),
.Y(n_777)
);

BUFx2_ASAP7_75t_L g778 ( 
.A(n_772),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_774),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_775),
.Y(n_780)
);

AND2x4_ASAP7_75t_L g781 ( 
.A(n_776),
.B(n_690),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_778),
.Y(n_782)
);

OAI21x1_ASAP7_75t_L g783 ( 
.A1(n_780),
.A2(n_779),
.B(n_777),
.Y(n_783)
);

NAND2x1_ASAP7_75t_SL g784 ( 
.A(n_781),
.B(n_604),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_778),
.Y(n_785)
);

AOI22xp33_ASAP7_75t_L g786 ( 
.A1(n_779),
.A2(n_585),
.B1(n_698),
.B2(n_602),
.Y(n_786)
);

OAI21xp5_ASAP7_75t_L g787 ( 
.A1(n_778),
.A2(n_602),
.B(n_588),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_782),
.Y(n_788)
);

AOI31xp33_ASAP7_75t_L g789 ( 
.A1(n_788),
.A2(n_785),
.A3(n_787),
.B(n_783),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_789),
.B(n_784),
.Y(n_790)
);

AOI22xp5_ASAP7_75t_L g791 ( 
.A1(n_790),
.A2(n_786),
.B1(n_588),
.B2(n_619),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_791),
.Y(n_792)
);

OAI221xp5_ASAP7_75t_R g793 ( 
.A1(n_792),
.A2(n_604),
.B1(n_592),
.B2(n_591),
.C(n_610),
.Y(n_793)
);

AOI211xp5_ASAP7_75t_L g794 ( 
.A1(n_793),
.A2(n_591),
.B(n_592),
.C(n_607),
.Y(n_794)
);


endmodule