module real_jpeg_7049_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g64 ( 
.A(n_0),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_1),
.Y(n_433)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_2),
.Y(n_77)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_2),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_2),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_3),
.A2(n_38),
.B1(n_54),
.B2(n_230),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_3),
.Y(n_230)
);

OAI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_3),
.A2(n_143),
.B1(n_230),
.B2(n_245),
.Y(n_244)
);

OAI22xp33_ASAP7_75t_SL g346 ( 
.A1(n_3),
.A2(n_230),
.B1(n_347),
.B2(n_348),
.Y(n_346)
);

AOI22xp33_ASAP7_75t_L g370 ( 
.A1(n_3),
.A2(n_171),
.B1(n_230),
.B2(n_371),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_4),
.A2(n_37),
.B1(n_42),
.B2(n_45),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_4),
.Y(n_45)
);

OAI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_4),
.A2(n_45),
.B1(n_124),
.B2(n_125),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_4),
.A2(n_45),
.B1(n_160),
.B2(n_162),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_4),
.A2(n_45),
.B1(n_219),
.B2(n_221),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_5),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_5),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_5),
.A2(n_39),
.B1(n_142),
.B2(n_143),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_5),
.A2(n_39),
.B1(n_184),
.B2(n_186),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_5),
.A2(n_39),
.B1(n_264),
.B2(n_266),
.Y(n_263)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_6),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_7),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_7),
.Y(n_176)
);

INVx8_ASAP7_75t_L g214 ( 
.A(n_7),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_7),
.Y(n_279)
);

BUFx5_ASAP7_75t_L g386 ( 
.A(n_7),
.Y(n_386)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_8),
.Y(n_261)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx3_ASAP7_75t_L g430 ( 
.A(n_10),
.Y(n_430)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_11),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_12),
.A2(n_85),
.B1(n_87),
.B2(n_88),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_12),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_12),
.A2(n_87),
.B1(n_104),
.B2(n_106),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_12),
.A2(n_87),
.B1(n_178),
.B2(n_181),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_12),
.B(n_25),
.Y(n_274)
);

O2A1O1Ixp33_ASAP7_75t_L g331 ( 
.A1(n_12),
.A2(n_93),
.B(n_332),
.C(n_339),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_12),
.B(n_361),
.C(n_362),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_12),
.B(n_147),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_12),
.B(n_279),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_12),
.B(n_71),
.Y(n_398)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_13),
.Y(n_66)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_13),
.Y(n_69)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_13),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g361 ( 
.A(n_13),
.Y(n_361)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_428),
.B(n_431),
.Y(n_14)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_196),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_195),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_148),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_19),
.B(n_148),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_138),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_131),
.B2(n_132),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_55),
.B1(n_56),
.B2(n_130),
.Y(n_22)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_23),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_36),
.B(n_40),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_24),
.A2(n_193),
.B(n_194),
.Y(n_192)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NOR2x1_ASAP7_75t_L g46 ( 
.A(n_25),
.B(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_25),
.B(n_41),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_25),
.B(n_135),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_25),
.B(n_229),
.Y(n_239)
);

AO22x2_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_28),
.B1(n_32),
.B2(n_34),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_31),
.Y(n_105)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_31),
.Y(n_109)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_31),
.Y(n_116)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_31),
.Y(n_128)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_33),
.Y(n_258)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx8_ASAP7_75t_L g137 ( 
.A(n_37),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_40),
.B(n_239),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_46),
.Y(n_40)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_46),
.B(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_46),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_46),
.B(n_229),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_50),
.B1(n_52),
.B2(n_54),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_48),
.A2(n_87),
.B(n_136),
.Y(n_135)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_51),
.Y(n_53)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_51),
.Y(n_251)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_57),
.A2(n_89),
.B1(n_90),
.B2(n_129),
.Y(n_56)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_57),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_57),
.A2(n_129),
.B1(n_139),
.B2(n_152),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_57),
.A2(n_129),
.B1(n_241),
.B2(n_247),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_57),
.B(n_238),
.C(n_241),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_82),
.B(n_83),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_58),
.A2(n_183),
.B(n_190),
.Y(n_182)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_59),
.B(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_59),
.B(n_84),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_59),
.B(n_346),
.Y(n_345)
);

NOR2x1_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_71),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_65),
.B1(n_67),
.B2(n_70),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_63),
.Y(n_97)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_63),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_63),
.Y(n_185)
);

INVx6_ASAP7_75t_L g338 ( 
.A(n_63),
.Y(n_338)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_64),
.Y(n_96)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_64),
.Y(n_164)
);

INVx3_ASAP7_75t_L g350 ( 
.A(n_64),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_64),
.Y(n_359)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

AO22x2_ASAP7_75t_L g71 ( 
.A1(n_68),
.A2(n_72),
.B1(n_74),
.B2(n_78),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_71),
.B(n_159),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_71),
.B(n_346),
.Y(n_365)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g220 ( 
.A(n_77),
.Y(n_220)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx5_ASAP7_75t_L g222 ( 
.A(n_80),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_81),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g363 ( 
.A(n_81),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_82),
.B(n_83),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_82),
.A2(n_158),
.B(n_183),
.Y(n_223)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_86),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_87),
.B(n_137),
.Y(n_136)
);

OAI21xp33_ASAP7_75t_L g332 ( 
.A1(n_87),
.A2(n_333),
.B(n_336),
.Y(n_332)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_110),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_91),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_102),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_92),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_95),
.B1(n_97),
.B2(n_98),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_94),
.Y(n_101)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_94),
.Y(n_114)
);

INVx5_ASAP7_75t_L g347 ( 
.A(n_95),
.Y(n_347)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_100),
.Y(n_118)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVxp67_ASAP7_75t_SL g102 ( 
.A(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_103),
.B(n_140),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_103),
.A2(n_140),
.B(n_147),
.Y(n_302)
);

INVx6_ASAP7_75t_SL g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_109),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_109),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g144 ( 
.A(n_109),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_109),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_110),
.A2(n_141),
.B(n_147),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_110),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_111),
.B(n_122),
.Y(n_110)
);

INVx1_ASAP7_75t_SL g140 ( 
.A(n_111),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_115),
.B1(n_117),
.B2(n_119),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx4_ASAP7_75t_L g335 ( 
.A(n_114),
.Y(n_335)
);

AOI32xp33_ASAP7_75t_L g250 ( 
.A1(n_115),
.A2(n_251),
.A3(n_252),
.B1(n_255),
.B2(n_256),
.Y(n_250)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_SL g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_120),
.Y(n_142)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_123),
.B(n_147),
.Y(n_146)
);

INVx6_ASAP7_75t_L g246 ( 
.A(n_124),
.Y(n_246)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_129),
.B(n_132),
.C(n_139),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_131),
.A2(n_132),
.B1(n_150),
.B2(n_151),
.Y(n_149)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_134),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_133),
.B(n_228),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_134),
.B(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_135),
.Y(n_194)
);

INVxp33_ASAP7_75t_L g255 ( 
.A(n_136),
.Y(n_255)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_139),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_141),
.B(n_145),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_140),
.B(n_244),
.Y(n_272)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_146),
.B(n_225),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_146),
.B(n_272),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_147),
.B(n_244),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_153),
.C(n_166),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_149),
.A2(n_153),
.B1(n_154),
.B2(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_149),
.Y(n_200)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_154),
.A2(n_155),
.B(n_165),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_155),
.B(n_165),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_157),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_156),
.Y(n_344)
);

INVxp67_ASAP7_75t_SL g157 ( 
.A(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_158),
.B(n_365),
.Y(n_407)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_164),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_166),
.B(n_199),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_191),
.B(n_192),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_167),
.A2(n_168),
.B1(n_203),
.B2(n_204),
.Y(n_202)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_182),
.Y(n_168)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_169),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_169),
.A2(n_191),
.B1(n_192),
.B2(n_205),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_169),
.A2(n_182),
.B1(n_191),
.B2(n_314),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_169),
.B(n_331),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_169),
.A2(n_191),
.B1(n_331),
.B2(n_410),
.Y(n_409)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_175),
.B(n_177),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_170),
.B(n_218),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_170),
.B(n_177),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_170),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_170),
.B(n_370),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_173),
.Y(n_170)
);

INVx8_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_172),
.Y(n_181)
);

INVx4_ASAP7_75t_L g372 ( 
.A(n_172),
.Y(n_372)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_177),
.Y(n_215)
);

INVx5_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

BUFx5_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_180),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_182),
.Y(n_314)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

AND2x2_ASAP7_75t_SL g286 ( 
.A(n_190),
.B(n_287),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_190),
.B(n_345),
.Y(n_374)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_192),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_231),
.B(n_427),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_198),
.B(n_201),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_198),
.B(n_201),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_206),
.C(n_208),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_202),
.A2(n_206),
.B1(n_207),
.B2(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_202),
.Y(n_318)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_208),
.B(n_317),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_224),
.C(n_226),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_209),
.A2(n_210),
.B1(n_311),
.B2(n_312),
.Y(n_310)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_223),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_211),
.B(n_223),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_216),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_212),
.B(n_368),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_215),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_214),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_216),
.B(n_383),
.Y(n_382)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_217),
.A2(n_263),
.B(n_268),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_218),
.B(n_278),
.Y(n_277)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_220),
.Y(n_265)
);

BUFx2_ASAP7_75t_L g267 ( 
.A(n_220),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_224),
.B(n_226),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_225),
.B(n_243),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_419),
.Y(n_232)
);

NAND3xp33_ASAP7_75t_SL g233 ( 
.A(n_234),
.B(n_307),
.C(n_321),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_294),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_280),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_236),
.B(n_280),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_248),
.C(n_270),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_237),
.B(n_324),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_238),
.B(n_240),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_241),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

INVx6_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_248),
.A2(n_249),
.B1(n_270),
.B2(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_262),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_250),
.B(n_262),
.Y(n_289)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx8_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

NAND2xp33_ASAP7_75t_SL g256 ( 
.A(n_257),
.B(n_259),
.Y(n_256)
);

INVx5_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_263),
.A2(n_277),
.B(n_285),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx8_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_270),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_273),
.C(n_275),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_271),
.B(n_328),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_272),
.B(n_293),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_273),
.A2(n_274),
.B1(n_275),
.B2(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_275),
.Y(n_329)
);

OR2x2_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_276),
.B(n_384),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_SL g397 ( 
.A(n_277),
.B(n_369),
.Y(n_397)
);

INVx4_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_288),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_282),
.B(n_283),
.C(n_288),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_286),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_284),
.B(n_286),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_287),
.B(n_365),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_SL g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_289),
.B(n_291),
.C(n_292),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g421 ( 
.A1(n_294),
.A2(n_422),
.B(n_423),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_295),
.B(n_306),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_295),
.B(n_306),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_296),
.B(n_298),
.C(n_299),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_301),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_300),
.B(n_303),
.C(n_304),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_302),
.A2(n_303),
.B1(n_304),
.B2(n_305),
.Y(n_301)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_302),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_303),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_319),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g425 ( 
.A(n_308),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_316),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_309),
.B(n_320),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_309),
.B(n_320),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_309),
.B(n_316),
.Y(n_426)
);

FAx1_ASAP7_75t_SL g309 ( 
.A(n_310),
.B(n_313),
.CI(n_315),
.CON(n_309),
.SN(n_309)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_319),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_322),
.A2(n_351),
.B(n_418),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_323),
.B(n_326),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_323),
.B(n_326),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_330),
.C(n_342),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_327),
.B(n_414),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_330),
.A2(n_342),
.B1(n_343),
.B2(n_415),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_330),
.Y(n_415)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_331),
.Y(n_410)
);

INVx4_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx8_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx3_ASAP7_75t_SL g336 ( 
.A(n_337),
.Y(n_336)
);

INVx8_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

BUFx12f_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_345),
.Y(n_343)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g351 ( 
.A1(n_352),
.A2(n_412),
.B(n_417),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_SL g352 ( 
.A1(n_353),
.A2(n_402),
.B(n_411),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_354),
.A2(n_378),
.B(n_401),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_366),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_355),
.B(n_366),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_364),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_356),
.A2(n_357),
.B1(n_364),
.B2(n_381),
.Y(n_380)
);

CKINVDCx16_ASAP7_75t_R g356 ( 
.A(n_357),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_360),
.Y(n_357)
);

INVx5_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_364),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_373),
.Y(n_366)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_367),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_370),
.B(n_385),
.Y(n_384)
);

INVx3_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_374),
.A2(n_375),
.B1(n_376),
.B2(n_377),
.Y(n_373)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_374),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_375),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_375),
.B(n_376),
.C(n_404),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_SL g378 ( 
.A1(n_379),
.A2(n_387),
.B(n_400),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_SL g379 ( 
.A(n_380),
.B(n_382),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_380),
.B(n_382),
.Y(n_400)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g387 ( 
.A1(n_388),
.A2(n_396),
.B(n_399),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_395),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_394),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVx6_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_397),
.B(n_398),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_397),
.B(n_398),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_405),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_403),
.B(n_405),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_409),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_408),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_407),
.B(n_408),
.C(n_409),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_413),
.B(n_416),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_413),
.B(n_416),
.Y(n_417)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g419 ( 
.A1(n_420),
.A2(n_421),
.B(n_424),
.C(n_425),
.D(n_426),
.Y(n_419)
);

BUFx4f_ASAP7_75t_SL g428 ( 
.A(n_429),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_429),
.Y(n_432)
);

INVx13_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_432),
.B(n_433),
.Y(n_431)
);


endmodule