module fake_jpeg_23742_n_59 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_59);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_59;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_27;
wire n_55;
wire n_51;
wire n_47;
wire n_40;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_36;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

INVx1_ASAP7_75t_L g26 ( 
.A(n_24),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_19),
.B(n_20),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx6_ASAP7_75t_SL g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_25),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_32),
.B(n_3),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_34),
.B(n_6),
.Y(n_43)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_36),
.Y(n_38)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_4),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_37),
.B(n_5),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_39),
.B(n_42),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_37),
.B(n_33),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_43),
.C(n_44),
.Y(n_48)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_41),
.A2(n_8),
.B1(n_12),
.B2(n_13),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_27),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_26),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_7),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_45),
.A2(n_31),
.B1(n_9),
.B2(n_11),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_46),
.B(n_14),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_49),
.A2(n_38),
.B(n_15),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_50),
.B(n_51),
.Y(n_53)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_51),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_52),
.B(n_47),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_54),
.B(n_53),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_55),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_56),
.B(n_48),
.C(n_17),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_16),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_58),
.A2(n_18),
.B1(n_21),
.B2(n_22),
.Y(n_59)
);


endmodule