module real_aes_8626_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_746;
wire n_153;
wire n_532;
wire n_284;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_504;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_754;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_527;
wire n_434;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_756;
wire n_288;
wire n_404;
wire n_598;
wire n_728;
wire n_713;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_749;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_762;
wire n_325;
wire n_575;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g109 ( .A(n_0), .Y(n_109) );
A2O1A1Ixp33_ASAP7_75t_L g224 ( .A1(n_1), .A2(n_147), .B(n_150), .C(n_225), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g174 ( .A1(n_2), .A2(n_175), .B(n_176), .Y(n_174) );
INVx1_ASAP7_75t_L g507 ( .A(n_3), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_4), .B(n_186), .Y(n_185) );
AOI21xp33_ASAP7_75t_L g484 ( .A1(n_5), .A2(n_175), .B(n_485), .Y(n_484) );
AND2x6_ASAP7_75t_L g147 ( .A(n_6), .B(n_148), .Y(n_147) );
INVx1_ASAP7_75t_L g250 ( .A(n_7), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_8), .B(n_115), .Y(n_114) );
NOR2xp33_ASAP7_75t_L g455 ( .A(n_8), .B(n_42), .Y(n_455) );
AOI21xp5_ASAP7_75t_L g547 ( .A1(n_9), .A2(n_274), .B(n_548), .Y(n_547) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_10), .B(n_159), .Y(n_227) );
INVx1_ASAP7_75t_L g489 ( .A(n_11), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_12), .B(n_180), .Y(n_540) );
INVx1_ASAP7_75t_L g139 ( .A(n_13), .Y(n_139) );
INVx1_ASAP7_75t_L g552 ( .A(n_14), .Y(n_552) );
A2O1A1Ixp33_ASAP7_75t_L g234 ( .A1(n_15), .A2(n_194), .B(n_235), .C(n_237), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_16), .B(n_186), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_17), .B(n_478), .Y(n_530) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_18), .B(n_175), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_19), .B(n_282), .Y(n_281) );
A2O1A1Ixp33_ASAP7_75t_L g210 ( .A1(n_20), .A2(n_180), .B(n_211), .C(n_214), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_21), .B(n_186), .Y(n_481) );
NAND2xp5_ASAP7_75t_SL g158 ( .A(n_22), .B(n_159), .Y(n_158) );
AOI22xp5_ASAP7_75t_L g103 ( .A1(n_23), .A2(n_104), .B1(n_116), .B2(n_763), .Y(n_103) );
A2O1A1Ixp33_ASAP7_75t_L g550 ( .A1(n_24), .A2(n_213), .B(n_237), .C(n_551), .Y(n_550) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_25), .B(n_159), .Y(n_195) );
CKINVDCx16_ASAP7_75t_R g141 ( .A(n_26), .Y(n_141) );
INVx1_ASAP7_75t_L g192 ( .A(n_27), .Y(n_192) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_28), .Y(n_146) );
CKINVDCx20_ASAP7_75t_R g223 ( .A(n_29), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_30), .B(n_159), .Y(n_508) );
INVx1_ASAP7_75t_L g279 ( .A(n_31), .Y(n_279) );
INVx1_ASAP7_75t_L g497 ( .A(n_32), .Y(n_497) );
AOI22xp5_ASAP7_75t_L g122 ( .A1(n_33), .A2(n_123), .B1(n_124), .B2(n_449), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g449 ( .A(n_33), .Y(n_449) );
INVx2_ASAP7_75t_L g145 ( .A(n_34), .Y(n_145) );
CKINVDCx20_ASAP7_75t_R g229 ( .A(n_35), .Y(n_229) );
NAND2xp5_ASAP7_75t_SL g456 ( .A(n_36), .B(n_457), .Y(n_456) );
A2O1A1Ixp33_ASAP7_75t_L g179 ( .A1(n_37), .A2(n_180), .B(n_181), .C(n_183), .Y(n_179) );
INVxp67_ASAP7_75t_L g280 ( .A(n_38), .Y(n_280) );
CKINVDCx14_ASAP7_75t_R g177 ( .A(n_39), .Y(n_177) );
A2O1A1Ixp33_ASAP7_75t_L g190 ( .A1(n_40), .A2(n_150), .B(n_191), .C(n_198), .Y(n_190) );
A2O1A1Ixp33_ASAP7_75t_L g518 ( .A1(n_41), .A2(n_147), .B(n_150), .C(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g115 ( .A(n_42), .Y(n_115) );
INVx1_ASAP7_75t_L g496 ( .A(n_43), .Y(n_496) );
OAI22xp5_ASAP7_75t_SL g446 ( .A1(n_44), .A2(n_52), .B1(n_447), .B2(n_448), .Y(n_446) );
CKINVDCx20_ASAP7_75t_R g448 ( .A(n_44), .Y(n_448) );
AOI22xp5_ASAP7_75t_L g752 ( .A1(n_45), .A2(n_65), .B1(n_753), .B2(n_754), .Y(n_752) );
CKINVDCx20_ASAP7_75t_R g754 ( .A(n_45), .Y(n_754) );
OAI22xp5_ASAP7_75t_SL g750 ( .A1(n_46), .A2(n_751), .B1(n_752), .B2(n_755), .Y(n_750) );
CKINVDCx20_ASAP7_75t_R g755 ( .A(n_46), .Y(n_755) );
A2O1A1Ixp33_ASAP7_75t_L g247 ( .A1(n_47), .A2(n_161), .B(n_248), .C(n_249), .Y(n_247) );
AOI222xp33_ASAP7_75t_L g459 ( .A1(n_48), .A2(n_460), .B1(n_749), .B2(n_750), .C1(n_756), .C2(n_759), .Y(n_459) );
NAND2xp5_ASAP7_75t_SL g529 ( .A(n_49), .B(n_159), .Y(n_529) );
CKINVDCx20_ASAP7_75t_R g200 ( .A(n_50), .Y(n_200) );
CKINVDCx20_ASAP7_75t_R g276 ( .A(n_51), .Y(n_276) );
CKINVDCx20_ASAP7_75t_R g447 ( .A(n_52), .Y(n_447) );
INVx1_ASAP7_75t_L g209 ( .A(n_53), .Y(n_209) );
CKINVDCx16_ASAP7_75t_R g498 ( .A(n_54), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_55), .B(n_175), .Y(n_542) );
AOI22xp5_ASAP7_75t_L g494 ( .A1(n_56), .A2(n_150), .B1(n_214), .B2(n_495), .Y(n_494) );
CKINVDCx20_ASAP7_75t_R g523 ( .A(n_57), .Y(n_523) );
CKINVDCx16_ASAP7_75t_R g504 ( .A(n_58), .Y(n_504) );
CKINVDCx14_ASAP7_75t_R g246 ( .A(n_59), .Y(n_246) );
A2O1A1Ixp33_ASAP7_75t_L g487 ( .A1(n_60), .A2(n_183), .B(n_248), .C(n_488), .Y(n_487) );
CKINVDCx20_ASAP7_75t_R g532 ( .A(n_61), .Y(n_532) );
INVx1_ASAP7_75t_L g486 ( .A(n_62), .Y(n_486) );
INVx1_ASAP7_75t_L g148 ( .A(n_63), .Y(n_148) );
INVx1_ASAP7_75t_L g138 ( .A(n_64), .Y(n_138) );
CKINVDCx20_ASAP7_75t_R g753 ( .A(n_65), .Y(n_753) );
INVx1_ASAP7_75t_SL g182 ( .A(n_66), .Y(n_182) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_67), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_68), .B(n_186), .Y(n_216) );
INVx1_ASAP7_75t_L g154 ( .A(n_69), .Y(n_154) );
A2O1A1Ixp33_ASAP7_75t_SL g477 ( .A1(n_70), .A2(n_183), .B(n_478), .C(n_479), .Y(n_477) );
INVxp67_ASAP7_75t_L g480 ( .A(n_71), .Y(n_480) );
INVx1_ASAP7_75t_L g112 ( .A(n_72), .Y(n_112) );
AOI21xp5_ASAP7_75t_L g244 ( .A1(n_73), .A2(n_175), .B(n_245), .Y(n_244) );
CKINVDCx20_ASAP7_75t_R g166 ( .A(n_74), .Y(n_166) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_75), .A2(n_175), .B(n_232), .Y(n_231) );
CKINVDCx20_ASAP7_75t_R g500 ( .A(n_76), .Y(n_500) );
INVx1_ASAP7_75t_L g526 ( .A(n_77), .Y(n_526) );
AOI21xp5_ASAP7_75t_L g273 ( .A1(n_78), .A2(n_274), .B(n_275), .Y(n_273) );
CKINVDCx16_ASAP7_75t_R g189 ( .A(n_79), .Y(n_189) );
INVx1_ASAP7_75t_L g233 ( .A(n_80), .Y(n_233) );
A2O1A1Ixp33_ASAP7_75t_L g527 ( .A1(n_81), .A2(n_147), .B(n_150), .C(n_528), .Y(n_527) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_82), .A2(n_175), .B(n_208), .Y(n_207) );
INVx1_ASAP7_75t_L g236 ( .A(n_83), .Y(n_236) );
NAND2xp5_ASAP7_75t_SL g520 ( .A(n_84), .B(n_193), .Y(n_520) );
INVx2_ASAP7_75t_L g136 ( .A(n_85), .Y(n_136) );
INVx1_ASAP7_75t_L g226 ( .A(n_86), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_87), .B(n_478), .Y(n_521) );
A2O1A1Ixp33_ASAP7_75t_L g505 ( .A1(n_88), .A2(n_147), .B(n_150), .C(n_506), .Y(n_505) );
NAND3xp33_ASAP7_75t_SL g108 ( .A(n_89), .B(n_109), .C(n_110), .Y(n_108) );
OR2x2_ASAP7_75t_L g452 ( .A(n_89), .B(n_453), .Y(n_452) );
INVx2_ASAP7_75t_L g464 ( .A(n_89), .Y(n_464) );
OR2x2_ASAP7_75t_L g747 ( .A(n_89), .B(n_454), .Y(n_747) );
A2O1A1Ixp33_ASAP7_75t_L g149 ( .A1(n_90), .A2(n_150), .B(n_153), .C(n_163), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_91), .B(n_168), .Y(n_490) );
CKINVDCx20_ASAP7_75t_R g511 ( .A(n_92), .Y(n_511) );
A2O1A1Ixp33_ASAP7_75t_L g537 ( .A1(n_93), .A2(n_147), .B(n_150), .C(n_538), .Y(n_537) );
CKINVDCx20_ASAP7_75t_R g544 ( .A(n_94), .Y(n_544) );
INVx1_ASAP7_75t_L g476 ( .A(n_95), .Y(n_476) );
CKINVDCx16_ASAP7_75t_R g549 ( .A(n_96), .Y(n_549) );
NAND2xp5_ASAP7_75t_SL g539 ( .A(n_97), .B(n_193), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_98), .B(n_134), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_99), .B(n_134), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_100), .B(n_112), .Y(n_111) );
INVx2_ASAP7_75t_L g212 ( .A(n_101), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g474 ( .A1(n_102), .A2(n_175), .B(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g763 ( .A(n_104), .Y(n_763) );
INVx1_ASAP7_75t_SL g104 ( .A(n_105), .Y(n_104) );
INVx2_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
AND2x2_ASAP7_75t_SL g106 ( .A(n_107), .B(n_113), .Y(n_106) );
CKINVDCx16_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
AND2x2_ASAP7_75t_L g454 ( .A(n_109), .B(n_455), .Y(n_454) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
INVxp67_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
AO21x2_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_121), .B(n_458), .Y(n_116) );
HB1xp67_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
BUFx3_ASAP7_75t_L g762 ( .A(n_118), .Y(n_762) );
INVx2_ASAP7_75t_SL g118 ( .A(n_119), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
OAI21xp5_ASAP7_75t_SL g121 ( .A1(n_122), .A2(n_450), .B(n_456), .Y(n_121) );
INVx1_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
XNOR2xp5_ASAP7_75t_L g124 ( .A(n_125), .B(n_446), .Y(n_124) );
INVx3_ASAP7_75t_L g748 ( .A(n_125), .Y(n_748) );
AOI22xp5_ASAP7_75t_L g760 ( .A1(n_125), .A2(n_462), .B1(n_746), .B2(n_761), .Y(n_760) );
AND2x2_ASAP7_75t_SL g125 ( .A(n_126), .B(n_401), .Y(n_125) );
NOR4xp25_ASAP7_75t_L g126 ( .A(n_127), .B(n_338), .C(n_372), .D(n_388), .Y(n_126) );
NAND4xp25_ASAP7_75t_SL g127 ( .A(n_128), .B(n_264), .C(n_302), .D(n_318), .Y(n_127) );
AOI222xp33_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_201), .B1(n_239), .B2(n_252), .C1(n_257), .C2(n_263), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
AOI31xp33_ASAP7_75t_L g434 ( .A1(n_130), .A2(n_435), .A3(n_436), .B(n_438), .Y(n_434) );
OR2x2_ASAP7_75t_L g130 ( .A(n_131), .B(n_169), .Y(n_130) );
AND2x2_ASAP7_75t_L g409 ( .A(n_131), .B(n_171), .Y(n_409) );
BUFx2_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx2_ASAP7_75t_SL g256 ( .A(n_132), .Y(n_256) );
AND2x2_ASAP7_75t_L g263 ( .A(n_132), .B(n_187), .Y(n_263) );
AND2x2_ASAP7_75t_L g323 ( .A(n_132), .B(n_172), .Y(n_323) );
AO21x2_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_140), .B(n_165), .Y(n_132) );
INVx3_ASAP7_75t_L g186 ( .A(n_133), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_133), .B(n_200), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_133), .B(n_229), .Y(n_228) );
NOR2xp33_ASAP7_75t_SL g522 ( .A(n_133), .B(n_523), .Y(n_522) );
INVx4_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
HB1xp67_ASAP7_75t_L g173 ( .A(n_134), .Y(n_173) );
OA21x2_ASAP7_75t_L g473 ( .A1(n_134), .A2(n_474), .B(n_481), .Y(n_473) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx1_ASAP7_75t_L g272 ( .A(n_135), .Y(n_272) );
AND2x2_ASAP7_75t_L g135 ( .A(n_136), .B(n_137), .Y(n_135) );
AND2x2_ASAP7_75t_SL g168 ( .A(n_136), .B(n_137), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_138), .B(n_139), .Y(n_137) );
OAI21xp5_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_142), .B(n_149), .Y(n_140) );
O2A1O1Ixp33_ASAP7_75t_L g188 ( .A1(n_142), .A2(n_168), .B(n_189), .C(n_190), .Y(n_188) );
OAI21xp5_ASAP7_75t_L g222 ( .A1(n_142), .A2(n_223), .B(n_224), .Y(n_222) );
OAI22xp33_ASAP7_75t_L g493 ( .A1(n_142), .A2(n_164), .B1(n_494), .B2(n_498), .Y(n_493) );
OAI21xp5_ASAP7_75t_L g503 ( .A1(n_142), .A2(n_504), .B(n_505), .Y(n_503) );
OAI21xp5_ASAP7_75t_L g525 ( .A1(n_142), .A2(n_526), .B(n_527), .Y(n_525) );
NAND2x1p5_ASAP7_75t_L g142 ( .A(n_143), .B(n_147), .Y(n_142) );
AND2x4_ASAP7_75t_L g175 ( .A(n_143), .B(n_147), .Y(n_175) );
AND2x2_ASAP7_75t_L g143 ( .A(n_144), .B(n_146), .Y(n_143) );
INVx1_ASAP7_75t_L g197 ( .A(n_144), .Y(n_197) );
INVx1_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx2_ASAP7_75t_L g151 ( .A(n_145), .Y(n_151) );
INVx1_ASAP7_75t_L g215 ( .A(n_145), .Y(n_215) );
INVx1_ASAP7_75t_L g152 ( .A(n_146), .Y(n_152) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_146), .Y(n_157) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_146), .Y(n_159) );
INVx3_ASAP7_75t_L g194 ( .A(n_146), .Y(n_194) );
INVx1_ASAP7_75t_L g478 ( .A(n_146), .Y(n_478) );
INVx4_ASAP7_75t_SL g164 ( .A(n_147), .Y(n_164) );
BUFx3_ASAP7_75t_L g198 ( .A(n_147), .Y(n_198) );
INVx5_ASAP7_75t_L g178 ( .A(n_150), .Y(n_178) );
AND2x6_ASAP7_75t_L g150 ( .A(n_151), .B(n_152), .Y(n_150) );
BUFx3_ASAP7_75t_L g162 ( .A(n_151), .Y(n_162) );
BUFx6f_ASAP7_75t_L g184 ( .A(n_151), .Y(n_184) );
O2A1O1Ixp33_ASAP7_75t_L g153 ( .A1(n_154), .A2(n_155), .B(n_158), .C(n_160), .Y(n_153) );
O2A1O1Ixp5_ASAP7_75t_L g225 ( .A1(n_155), .A2(n_160), .B(n_226), .C(n_227), .Y(n_225) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
OAI22xp5_ASAP7_75t_SL g495 ( .A1(n_156), .A2(n_157), .B1(n_496), .B2(n_497), .Y(n_495) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx4_ASAP7_75t_L g213 ( .A(n_157), .Y(n_213) );
INVx4_ASAP7_75t_L g180 ( .A(n_159), .Y(n_180) );
INVx2_ASAP7_75t_L g248 ( .A(n_159), .Y(n_248) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_160), .A2(n_520), .B(n_521), .Y(n_519) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_160), .A2(n_529), .B(n_530), .Y(n_528) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx1_ASAP7_75t_L g237 ( .A(n_162), .Y(n_237) );
INVx1_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
O2A1O1Ixp33_ASAP7_75t_L g176 ( .A1(n_164), .A2(n_177), .B(n_178), .C(n_179), .Y(n_176) );
O2A1O1Ixp33_ASAP7_75t_SL g208 ( .A1(n_164), .A2(n_178), .B(n_209), .C(n_210), .Y(n_208) );
O2A1O1Ixp33_ASAP7_75t_SL g232 ( .A1(n_164), .A2(n_178), .B(n_233), .C(n_234), .Y(n_232) );
O2A1O1Ixp33_ASAP7_75t_SL g245 ( .A1(n_164), .A2(n_178), .B(n_246), .C(n_247), .Y(n_245) );
O2A1O1Ixp33_ASAP7_75t_SL g275 ( .A1(n_164), .A2(n_178), .B(n_276), .C(n_277), .Y(n_275) );
O2A1O1Ixp33_ASAP7_75t_L g475 ( .A1(n_164), .A2(n_178), .B(n_476), .C(n_477), .Y(n_475) );
O2A1O1Ixp33_ASAP7_75t_L g485 ( .A1(n_164), .A2(n_178), .B(n_486), .C(n_487), .Y(n_485) );
O2A1O1Ixp33_ASAP7_75t_L g548 ( .A1(n_164), .A2(n_178), .B(n_549), .C(n_550), .Y(n_548) );
NOR2xp33_ASAP7_75t_L g165 ( .A(n_166), .B(n_167), .Y(n_165) );
INVx1_ASAP7_75t_L g282 ( .A(n_167), .Y(n_282) );
AO21x2_ASAP7_75t_L g535 ( .A1(n_167), .A2(n_536), .B(n_543), .Y(n_535) );
INVx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx1_ASAP7_75t_L g221 ( .A(n_168), .Y(n_221) );
OA21x2_ASAP7_75t_L g243 ( .A1(n_168), .A2(n_244), .B(n_251), .Y(n_243) );
OA21x2_ASAP7_75t_L g546 ( .A1(n_168), .A2(n_547), .B(n_553), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_169), .B(n_353), .Y(n_352) );
INVx3_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g286 ( .A(n_170), .B(n_287), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_170), .B(n_267), .Y(n_313) );
AND2x2_ASAP7_75t_L g406 ( .A(n_170), .B(n_346), .Y(n_406) );
OAI321xp33_ASAP7_75t_L g440 ( .A1(n_170), .A2(n_256), .A3(n_413), .B1(n_441), .B2(n_443), .C(n_444), .Y(n_440) );
NAND4xp25_ASAP7_75t_L g444 ( .A(n_170), .B(n_242), .C(n_353), .D(n_445), .Y(n_444) );
AND2x4_ASAP7_75t_L g170 ( .A(n_171), .B(n_187), .Y(n_170) );
AND2x2_ASAP7_75t_L g308 ( .A(n_171), .B(n_254), .Y(n_308) );
AND2x2_ASAP7_75t_L g327 ( .A(n_171), .B(n_256), .Y(n_327) );
INVx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
AND2x2_ASAP7_75t_L g255 ( .A(n_172), .B(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g283 ( .A(n_172), .B(n_187), .Y(n_283) );
AND2x2_ASAP7_75t_L g369 ( .A(n_172), .B(n_254), .Y(n_369) );
OA21x2_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_174), .B(n_185), .Y(n_172) );
OA21x2_ASAP7_75t_L g206 ( .A1(n_173), .A2(n_207), .B(n_216), .Y(n_206) );
OA21x2_ASAP7_75t_L g230 ( .A1(n_173), .A2(n_231), .B(n_238), .Y(n_230) );
BUFx2_ASAP7_75t_L g274 ( .A(n_175), .Y(n_274) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_180), .B(n_182), .Y(n_181) );
INVx3_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
HB1xp67_ASAP7_75t_L g541 ( .A(n_184), .Y(n_541) );
OA21x2_ASAP7_75t_L g483 ( .A1(n_186), .A2(n_484), .B(n_490), .Y(n_483) );
INVx3_ASAP7_75t_SL g254 ( .A(n_187), .Y(n_254) );
AND2x2_ASAP7_75t_L g301 ( .A(n_187), .B(n_288), .Y(n_301) );
OR2x2_ASAP7_75t_L g334 ( .A(n_187), .B(n_256), .Y(n_334) );
HB1xp67_ASAP7_75t_L g341 ( .A(n_187), .Y(n_341) );
AND2x2_ASAP7_75t_L g370 ( .A(n_187), .B(n_255), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_187), .B(n_343), .Y(n_385) );
AND2x2_ASAP7_75t_L g417 ( .A(n_187), .B(n_409), .Y(n_417) );
AND2x2_ASAP7_75t_L g426 ( .A(n_187), .B(n_268), .Y(n_426) );
OR2x6_ASAP7_75t_L g187 ( .A(n_188), .B(n_199), .Y(n_187) );
O2A1O1Ixp33_ASAP7_75t_L g191 ( .A1(n_192), .A2(n_193), .B(n_195), .C(n_196), .Y(n_191) );
OAI22xp33_ASAP7_75t_L g278 ( .A1(n_193), .A2(n_213), .B1(n_279), .B2(n_280), .Y(n_278) );
O2A1O1Ixp33_ASAP7_75t_L g506 ( .A1(n_193), .A2(n_507), .B(n_508), .C(n_509), .Y(n_506) );
INVx5_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g249 ( .A(n_194), .B(n_250), .Y(n_249) );
NOR2xp33_ASAP7_75t_L g479 ( .A(n_194), .B(n_480), .Y(n_479) );
NOR2xp33_ASAP7_75t_L g488 ( .A(n_194), .B(n_489), .Y(n_488) );
INVx2_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g277 ( .A(n_197), .B(n_278), .Y(n_277) );
INVx1_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_203), .B(n_217), .Y(n_202) );
INVx1_ASAP7_75t_SL g394 ( .A(n_203), .Y(n_394) );
INVx2_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
AND2x2_ASAP7_75t_L g259 ( .A(n_204), .B(n_260), .Y(n_259) );
INVx2_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
AND2x2_ASAP7_75t_L g241 ( .A(n_205), .B(n_219), .Y(n_241) );
AND2x2_ASAP7_75t_L g330 ( .A(n_205), .B(n_243), .Y(n_330) );
INVx2_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
AND2x2_ASAP7_75t_L g300 ( .A(n_206), .B(n_230), .Y(n_300) );
OR2x2_ASAP7_75t_L g311 ( .A(n_206), .B(n_243), .Y(n_311) );
AND2x2_ASAP7_75t_L g337 ( .A(n_206), .B(n_243), .Y(n_337) );
HB1xp67_ASAP7_75t_L g382 ( .A(n_206), .Y(n_382) );
NOR2xp33_ASAP7_75t_L g211 ( .A(n_212), .B(n_213), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_213), .B(n_236), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g551 ( .A(n_213), .B(n_552), .Y(n_551) );
INVx2_ASAP7_75t_L g509 ( .A(n_214), .Y(n_509) );
INVx3_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_217), .B(n_337), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_217), .B(n_394), .Y(n_393) );
INVx2_ASAP7_75t_SL g217 ( .A(n_218), .Y(n_217) );
OR2x2_ASAP7_75t_L g310 ( .A(n_218), .B(n_311), .Y(n_310) );
AOI322xp5_ASAP7_75t_L g396 ( .A1(n_218), .A2(n_300), .A3(n_306), .B1(n_337), .B2(n_387), .C1(n_397), .C2(n_399), .Y(n_396) );
OR2x2_ASAP7_75t_L g218 ( .A(n_219), .B(n_230), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_219), .B(n_242), .Y(n_262) );
NOR2xp33_ASAP7_75t_L g293 ( .A(n_219), .B(n_243), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_219), .B(n_260), .Y(n_317) );
AND2x2_ASAP7_75t_L g371 ( .A(n_219), .B(n_337), .Y(n_371) );
INVx1_ASAP7_75t_L g375 ( .A(n_219), .Y(n_375) );
AND2x2_ASAP7_75t_L g387 ( .A(n_219), .B(n_230), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_219), .B(n_259), .Y(n_419) );
INVx4_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
AND2x2_ASAP7_75t_L g284 ( .A(n_220), .B(n_230), .Y(n_284) );
BUFx3_ASAP7_75t_L g298 ( .A(n_220), .Y(n_298) );
AND3x2_ASAP7_75t_L g380 ( .A(n_220), .B(n_360), .C(n_381), .Y(n_380) );
AO21x2_ASAP7_75t_L g220 ( .A1(n_221), .A2(n_222), .B(n_228), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_221), .B(n_511), .Y(n_510) );
NOR2xp33_ASAP7_75t_L g531 ( .A(n_221), .B(n_532), .Y(n_531) );
NOR2xp33_ASAP7_75t_L g543 ( .A(n_221), .B(n_544), .Y(n_543) );
NAND3xp33_ASAP7_75t_L g240 ( .A(n_230), .B(n_241), .C(n_242), .Y(n_240) );
INVx1_ASAP7_75t_SL g260 ( .A(n_230), .Y(n_260) );
HB1xp67_ASAP7_75t_L g365 ( .A(n_230), .Y(n_365) );
INVx1_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
AND2x2_ASAP7_75t_L g359 ( .A(n_241), .B(n_360), .Y(n_359) );
INVxp67_ASAP7_75t_L g366 ( .A(n_241), .Y(n_366) );
AND2x2_ASAP7_75t_L g404 ( .A(n_242), .B(n_382), .Y(n_404) );
INVx2_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
BUFx3_ASAP7_75t_L g285 ( .A(n_243), .Y(n_285) );
AND2x2_ASAP7_75t_L g360 ( .A(n_243), .B(n_260), .Y(n_360) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
OR2x2_ASAP7_75t_L g304 ( .A(n_254), .B(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g423 ( .A(n_254), .B(n_323), .Y(n_423) );
AND2x2_ASAP7_75t_L g437 ( .A(n_254), .B(n_256), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_255), .B(n_268), .Y(n_378) );
AND2x2_ASAP7_75t_L g425 ( .A(n_255), .B(n_426), .Y(n_425) );
AND2x2_ASAP7_75t_L g288 ( .A(n_256), .B(n_289), .Y(n_288) );
OR2x2_ASAP7_75t_L g305 ( .A(n_256), .B(n_268), .Y(n_305) );
INVx1_ASAP7_75t_L g315 ( .A(n_256), .Y(n_315) );
AND2x2_ASAP7_75t_L g346 ( .A(n_256), .B(n_268), .Y(n_346) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
OAI221xp5_ASAP7_75t_L g388 ( .A1(n_258), .A2(n_389), .B1(n_393), .B2(n_395), .C(n_396), .Y(n_388) );
NAND2xp5_ASAP7_75t_SL g258 ( .A(n_259), .B(n_261), .Y(n_258) );
AND2x2_ASAP7_75t_L g292 ( .A(n_259), .B(n_293), .Y(n_292) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
NOR2xp33_ASAP7_75t_L g442 ( .A(n_262), .B(n_299), .Y(n_442) );
AOI322xp5_ASAP7_75t_L g264 ( .A1(n_265), .A2(n_284), .A3(n_285), .B1(n_286), .B2(n_292), .C1(n_294), .C2(n_301), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_267), .B(n_283), .Y(n_266) );
NAND2x1p5_ASAP7_75t_L g322 ( .A(n_267), .B(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_267), .B(n_333), .Y(n_332) );
O2A1O1Ixp33_ASAP7_75t_L g356 ( .A1(n_267), .A2(n_283), .B(n_357), .C(n_358), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_267), .B(n_369), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_267), .B(n_327), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_267), .B(n_409), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_267), .B(n_437), .Y(n_436) );
BUFx3_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_268), .B(n_308), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_268), .B(n_315), .Y(n_314) );
OR2x2_ASAP7_75t_L g398 ( .A(n_268), .B(n_285), .Y(n_398) );
OA21x2_ASAP7_75t_L g268 ( .A1(n_269), .A2(n_273), .B(n_281), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
AO21x2_ASAP7_75t_L g289 ( .A1(n_270), .A2(n_290), .B(n_291), .Y(n_289) );
AO21x2_ASAP7_75t_L g524 ( .A1(n_270), .A2(n_525), .B(n_531), .Y(n_524) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
AOI21xp5_ASAP7_75t_SL g516 ( .A1(n_271), .A2(n_517), .B(n_518), .Y(n_516) );
INVx2_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AO21x2_ASAP7_75t_L g492 ( .A1(n_272), .A2(n_493), .B(n_499), .Y(n_492) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_272), .B(n_500), .Y(n_499) );
AO21x2_ASAP7_75t_L g502 ( .A1(n_272), .A2(n_503), .B(n_510), .Y(n_502) );
INVx1_ASAP7_75t_L g290 ( .A(n_273), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_281), .Y(n_291) );
INVx1_ASAP7_75t_L g373 ( .A(n_283), .Y(n_373) );
OAI31xp33_ASAP7_75t_L g383 ( .A1(n_283), .A2(n_308), .A3(n_384), .B(n_386), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_283), .B(n_289), .Y(n_435) );
INVx1_ASAP7_75t_SL g296 ( .A(n_284), .Y(n_296) );
AND2x2_ASAP7_75t_L g329 ( .A(n_284), .B(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g410 ( .A(n_284), .B(n_411), .Y(n_410) );
OR2x2_ASAP7_75t_L g295 ( .A(n_285), .B(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g320 ( .A(n_285), .Y(n_320) );
AND2x2_ASAP7_75t_L g347 ( .A(n_285), .B(n_300), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_285), .B(n_365), .Y(n_364) );
AND2x2_ASAP7_75t_L g439 ( .A(n_285), .B(n_387), .Y(n_439) );
NOR2xp33_ASAP7_75t_L g430 ( .A(n_287), .B(n_357), .Y(n_430) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g326 ( .A(n_289), .B(n_327), .Y(n_326) );
INVx1_ASAP7_75t_SL g344 ( .A(n_289), .Y(n_344) );
NAND2xp33_ASAP7_75t_SL g294 ( .A(n_295), .B(n_297), .Y(n_294) );
OAI211xp5_ASAP7_75t_SL g338 ( .A1(n_296), .A2(n_339), .B(n_345), .C(n_361), .Y(n_338) );
OR2x2_ASAP7_75t_L g413 ( .A(n_296), .B(n_394), .Y(n_413) );
OR2x2_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
CKINVDCx16_ASAP7_75t_R g350 ( .A(n_298), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_298), .B(n_404), .Y(n_403) );
INVx1_ASAP7_75t_SL g299 ( .A(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g319 ( .A(n_300), .B(n_320), .Y(n_319) );
O2A1O1Ixp33_ASAP7_75t_L g302 ( .A1(n_303), .A2(n_306), .B(n_309), .C(n_312), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx1_ASAP7_75t_SL g353 ( .A(n_305), .Y(n_353) );
INVx1_ASAP7_75t_SL g306 ( .A(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_308), .B(n_346), .Y(n_351) );
INVx1_ASAP7_75t_L g357 ( .A(n_308), .Y(n_357) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
OR2x2_ASAP7_75t_L g316 ( .A(n_311), .B(n_317), .Y(n_316) );
OR2x2_ASAP7_75t_L g349 ( .A(n_311), .B(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g411 ( .A(n_311), .Y(n_411) );
AOI21xp33_ASAP7_75t_SL g312 ( .A1(n_313), .A2(n_314), .B(n_316), .Y(n_312) );
AOI21xp5_ASAP7_75t_L g324 ( .A1(n_314), .A2(n_325), .B(n_328), .Y(n_324) );
AOI211xp5_ASAP7_75t_L g318 ( .A1(n_319), .A2(n_321), .B(n_324), .C(n_331), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_319), .B(n_375), .Y(n_374) );
INVx1_ASAP7_75t_SL g321 ( .A(n_322), .Y(n_321) );
NOR2xp33_ASAP7_75t_L g412 ( .A(n_322), .B(n_413), .Y(n_412) );
INVx2_ASAP7_75t_SL g335 ( .A(n_323), .Y(n_335) );
OAI21xp5_ASAP7_75t_L g390 ( .A1(n_325), .A2(n_391), .B(n_392), .Y(n_390) );
INVx1_ASAP7_75t_SL g325 ( .A(n_326), .Y(n_325) );
INVx1_ASAP7_75t_SL g328 ( .A(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_330), .B(n_343), .Y(n_342) );
INVx1_ASAP7_75t_SL g355 ( .A(n_330), .Y(n_355) );
AOI21xp33_ASAP7_75t_SL g331 ( .A1(n_332), .A2(n_335), .B(n_336), .Y(n_331) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
AND2x2_ASAP7_75t_L g386 ( .A(n_337), .B(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
NOR2xp33_ASAP7_75t_L g340 ( .A(n_341), .B(n_342), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_343), .B(n_369), .Y(n_395) );
AND2x2_ASAP7_75t_L g408 ( .A(n_343), .B(n_409), .Y(n_408) );
AND2x2_ASAP7_75t_L g422 ( .A(n_343), .B(n_423), .Y(n_422) );
AND2x2_ASAP7_75t_L g432 ( .A(n_343), .B(n_370), .Y(n_432) );
INVx2_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
AOI211xp5_ASAP7_75t_L g345 ( .A1(n_346), .A2(n_347), .B(n_348), .C(n_356), .Y(n_345) );
INVx1_ASAP7_75t_L g392 ( .A(n_346), .Y(n_392) );
OAI22xp33_ASAP7_75t_L g348 ( .A1(n_349), .A2(n_351), .B1(n_352), .B2(n_354), .Y(n_348) );
OR2x2_ASAP7_75t_L g354 ( .A(n_350), .B(n_355), .Y(n_354) );
NAND2xp5_ASAP7_75t_SL g433 ( .A(n_350), .B(n_411), .Y(n_433) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g427 ( .A(n_360), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g361 ( .A1(n_362), .A2(n_367), .B1(n_370), .B2(n_371), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
OR2x2_ASAP7_75t_L g363 ( .A(n_364), .B(n_366), .Y(n_363) );
INVx1_ASAP7_75t_L g445 ( .A(n_365), .Y(n_445) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g391 ( .A(n_369), .Y(n_391) );
OAI211xp5_ASAP7_75t_SL g372 ( .A1(n_373), .A2(n_374), .B(n_376), .C(n_383), .Y(n_372) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
NOR2xp33_ASAP7_75t_L g377 ( .A(n_378), .B(n_379), .Y(n_377) );
INVx2_ASAP7_75t_SL g379 ( .A(n_380), .Y(n_379) );
INVxp67_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVxp67_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
NOR2xp33_ASAP7_75t_L g397 ( .A(n_391), .B(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
NOR5xp2_ASAP7_75t_L g401 ( .A(n_402), .B(n_420), .C(n_428), .D(n_434), .E(n_440), .Y(n_401) );
OAI211xp5_ASAP7_75t_SL g402 ( .A1(n_403), .A2(n_405), .B(n_407), .C(n_414), .Y(n_402) );
INVxp67_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
AOI21xp5_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_410), .B(n_412), .Y(n_407) );
OAI21xp33_ASAP7_75t_L g414 ( .A1(n_415), .A2(n_417), .B(n_418), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
NOR2xp33_ASAP7_75t_L g429 ( .A(n_417), .B(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
AOI21xp33_ASAP7_75t_L g420 ( .A1(n_421), .A2(n_424), .B(n_427), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_SL g443 ( .A(n_423), .Y(n_443) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
AOI21xp5_ASAP7_75t_L g428 ( .A1(n_429), .A2(n_431), .B(n_433), .Y(n_428) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
HB1xp67_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx2_ASAP7_75t_L g457 ( .A(n_452), .Y(n_457) );
NOR2x2_ASAP7_75t_L g758 ( .A(n_453), .B(n_464), .Y(n_758) );
INVx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
OR2x2_ASAP7_75t_L g463 ( .A(n_454), .B(n_464), .Y(n_463) );
AOI21xp33_ASAP7_75t_L g458 ( .A1(n_456), .A2(n_459), .B(n_762), .Y(n_458) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
AOI22xp5_ASAP7_75t_L g461 ( .A1(n_462), .A2(n_465), .B1(n_746), .B2(n_748), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx2_ASAP7_75t_L g761 ( .A(n_465), .Y(n_761) );
INVx3_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
AND4x1_ASAP7_75t_L g466 ( .A(n_467), .B(n_664), .C(n_711), .D(n_731), .Y(n_466) );
NOR3xp33_ASAP7_75t_SL g467 ( .A(n_468), .B(n_594), .C(n_619), .Y(n_467) );
OAI211xp5_ASAP7_75t_SL g468 ( .A1(n_469), .A2(n_512), .B(n_554), .C(n_584), .Y(n_468) );
INVxp67_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
NOR2xp33_ASAP7_75t_L g470 ( .A(n_471), .B(n_491), .Y(n_470) );
INVx3_ASAP7_75t_SL g636 ( .A(n_471), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_471), .B(n_567), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_471), .B(n_501), .Y(n_717) );
AND2x2_ASAP7_75t_L g740 ( .A(n_471), .B(n_606), .Y(n_740) );
AND2x4_ASAP7_75t_L g471 ( .A(n_472), .B(n_482), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
AND2x2_ASAP7_75t_L g558 ( .A(n_473), .B(n_483), .Y(n_558) );
INVx3_ASAP7_75t_L g571 ( .A(n_473), .Y(n_571) );
AND2x2_ASAP7_75t_L g576 ( .A(n_473), .B(n_482), .Y(n_576) );
OR2x2_ASAP7_75t_L g627 ( .A(n_473), .B(n_568), .Y(n_627) );
BUFx2_ASAP7_75t_L g647 ( .A(n_473), .Y(n_647) );
AND2x2_ASAP7_75t_L g657 ( .A(n_473), .B(n_568), .Y(n_657) );
AND2x2_ASAP7_75t_L g663 ( .A(n_473), .B(n_492), .Y(n_663) );
INVx1_ASAP7_75t_SL g482 ( .A(n_483), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_483), .B(n_568), .Y(n_582) );
INVx2_ASAP7_75t_L g592 ( .A(n_483), .Y(n_592) );
AND2x2_ASAP7_75t_L g605 ( .A(n_483), .B(n_571), .Y(n_605) );
OR2x2_ASAP7_75t_L g616 ( .A(n_483), .B(n_568), .Y(n_616) );
AND2x2_ASAP7_75t_SL g662 ( .A(n_483), .B(n_663), .Y(n_662) );
BUFx2_ASAP7_75t_L g674 ( .A(n_483), .Y(n_674) );
AND2x2_ASAP7_75t_L g720 ( .A(n_483), .B(n_492), .Y(n_720) );
INVx3_ASAP7_75t_SL g593 ( .A(n_491), .Y(n_593) );
OR2x2_ASAP7_75t_L g646 ( .A(n_491), .B(n_647), .Y(n_646) );
OR2x2_ASAP7_75t_L g491 ( .A(n_492), .B(n_501), .Y(n_491) );
INVx3_ASAP7_75t_L g568 ( .A(n_492), .Y(n_568) );
AND2x2_ASAP7_75t_L g635 ( .A(n_492), .B(n_502), .Y(n_635) );
HB1xp67_ASAP7_75t_L g703 ( .A(n_492), .Y(n_703) );
AOI33xp33_ASAP7_75t_L g707 ( .A1(n_492), .A2(n_636), .A3(n_643), .B1(n_652), .B2(n_708), .B3(n_709), .Y(n_707) );
INVx1_ASAP7_75t_L g556 ( .A(n_501), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_501), .B(n_571), .Y(n_570) );
NOR3xp33_ASAP7_75t_L g630 ( .A(n_501), .B(n_631), .C(n_633), .Y(n_630) );
AND2x2_ASAP7_75t_L g656 ( .A(n_501), .B(n_657), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_501), .B(n_663), .Y(n_666) );
AND2x2_ASAP7_75t_L g719 ( .A(n_501), .B(n_720), .Y(n_719) );
INVx3_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx3_ASAP7_75t_L g575 ( .A(n_502), .Y(n_575) );
OR2x2_ASAP7_75t_L g669 ( .A(n_502), .B(n_568), .Y(n_669) );
OR2x2_ASAP7_75t_L g512 ( .A(n_513), .B(n_533), .Y(n_512) );
AOI32xp33_ASAP7_75t_L g620 ( .A1(n_513), .A2(n_621), .A3(n_623), .B1(n_625), .B2(n_628), .Y(n_620) );
NOR2xp67_ASAP7_75t_L g693 ( .A(n_513), .B(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g723 ( .A(n_513), .Y(n_723) );
INVx4_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
AND2x2_ASAP7_75t_L g655 ( .A(n_514), .B(n_639), .Y(n_655) );
AND2x2_ASAP7_75t_L g675 ( .A(n_514), .B(n_601), .Y(n_675) );
AND2x2_ASAP7_75t_L g743 ( .A(n_514), .B(n_661), .Y(n_743) );
AND2x2_ASAP7_75t_L g514 ( .A(n_515), .B(n_524), .Y(n_514) );
INVx3_ASAP7_75t_L g564 ( .A(n_515), .Y(n_564) );
AND2x2_ASAP7_75t_L g578 ( .A(n_515), .B(n_562), .Y(n_578) );
OR2x2_ASAP7_75t_L g583 ( .A(n_515), .B(n_561), .Y(n_583) );
INVx1_ASAP7_75t_L g590 ( .A(n_515), .Y(n_590) );
AND2x2_ASAP7_75t_L g598 ( .A(n_515), .B(n_572), .Y(n_598) );
AND2x2_ASAP7_75t_L g600 ( .A(n_515), .B(n_601), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_515), .B(n_639), .Y(n_638) );
INVx2_ASAP7_75t_L g653 ( .A(n_515), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_515), .B(n_738), .Y(n_737) );
OR2x6_ASAP7_75t_L g515 ( .A(n_516), .B(n_522), .Y(n_515) );
INVx2_ASAP7_75t_L g562 ( .A(n_524), .Y(n_562) );
AND2x2_ASAP7_75t_L g608 ( .A(n_524), .B(n_534), .Y(n_608) );
AND2x2_ASAP7_75t_L g618 ( .A(n_524), .B(n_546), .Y(n_618) );
INVx2_ASAP7_75t_L g738 ( .A(n_533), .Y(n_738) );
OR2x2_ASAP7_75t_L g533 ( .A(n_534), .B(n_545), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_534), .B(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g579 ( .A(n_534), .Y(n_579) );
AND2x2_ASAP7_75t_L g623 ( .A(n_534), .B(n_624), .Y(n_623) );
AND2x2_ASAP7_75t_L g639 ( .A(n_534), .B(n_602), .Y(n_639) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g587 ( .A(n_535), .Y(n_587) );
AND2x2_ASAP7_75t_L g601 ( .A(n_535), .B(n_602), .Y(n_601) );
AND2x2_ASAP7_75t_L g652 ( .A(n_535), .B(n_653), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_535), .B(n_562), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_537), .B(n_542), .Y(n_536) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_539), .A2(n_540), .B(n_541), .Y(n_538) );
AND2x2_ASAP7_75t_L g563 ( .A(n_545), .B(n_564), .Y(n_563) );
INVx2_ASAP7_75t_L g624 ( .A(n_545), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_545), .B(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g661 ( .A(n_545), .Y(n_661) );
INVx1_ASAP7_75t_L g694 ( .A(n_545), .Y(n_694) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
AND2x2_ASAP7_75t_L g572 ( .A(n_546), .B(n_562), .Y(n_572) );
INVx1_ASAP7_75t_L g602 ( .A(n_546), .Y(n_602) );
AOI221xp5_ASAP7_75t_L g554 ( .A1(n_555), .A2(n_559), .B1(n_565), .B2(n_572), .C(n_573), .Y(n_554) );
NOR2xp33_ASAP7_75t_L g555 ( .A(n_556), .B(n_557), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_556), .B(n_576), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_556), .B(n_639), .Y(n_716) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_558), .B(n_606), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_558), .B(n_567), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_558), .B(n_581), .Y(n_710) );
AND2x2_ASAP7_75t_L g559 ( .A(n_560), .B(n_563), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx2_ASAP7_75t_L g632 ( .A(n_562), .Y(n_632) );
AND2x2_ASAP7_75t_L g607 ( .A(n_563), .B(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g685 ( .A(n_563), .Y(n_685) );
AND2x2_ASAP7_75t_L g617 ( .A(n_564), .B(n_618), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_564), .B(n_587), .Y(n_633) );
AND2x2_ASAP7_75t_L g697 ( .A(n_564), .B(n_623), .Y(n_697) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_567), .B(n_569), .Y(n_566) );
BUFx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g606 ( .A(n_568), .B(n_575), .Y(n_606) );
AND2x2_ASAP7_75t_L g702 ( .A(n_569), .B(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_571), .B(n_615), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_572), .B(n_590), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_572), .B(n_579), .Y(n_667) );
AND2x2_ASAP7_75t_L g687 ( .A(n_572), .B(n_587), .Y(n_687) );
AND2x2_ASAP7_75t_L g708 ( .A(n_572), .B(n_652), .Y(n_708) );
OAI32xp33_ASAP7_75t_L g573 ( .A1(n_574), .A2(n_577), .A3(n_579), .B1(n_580), .B2(n_583), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_575), .B(n_576), .Y(n_574) );
INVx1_ASAP7_75t_SL g581 ( .A(n_575), .Y(n_581) );
NAND2x1_ASAP7_75t_L g622 ( .A(n_575), .B(n_605), .Y(n_622) );
OR2x2_ASAP7_75t_L g626 ( .A(n_575), .B(n_627), .Y(n_626) );
NOR2xp33_ASAP7_75t_L g727 ( .A(n_575), .B(n_674), .Y(n_727) );
INVx1_ASAP7_75t_L g595 ( .A(n_576), .Y(n_595) );
OAI221xp5_ASAP7_75t_SL g713 ( .A1(n_577), .A2(n_668), .B1(n_714), .B2(n_717), .C(n_718), .Y(n_713) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_L g585 ( .A(n_578), .B(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g628 ( .A(n_578), .B(n_601), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_578), .B(n_660), .Y(n_659) );
AND2x2_ASAP7_75t_L g706 ( .A(n_578), .B(n_639), .Y(n_706) );
INVxp67_ASAP7_75t_L g642 ( .A(n_579), .Y(n_642) );
OR2x2_ASAP7_75t_L g580 ( .A(n_581), .B(n_582), .Y(n_580) );
AND2x2_ASAP7_75t_L g712 ( .A(n_581), .B(n_699), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_581), .B(n_662), .Y(n_735) );
INVx1_ASAP7_75t_L g610 ( .A(n_583), .Y(n_610) );
NAND2xp5_ASAP7_75t_SL g691 ( .A(n_583), .B(n_692), .Y(n_691) );
OR2x2_ASAP7_75t_L g728 ( .A(n_583), .B(n_729), .Y(n_728) );
OAI21xp5_ASAP7_75t_SL g584 ( .A1(n_585), .A2(n_588), .B(n_591), .Y(n_584) );
AND2x2_ASAP7_75t_L g597 ( .A(n_586), .B(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_L g681 ( .A(n_590), .B(n_601), .Y(n_681) );
AND2x2_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .Y(n_591) );
AND2x2_ASAP7_75t_L g699 ( .A(n_592), .B(n_657), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_592), .B(n_656), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_593), .B(n_605), .Y(n_679) );
OAI211xp5_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_596), .B(n_599), .C(n_609), .Y(n_594) );
AOI221xp5_ASAP7_75t_L g629 ( .A1(n_595), .A2(n_630), .B1(n_634), .B2(n_637), .C(n_640), .Y(n_629) );
AOI31xp33_ASAP7_75t_L g724 ( .A1(n_595), .A2(n_725), .A3(n_726), .B(n_728), .Y(n_724) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
AOI22xp5_ASAP7_75t_L g599 ( .A1(n_600), .A2(n_603), .B1(n_605), .B2(n_607), .Y(n_599) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_605), .B(n_606), .Y(n_604) );
INVx1_ASAP7_75t_L g725 ( .A(n_605), .Y(n_725) );
INVx1_ASAP7_75t_L g688 ( .A(n_606), .Y(n_688) );
O2A1O1Ixp33_ASAP7_75t_L g731 ( .A1(n_608), .A2(n_732), .B(n_734), .C(n_736), .Y(n_731) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_610), .A2(n_611), .B1(n_613), .B2(n_617), .Y(n_609) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_614), .B(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
OAI221xp5_ASAP7_75t_SL g704 ( .A1(n_616), .A2(n_650), .B1(n_669), .B2(n_705), .C(n_707), .Y(n_704) );
INVx1_ASAP7_75t_L g700 ( .A(n_617), .Y(n_700) );
INVx1_ASAP7_75t_L g654 ( .A(n_618), .Y(n_654) );
NAND3xp33_ASAP7_75t_SL g619 ( .A(n_620), .B(n_629), .C(n_644), .Y(n_619) );
OAI21xp33_ASAP7_75t_L g670 ( .A1(n_621), .A2(n_671), .B(n_675), .Y(n_670) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_623), .B(n_723), .Y(n_722) );
INVxp67_ASAP7_75t_L g730 ( .A(n_624), .Y(n_730) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
OR2x2_ASAP7_75t_L g668 ( .A(n_631), .B(n_651), .Y(n_668) );
INVx1_ASAP7_75t_L g643 ( .A(n_632), .Y(n_643) );
AND2x2_ASAP7_75t_L g634 ( .A(n_635), .B(n_636), .Y(n_634) );
INVx1_ASAP7_75t_L g641 ( .A(n_635), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_635), .B(n_673), .Y(n_672) );
NOR4xp25_ASAP7_75t_L g640 ( .A(n_636), .B(n_641), .C(n_642), .D(n_643), .Y(n_640) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
AOI222xp33_ASAP7_75t_L g644 ( .A1(n_645), .A2(n_649), .B1(n_655), .B2(n_656), .C1(n_658), .C2(n_662), .Y(n_644) );
NAND2xp5_ASAP7_75t_SL g645 ( .A(n_646), .B(n_648), .Y(n_645) );
INVx1_ASAP7_75t_L g742 ( .A(n_646), .Y(n_742) );
INVx1_ASAP7_75t_SL g649 ( .A(n_650), .Y(n_649) );
OR2x2_ASAP7_75t_L g650 ( .A(n_651), .B(n_654), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_658), .B(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
OAI21xp5_ASAP7_75t_SL g718 ( .A1(n_663), .A2(n_719), .B(n_721), .Y(n_718) );
NOR4xp25_ASAP7_75t_L g664 ( .A(n_665), .B(n_676), .C(n_689), .D(n_704), .Y(n_664) );
OAI221xp5_ASAP7_75t_SL g665 ( .A1(n_666), .A2(n_667), .B1(n_668), .B2(n_669), .C(n_670), .Y(n_665) );
INVx1_ASAP7_75t_L g745 ( .A(n_666), .Y(n_745) );
INVx1_ASAP7_75t_SL g671 ( .A(n_672), .Y(n_671) );
NOR2xp33_ASAP7_75t_L g715 ( .A(n_673), .B(n_716), .Y(n_715) );
INVx1_ASAP7_75t_SL g673 ( .A(n_674), .Y(n_673) );
OAI222xp33_ASAP7_75t_L g676 ( .A1(n_677), .A2(n_680), .B1(n_682), .B2(n_683), .C1(n_686), .C2(n_688), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
AOI211xp5_ASAP7_75t_L g711 ( .A1(n_681), .A2(n_712), .B(n_713), .C(n_724), .Y(n_711) );
OR2x2_ASAP7_75t_L g683 ( .A(n_684), .B(n_685), .Y(n_683) );
INVx1_ASAP7_75t_SL g686 ( .A(n_687), .Y(n_686) );
OAI222xp33_ASAP7_75t_L g689 ( .A1(n_690), .A2(n_695), .B1(n_696), .B2(n_698), .C1(n_700), .C2(n_701), .Y(n_689) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVxp67_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
AOI22xp5_ASAP7_75t_L g741 ( .A1(n_706), .A2(n_709), .B1(n_742), .B2(n_743), .Y(n_741) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
HB1xp67_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
OAI211xp5_ASAP7_75t_SL g736 ( .A1(n_737), .A2(n_739), .B(n_741), .C(n_744), .Y(n_736) );
INVx2_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
INVx1_ASAP7_75t_SL g756 ( .A(n_757), .Y(n_756) );
INVx3_ASAP7_75t_SL g757 ( .A(n_758), .Y(n_757) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
endmodule