module real_aes_8961_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_369;
wire n_343;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_656;
wire n_532;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_617;
wire n_552;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_717;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_241;
wire n_175;
wire n_168;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g110 ( .A(n_0), .B(n_111), .C(n_112), .Y(n_110) );
INVx1_ASAP7_75t_L g442 ( .A(n_0), .Y(n_442) );
A2O1A1Ixp33_ASAP7_75t_L g188 ( .A1(n_1), .A2(n_147), .B(n_152), .C(n_189), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_2), .A2(n_142), .B(n_212), .Y(n_211) );
INVx1_ASAP7_75t_L g460 ( .A(n_3), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_4), .B(n_166), .Y(n_219) );
AOI22xp5_ASAP7_75t_L g721 ( .A1(n_5), .A2(n_15), .B1(n_722), .B2(n_723), .Y(n_721) );
CKINVDCx20_ASAP7_75t_R g723 ( .A(n_5), .Y(n_723) );
AOI21xp33_ASAP7_75t_L g477 ( .A1(n_6), .A2(n_142), .B(n_478), .Y(n_477) );
AND2x6_ASAP7_75t_L g147 ( .A(n_7), .B(n_148), .Y(n_147) );
INVx1_ASAP7_75t_L g176 ( .A(n_8), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_9), .B(n_109), .Y(n_108) );
NOR2xp33_ASAP7_75t_L g443 ( .A(n_9), .B(n_43), .Y(n_443) );
AOI21xp5_ASAP7_75t_L g537 ( .A1(n_10), .A2(n_254), .B(n_538), .Y(n_537) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_11), .B(n_157), .Y(n_193) );
INVx1_ASAP7_75t_L g482 ( .A(n_12), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_13), .B(n_156), .Y(n_530) );
INVx1_ASAP7_75t_L g140 ( .A(n_14), .Y(n_140) );
CKINVDCx20_ASAP7_75t_R g722 ( .A(n_15), .Y(n_722) );
INVx1_ASAP7_75t_L g542 ( .A(n_16), .Y(n_542) );
A2O1A1Ixp33_ASAP7_75t_L g201 ( .A1(n_17), .A2(n_177), .B(n_202), .C(n_204), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_18), .B(n_166), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_19), .B(n_471), .Y(n_521) );
NAND2xp5_ASAP7_75t_SL g508 ( .A(n_20), .B(n_142), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_21), .B(n_262), .Y(n_261) );
A2O1A1Ixp33_ASAP7_75t_L g155 ( .A1(n_22), .A2(n_156), .B(n_158), .C(n_162), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_23), .B(n_166), .Y(n_474) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_24), .B(n_157), .Y(n_226) );
A2O1A1Ixp33_ASAP7_75t_L g540 ( .A1(n_25), .A2(n_160), .B(n_204), .C(n_541), .Y(n_540) );
NAND2xp5_ASAP7_75t_SL g238 ( .A(n_26), .B(n_157), .Y(n_238) );
CKINVDCx16_ASAP7_75t_R g222 ( .A(n_27), .Y(n_222) );
INVx1_ASAP7_75t_L g236 ( .A(n_28), .Y(n_236) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_29), .Y(n_146) );
CKINVDCx20_ASAP7_75t_R g186 ( .A(n_30), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_31), .B(n_157), .Y(n_461) );
INVx1_ASAP7_75t_L g259 ( .A(n_32), .Y(n_259) );
INVx1_ASAP7_75t_L g495 ( .A(n_33), .Y(n_495) );
NAND2xp5_ASAP7_75t_SL g444 ( .A(n_34), .B(n_445), .Y(n_444) );
INVx2_ASAP7_75t_L g145 ( .A(n_35), .Y(n_145) );
CKINVDCx20_ASAP7_75t_R g196 ( .A(n_36), .Y(n_196) );
A2O1A1Ixp33_ASAP7_75t_L g214 ( .A1(n_37), .A2(n_156), .B(n_215), .C(n_217), .Y(n_214) );
INVxp67_ASAP7_75t_L g260 ( .A(n_38), .Y(n_260) );
CKINVDCx14_ASAP7_75t_R g213 ( .A(n_39), .Y(n_213) );
A2O1A1Ixp33_ASAP7_75t_L g234 ( .A1(n_40), .A2(n_152), .B(n_235), .C(n_241), .Y(n_234) );
A2O1A1Ixp33_ASAP7_75t_L g509 ( .A1(n_41), .A2(n_147), .B(n_152), .C(n_510), .Y(n_509) );
OAI22xp5_ASAP7_75t_SL g124 ( .A1(n_42), .A2(n_91), .B1(n_125), .B2(n_126), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_42), .Y(n_126) );
INVx1_ASAP7_75t_L g109 ( .A(n_43), .Y(n_109) );
INVx1_ASAP7_75t_L g494 ( .A(n_44), .Y(n_494) );
A2O1A1Ixp33_ASAP7_75t_L g173 ( .A1(n_45), .A2(n_174), .B(n_175), .C(n_178), .Y(n_173) );
NAND2xp5_ASAP7_75t_SL g520 ( .A(n_46), .B(n_157), .Y(n_520) );
AOI22xp33_ASAP7_75t_L g122 ( .A1(n_47), .A2(n_123), .B1(n_435), .B2(n_436), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g435 ( .A(n_47), .Y(n_435) );
CKINVDCx20_ASAP7_75t_R g243 ( .A(n_48), .Y(n_243) );
CKINVDCx20_ASAP7_75t_R g256 ( .A(n_49), .Y(n_256) );
INVx1_ASAP7_75t_L g150 ( .A(n_50), .Y(n_150) );
CKINVDCx16_ASAP7_75t_R g496 ( .A(n_51), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_52), .B(n_142), .Y(n_532) );
AOI22xp5_ASAP7_75t_L g492 ( .A1(n_53), .A2(n_152), .B1(n_162), .B2(n_493), .Y(n_492) );
CKINVDCx20_ASAP7_75t_R g514 ( .A(n_54), .Y(n_514) );
CKINVDCx16_ASAP7_75t_R g457 ( .A(n_55), .Y(n_457) );
CKINVDCx14_ASAP7_75t_R g172 ( .A(n_56), .Y(n_172) );
A2O1A1Ixp33_ASAP7_75t_L g480 ( .A1(n_57), .A2(n_174), .B(n_217), .C(n_481), .Y(n_480) );
CKINVDCx20_ASAP7_75t_R g523 ( .A(n_58), .Y(n_523) );
INVx1_ASAP7_75t_L g479 ( .A(n_59), .Y(n_479) );
INVx1_ASAP7_75t_L g148 ( .A(n_60), .Y(n_148) );
INVx1_ASAP7_75t_L g139 ( .A(n_61), .Y(n_139) );
INVx1_ASAP7_75t_SL g216 ( .A(n_62), .Y(n_216) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_63), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_64), .B(n_166), .Y(n_165) );
INVx1_ASAP7_75t_L g225 ( .A(n_65), .Y(n_225) );
A2O1A1Ixp33_ASAP7_75t_SL g470 ( .A1(n_66), .A2(n_217), .B(n_471), .C(n_472), .Y(n_470) );
INVxp67_ASAP7_75t_L g473 ( .A(n_67), .Y(n_473) );
INVx1_ASAP7_75t_L g114 ( .A(n_68), .Y(n_114) );
AOI21xp5_ASAP7_75t_L g170 ( .A1(n_69), .A2(n_142), .B(n_171), .Y(n_170) );
CKINVDCx20_ASAP7_75t_R g229 ( .A(n_70), .Y(n_229) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_71), .A2(n_142), .B(n_199), .Y(n_198) );
CKINVDCx20_ASAP7_75t_R g498 ( .A(n_72), .Y(n_498) );
INVx1_ASAP7_75t_L g517 ( .A(n_73), .Y(n_517) );
AOI21xp5_ASAP7_75t_L g253 ( .A1(n_74), .A2(n_254), .B(n_255), .Y(n_253) );
INVx1_ASAP7_75t_L g200 ( .A(n_75), .Y(n_200) );
CKINVDCx16_ASAP7_75t_R g233 ( .A(n_76), .Y(n_233) );
AOI222xp33_ASAP7_75t_L g447 ( .A1(n_77), .A2(n_448), .B1(n_719), .B2(n_725), .C1(n_729), .C2(n_730), .Y(n_447) );
A2O1A1Ixp33_ASAP7_75t_L g518 ( .A1(n_78), .A2(n_147), .B(n_152), .C(n_519), .Y(n_518) );
AOI21xp5_ASAP7_75t_L g141 ( .A1(n_79), .A2(n_142), .B(n_149), .Y(n_141) );
INVx1_ASAP7_75t_L g203 ( .A(n_80), .Y(n_203) );
NAND2xp5_ASAP7_75t_SL g511 ( .A(n_81), .B(n_237), .Y(n_511) );
INVx2_ASAP7_75t_L g137 ( .A(n_82), .Y(n_137) );
INVx1_ASAP7_75t_L g190 ( .A(n_83), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_84), .B(n_471), .Y(n_512) );
A2O1A1Ixp33_ASAP7_75t_L g458 ( .A1(n_85), .A2(n_147), .B(n_152), .C(n_459), .Y(n_458) );
INVx2_ASAP7_75t_L g111 ( .A(n_86), .Y(n_111) );
OR2x2_ASAP7_75t_L g439 ( .A(n_86), .B(n_440), .Y(n_439) );
OR2x2_ASAP7_75t_L g718 ( .A(n_86), .B(n_441), .Y(n_718) );
A2O1A1Ixp33_ASAP7_75t_L g223 ( .A1(n_87), .A2(n_152), .B(n_224), .C(n_227), .Y(n_223) );
OAI22xp5_ASAP7_75t_SL g719 ( .A1(n_88), .A2(n_720), .B1(n_721), .B2(n_724), .Y(n_719) );
CKINVDCx20_ASAP7_75t_R g724 ( .A(n_88), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_89), .B(n_169), .Y(n_483) );
CKINVDCx20_ASAP7_75t_R g464 ( .A(n_90), .Y(n_464) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_91), .Y(n_125) );
A2O1A1Ixp33_ASAP7_75t_L g527 ( .A1(n_92), .A2(n_147), .B(n_152), .C(n_528), .Y(n_527) );
CKINVDCx20_ASAP7_75t_R g534 ( .A(n_93), .Y(n_534) );
INVx1_ASAP7_75t_L g469 ( .A(n_94), .Y(n_469) );
CKINVDCx16_ASAP7_75t_R g539 ( .A(n_95), .Y(n_539) );
NAND2xp5_ASAP7_75t_SL g529 ( .A(n_96), .B(n_237), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_97), .A2(n_104), .B1(n_115), .B2(n_734), .Y(n_103) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_98), .B(n_135), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_99), .B(n_135), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_100), .B(n_114), .Y(n_113) );
INVx2_ASAP7_75t_L g159 ( .A(n_101), .Y(n_159) );
AOI21xp5_ASAP7_75t_L g467 ( .A1(n_102), .A2(n_142), .B(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
CKINVDCx12_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_SL g735 ( .A(n_107), .Y(n_735) );
OR2x2_ASAP7_75t_L g107 ( .A(n_108), .B(n_110), .Y(n_107) );
OR2x2_ASAP7_75t_L g717 ( .A(n_111), .B(n_441), .Y(n_717) );
NOR2x2_ASAP7_75t_L g732 ( .A(n_111), .B(n_440), .Y(n_732) );
INVx1_ASAP7_75t_SL g112 ( .A(n_113), .Y(n_112) );
AO21x1_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_121), .B(n_446), .Y(n_115) );
INVx1_ASAP7_75t_SL g116 ( .A(n_117), .Y(n_116) );
BUFx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx2_ASAP7_75t_SL g733 ( .A(n_118), .Y(n_733) );
BUFx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
OAI21xp5_ASAP7_75t_SL g121 ( .A1(n_122), .A2(n_437), .B(n_444), .Y(n_121) );
INVx1_ASAP7_75t_L g436 ( .A(n_123), .Y(n_436) );
AOI22xp5_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_127), .B1(n_433), .B2(n_434), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g433 ( .A(n_124), .Y(n_433) );
OAI22xp5_ASAP7_75t_L g725 ( .A1(n_127), .A2(n_717), .B1(n_726), .B2(n_727), .Y(n_725) );
BUFx2_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx1_ASAP7_75t_L g434 ( .A(n_128), .Y(n_434) );
AND2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_359), .Y(n_128) );
NOR4xp25_ASAP7_75t_L g129 ( .A(n_130), .B(n_301), .C(n_331), .D(n_341), .Y(n_129) );
OAI211xp5_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_206), .B(n_264), .C(n_291), .Y(n_130) );
OAI222xp33_ASAP7_75t_L g386 ( .A1(n_131), .A2(n_306), .B1(n_387), .B2(n_388), .C1(n_389), .C2(n_390), .Y(n_386) );
OR2x2_ASAP7_75t_L g131 ( .A(n_132), .B(n_181), .Y(n_131) );
AOI33xp33_ASAP7_75t_L g312 ( .A1(n_132), .A2(n_299), .A3(n_300), .B1(n_313), .B2(n_318), .B3(n_320), .Y(n_312) );
OAI211xp5_ASAP7_75t_SL g369 ( .A1(n_132), .A2(n_370), .B(n_372), .C(n_374), .Y(n_369) );
OR2x2_ASAP7_75t_L g385 ( .A(n_132), .B(n_371), .Y(n_385) );
INVx1_ASAP7_75t_L g418 ( .A(n_132), .Y(n_418) );
OR2x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_168), .Y(n_132) );
INVx2_ASAP7_75t_L g295 ( .A(n_133), .Y(n_295) );
AND2x2_ASAP7_75t_L g311 ( .A(n_133), .B(n_197), .Y(n_311) );
HB1xp67_ASAP7_75t_L g346 ( .A(n_133), .Y(n_346) );
AND2x2_ASAP7_75t_L g375 ( .A(n_133), .B(n_168), .Y(n_375) );
OA21x2_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_141), .B(n_165), .Y(n_133) );
OA21x2_ASAP7_75t_L g197 ( .A1(n_134), .A2(n_198), .B(n_205), .Y(n_197) );
OA21x2_ASAP7_75t_L g210 ( .A1(n_134), .A2(n_211), .B(n_219), .Y(n_210) );
HB1xp67_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx4_ASAP7_75t_L g167 ( .A(n_135), .Y(n_167) );
OA21x2_ASAP7_75t_L g466 ( .A1(n_135), .A2(n_467), .B(n_474), .Y(n_466) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx1_ASAP7_75t_L g252 ( .A(n_136), .Y(n_252) );
AND2x2_ASAP7_75t_L g136 ( .A(n_137), .B(n_138), .Y(n_136) );
AND2x2_ASAP7_75t_SL g169 ( .A(n_137), .B(n_138), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_139), .B(n_140), .Y(n_138) );
BUFx2_ASAP7_75t_L g254 ( .A(n_142), .Y(n_254) );
AND2x4_ASAP7_75t_L g142 ( .A(n_143), .B(n_147), .Y(n_142) );
NAND2x1p5_ASAP7_75t_L g187 ( .A(n_143), .B(n_147), .Y(n_187) );
AND2x2_ASAP7_75t_L g143 ( .A(n_144), .B(n_146), .Y(n_143) );
INVx1_ASAP7_75t_L g240 ( .A(n_144), .Y(n_240) );
INVx1_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx2_ASAP7_75t_L g153 ( .A(n_145), .Y(n_153) );
INVx1_ASAP7_75t_L g163 ( .A(n_145), .Y(n_163) );
INVx1_ASAP7_75t_L g154 ( .A(n_146), .Y(n_154) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_146), .Y(n_157) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_146), .Y(n_161) );
INVx3_ASAP7_75t_L g177 ( .A(n_146), .Y(n_177) );
INVx1_ASAP7_75t_L g471 ( .A(n_146), .Y(n_471) );
INVx4_ASAP7_75t_SL g164 ( .A(n_147), .Y(n_164) );
BUFx3_ASAP7_75t_L g241 ( .A(n_147), .Y(n_241) );
O2A1O1Ixp33_ASAP7_75t_SL g149 ( .A1(n_150), .A2(n_151), .B(n_155), .C(n_164), .Y(n_149) );
O2A1O1Ixp33_ASAP7_75t_SL g171 ( .A1(n_151), .A2(n_164), .B(n_172), .C(n_173), .Y(n_171) );
O2A1O1Ixp33_ASAP7_75t_SL g199 ( .A1(n_151), .A2(n_164), .B(n_200), .C(n_201), .Y(n_199) );
O2A1O1Ixp33_ASAP7_75t_L g212 ( .A1(n_151), .A2(n_164), .B(n_213), .C(n_214), .Y(n_212) );
O2A1O1Ixp33_ASAP7_75t_SL g255 ( .A1(n_151), .A2(n_164), .B(n_256), .C(n_257), .Y(n_255) );
O2A1O1Ixp33_ASAP7_75t_L g468 ( .A1(n_151), .A2(n_164), .B(n_469), .C(n_470), .Y(n_468) );
O2A1O1Ixp33_ASAP7_75t_L g478 ( .A1(n_151), .A2(n_164), .B(n_479), .C(n_480), .Y(n_478) );
O2A1O1Ixp33_ASAP7_75t_L g538 ( .A1(n_151), .A2(n_164), .B(n_539), .C(n_540), .Y(n_538) );
INVx5_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
AND2x6_ASAP7_75t_L g152 ( .A(n_153), .B(n_154), .Y(n_152) );
BUFx3_ASAP7_75t_L g179 ( .A(n_153), .Y(n_179) );
BUFx6f_ASAP7_75t_L g218 ( .A(n_153), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g215 ( .A(n_156), .B(n_216), .Y(n_215) );
INVx4_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx2_ASAP7_75t_L g174 ( .A(n_157), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g158 ( .A(n_159), .B(n_160), .Y(n_158) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_160), .B(n_203), .Y(n_202) );
OAI22xp33_ASAP7_75t_L g258 ( .A1(n_160), .A2(n_237), .B1(n_259), .B2(n_260), .Y(n_258) );
NOR2xp33_ASAP7_75t_L g541 ( .A(n_160), .B(n_542), .Y(n_541) );
INVx4_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx2_ASAP7_75t_L g192 ( .A(n_161), .Y(n_192) );
OAI22xp5_ASAP7_75t_SL g493 ( .A1(n_161), .A2(n_192), .B1(n_494), .B2(n_495), .Y(n_493) );
INVx2_ASAP7_75t_L g462 ( .A(n_162), .Y(n_462) );
INVx3_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx1_ASAP7_75t_L g227 ( .A(n_164), .Y(n_227) );
OAI22xp33_ASAP7_75t_L g491 ( .A1(n_164), .A2(n_187), .B1(n_492), .B2(n_496), .Y(n_491) );
OA21x2_ASAP7_75t_L g476 ( .A1(n_166), .A2(n_477), .B(n_483), .Y(n_476) );
INVx3_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g195 ( .A(n_167), .B(n_196), .Y(n_195) );
AO21x2_ASAP7_75t_L g220 ( .A1(n_167), .A2(n_221), .B(n_228), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_167), .B(n_243), .Y(n_242) );
NOR2xp33_ASAP7_75t_SL g513 ( .A(n_167), .B(n_514), .Y(n_513) );
INVx2_ASAP7_75t_L g275 ( .A(n_168), .Y(n_275) );
BUFx3_ASAP7_75t_L g283 ( .A(n_168), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_168), .B(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g294 ( .A(n_168), .B(n_295), .Y(n_294) );
NOR2xp33_ASAP7_75t_L g323 ( .A(n_168), .B(n_182), .Y(n_323) );
AND2x2_ASAP7_75t_L g392 ( .A(n_168), .B(n_326), .Y(n_392) );
OA21x2_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_170), .B(n_180), .Y(n_168) );
INVx1_ASAP7_75t_L g184 ( .A(n_169), .Y(n_184) );
INVx2_ASAP7_75t_L g230 ( .A(n_169), .Y(n_230) );
O2A1O1Ixp33_ASAP7_75t_L g232 ( .A1(n_169), .A2(n_187), .B(n_233), .C(n_234), .Y(n_232) );
OA21x2_ASAP7_75t_L g536 ( .A1(n_169), .A2(n_537), .B(n_543), .Y(n_536) );
NOR2xp33_ASAP7_75t_L g175 ( .A(n_176), .B(n_177), .Y(n_175) );
INVx5_ASAP7_75t_L g237 ( .A(n_177), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g472 ( .A(n_177), .B(n_473), .Y(n_472) );
NOR2xp33_ASAP7_75t_L g481 ( .A(n_177), .B(n_482), .Y(n_481) );
INVx2_ASAP7_75t_L g194 ( .A(n_178), .Y(n_194) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
INVx1_ASAP7_75t_L g204 ( .A(n_179), .Y(n_204) );
INVx2_ASAP7_75t_SL g286 ( .A(n_181), .Y(n_286) );
OR2x2_ASAP7_75t_L g181 ( .A(n_182), .B(n_197), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_182), .B(n_275), .Y(n_274) );
INVx1_ASAP7_75t_L g328 ( .A(n_182), .Y(n_328) );
AND2x2_ASAP7_75t_L g339 ( .A(n_182), .B(n_295), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_182), .B(n_324), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_182), .B(n_326), .Y(n_371) );
AND2x2_ASAP7_75t_L g430 ( .A(n_182), .B(n_375), .Y(n_430) );
INVx4_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
AND2x2_ASAP7_75t_L g300 ( .A(n_183), .B(n_197), .Y(n_300) );
AND2x2_ASAP7_75t_L g310 ( .A(n_183), .B(n_311), .Y(n_310) );
BUFx3_ASAP7_75t_L g332 ( .A(n_183), .Y(n_332) );
AND3x2_ASAP7_75t_L g391 ( .A(n_183), .B(n_392), .C(n_393), .Y(n_391) );
AO21x2_ASAP7_75t_L g183 ( .A1(n_184), .A2(n_185), .B(n_195), .Y(n_183) );
NOR2xp33_ASAP7_75t_L g463 ( .A(n_184), .B(n_464), .Y(n_463) );
NOR2xp33_ASAP7_75t_L g522 ( .A(n_184), .B(n_523), .Y(n_522) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_184), .B(n_534), .Y(n_533) );
OAI21xp5_ASAP7_75t_L g185 ( .A1(n_186), .A2(n_187), .B(n_188), .Y(n_185) );
OAI21xp5_ASAP7_75t_L g221 ( .A1(n_187), .A2(n_222), .B(n_223), .Y(n_221) );
OAI21xp5_ASAP7_75t_L g456 ( .A1(n_187), .A2(n_457), .B(n_458), .Y(n_456) );
OAI21xp5_ASAP7_75t_L g516 ( .A1(n_187), .A2(n_517), .B(n_518), .Y(n_516) );
O2A1O1Ixp5_ASAP7_75t_L g189 ( .A1(n_190), .A2(n_191), .B(n_193), .C(n_194), .Y(n_189) );
O2A1O1Ixp33_ASAP7_75t_L g224 ( .A1(n_191), .A2(n_194), .B(n_225), .C(n_226), .Y(n_224) );
INVx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_194), .A2(n_511), .B(n_512), .Y(n_510) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_194), .A2(n_520), .B(n_521), .Y(n_519) );
HB1xp67_ASAP7_75t_L g282 ( .A(n_197), .Y(n_282) );
INVx1_ASAP7_75t_SL g326 ( .A(n_197), .Y(n_326) );
NAND3xp33_ASAP7_75t_L g338 ( .A(n_197), .B(n_275), .C(n_339), .Y(n_338) );
NOR2xp33_ASAP7_75t_L g206 ( .A(n_207), .B(n_244), .Y(n_206) );
A2O1A1Ixp33_ASAP7_75t_L g361 ( .A1(n_207), .A2(n_310), .B(n_362), .C(n_364), .Y(n_361) );
INVx1_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_209), .B(n_231), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_209), .B(n_368), .Y(n_367) );
INVx2_ASAP7_75t_SL g378 ( .A(n_209), .Y(n_378) );
AND2x2_ASAP7_75t_L g399 ( .A(n_209), .B(n_246), .Y(n_399) );
NOR2xp33_ASAP7_75t_L g427 ( .A(n_209), .B(n_308), .Y(n_427) );
AND2x2_ASAP7_75t_L g209 ( .A(n_210), .B(n_220), .Y(n_209) );
AND2x2_ASAP7_75t_L g272 ( .A(n_210), .B(n_263), .Y(n_272) );
INVx2_ASAP7_75t_L g279 ( .A(n_210), .Y(n_279) );
AND2x2_ASAP7_75t_L g299 ( .A(n_210), .B(n_246), .Y(n_299) );
AND2x2_ASAP7_75t_L g349 ( .A(n_210), .B(n_231), .Y(n_349) );
INVx1_ASAP7_75t_L g353 ( .A(n_210), .Y(n_353) );
INVx3_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
HB1xp67_ASAP7_75t_L g531 ( .A(n_218), .Y(n_531) );
INVx2_ASAP7_75t_SL g263 ( .A(n_220), .Y(n_263) );
BUFx2_ASAP7_75t_L g289 ( .A(n_220), .Y(n_289) );
AND2x2_ASAP7_75t_L g416 ( .A(n_220), .B(n_231), .Y(n_416) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_229), .B(n_230), .Y(n_228) );
INVx1_ASAP7_75t_L g262 ( .A(n_230), .Y(n_262) );
AO21x2_ASAP7_75t_L g525 ( .A1(n_230), .A2(n_526), .B(n_533), .Y(n_525) );
INVx3_ASAP7_75t_SL g246 ( .A(n_231), .Y(n_246) );
AND2x2_ASAP7_75t_L g271 ( .A(n_231), .B(n_272), .Y(n_271) );
AND2x4_ASAP7_75t_L g278 ( .A(n_231), .B(n_279), .Y(n_278) );
OR2x2_ASAP7_75t_L g308 ( .A(n_231), .B(n_268), .Y(n_308) );
OR2x2_ASAP7_75t_L g317 ( .A(n_231), .B(n_263), .Y(n_317) );
HB1xp67_ASAP7_75t_L g335 ( .A(n_231), .Y(n_335) );
AND2x2_ASAP7_75t_L g340 ( .A(n_231), .B(n_293), .Y(n_340) );
AND2x2_ASAP7_75t_L g368 ( .A(n_231), .B(n_248), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_231), .B(n_404), .Y(n_403) );
OR2x2_ASAP7_75t_L g406 ( .A(n_231), .B(n_247), .Y(n_406) );
OR2x6_ASAP7_75t_L g231 ( .A(n_232), .B(n_242), .Y(n_231) );
O2A1O1Ixp33_ASAP7_75t_L g235 ( .A1(n_236), .A2(n_237), .B(n_238), .C(n_239), .Y(n_235) );
O2A1O1Ixp33_ASAP7_75t_L g459 ( .A1(n_237), .A2(n_460), .B(n_461), .C(n_462), .Y(n_459) );
INVx2_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
NAND2xp5_ASAP7_75t_SL g257 ( .A(n_240), .B(n_258), .Y(n_257) );
INVx1_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
OR2x2_ASAP7_75t_L g245 ( .A(n_246), .B(n_247), .Y(n_245) );
AND2x2_ASAP7_75t_L g330 ( .A(n_246), .B(n_279), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_246), .B(n_272), .Y(n_358) );
AND2x2_ASAP7_75t_L g376 ( .A(n_246), .B(n_293), .Y(n_376) );
OR2x2_ASAP7_75t_L g247 ( .A(n_248), .B(n_263), .Y(n_247) );
AND2x2_ASAP7_75t_L g277 ( .A(n_248), .B(n_263), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_248), .B(n_306), .Y(n_305) );
BUFx3_ASAP7_75t_L g315 ( .A(n_248), .Y(n_315) );
OR2x2_ASAP7_75t_L g363 ( .A(n_248), .B(n_283), .Y(n_363) );
OA21x2_ASAP7_75t_L g248 ( .A1(n_249), .A2(n_253), .B(n_261), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
AO21x2_ASAP7_75t_L g268 ( .A1(n_250), .A2(n_269), .B(n_270), .Y(n_268) );
AO21x2_ASAP7_75t_L g515 ( .A1(n_250), .A2(n_516), .B(n_522), .Y(n_515) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
AOI21xp5_ASAP7_75t_SL g507 ( .A1(n_251), .A2(n_508), .B(n_509), .Y(n_507) );
INVx2_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
AO21x2_ASAP7_75t_L g455 ( .A1(n_252), .A2(n_456), .B(n_463), .Y(n_455) );
AO21x2_ASAP7_75t_L g490 ( .A1(n_252), .A2(n_491), .B(n_497), .Y(n_490) );
NOR2xp33_ASAP7_75t_L g497 ( .A(n_252), .B(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g269 ( .A(n_253), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_261), .Y(n_270) );
AND2x2_ASAP7_75t_L g298 ( .A(n_263), .B(n_268), .Y(n_298) );
INVx1_ASAP7_75t_L g306 ( .A(n_263), .Y(n_306) );
AND2x2_ASAP7_75t_L g401 ( .A(n_263), .B(n_279), .Y(n_401) );
AOI222xp33_ASAP7_75t_L g264 ( .A1(n_265), .A2(n_273), .B1(n_276), .B2(n_280), .C1(n_284), .C2(n_287), .Y(n_264) );
INVx1_ASAP7_75t_L g396 ( .A(n_265), .Y(n_396) );
AND2x2_ASAP7_75t_L g265 ( .A(n_266), .B(n_271), .Y(n_265) );
AND2x2_ASAP7_75t_L g292 ( .A(n_266), .B(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g303 ( .A(n_266), .B(n_272), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_266), .B(n_294), .Y(n_319) );
OAI222xp33_ASAP7_75t_L g341 ( .A1(n_266), .A2(n_342), .B1(n_347), .B2(n_348), .C1(n_356), .C2(n_358), .Y(n_341) );
INVx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
INVx1_ASAP7_75t_SL g267 ( .A(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g329 ( .A(n_268), .B(n_330), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_268), .B(n_349), .Y(n_389) );
AND2x2_ASAP7_75t_L g400 ( .A(n_268), .B(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g408 ( .A(n_271), .Y(n_408) );
NAND2xp5_ASAP7_75t_SL g387 ( .A(n_273), .B(n_324), .Y(n_387) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
NOR2xp33_ASAP7_75t_L g327 ( .A(n_275), .B(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g345 ( .A(n_275), .B(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
INVx3_ASAP7_75t_L g290 ( .A(n_278), .Y(n_290) );
O2A1O1Ixp33_ASAP7_75t_L g380 ( .A1(n_278), .A2(n_381), .B(n_384), .C(n_386), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_278), .B(n_315), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_278), .B(n_298), .Y(n_420) );
AND2x2_ASAP7_75t_L g293 ( .A(n_279), .B(n_289), .Y(n_293) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
INVx1_ASAP7_75t_L g320 ( .A(n_282), .Y(n_320) );
NAND2xp5_ASAP7_75t_SL g309 ( .A(n_283), .B(n_310), .Y(n_309) );
OR2x2_ASAP7_75t_L g372 ( .A(n_283), .B(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g411 ( .A(n_283), .B(n_311), .Y(n_411) );
INVx1_ASAP7_75t_L g423 ( .A(n_283), .Y(n_423) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_286), .B(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
OR2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_290), .Y(n_288) );
INVx1_ASAP7_75t_L g404 ( .A(n_289), .Y(n_404) );
A2O1A1Ixp33_ASAP7_75t_SL g291 ( .A1(n_292), .A2(n_294), .B(n_296), .C(n_300), .Y(n_291) );
AOI22xp33_ASAP7_75t_L g336 ( .A1(n_292), .A2(n_322), .B1(n_337), .B2(n_340), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_293), .B(n_307), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_293), .B(n_315), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_294), .B(n_352), .Y(n_351) );
INVx1_ASAP7_75t_SL g357 ( .A(n_294), .Y(n_357) );
AND2x2_ASAP7_75t_L g364 ( .A(n_294), .B(n_344), .Y(n_364) );
INVx2_ASAP7_75t_L g325 ( .A(n_295), .Y(n_325) );
INVxp67_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
NOR4xp25_ASAP7_75t_L g302 ( .A(n_299), .B(n_303), .C(n_304), .D(n_307), .Y(n_302) );
INVx1_ASAP7_75t_SL g373 ( .A(n_300), .Y(n_373) );
AND2x2_ASAP7_75t_L g417 ( .A(n_300), .B(n_418), .Y(n_417) );
OAI211xp5_ASAP7_75t_SL g301 ( .A1(n_302), .A2(n_309), .B(n_312), .C(n_321), .Y(n_301) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx1_ASAP7_75t_SL g307 ( .A(n_308), .Y(n_307) );
NOR2xp33_ASAP7_75t_L g429 ( .A(n_308), .B(n_378), .Y(n_429) );
AOI22xp5_ASAP7_75t_L g428 ( .A1(n_310), .A2(n_429), .B1(n_430), .B2(n_431), .Y(n_428) );
INVx1_ASAP7_75t_SL g383 ( .A(n_311), .Y(n_383) );
AND2x2_ASAP7_75t_L g422 ( .A(n_311), .B(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
NAND2xp5_ASAP7_75t_SL g415 ( .A(n_315), .B(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
NOR2xp33_ASAP7_75t_L g334 ( .A(n_319), .B(n_335), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_320), .B(n_345), .Y(n_405) );
OAI21xp5_ASAP7_75t_SL g321 ( .A1(n_322), .A2(n_327), .B(n_329), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
INVx1_ASAP7_75t_L g397 ( .A(n_324), .Y(n_397) );
AND2x2_ASAP7_75t_L g324 ( .A(n_325), .B(n_326), .Y(n_324) );
INVx2_ASAP7_75t_L g425 ( .A(n_325), .Y(n_425) );
HB1xp67_ASAP7_75t_L g352 ( .A(n_326), .Y(n_352) );
OAI21xp33_ASAP7_75t_L g331 ( .A1(n_332), .A2(n_333), .B(n_336), .Y(n_331) );
CKINVDCx16_ASAP7_75t_R g344 ( .A(n_332), .Y(n_344) );
OR2x2_ASAP7_75t_L g382 ( .A(n_332), .B(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
AOI21xp33_ASAP7_75t_SL g377 ( .A1(n_335), .A2(n_378), .B(n_379), .Y(n_377) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
AOI221xp5_ASAP7_75t_L g365 ( .A1(n_339), .A2(n_366), .B1(n_369), .B2(n_376), .C(n_377), .Y(n_365) );
INVx1_ASAP7_75t_SL g409 ( .A(n_340), .Y(n_409) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
OR2x2_ASAP7_75t_L g356 ( .A(n_344), .B(n_357), .Y(n_356) );
INVxp67_ASAP7_75t_L g393 ( .A(n_346), .Y(n_393) );
AOI22xp5_ASAP7_75t_L g348 ( .A1(n_349), .A2(n_350), .B1(n_353), .B2(n_354), .Y(n_348) );
INVx1_ASAP7_75t_L g388 ( .A(n_349), .Y(n_388) );
INVxp67_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_352), .B(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
NOR4xp25_ASAP7_75t_L g359 ( .A(n_360), .B(n_394), .C(n_407), .D(n_419), .Y(n_359) );
NAND3xp33_ASAP7_75t_SL g360 ( .A(n_361), .B(n_365), .C(n_380), .Y(n_360) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
NOR2xp33_ASAP7_75t_L g381 ( .A(n_363), .B(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_370), .B(n_375), .Y(n_379) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
OAI221xp5_ASAP7_75t_SL g407 ( .A1(n_382), .A2(n_408), .B1(n_409), .B2(n_410), .C(n_412), .Y(n_407) );
O2A1O1Ixp33_ASAP7_75t_L g398 ( .A1(n_384), .A2(n_399), .B(n_400), .C(n_402), .Y(n_398) );
INVx2_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
OAI22xp5_ASAP7_75t_L g402 ( .A1(n_385), .A2(n_403), .B1(n_405), .B2(n_406), .Y(n_402) );
INVx2_ASAP7_75t_SL g390 ( .A(n_391), .Y(n_390) );
A2O1A1Ixp33_ASAP7_75t_L g394 ( .A1(n_395), .A2(n_396), .B(n_397), .C(n_398), .Y(n_394) );
INVx1_ASAP7_75t_L g413 ( .A(n_406), .Y(n_413) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
OAI21xp5_ASAP7_75t_SL g412 ( .A1(n_413), .A2(n_414), .B(n_417), .Y(n_412) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
OAI221xp5_ASAP7_75t_SL g419 ( .A1(n_420), .A2(n_421), .B1(n_424), .B2(n_426), .C(n_428), .Y(n_419) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVxp67_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
OAI22xp5_ASAP7_75t_SL g448 ( .A1(n_434), .A2(n_449), .B1(n_717), .B2(n_718), .Y(n_448) );
INVx1_ASAP7_75t_SL g437 ( .A(n_438), .Y(n_437) );
HB1xp67_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_SL g445 ( .A(n_439), .Y(n_445) );
INVx2_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_442), .B(n_443), .Y(n_441) );
AOI21xp33_ASAP7_75t_SL g446 ( .A1(n_444), .A2(n_447), .B(n_733), .Y(n_446) );
INVx1_ASAP7_75t_L g726 ( .A(n_449), .Y(n_726) );
NAND2x1_ASAP7_75t_L g449 ( .A(n_450), .B(n_633), .Y(n_449) );
NOR5xp2_ASAP7_75t_L g450 ( .A(n_451), .B(n_556), .C(n_588), .D(n_603), .E(n_620), .Y(n_450) );
A2O1A1Ixp33_ASAP7_75t_L g451 ( .A1(n_452), .A2(n_484), .B(n_503), .C(n_544), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_453), .B(n_465), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_453), .B(n_656), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_453), .B(n_608), .Y(n_671) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_454), .B(n_553), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_454), .B(n_500), .Y(n_557) );
AND2x2_ASAP7_75t_L g598 ( .A(n_454), .B(n_599), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_454), .B(n_567), .Y(n_602) );
OR2x2_ASAP7_75t_L g639 ( .A(n_454), .B(n_490), .Y(n_639) );
INVx3_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
AND2x2_ASAP7_75t_L g489 ( .A(n_455), .B(n_490), .Y(n_489) );
INVx3_ASAP7_75t_L g547 ( .A(n_455), .Y(n_547) );
OR2x2_ASAP7_75t_L g710 ( .A(n_455), .B(n_550), .Y(n_710) );
AOI22xp5_ASAP7_75t_L g612 ( .A1(n_465), .A2(n_613), .B1(n_614), .B2(n_617), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_465), .B(n_547), .Y(n_696) );
AND2x2_ASAP7_75t_L g465 ( .A(n_466), .B(n_475), .Y(n_465) );
AND2x2_ASAP7_75t_L g502 ( .A(n_466), .B(n_490), .Y(n_502) );
AND2x2_ASAP7_75t_L g549 ( .A(n_466), .B(n_550), .Y(n_549) );
INVx1_ASAP7_75t_L g554 ( .A(n_466), .Y(n_554) );
INVx3_ASAP7_75t_L g567 ( .A(n_466), .Y(n_567) );
OR2x2_ASAP7_75t_L g587 ( .A(n_466), .B(n_550), .Y(n_587) );
AND2x2_ASAP7_75t_L g606 ( .A(n_466), .B(n_476), .Y(n_606) );
BUFx2_ASAP7_75t_L g638 ( .A(n_466), .Y(n_638) );
AND2x4_ASAP7_75t_L g553 ( .A(n_475), .B(n_554), .Y(n_553) );
INVx1_ASAP7_75t_SL g475 ( .A(n_476), .Y(n_475) );
BUFx2_ASAP7_75t_L g488 ( .A(n_476), .Y(n_488) );
INVx2_ASAP7_75t_L g501 ( .A(n_476), .Y(n_501) );
OR2x2_ASAP7_75t_L g569 ( .A(n_476), .B(n_550), .Y(n_569) );
AND2x2_ASAP7_75t_L g599 ( .A(n_476), .B(n_490), .Y(n_599) );
AND2x2_ASAP7_75t_L g616 ( .A(n_476), .B(n_547), .Y(n_616) );
AND2x2_ASAP7_75t_L g656 ( .A(n_476), .B(n_567), .Y(n_656) );
AND2x2_ASAP7_75t_SL g692 ( .A(n_476), .B(n_502), .Y(n_692) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
NAND2xp33_ASAP7_75t_SL g485 ( .A(n_486), .B(n_499), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_487), .B(n_489), .Y(n_486) );
NOR2xp33_ASAP7_75t_L g670 ( .A(n_487), .B(n_671), .Y(n_670) );
INVx1_ASAP7_75t_SL g487 ( .A(n_488), .Y(n_487) );
OAI21xp33_ASAP7_75t_L g630 ( .A1(n_488), .A2(n_502), .B(n_631), .Y(n_630) );
NOR2xp33_ASAP7_75t_L g686 ( .A(n_488), .B(n_490), .Y(n_686) );
AND2x2_ASAP7_75t_L g622 ( .A(n_489), .B(n_623), .Y(n_622) );
INVx3_ASAP7_75t_L g550 ( .A(n_490), .Y(n_550) );
HB1xp67_ASAP7_75t_L g648 ( .A(n_490), .Y(n_648) );
NOR2xp33_ASAP7_75t_L g715 ( .A(n_499), .B(n_547), .Y(n_715) );
INVx2_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
AOI22xp33_ASAP7_75t_L g657 ( .A1(n_500), .A2(n_658), .B1(n_659), .B2(n_664), .Y(n_657) );
AND2x2_ASAP7_75t_L g500 ( .A(n_501), .B(n_502), .Y(n_500) );
AND2x2_ASAP7_75t_L g548 ( .A(n_501), .B(n_549), .Y(n_548) );
OR2x2_ASAP7_75t_L g586 ( .A(n_501), .B(n_587), .Y(n_586) );
INVx1_ASAP7_75t_SL g623 ( .A(n_501), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_502), .B(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g677 ( .A(n_502), .Y(n_677) );
CKINVDCx16_ASAP7_75t_R g503 ( .A(n_504), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_505), .B(n_524), .Y(n_504) );
INVx4_ASAP7_75t_L g563 ( .A(n_505), .Y(n_563) );
AND2x2_ASAP7_75t_L g641 ( .A(n_505), .B(n_608), .Y(n_641) );
AND2x2_ASAP7_75t_L g505 ( .A(n_506), .B(n_515), .Y(n_505) );
INVx3_ASAP7_75t_L g560 ( .A(n_506), .Y(n_560) );
AND2x2_ASAP7_75t_L g574 ( .A(n_506), .B(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g578 ( .A(n_506), .Y(n_578) );
INVx2_ASAP7_75t_L g592 ( .A(n_506), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_506), .B(n_608), .Y(n_607) );
AND2x2_ASAP7_75t_L g649 ( .A(n_506), .B(n_644), .Y(n_649) );
AND2x2_ASAP7_75t_L g714 ( .A(n_506), .B(n_684), .Y(n_714) );
OR2x6_ASAP7_75t_L g506 ( .A(n_507), .B(n_513), .Y(n_506) );
AND2x2_ASAP7_75t_L g555 ( .A(n_515), .B(n_536), .Y(n_555) );
INVx2_ASAP7_75t_L g575 ( .A(n_515), .Y(n_575) );
INVx1_ASAP7_75t_L g580 ( .A(n_524), .Y(n_580) );
AND2x2_ASAP7_75t_L g626 ( .A(n_524), .B(n_574), .Y(n_626) );
AND2x2_ASAP7_75t_L g524 ( .A(n_525), .B(n_535), .Y(n_524) );
INVx2_ASAP7_75t_L g565 ( .A(n_525), .Y(n_565) );
INVx1_ASAP7_75t_L g573 ( .A(n_525), .Y(n_573) );
AND2x2_ASAP7_75t_L g591 ( .A(n_525), .B(n_592), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_525), .B(n_575), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_527), .B(n_532), .Y(n_526) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_529), .A2(n_530), .B(n_531), .Y(n_528) );
AND2x2_ASAP7_75t_L g608 ( .A(n_535), .B(n_565), .Y(n_608) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx2_ASAP7_75t_L g561 ( .A(n_536), .Y(n_561) );
AND2x2_ASAP7_75t_L g644 ( .A(n_536), .B(n_575), .Y(n_644) );
OAI21xp5_ASAP7_75t_SL g544 ( .A1(n_545), .A2(n_551), .B(n_555), .Y(n_544) );
INVx1_ASAP7_75t_SL g589 ( .A(n_545), .Y(n_589) );
AND2x2_ASAP7_75t_L g545 ( .A(n_546), .B(n_548), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_546), .B(n_553), .Y(n_646) );
INVx1_ASAP7_75t_SL g546 ( .A(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g595 ( .A(n_547), .B(n_550), .Y(n_595) );
AND2x2_ASAP7_75t_L g624 ( .A(n_547), .B(n_568), .Y(n_624) );
OR2x2_ASAP7_75t_L g627 ( .A(n_547), .B(n_587), .Y(n_627) );
AOI222xp33_ASAP7_75t_L g691 ( .A1(n_548), .A2(n_640), .B1(n_692), .B2(n_693), .C1(n_695), .C2(n_697), .Y(n_691) );
BUFx2_ASAP7_75t_L g605 ( .A(n_550), .Y(n_605) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g594 ( .A(n_553), .B(n_595), .Y(n_594) );
INVx3_ASAP7_75t_SL g611 ( .A(n_553), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_553), .B(n_605), .Y(n_665) );
AND2x2_ASAP7_75t_L g600 ( .A(n_555), .B(n_560), .Y(n_600) );
INVx1_ASAP7_75t_L g619 ( .A(n_555), .Y(n_619) );
OAI221xp5_ASAP7_75t_SL g556 ( .A1(n_557), .A2(n_558), .B1(n_562), .B2(n_566), .C(n_570), .Y(n_556) );
OR2x2_ASAP7_75t_L g628 ( .A(n_558), .B(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_560), .B(n_561), .Y(n_559) );
AND2x2_ASAP7_75t_L g613 ( .A(n_560), .B(n_583), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_560), .B(n_573), .Y(n_653) );
AND2x2_ASAP7_75t_L g658 ( .A(n_560), .B(n_608), .Y(n_658) );
HB1xp67_ASAP7_75t_L g668 ( .A(n_560), .Y(n_668) );
NAND2x1_ASAP7_75t_SL g679 ( .A(n_560), .B(n_680), .Y(n_679) );
OR2x2_ASAP7_75t_L g564 ( .A(n_561), .B(n_565), .Y(n_564) );
INVx2_ASAP7_75t_L g584 ( .A(n_561), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_561), .B(n_579), .Y(n_610) );
INVx1_ASAP7_75t_L g676 ( .A(n_561), .Y(n_676) );
INVx1_ASAP7_75t_L g651 ( .A(n_562), .Y(n_651) );
OR2x2_ASAP7_75t_L g562 ( .A(n_563), .B(n_564), .Y(n_562) );
INVx1_ASAP7_75t_L g663 ( .A(n_563), .Y(n_663) );
NOR2xp67_ASAP7_75t_L g675 ( .A(n_563), .B(n_676), .Y(n_675) );
INVx2_ASAP7_75t_L g680 ( .A(n_564), .Y(n_680) );
NOR2xp33_ASAP7_75t_L g687 ( .A(n_564), .B(n_688), .Y(n_687) );
AND2x2_ASAP7_75t_L g583 ( .A(n_565), .B(n_584), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_565), .B(n_575), .Y(n_596) );
INVx1_ASAP7_75t_L g662 ( .A(n_565), .Y(n_662) );
INVx1_ASAP7_75t_L g683 ( .A(n_566), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .Y(n_566) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
OAI21xp5_ASAP7_75t_SL g570 ( .A1(n_571), .A2(n_576), .B(n_585), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_572), .B(n_574), .Y(n_571) );
AND2x2_ASAP7_75t_L g716 ( .A(n_572), .B(n_649), .Y(n_716) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g684 ( .A(n_573), .B(n_644), .Y(n_684) );
AOI32xp33_ASAP7_75t_L g597 ( .A1(n_574), .A2(n_580), .A3(n_598), .B1(n_600), .B2(n_601), .Y(n_597) );
AOI322xp5_ASAP7_75t_L g699 ( .A1(n_574), .A2(n_606), .A3(n_689), .B1(n_700), .B2(n_701), .C1(n_702), .C2(n_704), .Y(n_699) );
INVx2_ASAP7_75t_L g579 ( .A(n_575), .Y(n_579) );
INVx1_ASAP7_75t_L g689 ( .A(n_575), .Y(n_689) );
OAI22xp5_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_580), .B1(n_581), .B2(n_582), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_577), .B(n_583), .Y(n_632) );
AND2x2_ASAP7_75t_L g577 ( .A(n_578), .B(n_579), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_578), .B(n_644), .Y(n_694) );
INVx1_ASAP7_75t_L g581 ( .A(n_579), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_579), .B(n_608), .Y(n_698) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx1_ASAP7_75t_SL g585 ( .A(n_586), .Y(n_585) );
NOR2xp33_ASAP7_75t_L g681 ( .A(n_587), .B(n_682), .Y(n_681) );
OAI221xp5_ASAP7_75t_SL g588 ( .A1(n_589), .A2(n_590), .B1(n_593), .B2(n_596), .C(n_597), .Y(n_588) );
OR2x2_ASAP7_75t_L g609 ( .A(n_590), .B(n_610), .Y(n_609) );
OR2x2_ASAP7_75t_L g618 ( .A(n_590), .B(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g643 ( .A(n_591), .B(n_644), .Y(n_643) );
INVx2_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
AND2x2_ASAP7_75t_L g647 ( .A(n_601), .B(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
OAI221xp5_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_607), .B1(n_609), .B2(n_611), .C(n_612), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_605), .B(n_606), .Y(n_604) );
AOI22xp5_ASAP7_75t_L g635 ( .A1(n_605), .A2(n_636), .B1(n_640), .B2(n_641), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_606), .B(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g711 ( .A(n_606), .Y(n_711) );
INVx1_ASAP7_75t_L g705 ( .A(n_608), .Y(n_705) );
INVx1_ASAP7_75t_SL g640 ( .A(n_609), .Y(n_640) );
NOR2xp33_ASAP7_75t_L g701 ( .A(n_611), .B(n_639), .Y(n_701) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_616), .B(n_675), .Y(n_674) );
INVx1_ASAP7_75t_SL g682 ( .A(n_616), .Y(n_682) );
INVx1_ASAP7_75t_SL g617 ( .A(n_618), .Y(n_617) );
OAI221xp5_ASAP7_75t_SL g620 ( .A1(n_621), .A2(n_625), .B1(n_627), .B2(n_628), .C(n_630), .Y(n_620) );
NOR2xp33_ASAP7_75t_SL g621 ( .A(n_622), .B(n_624), .Y(n_621) );
AOI22xp5_ASAP7_75t_L g685 ( .A1(n_622), .A2(n_640), .B1(n_686), .B2(n_687), .Y(n_685) );
CKINVDCx14_ASAP7_75t_R g625 ( .A(n_626), .Y(n_625) );
OAI21xp33_ASAP7_75t_L g704 ( .A1(n_627), .A2(n_705), .B(n_706), .Y(n_704) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
NOR3xp33_ASAP7_75t_SL g633 ( .A(n_634), .B(n_666), .C(n_690), .Y(n_633) );
NAND4xp25_ASAP7_75t_L g634 ( .A(n_635), .B(n_642), .C(n_650), .D(n_657), .Y(n_634) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
OR2x2_ASAP7_75t_L g637 ( .A(n_638), .B(n_639), .Y(n_637) );
INVx1_ASAP7_75t_L g713 ( .A(n_638), .Y(n_713) );
INVx3_ASAP7_75t_SL g707 ( .A(n_639), .Y(n_707) );
OR2x2_ASAP7_75t_L g712 ( .A(n_639), .B(n_713), .Y(n_712) );
AOI22xp5_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_645), .B1(n_647), .B2(n_649), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_644), .B(n_662), .Y(n_703) );
INVxp67_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
OAI21xp5_ASAP7_75t_SL g650 ( .A1(n_651), .A2(n_652), .B(n_654), .Y(n_650) );
INVxp67_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_661), .B(n_663), .Y(n_660) );
INVxp67_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
OAI211xp5_ASAP7_75t_SL g666 ( .A1(n_667), .A2(n_669), .B(n_672), .C(n_685), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g700 ( .A(n_671), .Y(n_700) );
AOI222xp33_ASAP7_75t_L g672 ( .A1(n_673), .A2(n_677), .B1(n_678), .B2(n_681), .C1(n_683), .C2(n_684), .Y(n_672) );
INVxp67_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
NAND4xp25_ASAP7_75t_SL g709 ( .A(n_682), .B(n_710), .C(n_711), .D(n_712), .Y(n_709) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
NAND3xp33_ASAP7_75t_SL g690 ( .A(n_691), .B(n_699), .C(n_708), .Y(n_690) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
AOI22xp33_ASAP7_75t_L g708 ( .A1(n_709), .A2(n_714), .B1(n_715), .B2(n_716), .Y(n_708) );
INVx1_ASAP7_75t_L g728 ( .A(n_718), .Y(n_728) );
INVx1_ASAP7_75t_L g729 ( .A(n_719), .Y(n_729) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx2_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_SL g730 ( .A(n_731), .Y(n_730) );
INVx2_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
endmodule