module fake_jpeg_14623_n_147 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_147);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_147;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_28),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_9),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_3),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_3),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_27),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_2),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_59),
.B(n_0),
.Y(n_60)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_64),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_53),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_42),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_65),
.B(n_54),
.Y(n_83)
);

INVx2_ASAP7_75t_R g66 ( 
.A(n_55),
.Y(n_66)
);

NAND2xp33_ASAP7_75t_SL g81 ( 
.A(n_66),
.B(n_67),
.Y(n_81)
);

AOI21xp33_ASAP7_75t_L g67 ( 
.A1(n_43),
.A2(n_0),
.B(n_1),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_62),
.A2(n_51),
.B1(n_44),
.B2(n_45),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_68),
.A2(n_70),
.B1(n_56),
.B2(n_4),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_66),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_64),
.A2(n_41),
.B1(n_47),
.B2(n_51),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_61),
.A2(n_45),
.B1(n_48),
.B2(n_58),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_71),
.A2(n_75),
.B1(n_52),
.B2(n_50),
.Y(n_84)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

INVx3_ASAP7_75t_SL g93 ( 
.A(n_73),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_61),
.A2(n_48),
.B1(n_58),
.B2(n_50),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_64),
.B(n_57),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_76),
.B(n_49),
.Y(n_85)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_77),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_82),
.B(n_83),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_84),
.A2(n_96),
.B1(n_71),
.B2(n_9),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_85),
.B(n_86),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_SL g86 ( 
.A(n_81),
.B(n_56),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_78),
.B(n_1),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_88),
.B(n_92),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_90),
.A2(n_97),
.B1(n_98),
.B2(n_100),
.Y(n_108)
);

NAND2xp33_ASAP7_75t_SL g91 ( 
.A(n_68),
.B(n_2),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_91),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_4),
.Y(n_92)
);

NAND2xp33_ASAP7_75t_SL g96 ( 
.A(n_79),
.B(n_5),
.Y(n_96)
);

HAxp5_ASAP7_75t_SL g97 ( 
.A(n_69),
.B(n_5),
.CON(n_97),
.SN(n_97)
);

OA22x2_ASAP7_75t_L g98 ( 
.A1(n_80),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_73),
.B(n_6),
.Y(n_99)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_99),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_75),
.A2(n_22),
.B1(n_38),
.B2(n_36),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_82),
.B(n_7),
.Y(n_101)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_101),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_89),
.Y(n_104)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_104),
.Y(n_115)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_105),
.Y(n_116)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_95),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_107),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_110),
.A2(n_98),
.B1(n_97),
.B2(n_84),
.Y(n_113)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_94),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_112),
.B(n_87),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_R g122 ( 
.A(n_113),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_111),
.B(n_86),
.C(n_93),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_114),
.B(n_109),
.Y(n_120)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_117),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_120),
.B(n_121),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_115),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_113),
.A2(n_109),
.B(n_108),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_123),
.A2(n_108),
.B(n_98),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_119),
.B(n_106),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_124),
.B(n_125),
.Y(n_130)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_123),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_122),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_127),
.B(n_129),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_128),
.A2(n_118),
.B1(n_116),
.B2(n_102),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_119),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_126),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_132),
.B(n_103),
.C(n_128),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_133),
.B(n_93),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_134),
.B(n_135),
.C(n_133),
.Y(n_137)
);

OAI21xp33_ASAP7_75t_L g136 ( 
.A1(n_134),
.A2(n_130),
.B(n_131),
.Y(n_136)
);

HB1xp67_ASAP7_75t_L g138 ( 
.A(n_136),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_137),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_139),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_23),
.Y(n_141)
);

CKINVDCx14_ASAP7_75t_R g142 ( 
.A(n_141),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_142),
.A2(n_20),
.B(n_34),
.Y(n_143)
);

AO221x1_ASAP7_75t_L g144 ( 
.A1(n_143),
.A2(n_19),
.B1(n_33),
.B2(n_11),
.C(n_13),
.Y(n_144)
);

OAI321xp33_ASAP7_75t_L g145 ( 
.A1(n_144),
.A2(n_26),
.A3(n_32),
.B1(n_14),
.B2(n_16),
.C(n_17),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_145),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_30),
.Y(n_147)
);


endmodule