module fake_jpeg_18972_n_378 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_378);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_378;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_377;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_1),
.B(n_7),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_2),
.B(n_4),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_2),
.B(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx14_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_4),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_24),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_38),
.B(n_39),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_24),
.B(n_25),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

BUFx10_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g96 ( 
.A(n_41),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx4_ASAP7_75t_SL g98 ( 
.A(n_44),
.Y(n_98)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_45),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_25),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_46),
.B(n_55),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_17),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_50),
.A2(n_35),
.B1(n_20),
.B2(n_31),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_51),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_27),
.B(n_36),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_53),
.B(n_34),
.Y(n_87)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_27),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

CKINVDCx9p33_ASAP7_75t_R g57 ( 
.A(n_34),
.Y(n_57)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_58),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_16),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_59),
.B(n_40),
.Y(n_82)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_16),
.Y(n_61)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_61),
.Y(n_100)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_17),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_38),
.A2(n_17),
.B1(n_32),
.B2(n_36),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_72),
.A2(n_73),
.B1(n_80),
.B2(n_99),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_46),
.A2(n_36),
.B1(n_32),
.B2(n_18),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_78),
.A2(n_88),
.B1(n_92),
.B2(n_97),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_55),
.A2(n_32),
.B1(n_18),
.B2(n_26),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_82),
.B(n_94),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_87),
.B(n_91),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_50),
.A2(n_19),
.B1(n_26),
.B2(n_28),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_53),
.B(n_35),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_89),
.B(n_102),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_61),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_45),
.A2(n_19),
.B1(n_28),
.B2(n_29),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_39),
.B(n_29),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_59),
.B(n_21),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_95),
.B(n_41),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_49),
.A2(n_19),
.B1(n_21),
.B2(n_30),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_43),
.A2(n_35),
.B1(n_31),
.B2(n_30),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_54),
.A2(n_31),
.B1(n_30),
.B2(n_20),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_101),
.A2(n_47),
.B1(n_42),
.B2(n_48),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_65),
.B(n_20),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_101),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g145 ( 
.A(n_107),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_108),
.B(n_114),
.Y(n_154)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_67),
.Y(n_110)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_110),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_65),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_111),
.B(n_112),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_87),
.B(n_42),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_102),
.Y(n_113)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_113),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_77),
.B(n_44),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_69),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_115),
.Y(n_170)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_85),
.Y(n_116)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_116),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_83),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_117),
.B(n_127),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_76),
.Y(n_118)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_118),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_74),
.A2(n_62),
.B1(n_60),
.B2(n_57),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_119),
.A2(n_120),
.B1(n_141),
.B2(n_142),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_74),
.A2(n_64),
.B1(n_56),
.B2(n_41),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_69),
.Y(n_122)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_122),
.Y(n_150)
);

OAI21xp33_ASAP7_75t_L g123 ( 
.A1(n_91),
.A2(n_0),
.B(n_1),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_123),
.B(n_134),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_66),
.B(n_51),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_124),
.B(n_144),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_66),
.B(n_41),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_125),
.B(n_126),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_100),
.B(n_41),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_85),
.Y(n_127)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_67),
.Y(n_128)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_128),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_88),
.A2(n_64),
.B1(n_63),
.B2(n_58),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_129),
.A2(n_90),
.B1(n_75),
.B2(n_79),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_100),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_130),
.B(n_132),
.Y(n_175)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_68),
.Y(n_131)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_131),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_78),
.B(n_63),
.Y(n_132)
);

OAI32xp33_ASAP7_75t_L g133 ( 
.A1(n_81),
.A2(n_58),
.A3(n_52),
.B1(n_51),
.B2(n_48),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_133),
.B(n_104),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_81),
.B(n_52),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_68),
.Y(n_135)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_135),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_137),
.A2(n_107),
.B1(n_113),
.B2(n_136),
.Y(n_146)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_71),
.Y(n_138)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_138),
.Y(n_173)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_83),
.Y(n_139)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_139),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_76),
.Y(n_140)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_140),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_98),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_98),
.B(n_3),
.Y(n_142)
);

BUFx8_ASAP7_75t_L g143 ( 
.A(n_96),
.Y(n_143)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_143),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_103),
.B(n_47),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_146),
.A2(n_160),
.B1(n_166),
.B2(n_179),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_121),
.A2(n_71),
.B1(n_93),
.B2(n_86),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_162),
.A2(n_172),
.B1(n_174),
.B2(n_135),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_115),
.A2(n_104),
.B(n_93),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_163),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_130),
.A2(n_98),
.B1(n_70),
.B2(n_79),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_164),
.A2(n_165),
.B1(n_168),
.B2(n_151),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_106),
.A2(n_84),
.B1(n_86),
.B2(n_90),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_106),
.B(n_103),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_167),
.B(n_171),
.Y(n_199)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_124),
.Y(n_169)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_169),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_111),
.B(n_103),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_121),
.A2(n_84),
.B1(n_70),
.B2(n_75),
.Y(n_172)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_144),
.Y(n_176)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_176),
.Y(n_189)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_131),
.Y(n_178)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_178),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_112),
.A2(n_76),
.B1(n_96),
.B2(n_6),
.Y(n_179)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_173),
.Y(n_181)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_181),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_152),
.B(n_109),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_182),
.B(n_191),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_152),
.B(n_109),
.C(n_126),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_183),
.B(n_185),
.C(n_13),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_148),
.B(n_125),
.C(n_126),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_145),
.A2(n_133),
.B1(n_129),
.B2(n_127),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_186),
.A2(n_190),
.B1(n_217),
.B2(n_11),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_159),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_187),
.B(n_194),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_147),
.B(n_125),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_188),
.A2(n_197),
.B(n_207),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_167),
.B(n_122),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_150),
.B(n_105),
.Y(n_193)
);

CKINVDCx14_ASAP7_75t_R g225 ( 
.A(n_193),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_158),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_150),
.B(n_110),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_195),
.B(n_204),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_160),
.A2(n_139),
.B(n_142),
.Y(n_197)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_156),
.Y(n_200)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_200),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_180),
.B(n_140),
.Y(n_201)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_201),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_180),
.B(n_138),
.Y(n_202)
);

OAI21xp33_ASAP7_75t_L g229 ( 
.A1(n_202),
.A2(n_206),
.B(n_178),
.Y(n_229)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_156),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_203),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_154),
.B(n_128),
.Y(n_204)
);

FAx1_ASAP7_75t_SL g205 ( 
.A(n_147),
.B(n_96),
.CI(n_143),
.CON(n_205),
.SN(n_205)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_205),
.B(n_12),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_148),
.B(n_116),
.Y(n_206)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_157),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_208),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_174),
.A2(n_140),
.B1(n_118),
.B2(n_6),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_209),
.A2(n_218),
.B1(n_179),
.B2(n_169),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_146),
.A2(n_118),
.B1(n_143),
.B2(n_8),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_210),
.A2(n_153),
.B1(n_161),
.B2(n_149),
.Y(n_227)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_168),
.Y(n_211)
);

INVx2_ASAP7_75t_SL g240 ( 
.A(n_211),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_173),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_212),
.Y(n_223)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_157),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_213),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_163),
.B(n_3),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_214),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_175),
.B(n_3),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_215),
.Y(n_252)
);

INVx8_ASAP7_75t_L g216 ( 
.A(n_155),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_216),
.A2(n_165),
.B1(n_149),
.B2(n_161),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_166),
.B(n_3),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_176),
.A2(n_5),
.B1(n_9),
.B2(n_10),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_220),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_183),
.B(n_171),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_221),
.B(n_239),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_222),
.A2(n_231),
.B1(n_235),
.B2(n_237),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_227),
.A2(n_234),
.B1(n_207),
.B2(n_209),
.Y(n_260)
);

CKINVDCx14_ASAP7_75t_R g271 ( 
.A(n_229),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_192),
.A2(n_170),
.B1(n_177),
.B2(n_159),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_198),
.A2(n_177),
.B1(n_170),
.B2(n_151),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_192),
.A2(n_177),
.B1(n_155),
.B2(n_143),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_197),
.A2(n_5),
.B1(n_9),
.B2(n_10),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_191),
.B(n_5),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_188),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_241)
);

NAND2xp33_ASAP7_75t_R g254 ( 
.A(n_241),
.B(n_242),
.Y(n_254)
);

MAJx2_ASAP7_75t_L g242 ( 
.A(n_188),
.B(n_11),
.C(n_12),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_244),
.A2(n_246),
.B1(n_247),
.B2(n_187),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_185),
.B(n_11),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_245),
.B(n_249),
.C(n_205),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_190),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_198),
.A2(n_201),
.B1(n_199),
.B2(n_184),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_248),
.B(n_218),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_182),
.B(n_13),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_250),
.B(n_15),
.C(n_245),
.Y(n_280)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_224),
.Y(n_253)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_253),
.Y(n_282)
);

INVxp33_ASAP7_75t_SL g255 ( 
.A(n_238),
.Y(n_255)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_255),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_256),
.B(n_257),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_226),
.B(n_194),
.Y(n_257)
);

A2O1A1Ixp33_ASAP7_75t_L g258 ( 
.A1(n_251),
.A2(n_199),
.B(n_184),
.C(n_189),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_258),
.B(n_262),
.Y(n_298)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_224),
.Y(n_259)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_259),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_260),
.A2(n_272),
.B1(n_276),
.B2(n_278),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_251),
.B(n_202),
.Y(n_262)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_233),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_264),
.B(n_275),
.Y(n_299)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_228),
.Y(n_265)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_265),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_225),
.B(n_247),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_266),
.B(n_267),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_237),
.B(n_206),
.Y(n_267)
);

NAND3xp33_ASAP7_75t_SL g268 ( 
.A(n_234),
.B(n_189),
.C(n_208),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_268),
.B(n_269),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_270),
.B(n_280),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_227),
.A2(n_210),
.B1(n_213),
.B2(n_196),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_273),
.A2(n_230),
.B1(n_252),
.B2(n_239),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_221),
.B(n_205),
.C(n_196),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_249),
.C(n_231),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_228),
.B(n_200),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_219),
.A2(n_203),
.B1(n_216),
.B2(n_181),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_232),
.Y(n_277)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_277),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_219),
.A2(n_216),
.B1(n_211),
.B2(n_212),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_222),
.A2(n_15),
.B1(n_212),
.B2(n_246),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_279),
.A2(n_223),
.B1(n_236),
.B2(n_243),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_281),
.A2(n_280),
.B1(n_240),
.B2(n_15),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_274),
.B(n_248),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_284),
.B(n_287),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_285),
.A2(n_292),
.B1(n_301),
.B2(n_260),
.Y(n_305)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_275),
.Y(n_286)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_286),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_261),
.A2(n_235),
.B(n_230),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_288),
.B(n_291),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_271),
.B(n_241),
.Y(n_291)
);

HB1xp67_ASAP7_75t_L g293 ( 
.A(n_262),
.Y(n_293)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_293),
.Y(n_306)
);

A2O1A1Ixp33_ASAP7_75t_L g300 ( 
.A1(n_258),
.A2(n_242),
.B(n_252),
.C(n_250),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_300),
.B(n_291),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_273),
.A2(n_223),
.B1(n_240),
.B2(n_233),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_263),
.B(n_240),
.C(n_15),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_302),
.B(n_296),
.C(n_283),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_287),
.B(n_263),
.C(n_270),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_304),
.B(n_296),
.C(n_302),
.Y(n_326)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_305),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_294),
.A2(n_261),
.B1(n_269),
.B2(n_279),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_307),
.A2(n_310),
.B1(n_317),
.B2(n_285),
.Y(n_327)
);

HB1xp67_ASAP7_75t_L g309 ( 
.A(n_298),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_309),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_294),
.A2(n_265),
.B1(n_272),
.B2(n_277),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_284),
.B(n_276),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_312),
.B(n_313),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_SL g313 ( 
.A(n_298),
.B(n_254),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_299),
.Y(n_314)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_314),
.Y(n_336)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_299),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_315),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_301),
.A2(n_278),
.B1(n_256),
.B2(n_253),
.Y(n_317)
);

OA21x2_ASAP7_75t_L g318 ( 
.A1(n_281),
.A2(n_259),
.B(n_256),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_318),
.B(n_288),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_283),
.B(n_264),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_319),
.B(n_320),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_321),
.B(n_322),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_326),
.B(n_332),
.C(n_334),
.Y(n_338)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_327),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_321),
.B(n_303),
.Y(n_328)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_328),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_307),
.A2(n_290),
.B1(n_295),
.B2(n_289),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_330),
.A2(n_315),
.B1(n_314),
.B2(n_306),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_322),
.B(n_295),
.C(n_289),
.Y(n_332)
);

XOR2x2_ASAP7_75t_L g333 ( 
.A(n_313),
.B(n_318),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_333),
.A2(n_337),
.B(n_316),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_312),
.B(n_282),
.C(n_297),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_330),
.B(n_318),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_339),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_340),
.B(n_348),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_332),
.B(n_310),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_342),
.B(n_343),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_329),
.B(n_334),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_324),
.A2(n_317),
.B(n_333),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_344),
.A2(n_349),
.B1(n_336),
.B2(n_306),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_323),
.Y(n_345)
);

OR2x2_ASAP7_75t_L g354 ( 
.A(n_345),
.B(n_329),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_326),
.B(n_311),
.C(n_304),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_347),
.B(n_325),
.C(n_335),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_335),
.B(n_311),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_SL g364 ( 
.A(n_350),
.B(n_308),
.Y(n_364)
);

HB1xp67_ASAP7_75t_L g352 ( 
.A(n_344),
.Y(n_352)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_352),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_354),
.B(n_356),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_338),
.B(n_305),
.C(n_331),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_338),
.B(n_331),
.C(n_297),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_357),
.B(n_358),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_SL g358 ( 
.A(n_348),
.B(n_327),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_359),
.B(n_349),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_351),
.B(n_347),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_361),
.B(n_362),
.Y(n_367)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_355),
.B(n_346),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_SL g369 ( 
.A1(n_363),
.A2(n_345),
.B(n_352),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_SL g368 ( 
.A(n_364),
.B(n_353),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_368),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g372 ( 
.A1(n_369),
.A2(n_370),
.B(n_371),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_SL g370 ( 
.A1(n_366),
.A2(n_340),
.B(n_336),
.Y(n_370)
);

AO21x1_ASAP7_75t_L g371 ( 
.A1(n_363),
.A2(n_354),
.B(n_358),
.Y(n_371)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_373),
.A2(n_367),
.B(n_360),
.Y(n_374)
);

OA21x2_ASAP7_75t_SL g375 ( 
.A1(n_374),
.A2(n_372),
.B(n_365),
.Y(n_375)
);

HB1xp67_ASAP7_75t_L g376 ( 
.A(n_375),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_376),
.A2(n_362),
.B1(n_341),
.B2(n_282),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_377),
.B(n_341),
.C(n_300),
.Y(n_378)
);


endmodule