module fake_netlist_6_921_n_2044 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_2044);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_2044;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1371;
wire n_1285;
wire n_200;
wire n_1985;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_2018;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_405;
wire n_213;
wire n_538;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_1970;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_1413;
wire n_1330;
wire n_1605;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_210;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1886;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_701;
wire n_295;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_527;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_2037;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_2017;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2026;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1373;
wire n_1292;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_2020;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1848;
wire n_763;
wire n_1147;
wire n_1785;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_2022;
wire n_1945;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_390;
wire n_1148;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_2001;
wire n_1884;
wire n_206;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_187),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_68),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_114),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_48),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_126),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_65),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g204 ( 
.A(n_56),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_196),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_158),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_48),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_113),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_109),
.Y(n_209)
);

BUFx5_ASAP7_75t_L g210 ( 
.A(n_150),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_74),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_86),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_17),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_2),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_134),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_184),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_82),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_50),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_9),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_32),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_183),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_21),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_29),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_26),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_154),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_174),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_136),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_135),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_8),
.Y(n_229)
);

BUFx10_ASAP7_75t_L g230 ( 
.A(n_102),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_189),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_4),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_67),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_6),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_115),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_119),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_148),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_74),
.Y(n_238)
);

BUFx2_ASAP7_75t_L g239 ( 
.A(n_77),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_10),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_29),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_123),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_2),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_169),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_139),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_144),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_14),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_73),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_170),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_163),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_122),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_42),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_161),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_54),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_15),
.Y(n_255)
);

INVx1_ASAP7_75t_SL g256 ( 
.A(n_142),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_5),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_173),
.Y(n_258)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_15),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_116),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_147),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_172),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g263 ( 
.A(n_54),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_101),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_177),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_25),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_180),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_76),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_73),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_108),
.Y(n_270)
);

INVx4_ASAP7_75t_R g271 ( 
.A(n_194),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_43),
.Y(n_272)
);

CKINVDCx14_ASAP7_75t_R g273 ( 
.A(n_192),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_138),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_35),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_44),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_121),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_83),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_47),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_131),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_84),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_157),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_124),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_165),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_190),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_6),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_120),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_64),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_21),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_28),
.Y(n_290)
);

CKINVDCx14_ASAP7_75t_R g291 ( 
.A(n_68),
.Y(n_291)
);

INVx1_ASAP7_75t_SL g292 ( 
.A(n_67),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_40),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_96),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_36),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_7),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_37),
.Y(n_297)
);

INVxp33_ASAP7_75t_SL g298 ( 
.A(n_43),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_23),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_75),
.Y(n_300)
);

BUFx5_ASAP7_75t_L g301 ( 
.A(n_88),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_31),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_129),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_149),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_4),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_56),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_91),
.Y(n_307)
);

BUFx5_ASAP7_75t_L g308 ( 
.A(n_39),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_98),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_85),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_151),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_127),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_145),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_66),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_72),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_133),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_63),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_153),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_156),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_143),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_51),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_5),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_167),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_40),
.Y(n_324)
);

INVx2_ASAP7_75t_SL g325 ( 
.A(n_99),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_162),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_107),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_181),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_9),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_50),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_16),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_155),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_17),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_16),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_10),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_185),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_61),
.Y(n_337)
);

BUFx2_ASAP7_75t_L g338 ( 
.A(n_171),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_118),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_58),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_65),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_97),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_137),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_27),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_63),
.Y(n_345)
);

BUFx3_ASAP7_75t_L g346 ( 
.A(n_110),
.Y(n_346)
);

BUFx3_ASAP7_75t_L g347 ( 
.A(n_44),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_42),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_175),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_182),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_60),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_35),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_130),
.Y(n_353)
);

BUFx2_ASAP7_75t_L g354 ( 
.A(n_81),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_76),
.Y(n_355)
);

CKINVDCx16_ASAP7_75t_R g356 ( 
.A(n_89),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_47),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_58),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_1),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_26),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_62),
.Y(n_361)
);

BUFx10_ASAP7_75t_L g362 ( 
.A(n_193),
.Y(n_362)
);

BUFx2_ASAP7_75t_SL g363 ( 
.A(n_28),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_62),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_51),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_61),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_72),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_128),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_66),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_38),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_38),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_93),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_52),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_31),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_19),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_179),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_11),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_57),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_103),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_59),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_64),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_166),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_188),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_57),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_39),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_69),
.Y(n_386)
);

HB1xp67_ASAP7_75t_L g387 ( 
.A(n_117),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_25),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_92),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_1),
.Y(n_390)
);

BUFx3_ASAP7_75t_L g391 ( 
.A(n_19),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_104),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_7),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_195),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_239),
.B(n_338),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_308),
.Y(n_396)
);

BUFx2_ASAP7_75t_L g397 ( 
.A(n_204),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_236),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_200),
.Y(n_399)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_199),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_251),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_258),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_202),
.Y(n_403)
);

NOR2xp67_ASAP7_75t_L g404 ( 
.A(n_248),
.B(n_0),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_262),
.Y(n_405)
);

CKINVDCx16_ASAP7_75t_R g406 ( 
.A(n_291),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_308),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_208),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_226),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_308),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_308),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_249),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_253),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_308),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_265),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_308),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_247),
.B(n_0),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_274),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_343),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_308),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_308),
.Y(n_421)
);

INVxp67_ASAP7_75t_SL g422 ( 
.A(n_387),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_272),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_277),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_272),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_272),
.Y(n_426)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_363),
.Y(n_427)
);

INVxp67_ASAP7_75t_SL g428 ( 
.A(n_354),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_282),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_272),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_319),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_356),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_272),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_284),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_273),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_211),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_222),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_222),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_325),
.B(n_298),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_330),
.Y(n_440)
);

INVxp67_ASAP7_75t_SL g441 ( 
.A(n_346),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_330),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_210),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_199),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_247),
.Y(n_445)
);

INVxp33_ASAP7_75t_SL g446 ( 
.A(n_201),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_259),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_259),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_303),
.Y(n_449)
);

INVxp67_ASAP7_75t_SL g450 ( 
.A(n_346),
.Y(n_450)
);

BUFx2_ASAP7_75t_L g451 ( 
.A(n_347),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_307),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_347),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_309),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_312),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_391),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_316),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_320),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_323),
.Y(n_459)
);

NOR2xp67_ASAP7_75t_L g460 ( 
.A(n_214),
.B(n_3),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_327),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_391),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_328),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_219),
.Y(n_464)
);

NOR2xp67_ASAP7_75t_L g465 ( 
.A(n_325),
.B(n_3),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_294),
.B(n_8),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_254),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_224),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_210),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_318),
.B(n_11),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_255),
.Y(n_471)
);

HB1xp67_ASAP7_75t_L g472 ( 
.A(n_201),
.Y(n_472)
);

HB1xp67_ASAP7_75t_L g473 ( 
.A(n_203),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_257),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_232),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_268),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_252),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_266),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_279),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_198),
.Y(n_480)
);

HB1xp67_ASAP7_75t_L g481 ( 
.A(n_203),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_205),
.B(n_12),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_289),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_198),
.Y(n_484)
);

INVxp33_ASAP7_75t_L g485 ( 
.A(n_293),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_317),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_269),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_322),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_210),
.Y(n_489)
);

CKINVDCx16_ASAP7_75t_R g490 ( 
.A(n_230),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_205),
.B(n_12),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_344),
.Y(n_492)
);

CKINVDCx16_ASAP7_75t_R g493 ( 
.A(n_230),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_276),
.Y(n_494)
);

CKINVDCx16_ASAP7_75t_R g495 ( 
.A(n_230),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_236),
.Y(n_496)
);

HB1xp67_ASAP7_75t_L g497 ( 
.A(n_400),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_423),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_423),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_425),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_420),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_420),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_398),
.Y(n_503)
);

BUFx2_ASAP7_75t_L g504 ( 
.A(n_467),
.Y(n_504)
);

HB1xp67_ASAP7_75t_L g505 ( 
.A(n_444),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_441),
.B(n_209),
.Y(n_506)
);

OAI21x1_ASAP7_75t_L g507 ( 
.A1(n_396),
.A2(n_267),
.B(n_245),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_398),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_450),
.B(n_209),
.Y(n_509)
);

HB1xp67_ASAP7_75t_L g510 ( 
.A(n_472),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_398),
.Y(n_511)
);

AND2x4_ASAP7_75t_L g512 ( 
.A(n_417),
.B(n_245),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_425),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_398),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_426),
.Y(n_515)
);

BUFx2_ASAP7_75t_L g516 ( 
.A(n_471),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_426),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_398),
.Y(n_518)
);

BUFx6f_ASAP7_75t_L g519 ( 
.A(n_398),
.Y(n_519)
);

INVx3_ASAP7_75t_L g520 ( 
.A(n_496),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_406),
.B(n_362),
.Y(n_521)
);

HB1xp67_ASAP7_75t_L g522 ( 
.A(n_473),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_430),
.Y(n_523)
);

NAND2x1p5_ASAP7_75t_L g524 ( 
.A(n_465),
.B(n_236),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_496),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_496),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_496),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_496),
.Y(n_528)
);

HB1xp67_ASAP7_75t_L g529 ( 
.A(n_481),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_496),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_430),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_396),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_433),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_433),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_407),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_407),
.Y(n_536)
);

AND2x6_ASAP7_75t_L g537 ( 
.A(n_417),
.B(n_267),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_410),
.Y(n_538)
);

INVx3_ASAP7_75t_L g539 ( 
.A(n_443),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_410),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_443),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_411),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_445),
.B(n_283),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_SL g544 ( 
.A(n_406),
.B(n_263),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_411),
.Y(n_545)
);

AND2x4_ASAP7_75t_L g546 ( 
.A(n_414),
.B(n_283),
.Y(n_546)
);

NAND3xp33_ASAP7_75t_L g547 ( 
.A(n_439),
.B(n_288),
.C(n_286),
.Y(n_547)
);

INVx3_ASAP7_75t_L g548 ( 
.A(n_469),
.Y(n_548)
);

INVx5_ASAP7_75t_L g549 ( 
.A(n_469),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_414),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_416),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_416),
.B(n_215),
.Y(n_552)
);

CKINVDCx8_ASAP7_75t_R g553 ( 
.A(n_490),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_421),
.Y(n_554)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_489),
.Y(n_555)
);

BUFx6f_ASAP7_75t_L g556 ( 
.A(n_489),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_421),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_437),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_464),
.Y(n_559)
);

AND2x4_ASAP7_75t_L g560 ( 
.A(n_465),
.B(n_313),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_437),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_482),
.B(n_215),
.Y(n_562)
);

CKINVDCx16_ASAP7_75t_R g563 ( 
.A(n_490),
.Y(n_563)
);

AND2x4_ASAP7_75t_L g564 ( 
.A(n_460),
.B(n_313),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_464),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_468),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_468),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_475),
.Y(n_568)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_438),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_475),
.Y(n_570)
);

INVx3_ASAP7_75t_L g571 ( 
.A(n_438),
.Y(n_571)
);

HB1xp67_ASAP7_75t_L g572 ( 
.A(n_451),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_477),
.Y(n_573)
);

OA21x2_ASAP7_75t_L g574 ( 
.A1(n_440),
.A2(n_373),
.B(n_348),
.Y(n_574)
);

OR2x2_ASAP7_75t_SL g575 ( 
.A(n_493),
.B(n_495),
.Y(n_575)
);

AND2x6_ASAP7_75t_L g576 ( 
.A(n_491),
.B(n_236),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_512),
.B(n_401),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_512),
.B(n_402),
.Y(n_578)
);

CKINVDCx20_ASAP7_75t_R g579 ( 
.A(n_563),
.Y(n_579)
);

AOI22xp33_ASAP7_75t_L g580 ( 
.A1(n_512),
.A2(n_395),
.B1(n_422),
.B2(n_397),
.Y(n_580)
);

NOR3xp33_ASAP7_75t_L g581 ( 
.A(n_547),
.B(n_495),
.C(n_493),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_538),
.Y(n_582)
);

HB1xp67_ASAP7_75t_L g583 ( 
.A(n_572),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_512),
.B(n_552),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_503),
.Y(n_585)
);

BUFx10_ASAP7_75t_L g586 ( 
.A(n_537),
.Y(n_586)
);

AND3x2_ASAP7_75t_L g587 ( 
.A(n_544),
.B(n_397),
.C(n_466),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_501),
.Y(n_588)
);

INVx1_ASAP7_75t_SL g589 ( 
.A(n_504),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_538),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_544),
.B(n_405),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_501),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_543),
.B(n_445),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_512),
.B(n_415),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_SL g595 ( 
.A(n_553),
.B(n_431),
.Y(n_595)
);

INVx5_ASAP7_75t_L g596 ( 
.A(n_537),
.Y(n_596)
);

OAI22xp5_ASAP7_75t_L g597 ( 
.A1(n_547),
.A2(n_562),
.B1(n_428),
.B2(n_435),
.Y(n_597)
);

INVx4_ASAP7_75t_L g598 ( 
.A(n_541),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_506),
.B(n_418),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_501),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_552),
.B(n_424),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_540),
.Y(n_602)
);

INVxp33_ASAP7_75t_L g603 ( 
.A(n_572),
.Y(n_603)
);

AND2x6_ASAP7_75t_L g604 ( 
.A(n_560),
.B(n_236),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_506),
.B(n_429),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_501),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_560),
.B(n_434),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_543),
.B(n_447),
.Y(n_608)
);

OR2x2_ASAP7_75t_L g609 ( 
.A(n_509),
.B(n_451),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_560),
.B(n_449),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_560),
.B(n_452),
.Y(n_611)
);

BUFx3_ASAP7_75t_L g612 ( 
.A(n_574),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_509),
.B(n_455),
.Y(n_613)
);

NAND2xp33_ASAP7_75t_L g614 ( 
.A(n_576),
.B(n_210),
.Y(n_614)
);

INVxp33_ASAP7_75t_L g615 ( 
.A(n_497),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_504),
.B(n_457),
.Y(n_616)
);

AO22x2_ASAP7_75t_L g617 ( 
.A1(n_521),
.A2(n_377),
.B1(n_384),
.B2(n_378),
.Y(n_617)
);

AOI22xp5_ASAP7_75t_L g618 ( 
.A1(n_521),
.A2(n_234),
.B1(n_275),
.B2(n_233),
.Y(n_618)
);

INVx4_ASAP7_75t_L g619 ( 
.A(n_541),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_540),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_542),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_560),
.B(n_459),
.Y(n_622)
);

OR2x6_ASAP7_75t_L g623 ( 
.A(n_504),
.B(n_404),
.Y(n_623)
);

AOI22xp33_ASAP7_75t_L g624 ( 
.A1(n_576),
.A2(n_470),
.B1(n_446),
.B2(n_390),
.Y(n_624)
);

INVx3_ASAP7_75t_L g625 ( 
.A(n_503),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_553),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_502),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_516),
.B(n_474),
.Y(n_628)
);

AOI22xp33_ASAP7_75t_L g629 ( 
.A1(n_576),
.A2(n_385),
.B1(n_436),
.B2(n_485),
.Y(n_629)
);

AOI22xp5_ASAP7_75t_L g630 ( 
.A1(n_516),
.A2(n_463),
.B1(n_454),
.B2(n_458),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_502),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_542),
.Y(n_632)
);

NAND3xp33_ASAP7_75t_L g633 ( 
.A(n_497),
.B(n_487),
.C(n_476),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_502),
.Y(n_634)
);

INVx4_ASAP7_75t_L g635 ( 
.A(n_541),
.Y(n_635)
);

AO22x2_ASAP7_75t_L g636 ( 
.A1(n_564),
.A2(n_292),
.B1(n_332),
.B2(n_326),
.Y(n_636)
);

XOR2xp5_ASAP7_75t_L g637 ( 
.A(n_563),
.B(n_399),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_502),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_553),
.Y(n_639)
);

AOI22xp33_ASAP7_75t_L g640 ( 
.A1(n_576),
.A2(n_447),
.B1(n_453),
.B2(n_456),
.Y(n_640)
);

BUFx3_ASAP7_75t_L g641 ( 
.A(n_574),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_532),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_516),
.B(n_494),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_505),
.B(n_461),
.Y(n_644)
);

AOI22xp33_ASAP7_75t_L g645 ( 
.A1(n_576),
.A2(n_448),
.B1(n_453),
.B2(n_456),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_545),
.B(n_227),
.Y(n_646)
);

OR2x6_ASAP7_75t_L g647 ( 
.A(n_505),
.B(n_448),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_532),
.Y(n_648)
);

BUFx6f_ASAP7_75t_L g649 ( 
.A(n_503),
.Y(n_649)
);

INVx2_ASAP7_75t_SL g650 ( 
.A(n_510),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_545),
.B(n_256),
.Y(n_651)
);

AOI22xp33_ASAP7_75t_L g652 ( 
.A1(n_576),
.A2(n_462),
.B1(n_492),
.B2(n_486),
.Y(n_652)
);

INVx4_ASAP7_75t_L g653 ( 
.A(n_541),
.Y(n_653)
);

AND2x6_ASAP7_75t_L g654 ( 
.A(n_546),
.B(n_206),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_510),
.B(n_480),
.Y(n_655)
);

BUFx6f_ASAP7_75t_L g656 ( 
.A(n_503),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_543),
.B(n_462),
.Y(n_657)
);

BUFx3_ASAP7_75t_L g658 ( 
.A(n_574),
.Y(n_658)
);

INVx2_ASAP7_75t_SL g659 ( 
.A(n_522),
.Y(n_659)
);

AND2x2_ASAP7_75t_SL g660 ( 
.A(n_564),
.B(n_212),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_522),
.B(n_484),
.Y(n_661)
);

INVxp33_ASAP7_75t_L g662 ( 
.A(n_529),
.Y(n_662)
);

AOI22xp33_ASAP7_75t_L g663 ( 
.A1(n_576),
.A2(n_492),
.B1(n_488),
.B2(n_486),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_559),
.B(n_440),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_564),
.B(n_432),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_529),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_564),
.B(n_427),
.Y(n_667)
);

BUFx3_ASAP7_75t_L g668 ( 
.A(n_574),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_550),
.Y(n_669)
);

INVx1_ASAP7_75t_SL g670 ( 
.A(n_575),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_532),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_532),
.Y(n_672)
);

AND3x2_ASAP7_75t_L g673 ( 
.A(n_564),
.B(n_228),
.C(n_216),
.Y(n_673)
);

BUFx3_ASAP7_75t_L g674 ( 
.A(n_574),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_576),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_546),
.B(n_362),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_550),
.B(n_270),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_536),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_536),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_546),
.B(n_362),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_559),
.B(n_442),
.Y(n_681)
);

NAND2xp33_ASAP7_75t_R g682 ( 
.A(n_574),
.B(n_217),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_557),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_557),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_565),
.B(n_442),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_535),
.Y(n_686)
);

BUFx3_ASAP7_75t_L g687 ( 
.A(n_537),
.Y(n_687)
);

BUFx10_ASAP7_75t_L g688 ( 
.A(n_537),
.Y(n_688)
);

OAI22xp33_ASAP7_75t_L g689 ( 
.A1(n_524),
.A2(n_331),
.B1(n_299),
.B2(n_297),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_535),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_546),
.B(n_217),
.Y(n_691)
);

AOI22xp33_ASAP7_75t_L g692 ( 
.A1(n_576),
.A2(n_488),
.B1(n_483),
.B2(n_479),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_535),
.B(n_231),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_546),
.B(n_221),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_536),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_536),
.Y(n_696)
);

OR2x2_ASAP7_75t_L g697 ( 
.A(n_575),
.B(n_477),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_551),
.Y(n_698)
);

AND2x6_ASAP7_75t_L g699 ( 
.A(n_551),
.B(n_235),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_551),
.Y(n_700)
);

INVx1_ASAP7_75t_SL g701 ( 
.A(n_575),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_551),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_537),
.B(n_237),
.Y(n_703)
);

INVx5_ASAP7_75t_L g704 ( 
.A(n_537),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_565),
.B(n_403),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_554),
.Y(n_706)
);

AND3x2_ASAP7_75t_L g707 ( 
.A(n_566),
.B(n_250),
.C(n_242),
.Y(n_707)
);

BUFx4f_ASAP7_75t_L g708 ( 
.A(n_576),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_554),
.Y(n_709)
);

INVxp33_ASAP7_75t_L g710 ( 
.A(n_566),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_554),
.Y(n_711)
);

HB1xp67_ASAP7_75t_L g712 ( 
.A(n_567),
.Y(n_712)
);

AND2x4_ASAP7_75t_L g713 ( 
.A(n_567),
.B(n_478),
.Y(n_713)
);

BUFx6f_ASAP7_75t_L g714 ( 
.A(n_503),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_554),
.Y(n_715)
);

BUFx10_ASAP7_75t_L g716 ( 
.A(n_537),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_498),
.Y(n_717)
);

NAND2xp33_ASAP7_75t_L g718 ( 
.A(n_576),
.B(n_210),
.Y(n_718)
);

CKINVDCx14_ASAP7_75t_R g719 ( 
.A(n_537),
.Y(n_719)
);

OR2x6_ASAP7_75t_L g720 ( 
.A(n_568),
.B(n_478),
.Y(n_720)
);

BUFx6f_ASAP7_75t_L g721 ( 
.A(n_503),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_533),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_533),
.Y(n_723)
);

AOI22xp33_ASAP7_75t_L g724 ( 
.A1(n_537),
.A2(n_483),
.B1(n_479),
.B2(n_339),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_524),
.B(n_221),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_498),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_524),
.B(n_225),
.Y(n_727)
);

AOI22xp33_ASAP7_75t_L g728 ( 
.A1(n_537),
.A2(n_264),
.B1(n_287),
.B2(n_310),
.Y(n_728)
);

AND2x4_ASAP7_75t_L g729 ( 
.A(n_720),
.B(n_568),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_722),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_601),
.B(n_225),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_712),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_597),
.B(n_244),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_584),
.B(n_524),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_660),
.B(n_541),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_609),
.B(n_244),
.Y(n_736)
);

INVx2_ASAP7_75t_SL g737 ( 
.A(n_593),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_577),
.B(n_408),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_660),
.B(n_541),
.Y(n_739)
);

AOI22x1_ASAP7_75t_L g740 ( 
.A1(n_636),
.A2(n_617),
.B1(n_675),
.B2(n_686),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_660),
.B(n_541),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_722),
.Y(n_742)
);

AOI22xp5_ASAP7_75t_L g743 ( 
.A1(n_670),
.A2(n_409),
.B1(n_412),
.B2(n_413),
.Y(n_743)
);

NOR2xp67_ASAP7_75t_SL g744 ( 
.A(n_612),
.B(n_503),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_609),
.B(n_246),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_582),
.B(n_541),
.Y(n_746)
);

NOR2x1_ASAP7_75t_L g747 ( 
.A(n_633),
.B(n_260),
.Y(n_747)
);

INVx3_ASAP7_75t_L g748 ( 
.A(n_612),
.Y(n_748)
);

NAND2xp33_ASAP7_75t_L g749 ( 
.A(n_675),
.B(n_210),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_590),
.B(n_555),
.Y(n_750)
);

AND2x2_ASAP7_75t_L g751 ( 
.A(n_593),
.B(n_570),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_710),
.B(n_246),
.Y(n_752)
);

HB1xp67_ASAP7_75t_L g753 ( 
.A(n_583),
.Y(n_753)
);

NAND3xp33_ASAP7_75t_L g754 ( 
.A(n_580),
.B(n_624),
.C(n_628),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_607),
.B(n_336),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_590),
.B(n_555),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_723),
.Y(n_757)
);

NOR2x1p5_ASAP7_75t_L g758 ( 
.A(n_626),
.B(n_207),
.Y(n_758)
);

AND2x2_ASAP7_75t_L g759 ( 
.A(n_608),
.B(n_570),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_578),
.B(n_419),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_602),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_602),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_620),
.Y(n_763)
);

NOR2xp67_ASAP7_75t_L g764 ( 
.A(n_630),
.B(n_573),
.Y(n_764)
);

BUFx8_ASAP7_75t_L g765 ( 
.A(n_650),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_620),
.B(n_555),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_664),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_610),
.B(n_336),
.Y(n_768)
);

OAI22xp5_ASAP7_75t_SL g769 ( 
.A1(n_618),
.A2(n_360),
.B1(n_337),
.B2(n_352),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_611),
.B(n_349),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_664),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_621),
.B(n_555),
.Y(n_772)
);

NAND2xp33_ASAP7_75t_SL g773 ( 
.A(n_697),
.B(n_357),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_681),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_621),
.B(n_632),
.Y(n_775)
);

INVx2_ASAP7_75t_SL g776 ( 
.A(n_608),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_657),
.B(n_573),
.Y(n_777)
);

AOI22xp33_ASAP7_75t_L g778 ( 
.A1(n_641),
.A2(n_507),
.B1(n_304),
.B2(n_392),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_632),
.B(n_555),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_622),
.B(n_349),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_669),
.B(n_555),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_669),
.B(n_683),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_594),
.B(n_350),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_723),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_641),
.Y(n_785)
);

BUFx3_ASAP7_75t_L g786 ( 
.A(n_687),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_689),
.B(n_350),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_658),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_697),
.B(n_353),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_683),
.Y(n_790)
);

BUFx2_ASAP7_75t_L g791 ( 
.A(n_650),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_658),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_603),
.B(n_599),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_684),
.B(n_555),
.Y(n_794)
);

AOI22xp5_ASAP7_75t_L g795 ( 
.A1(n_701),
.A2(n_682),
.B1(n_605),
.B2(n_613),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_684),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_686),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_681),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_690),
.B(n_555),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_L g800 ( 
.A(n_615),
.B(n_353),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_668),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_690),
.B(n_556),
.Y(n_802)
);

A2O1A1Ixp33_ASAP7_75t_L g803 ( 
.A1(n_668),
.A2(n_507),
.B(n_278),
.C(n_280),
.Y(n_803)
);

NAND2xp33_ASAP7_75t_L g804 ( 
.A(n_604),
.B(n_210),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_L g805 ( 
.A(n_662),
.B(n_376),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_717),
.B(n_556),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_685),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_674),
.Y(n_808)
);

OAI22xp33_ASAP7_75t_L g809 ( 
.A1(n_623),
.A2(n_342),
.B1(n_311),
.B2(n_285),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_SL g810 ( 
.A(n_646),
.B(n_376),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_674),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_685),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_717),
.B(n_726),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_726),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_651),
.B(n_389),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_588),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_588),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_677),
.B(n_556),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_698),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_698),
.Y(n_820)
);

INVxp67_ASAP7_75t_L g821 ( 
.A(n_655),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_581),
.B(n_389),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_657),
.B(n_629),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_706),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_592),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_705),
.B(n_394),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_591),
.B(n_616),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_706),
.Y(n_828)
);

INVx3_ASAP7_75t_L g829 ( 
.A(n_687),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_665),
.B(n_394),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_659),
.B(n_261),
.Y(n_831)
);

O2A1O1Ixp33_ASAP7_75t_L g832 ( 
.A1(n_614),
.A2(n_531),
.B(n_523),
.C(n_515),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_626),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_709),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_667),
.B(n_556),
.Y(n_835)
);

O2A1O1Ixp33_ASAP7_75t_L g836 ( 
.A1(n_614),
.A2(n_531),
.B(n_523),
.C(n_515),
.Y(n_836)
);

OAI22xp33_ASAP7_75t_L g837 ( 
.A1(n_623),
.A2(n_281),
.B1(n_368),
.B2(n_372),
.Y(n_837)
);

HB1xp67_ASAP7_75t_L g838 ( 
.A(n_659),
.Y(n_838)
);

BUFx5_ASAP7_75t_L g839 ( 
.A(n_586),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_639),
.Y(n_840)
);

OAI22xp33_ASAP7_75t_L g841 ( 
.A1(n_623),
.A2(n_379),
.B1(n_382),
.B2(n_383),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_L g842 ( 
.A(n_643),
.B(n_290),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_592),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_709),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_587),
.B(n_295),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_L g846 ( 
.A(n_589),
.B(n_296),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_SL g847 ( 
.A(n_708),
.B(n_300),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_600),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_625),
.B(n_556),
.Y(n_849)
);

INVx2_ASAP7_75t_SL g850 ( 
.A(n_720),
.Y(n_850)
);

NOR2xp33_ASAP7_75t_L g851 ( 
.A(n_623),
.B(n_302),
.Y(n_851)
);

AO221x1_ASAP7_75t_L g852 ( 
.A1(n_636),
.A2(n_569),
.B1(n_571),
.B2(n_517),
.C(n_513),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_625),
.B(n_556),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_711),
.Y(n_854)
);

OR2x2_ASAP7_75t_L g855 ( 
.A(n_647),
.B(n_666),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_708),
.B(n_305),
.Y(n_856)
);

AND2x6_ASAP7_75t_L g857 ( 
.A(n_703),
.B(n_711),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_600),
.Y(n_858)
);

INVxp67_ASAP7_75t_L g859 ( 
.A(n_661),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_625),
.B(n_693),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_642),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_606),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_606),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_642),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_713),
.B(n_556),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_713),
.B(n_556),
.Y(n_866)
);

INVx4_ASAP7_75t_L g867 ( 
.A(n_596),
.Y(n_867)
);

INVx4_ASAP7_75t_L g868 ( 
.A(n_596),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_L g869 ( 
.A(n_666),
.B(n_306),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_648),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_627),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_648),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_L g873 ( 
.A(n_647),
.B(n_314),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_627),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_671),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_671),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_631),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_631),
.Y(n_878)
);

AOI22x1_ASAP7_75t_L g879 ( 
.A1(n_636),
.A2(n_617),
.B1(n_672),
.B2(n_700),
.Y(n_879)
);

OAI21xp5_ASAP7_75t_L g880 ( 
.A1(n_708),
.A2(n_507),
.B(n_539),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_SL g881 ( 
.A(n_639),
.B(n_713),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_634),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_634),
.Y(n_883)
);

NAND3xp33_ASAP7_75t_L g884 ( 
.A(n_647),
.B(n_315),
.C(n_321),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_SL g885 ( 
.A(n_676),
.B(n_324),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_638),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_672),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_678),
.B(n_539),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_678),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_680),
.B(n_329),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_720),
.B(n_569),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_725),
.B(n_333),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_SL g893 ( 
.A(n_727),
.B(n_210),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_595),
.B(n_301),
.Y(n_894)
);

NOR3xp33_ASAP7_75t_L g895 ( 
.A(n_644),
.B(n_220),
.C(n_393),
.Y(n_895)
);

NOR3xp33_ASAP7_75t_L g896 ( 
.A(n_618),
.B(n_220),
.C(n_393),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_596),
.B(n_301),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_638),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_679),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_797),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_734),
.A2(n_619),
.B(n_598),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_735),
.A2(n_619),
.B(n_598),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_737),
.B(n_617),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_737),
.B(n_617),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_776),
.B(n_720),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_739),
.A2(n_619),
.B(n_598),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_776),
.B(n_636),
.Y(n_907)
);

BUFx3_ASAP7_75t_L g908 ( 
.A(n_791),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_741),
.A2(n_653),
.B(n_635),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_814),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_761),
.B(n_691),
.Y(n_911)
);

INVx3_ASAP7_75t_L g912 ( 
.A(n_786),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_761),
.B(n_694),
.Y(n_913)
);

NOR2xp67_ASAP7_75t_L g914 ( 
.A(n_821),
.B(n_569),
.Y(n_914)
);

AND2x2_ASAP7_75t_L g915 ( 
.A(n_791),
.B(n_647),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_880),
.A2(n_653),
.B(n_635),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_762),
.B(n_679),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_818),
.A2(n_653),
.B(n_635),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_762),
.B(n_695),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_SL g920 ( 
.A(n_795),
.B(n_596),
.Y(n_920)
);

A2O1A1Ixp33_ASAP7_75t_L g921 ( 
.A1(n_754),
.A2(n_719),
.B(n_718),
.C(n_640),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_763),
.B(n_695),
.Y(n_922)
);

BUFx6f_ASAP7_75t_L g923 ( 
.A(n_786),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_763),
.B(n_696),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_829),
.A2(n_704),
.B(n_596),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_L g926 ( 
.A(n_859),
.B(n_738),
.Y(n_926)
);

AOI22xp5_ASAP7_75t_L g927 ( 
.A1(n_827),
.A2(n_654),
.B1(n_718),
.B2(n_604),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_829),
.A2(n_704),
.B(n_692),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_790),
.B(n_696),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_829),
.A2(n_704),
.B(n_663),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_867),
.A2(n_704),
.B(n_652),
.Y(n_931)
);

HB1xp67_ASAP7_75t_L g932 ( 
.A(n_838),
.Y(n_932)
);

AND2x2_ASAP7_75t_L g933 ( 
.A(n_846),
.B(n_637),
.Y(n_933)
);

OAI21xp33_ASAP7_75t_L g934 ( 
.A1(n_842),
.A2(n_213),
.B(n_207),
.Y(n_934)
);

O2A1O1Ixp33_ASAP7_75t_L g935 ( 
.A1(n_733),
.A2(n_702),
.B(n_700),
.C(n_715),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_760),
.B(n_579),
.Y(n_936)
);

CKINVDCx8_ASAP7_75t_R g937 ( 
.A(n_833),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_SL g938 ( 
.A(n_833),
.B(n_579),
.Y(n_938)
);

AOI22xp5_ASAP7_75t_L g939 ( 
.A1(n_891),
.A2(n_654),
.B1(n_604),
.B2(n_586),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_797),
.Y(n_940)
);

INVx1_ASAP7_75t_SL g941 ( 
.A(n_753),
.Y(n_941)
);

AND2x4_ASAP7_75t_L g942 ( 
.A(n_729),
.B(n_673),
.Y(n_942)
);

BUFx12f_ASAP7_75t_L g943 ( 
.A(n_765),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_840),
.Y(n_944)
);

A2O1A1Ixp33_ASAP7_75t_L g945 ( 
.A1(n_830),
.A2(n_645),
.B(n_724),
.C(n_728),
.Y(n_945)
);

BUFx3_ASAP7_75t_L g946 ( 
.A(n_732),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_867),
.A2(n_704),
.B(n_649),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_881),
.B(n_637),
.Y(n_948)
);

NOR3xp33_ASAP7_75t_L g949 ( 
.A(n_773),
.B(n_243),
.C(n_218),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_751),
.B(n_213),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_790),
.B(n_654),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_729),
.B(n_586),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_867),
.A2(n_656),
.B(n_649),
.Y(n_953)
);

NAND2x1p5_ASAP7_75t_L g954 ( 
.A(n_748),
.B(n_585),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_796),
.B(n_654),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_796),
.B(n_654),
.Y(n_956)
);

A2O1A1Ixp33_ASAP7_75t_L g957 ( 
.A1(n_823),
.A2(n_569),
.B(n_571),
.C(n_499),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_814),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_868),
.A2(n_656),
.B(n_649),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_868),
.A2(n_656),
.B(n_649),
.Y(n_960)
);

OAI21xp5_ASAP7_75t_L g961 ( 
.A1(n_803),
.A2(n_654),
.B(n_699),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_868),
.A2(n_656),
.B(n_649),
.Y(n_962)
);

O2A1O1Ixp5_ASAP7_75t_L g963 ( 
.A1(n_893),
.A2(n_571),
.B(n_569),
.C(n_534),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_751),
.B(n_654),
.Y(n_964)
);

AOI22xp5_ASAP7_75t_L g965 ( 
.A1(n_891),
.A2(n_604),
.B1(n_716),
.B2(n_688),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_730),
.Y(n_966)
);

OR2x6_ASAP7_75t_L g967 ( 
.A(n_855),
.B(n_585),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_759),
.B(n_585),
.Y(n_968)
);

BUFx6f_ASAP7_75t_L g969 ( 
.A(n_785),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_L g970 ( 
.A(n_793),
.B(n_365),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_730),
.Y(n_971)
);

BUFx6f_ASAP7_75t_L g972 ( 
.A(n_785),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_L g973 ( 
.A(n_736),
.B(n_218),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_742),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_865),
.A2(n_866),
.B(n_860),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_819),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_759),
.B(n_585),
.Y(n_977)
);

HB1xp67_ASAP7_75t_L g978 ( 
.A(n_777),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_777),
.B(n_585),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_L g980 ( 
.A(n_745),
.B(n_223),
.Y(n_980)
);

AOI22x1_ASAP7_75t_L g981 ( 
.A1(n_788),
.A2(n_801),
.B1(n_808),
.B2(n_792),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_788),
.B(n_656),
.Y(n_982)
);

A2O1A1Ixp33_ASAP7_75t_L g983 ( 
.A1(n_748),
.A2(n_571),
.B(n_499),
.C(n_500),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_L g984 ( 
.A(n_869),
.B(n_223),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_748),
.A2(n_714),
.B(n_721),
.Y(n_985)
);

BUFx3_ASAP7_75t_L g986 ( 
.A(n_765),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_SL g987 ( 
.A(n_839),
.B(n_688),
.Y(n_987)
);

INVx4_ASAP7_75t_L g988 ( 
.A(n_729),
.Y(n_988)
);

A2O1A1Ixp33_ASAP7_75t_L g989 ( 
.A1(n_792),
.A2(n_571),
.B(n_513),
.C(n_517),
.Y(n_989)
);

AOI21xp33_ASAP7_75t_L g990 ( 
.A1(n_845),
.A2(n_229),
.B(n_388),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_819),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_742),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_L g993 ( 
.A(n_826),
.B(n_855),
.Y(n_993)
);

OAI22xp5_ASAP7_75t_L g994 ( 
.A1(n_801),
.A2(n_721),
.B1(n_714),
.B2(n_534),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_808),
.B(n_714),
.Y(n_995)
);

INVxp67_ASAP7_75t_L g996 ( 
.A(n_800),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_835),
.A2(n_714),
.B(n_721),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_778),
.A2(n_714),
.B(n_721),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_849),
.A2(n_721),
.B(n_549),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_853),
.A2(n_549),
.B(n_539),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_775),
.A2(n_549),
.B(n_539),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_811),
.B(n_782),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_820),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_811),
.B(n_604),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_L g1005 ( 
.A(n_767),
.B(n_771),
.Y(n_1005)
);

AND2x2_ASAP7_75t_L g1006 ( 
.A(n_774),
.B(n_229),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_813),
.A2(n_549),
.B(n_539),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_820),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_798),
.B(n_604),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_746),
.A2(n_549),
.B(n_548),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_750),
.A2(n_549),
.B(n_548),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_824),
.Y(n_1012)
);

O2A1O1Ixp33_ASAP7_75t_L g1013 ( 
.A1(n_787),
.A2(n_548),
.B(n_558),
.C(n_561),
.Y(n_1013)
);

BUFx2_ASAP7_75t_L g1014 ( 
.A(n_765),
.Y(n_1014)
);

OAI22xp5_ASAP7_75t_L g1015 ( 
.A1(n_807),
.A2(n_380),
.B1(n_240),
.B2(n_241),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_756),
.A2(n_549),
.B(n_548),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_757),
.Y(n_1017)
);

INVxp67_ASAP7_75t_L g1018 ( 
.A(n_805),
.Y(n_1018)
);

NAND2x1p5_ASAP7_75t_L g1019 ( 
.A(n_744),
.B(n_548),
.Y(n_1019)
);

BUFx3_ASAP7_75t_L g1020 ( 
.A(n_840),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_766),
.A2(n_549),
.B(n_716),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_757),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_772),
.A2(n_549),
.B(n_716),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_812),
.B(n_604),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_824),
.B(n_828),
.Y(n_1025)
);

INVx3_ASAP7_75t_L g1026 ( 
.A(n_784),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_779),
.A2(n_688),
.B(n_508),
.Y(n_1027)
);

OR2x2_ASAP7_75t_L g1028 ( 
.A(n_743),
.B(n_238),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_781),
.A2(n_503),
.B(n_508),
.Y(n_1029)
);

A2O1A1Ixp33_ASAP7_75t_L g1030 ( 
.A1(n_851),
.A2(n_558),
.B(n_561),
.C(n_238),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_873),
.B(n_240),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_794),
.A2(n_508),
.B(n_511),
.Y(n_1032)
);

AND2x4_ASAP7_75t_L g1033 ( 
.A(n_850),
.B(n_707),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_806),
.A2(n_511),
.B(n_518),
.Y(n_1034)
);

OAI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_799),
.A2(n_699),
.B(n_528),
.Y(n_1035)
);

NAND2xp33_ASAP7_75t_L g1036 ( 
.A(n_839),
.B(n_301),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_SL g1037 ( 
.A(n_839),
.B(n_301),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_802),
.A2(n_511),
.B(n_518),
.Y(n_1038)
);

AOI21xp33_ASAP7_75t_L g1039 ( 
.A1(n_731),
.A2(n_241),
.B(n_243),
.Y(n_1039)
);

O2A1O1Ixp33_ASAP7_75t_L g1040 ( 
.A1(n_894),
.A2(n_558),
.B(n_561),
.C(n_527),
.Y(n_1040)
);

AND2x4_ASAP7_75t_L g1041 ( 
.A(n_850),
.B(n_558),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_828),
.B(n_699),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_834),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_749),
.A2(n_508),
.B(n_511),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_SL g1045 ( 
.A(n_839),
.B(n_301),
.Y(n_1045)
);

INVx4_ASAP7_75t_L g1046 ( 
.A(n_857),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_L g1047 ( 
.A(n_789),
.B(n_334),
.Y(n_1047)
);

BUFx6f_ASAP7_75t_L g1048 ( 
.A(n_857),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_834),
.B(n_699),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_844),
.B(n_699),
.Y(n_1050)
);

NOR2xp33_ASAP7_75t_L g1051 ( 
.A(n_773),
.B(n_334),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_844),
.B(n_699),
.Y(n_1052)
);

NOR2xp33_ASAP7_75t_SL g1053 ( 
.A(n_769),
.B(n_335),
.Y(n_1053)
);

INVx3_ASAP7_75t_L g1054 ( 
.A(n_784),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_L g1055 ( 
.A(n_783),
.B(n_335),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_749),
.A2(n_508),
.B(n_530),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_SL g1057 ( 
.A(n_839),
.B(n_301),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_847),
.A2(n_508),
.B(n_530),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_854),
.B(n_699),
.Y(n_1059)
);

INVxp67_ASAP7_75t_L g1060 ( 
.A(n_831),
.Y(n_1060)
);

OAI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_857),
.A2(n_514),
.B(n_528),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_854),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_856),
.A2(n_530),
.B(n_511),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_888),
.A2(n_530),
.B(n_511),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_744),
.B(n_520),
.Y(n_1065)
);

OAI21xp33_ASAP7_75t_L g1066 ( 
.A1(n_896),
.A2(n_370),
.B(n_340),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_897),
.A2(n_530),
.B(n_511),
.Y(n_1067)
);

AOI22xp33_ASAP7_75t_L g1068 ( 
.A1(n_740),
.A2(n_301),
.B1(n_381),
.B2(n_380),
.Y(n_1068)
);

AOI22xp33_ASAP7_75t_L g1069 ( 
.A1(n_740),
.A2(n_301),
.B1(n_381),
.B2(n_375),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_861),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_804),
.A2(n_530),
.B(n_511),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_804),
.A2(n_530),
.B(n_518),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_899),
.A2(n_530),
.B(n_518),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_899),
.A2(n_508),
.B(n_518),
.Y(n_1074)
);

AO21x1_ASAP7_75t_L g1075 ( 
.A1(n_822),
.A2(n_528),
.B(n_527),
.Y(n_1075)
);

O2A1O1Ixp33_ASAP7_75t_L g1076 ( 
.A1(n_755),
.A2(n_768),
.B(n_780),
.C(n_770),
.Y(n_1076)
);

HB1xp67_ASAP7_75t_L g1077 ( 
.A(n_764),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_758),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_861),
.A2(n_519),
.B(n_518),
.Y(n_1079)
);

INVx3_ASAP7_75t_L g1080 ( 
.A(n_898),
.Y(n_1080)
);

OAI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_857),
.A2(n_527),
.B(n_526),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_864),
.A2(n_519),
.B(n_518),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_864),
.B(n_520),
.Y(n_1083)
);

A2O1A1Ixp33_ASAP7_75t_L g1084 ( 
.A1(n_884),
.A2(n_370),
.B(n_340),
.C(n_341),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_870),
.A2(n_519),
.B(n_518),
.Y(n_1085)
);

O2A1O1Ixp33_ASAP7_75t_L g1086 ( 
.A1(n_892),
.A2(n_527),
.B(n_526),
.C(n_525),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_816),
.Y(n_1087)
);

AOI22xp5_ASAP7_75t_L g1088 ( 
.A1(n_857),
.A2(n_520),
.B1(n_526),
.B2(n_525),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_870),
.B(n_872),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_872),
.B(n_520),
.Y(n_1090)
);

BUFx4f_ASAP7_75t_L g1091 ( 
.A(n_857),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_916),
.A2(n_1036),
.B(n_975),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_976),
.Y(n_1093)
);

OAI21xp33_ASAP7_75t_L g1094 ( 
.A1(n_984),
.A2(n_895),
.B(n_752),
.Y(n_1094)
);

O2A1O1Ixp33_ASAP7_75t_L g1095 ( 
.A1(n_984),
.A2(n_815),
.B(n_810),
.C(n_841),
.Y(n_1095)
);

OAI22xp5_ASAP7_75t_SL g1096 ( 
.A1(n_970),
.A2(n_341),
.B1(n_388),
.B2(n_386),
.Y(n_1096)
);

INVx3_ASAP7_75t_L g1097 ( 
.A(n_923),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_1026),
.Y(n_1098)
);

OR2x6_ASAP7_75t_SL g1099 ( 
.A(n_944),
.B(n_345),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_991),
.Y(n_1100)
);

INVx3_ASAP7_75t_L g1101 ( 
.A(n_923),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_1054),
.Y(n_1102)
);

AND2x4_ASAP7_75t_L g1103 ( 
.A(n_988),
.B(n_747),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_1002),
.A2(n_839),
.B(n_889),
.Y(n_1104)
);

AND2x2_ASAP7_75t_L g1105 ( 
.A(n_970),
.B(n_885),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_901),
.A2(n_839),
.B(n_889),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_937),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_902),
.A2(n_909),
.B(n_906),
.Y(n_1108)
);

A2O1A1Ixp33_ASAP7_75t_SL g1109 ( 
.A1(n_926),
.A2(n_832),
.B(n_836),
.C(n_887),
.Y(n_1109)
);

A2O1A1Ixp33_ASAP7_75t_L g1110 ( 
.A1(n_926),
.A2(n_890),
.B(n_875),
.C(n_887),
.Y(n_1110)
);

NOR2xp33_ASAP7_75t_L g1111 ( 
.A(n_996),
.B(n_809),
.Y(n_1111)
);

NOR2xp33_ASAP7_75t_L g1112 ( 
.A(n_996),
.B(n_837),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_978),
.B(n_852),
.Y(n_1113)
);

INVx1_ASAP7_75t_SL g1114 ( 
.A(n_941),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_978),
.B(n_852),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_1054),
.Y(n_1116)
);

OR2x2_ASAP7_75t_L g1117 ( 
.A(n_1028),
.B(n_875),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_1018),
.B(n_879),
.Y(n_1118)
);

A2O1A1Ixp33_ASAP7_75t_L g1119 ( 
.A1(n_1076),
.A2(n_876),
.B(n_886),
.C(n_883),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_1003),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1008),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_1018),
.B(n_879),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_987),
.A2(n_839),
.B(n_876),
.Y(n_1123)
);

INVx5_ASAP7_75t_L g1124 ( 
.A(n_1048),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_1005),
.B(n_816),
.Y(n_1125)
);

OAI21xp33_ASAP7_75t_L g1126 ( 
.A1(n_934),
.A2(n_351),
.B(n_355),
.Y(n_1126)
);

BUFx6f_ASAP7_75t_SL g1127 ( 
.A(n_1020),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1012),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1043),
.Y(n_1129)
);

AOI22xp5_ASAP7_75t_L g1130 ( 
.A1(n_993),
.A2(n_898),
.B1(n_886),
.B2(n_883),
.Y(n_1130)
);

INVx3_ASAP7_75t_L g1131 ( 
.A(n_923),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_987),
.A2(n_882),
.B(n_878),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_SL g1133 ( 
.A(n_988),
.B(n_817),
.Y(n_1133)
);

NOR2xp33_ASAP7_75t_R g1134 ( 
.A(n_1078),
.B(n_938),
.Y(n_1134)
);

NOR3xp33_ASAP7_75t_L g1135 ( 
.A(n_990),
.B(n_386),
.C(n_345),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_SL g1136 ( 
.A(n_923),
.B(n_817),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_943),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_918),
.A2(n_882),
.B(n_878),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_998),
.A2(n_877),
.B(n_874),
.Y(n_1139)
);

BUFx6f_ASAP7_75t_L g1140 ( 
.A(n_967),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_1027),
.A2(n_877),
.B(n_874),
.Y(n_1141)
);

HB1xp67_ASAP7_75t_L g1142 ( 
.A(n_908),
.Y(n_1142)
);

OAI22xp5_ASAP7_75t_L g1143 ( 
.A1(n_912),
.A2(n_863),
.B1(n_862),
.B2(n_858),
.Y(n_1143)
);

OAI22xp5_ASAP7_75t_SL g1144 ( 
.A1(n_936),
.A2(n_369),
.B1(n_351),
.B2(n_355),
.Y(n_1144)
);

NAND3xp33_ASAP7_75t_SL g1145 ( 
.A(n_1053),
.B(n_374),
.C(n_358),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_SL g1146 ( 
.A(n_915),
.B(n_825),
.Y(n_1146)
);

O2A1O1Ixp33_ASAP7_75t_L g1147 ( 
.A1(n_1051),
.A2(n_871),
.B(n_863),
.C(n_862),
.Y(n_1147)
);

AOI22xp33_ASAP7_75t_L g1148 ( 
.A1(n_949),
.A2(n_871),
.B1(n_858),
.B2(n_848),
.Y(n_1148)
);

AOI22xp5_ASAP7_75t_L g1149 ( 
.A1(n_993),
.A2(n_848),
.B1(n_843),
.B2(n_825),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1062),
.Y(n_1150)
);

A2O1A1Ixp33_ASAP7_75t_L g1151 ( 
.A1(n_1051),
.A2(n_843),
.B(n_371),
.C(n_369),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1005),
.B(n_358),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_968),
.A2(n_519),
.B(n_508),
.Y(n_1153)
);

INVx2_ASAP7_75t_SL g1154 ( 
.A(n_946),
.Y(n_1154)
);

NOR2xp33_ASAP7_75t_SL g1155 ( 
.A(n_933),
.B(n_359),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_1080),
.Y(n_1156)
);

AOI22xp33_ASAP7_75t_L g1157 ( 
.A1(n_949),
.A2(n_371),
.B1(n_366),
.B2(n_359),
.Y(n_1157)
);

AOI33xp33_ASAP7_75t_L g1158 ( 
.A1(n_950),
.A2(n_361),
.A3(n_364),
.B1(n_366),
.B2(n_367),
.B3(n_374),
.Y(n_1158)
);

AO32x1_ASAP7_75t_L g1159 ( 
.A1(n_994),
.A2(n_514),
.A3(n_525),
.B1(n_271),
.B2(n_20),
.Y(n_1159)
);

O2A1O1Ixp33_ASAP7_75t_L g1160 ( 
.A1(n_1077),
.A2(n_525),
.B(n_514),
.C(n_520),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_914),
.B(n_361),
.Y(n_1161)
);

OAI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_921),
.A2(n_514),
.B(n_364),
.Y(n_1162)
);

NAND2xp33_ASAP7_75t_L g1163 ( 
.A(n_1048),
.B(n_375),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_977),
.A2(n_519),
.B(n_367),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_979),
.A2(n_519),
.B(n_78),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_964),
.A2(n_519),
.B(n_79),
.Y(n_1166)
);

INVx4_ASAP7_75t_L g1167 ( 
.A(n_912),
.Y(n_1167)
);

O2A1O1Ixp33_ASAP7_75t_L g1168 ( 
.A1(n_1077),
.A2(n_13),
.B(n_14),
.C(n_18),
.Y(n_1168)
);

O2A1O1Ixp33_ASAP7_75t_L g1169 ( 
.A1(n_1084),
.A2(n_13),
.B(n_18),
.C(n_20),
.Y(n_1169)
);

OAI21xp33_ASAP7_75t_L g1170 ( 
.A1(n_973),
.A2(n_22),
.B(n_23),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_1025),
.A2(n_519),
.B(n_90),
.Y(n_1171)
);

NOR2xp33_ASAP7_75t_L g1172 ( 
.A(n_936),
.B(n_932),
.Y(n_1172)
);

O2A1O1Ixp5_ASAP7_75t_L g1173 ( 
.A1(n_1075),
.A2(n_87),
.B(n_191),
.C(n_186),
.Y(n_1173)
);

NOR2xp33_ASAP7_75t_L g1174 ( 
.A(n_932),
.B(n_22),
.Y(n_1174)
);

O2A1O1Ixp33_ASAP7_75t_L g1175 ( 
.A1(n_1039),
.A2(n_24),
.B(n_27),
.C(n_30),
.Y(n_1175)
);

AND2x2_ASAP7_75t_L g1176 ( 
.A(n_1031),
.B(n_24),
.Y(n_1176)
);

OAI21xp33_ASAP7_75t_L g1177 ( 
.A1(n_973),
.A2(n_30),
.B(n_32),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_900),
.B(n_33),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_1080),
.Y(n_1179)
);

AOI33xp33_ASAP7_75t_L g1180 ( 
.A1(n_1006),
.A2(n_33),
.A3(n_34),
.B1(n_36),
.B2(n_37),
.B3(n_41),
.Y(n_1180)
);

O2A1O1Ixp33_ASAP7_75t_L g1181 ( 
.A1(n_1030),
.A2(n_34),
.B(n_41),
.C(n_45),
.Y(n_1181)
);

AOI22xp33_ASAP7_75t_L g1182 ( 
.A1(n_1047),
.A2(n_45),
.B1(n_46),
.B2(n_49),
.Y(n_1182)
);

NOR2x1_ASAP7_75t_L g1183 ( 
.A(n_986),
.B(n_106),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_940),
.B(n_46),
.Y(n_1184)
);

OAI22xp5_ASAP7_75t_L g1185 ( 
.A1(n_911),
.A2(n_111),
.B1(n_178),
.B2(n_176),
.Y(n_1185)
);

OAI22xp5_ASAP7_75t_L g1186 ( 
.A1(n_913),
.A2(n_100),
.B1(n_168),
.B2(n_164),
.Y(n_1186)
);

AOI22xp33_ASAP7_75t_L g1187 ( 
.A1(n_1047),
.A2(n_49),
.B1(n_52),
.B2(n_53),
.Y(n_1187)
);

NOR2xp33_ASAP7_75t_L g1188 ( 
.A(n_1060),
.B(n_53),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_905),
.B(n_55),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_910),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_958),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_903),
.B(n_55),
.Y(n_1192)
);

AND2x2_ASAP7_75t_SL g1193 ( 
.A(n_1014),
.B(n_59),
.Y(n_1193)
);

AND2x2_ASAP7_75t_L g1194 ( 
.A(n_980),
.B(n_60),
.Y(n_1194)
);

AND2x2_ASAP7_75t_L g1195 ( 
.A(n_980),
.B(n_69),
.Y(n_1195)
);

INVx4_ASAP7_75t_L g1196 ( 
.A(n_967),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_SL g1197 ( 
.A(n_1060),
.B(n_125),
.Y(n_1197)
);

AOI21xp33_ASAP7_75t_L g1198 ( 
.A1(n_1055),
.A2(n_70),
.B(n_71),
.Y(n_1198)
);

A2O1A1Ixp33_ASAP7_75t_SL g1199 ( 
.A1(n_1055),
.A2(n_132),
.B(n_160),
.C(n_159),
.Y(n_1199)
);

NOR3xp33_ASAP7_75t_L g1200 ( 
.A(n_948),
.B(n_1066),
.C(n_1015),
.Y(n_1200)
);

HB1xp67_ASAP7_75t_L g1201 ( 
.A(n_967),
.Y(n_1201)
);

INVxp67_ASAP7_75t_L g1202 ( 
.A(n_948),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_904),
.B(n_70),
.Y(n_1203)
);

NOR2xp33_ASAP7_75t_L g1204 ( 
.A(n_907),
.B(n_71),
.Y(n_1204)
);

AOI22xp5_ASAP7_75t_L g1205 ( 
.A1(n_952),
.A2(n_112),
.B1(n_80),
.B2(n_94),
.Y(n_1205)
);

INVx3_ASAP7_75t_L g1206 ( 
.A(n_969),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_951),
.A2(n_141),
.B(n_95),
.Y(n_1207)
);

A2O1A1Ixp33_ASAP7_75t_L g1208 ( 
.A1(n_945),
.A2(n_75),
.B(n_105),
.C(n_140),
.Y(n_1208)
);

CKINVDCx16_ASAP7_75t_R g1209 ( 
.A(n_942),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_SL g1210 ( 
.A(n_942),
.B(n_146),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1070),
.B(n_152),
.Y(n_1211)
);

AO32x1_ASAP7_75t_L g1212 ( 
.A1(n_1046),
.A2(n_1022),
.A3(n_974),
.B1(n_992),
.B2(n_966),
.Y(n_1212)
);

OAI22xp5_ASAP7_75t_L g1213 ( 
.A1(n_927),
.A2(n_197),
.B1(n_1091),
.B2(n_1046),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_1087),
.Y(n_1214)
);

O2A1O1Ixp33_ASAP7_75t_L g1215 ( 
.A1(n_957),
.A2(n_989),
.B(n_983),
.C(n_920),
.Y(n_1215)
);

OAI22xp5_ASAP7_75t_L g1216 ( 
.A1(n_1091),
.A2(n_972),
.B1(n_969),
.B2(n_965),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_971),
.Y(n_1217)
);

OAI22xp5_ASAP7_75t_L g1218 ( 
.A1(n_969),
.A2(n_972),
.B1(n_954),
.B2(n_939),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_969),
.B(n_972),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_972),
.B(n_1041),
.Y(n_1220)
);

OAI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_954),
.A2(n_1009),
.B1(n_1024),
.B2(n_1069),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_SL g1222 ( 
.A(n_1033),
.B(n_1041),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_955),
.A2(n_956),
.B(n_995),
.Y(n_1223)
);

BUFx6f_ASAP7_75t_L g1224 ( 
.A(n_1048),
.Y(n_1224)
);

CKINVDCx14_ASAP7_75t_R g1225 ( 
.A(n_1033),
.Y(n_1225)
);

BUFx2_ASAP7_75t_L g1226 ( 
.A(n_1048),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1017),
.B(n_1089),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_982),
.A2(n_961),
.B(n_985),
.Y(n_1228)
);

INVxp67_ASAP7_75t_SL g1229 ( 
.A(n_1019),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_1088),
.Y(n_1230)
);

INVx4_ASAP7_75t_L g1231 ( 
.A(n_1019),
.Y(n_1231)
);

A2O1A1Ixp33_ASAP7_75t_L g1232 ( 
.A1(n_1068),
.A2(n_1069),
.B(n_935),
.C(n_1042),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_917),
.Y(n_1233)
);

INVx4_ASAP7_75t_L g1234 ( 
.A(n_981),
.Y(n_1234)
);

BUFx12f_ASAP7_75t_L g1235 ( 
.A(n_1086),
.Y(n_1235)
);

BUFx6f_ASAP7_75t_L g1236 ( 
.A(n_919),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_922),
.Y(n_1237)
);

OAI22xp5_ASAP7_75t_L g1238 ( 
.A1(n_1068),
.A2(n_924),
.B1(n_929),
.B2(n_1004),
.Y(n_1238)
);

AOI221xp5_ASAP7_75t_L g1239 ( 
.A1(n_1013),
.A2(n_1049),
.B1(n_1059),
.B2(n_1050),
.C(n_1052),
.Y(n_1239)
);

BUFx6f_ASAP7_75t_L g1240 ( 
.A(n_1083),
.Y(n_1240)
);

O2A1O1Ixp33_ASAP7_75t_L g1241 ( 
.A1(n_1037),
.A2(n_1045),
.B(n_963),
.C(n_1090),
.Y(n_1241)
);

OAI22xp5_ASAP7_75t_L g1242 ( 
.A1(n_928),
.A2(n_930),
.B1(n_1065),
.B2(n_931),
.Y(n_1242)
);

A2O1A1Ixp33_ASAP7_75t_SL g1243 ( 
.A1(n_1061),
.A2(n_1081),
.B(n_1035),
.C(n_1040),
.Y(n_1243)
);

NOR2xp33_ASAP7_75t_L g1244 ( 
.A(n_1037),
.B(n_1045),
.Y(n_1244)
);

CKINVDCx11_ASAP7_75t_R g1245 ( 
.A(n_963),
.Y(n_1245)
);

AOI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_997),
.A2(n_1057),
.B(n_1023),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1085),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_1001),
.Y(n_1248)
);

INVx1_ASAP7_75t_SL g1249 ( 
.A(n_1079),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_1038),
.Y(n_1250)
);

NOR2xp33_ASAP7_75t_R g1251 ( 
.A(n_1007),
.B(n_1072),
.Y(n_1251)
);

A2O1A1Ixp33_ASAP7_75t_L g1252 ( 
.A1(n_1021),
.A2(n_1056),
.B(n_1044),
.C(n_1010),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1029),
.B(n_1032),
.Y(n_1253)
);

BUFx6f_ASAP7_75t_L g1254 ( 
.A(n_1140),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1105),
.B(n_1233),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1237),
.B(n_1111),
.Y(n_1256)
);

NOR4xp25_ASAP7_75t_L g1257 ( 
.A(n_1170),
.B(n_1034),
.C(n_1082),
.D(n_1016),
.Y(n_1257)
);

OAI21x1_ASAP7_75t_L g1258 ( 
.A1(n_1132),
.A2(n_1058),
.B(n_1063),
.Y(n_1258)
);

AO32x2_ASAP7_75t_L g1259 ( 
.A1(n_1238),
.A2(n_1064),
.A3(n_1071),
.B1(n_1011),
.B2(n_1000),
.Y(n_1259)
);

NOR2xp33_ASAP7_75t_L g1260 ( 
.A(n_1202),
.B(n_1074),
.Y(n_1260)
);

OAI21x1_ASAP7_75t_L g1261 ( 
.A1(n_1132),
.A2(n_999),
.B(n_960),
.Y(n_1261)
);

OAI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1244),
.A2(n_925),
.B(n_1067),
.Y(n_1262)
);

AOI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1092),
.A2(n_953),
.B(n_959),
.Y(n_1263)
);

INVxp67_ASAP7_75t_L g1264 ( 
.A(n_1114),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1112),
.B(n_1073),
.Y(n_1265)
);

AO32x2_ASAP7_75t_L g1266 ( 
.A1(n_1234),
.A2(n_947),
.A3(n_962),
.B1(n_1221),
.B2(n_1242),
.Y(n_1266)
);

OAI22xp5_ASAP7_75t_L g1267 ( 
.A1(n_1230),
.A2(n_1172),
.B1(n_1125),
.B2(n_1117),
.Y(n_1267)
);

BUFx12f_ASAP7_75t_L g1268 ( 
.A(n_1137),
.Y(n_1268)
);

BUFx6f_ASAP7_75t_L g1269 ( 
.A(n_1140),
.Y(n_1269)
);

OAI21x1_ASAP7_75t_L g1270 ( 
.A1(n_1139),
.A2(n_1138),
.B(n_1141),
.Y(n_1270)
);

O2A1O1Ixp33_ASAP7_75t_SL g1271 ( 
.A1(n_1208),
.A2(n_1118),
.B(n_1122),
.C(n_1197),
.Y(n_1271)
);

O2A1O1Ixp33_ASAP7_75t_L g1272 ( 
.A1(n_1094),
.A2(n_1095),
.B(n_1200),
.C(n_1198),
.Y(n_1272)
);

NOR2xp33_ASAP7_75t_L g1273 ( 
.A(n_1155),
.B(n_1152),
.Y(n_1273)
);

INVx3_ASAP7_75t_L g1274 ( 
.A(n_1167),
.Y(n_1274)
);

AOI22xp5_ASAP7_75t_L g1275 ( 
.A1(n_1194),
.A2(n_1195),
.B1(n_1210),
.B2(n_1145),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1093),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1176),
.B(n_1204),
.Y(n_1277)
);

OR2x6_ASAP7_75t_L g1278 ( 
.A(n_1154),
.B(n_1140),
.Y(n_1278)
);

AOI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1092),
.A2(n_1108),
.B(n_1253),
.Y(n_1279)
);

INVx3_ASAP7_75t_SL g1280 ( 
.A(n_1107),
.Y(n_1280)
);

CKINVDCx11_ASAP7_75t_R g1281 ( 
.A(n_1099),
.Y(n_1281)
);

AO31x2_ASAP7_75t_L g1282 ( 
.A1(n_1234),
.A2(n_1252),
.A3(n_1108),
.B(n_1232),
.Y(n_1282)
);

A2O1A1Ixp33_ASAP7_75t_L g1283 ( 
.A1(n_1177),
.A2(n_1151),
.B(n_1188),
.C(n_1110),
.Y(n_1283)
);

AO21x2_ASAP7_75t_L g1284 ( 
.A1(n_1228),
.A2(n_1106),
.B(n_1246),
.Y(n_1284)
);

AO21x2_ASAP7_75t_L g1285 ( 
.A1(n_1228),
.A2(n_1106),
.B(n_1246),
.Y(n_1285)
);

CKINVDCx6p67_ASAP7_75t_R g1286 ( 
.A(n_1127),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1100),
.B(n_1120),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_1134),
.Y(n_1288)
);

NOR2xp33_ASAP7_75t_L g1289 ( 
.A(n_1222),
.B(n_1142),
.Y(n_1289)
);

AND2x4_ASAP7_75t_L g1290 ( 
.A(n_1196),
.B(n_1201),
.Y(n_1290)
);

AND2x4_ASAP7_75t_L g1291 ( 
.A(n_1196),
.B(n_1103),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_SL g1292 ( 
.A(n_1209),
.B(n_1236),
.Y(n_1292)
);

OR2x2_ASAP7_75t_L g1293 ( 
.A(n_1161),
.B(n_1189),
.Y(n_1293)
);

OAI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_1223),
.A2(n_1164),
.B(n_1162),
.Y(n_1294)
);

OAI21x1_ASAP7_75t_L g1295 ( 
.A1(n_1139),
.A2(n_1138),
.B(n_1141),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1121),
.B(n_1128),
.Y(n_1296)
);

BUFx10_ASAP7_75t_L g1297 ( 
.A(n_1127),
.Y(n_1297)
);

A2O1A1Ixp33_ASAP7_75t_L g1298 ( 
.A1(n_1215),
.A2(n_1181),
.B(n_1175),
.C(n_1169),
.Y(n_1298)
);

AO21x2_ASAP7_75t_L g1299 ( 
.A1(n_1104),
.A2(n_1251),
.B(n_1166),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1129),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1150),
.Y(n_1301)
);

AOI22xp5_ASAP7_75t_L g1302 ( 
.A1(n_1096),
.A2(n_1103),
.B1(n_1135),
.B2(n_1144),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1214),
.Y(n_1303)
);

AOI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1243),
.A2(n_1223),
.B(n_1123),
.Y(n_1304)
);

AO31x2_ASAP7_75t_L g1305 ( 
.A1(n_1166),
.A2(n_1165),
.A3(n_1119),
.B(n_1171),
.Y(n_1305)
);

AOI21xp5_ASAP7_75t_L g1306 ( 
.A1(n_1123),
.A2(n_1109),
.B(n_1241),
.Y(n_1306)
);

AOI21xp5_ASAP7_75t_L g1307 ( 
.A1(n_1249),
.A2(n_1250),
.B(n_1216),
.Y(n_1307)
);

INVx2_ASAP7_75t_L g1308 ( 
.A(n_1190),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1227),
.B(n_1236),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1217),
.Y(n_1310)
);

O2A1O1Ixp33_ASAP7_75t_L g1311 ( 
.A1(n_1168),
.A2(n_1181),
.B(n_1178),
.C(n_1184),
.Y(n_1311)
);

OAI21xp5_ASAP7_75t_L g1312 ( 
.A1(n_1164),
.A2(n_1203),
.B(n_1192),
.Y(n_1312)
);

A2O1A1Ixp33_ASAP7_75t_L g1313 ( 
.A1(n_1171),
.A2(n_1126),
.B(n_1165),
.C(n_1147),
.Y(n_1313)
);

CKINVDCx6p67_ASAP7_75t_R g1314 ( 
.A(n_1124),
.Y(n_1314)
);

A2O1A1Ixp33_ASAP7_75t_L g1315 ( 
.A1(n_1211),
.A2(n_1160),
.B(n_1207),
.C(n_1213),
.Y(n_1315)
);

AO32x2_ASAP7_75t_L g1316 ( 
.A1(n_1218),
.A2(n_1143),
.A3(n_1185),
.B1(n_1186),
.B2(n_1159),
.Y(n_1316)
);

AO32x2_ASAP7_75t_L g1317 ( 
.A1(n_1159),
.A2(n_1212),
.A3(n_1180),
.B1(n_1231),
.B2(n_1245),
.Y(n_1317)
);

AOI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1247),
.A2(n_1229),
.B(n_1219),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1236),
.B(n_1220),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1191),
.Y(n_1320)
);

O2A1O1Ixp33_ASAP7_75t_L g1321 ( 
.A1(n_1199),
.A2(n_1174),
.B(n_1163),
.C(n_1115),
.Y(n_1321)
);

AO31x2_ASAP7_75t_L g1322 ( 
.A1(n_1113),
.A2(n_1207),
.A3(n_1153),
.B(n_1212),
.Y(n_1322)
);

OAI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1239),
.A2(n_1148),
.B(n_1146),
.Y(n_1323)
);

AOI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1248),
.A2(n_1239),
.B(n_1212),
.Y(n_1324)
);

OAI21x1_ASAP7_75t_L g1325 ( 
.A1(n_1153),
.A2(n_1173),
.B(n_1136),
.Y(n_1325)
);

O2A1O1Ixp33_ASAP7_75t_SL g1326 ( 
.A1(n_1133),
.A2(n_1205),
.B(n_1098),
.C(n_1179),
.Y(n_1326)
);

AOI221x1_ASAP7_75t_L g1327 ( 
.A1(n_1240),
.A2(n_1159),
.B1(n_1206),
.B2(n_1224),
.C(n_1102),
.Y(n_1327)
);

O2A1O1Ixp33_ASAP7_75t_L g1328 ( 
.A1(n_1182),
.A2(n_1187),
.B(n_1157),
.C(n_1225),
.Y(n_1328)
);

NOR2xp33_ASAP7_75t_L g1329 ( 
.A(n_1193),
.B(n_1240),
.Y(n_1329)
);

OAI21x1_ASAP7_75t_L g1330 ( 
.A1(n_1130),
.A2(n_1149),
.B(n_1206),
.Y(n_1330)
);

AOI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1240),
.A2(n_1124),
.B(n_1226),
.Y(n_1331)
);

BUFx3_ASAP7_75t_L g1332 ( 
.A(n_1097),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1158),
.B(n_1097),
.Y(n_1333)
);

O2A1O1Ixp33_ASAP7_75t_SL g1334 ( 
.A1(n_1116),
.A2(n_1156),
.B(n_1131),
.C(n_1101),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_1101),
.Y(n_1335)
);

AOI21xp5_ASAP7_75t_L g1336 ( 
.A1(n_1124),
.A2(n_1131),
.B(n_1224),
.Y(n_1336)
);

AOI21x1_ASAP7_75t_L g1337 ( 
.A1(n_1183),
.A2(n_1235),
.B(n_1124),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1224),
.Y(n_1338)
);

AND2x4_ASAP7_75t_L g1339 ( 
.A(n_1222),
.B(n_988),
.Y(n_1339)
);

INVx5_ASAP7_75t_L g1340 ( 
.A(n_1140),
.Y(n_1340)
);

AO31x2_ASAP7_75t_L g1341 ( 
.A1(n_1092),
.A2(n_1234),
.A3(n_1252),
.B(n_1108),
.Y(n_1341)
);

AOI21xp33_ASAP7_75t_L g1342 ( 
.A1(n_1095),
.A2(n_970),
.B(n_984),
.Y(n_1342)
);

AOI21xp5_ASAP7_75t_L g1343 ( 
.A1(n_1092),
.A2(n_708),
.B(n_1036),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1202),
.B(n_1031),
.Y(n_1344)
);

AOI21xp5_ASAP7_75t_L g1345 ( 
.A1(n_1092),
.A2(n_708),
.B(n_1036),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1202),
.B(n_1031),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1105),
.B(n_926),
.Y(n_1347)
);

INVx4_ASAP7_75t_L g1348 ( 
.A(n_1140),
.Y(n_1348)
);

AOI21xp5_ASAP7_75t_L g1349 ( 
.A1(n_1092),
.A2(n_708),
.B(n_1036),
.Y(n_1349)
);

CKINVDCx6p67_ASAP7_75t_R g1350 ( 
.A(n_1127),
.Y(n_1350)
);

AOI21xp5_ASAP7_75t_L g1351 ( 
.A1(n_1092),
.A2(n_708),
.B(n_1036),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1105),
.B(n_926),
.Y(n_1352)
);

AOI21xp5_ASAP7_75t_L g1353 ( 
.A1(n_1092),
.A2(n_708),
.B(n_1036),
.Y(n_1353)
);

INVxp67_ASAP7_75t_L g1354 ( 
.A(n_1114),
.Y(n_1354)
);

AO31x2_ASAP7_75t_L g1355 ( 
.A1(n_1092),
.A2(n_1234),
.A3(n_1252),
.B(n_1108),
.Y(n_1355)
);

AND2x6_ASAP7_75t_L g1356 ( 
.A(n_1224),
.B(n_1048),
.Y(n_1356)
);

OAI22x1_ASAP7_75t_L g1357 ( 
.A1(n_1194),
.A2(n_618),
.B1(n_970),
.B2(n_740),
.Y(n_1357)
);

OAI21x1_ASAP7_75t_L g1358 ( 
.A1(n_1132),
.A2(n_1139),
.B(n_1138),
.Y(n_1358)
);

CKINVDCx5p33_ASAP7_75t_R g1359 ( 
.A(n_1107),
.Y(n_1359)
);

OAI21x1_ASAP7_75t_L g1360 ( 
.A1(n_1132),
.A2(n_1139),
.B(n_1138),
.Y(n_1360)
);

BUFx2_ASAP7_75t_L g1361 ( 
.A(n_1142),
.Y(n_1361)
);

INVx3_ASAP7_75t_L g1362 ( 
.A(n_1167),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_SL g1363 ( 
.A(n_1172),
.B(n_589),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1202),
.B(n_1031),
.Y(n_1364)
);

INVxp67_ASAP7_75t_L g1365 ( 
.A(n_1114),
.Y(n_1365)
);

AO31x2_ASAP7_75t_L g1366 ( 
.A1(n_1092),
.A2(n_1234),
.A3(n_1252),
.B(n_1108),
.Y(n_1366)
);

AOI21x1_ASAP7_75t_L g1367 ( 
.A1(n_1106),
.A2(n_1104),
.B(n_1092),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_1093),
.Y(n_1368)
);

OAI21x1_ASAP7_75t_L g1369 ( 
.A1(n_1132),
.A2(n_1139),
.B(n_1138),
.Y(n_1369)
);

OR2x2_ASAP7_75t_L g1370 ( 
.A(n_1202),
.B(n_1117),
.Y(n_1370)
);

AOI221xp5_ASAP7_75t_SL g1371 ( 
.A1(n_1096),
.A2(n_934),
.B1(n_1195),
.B2(n_1194),
.C(n_1144),
.Y(n_1371)
);

OAI21xp5_ASAP7_75t_L g1372 ( 
.A1(n_1244),
.A2(n_754),
.B(n_921),
.Y(n_1372)
);

AND2x4_ASAP7_75t_L g1373 ( 
.A(n_1222),
.B(n_988),
.Y(n_1373)
);

OAI22xp5_ASAP7_75t_L g1374 ( 
.A1(n_1230),
.A2(n_754),
.B1(n_926),
.B2(n_795),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1202),
.B(n_1031),
.Y(n_1375)
);

AND2x4_ASAP7_75t_L g1376 ( 
.A(n_1222),
.B(n_988),
.Y(n_1376)
);

AOI21xp5_ASAP7_75t_L g1377 ( 
.A1(n_1092),
.A2(n_708),
.B(n_1036),
.Y(n_1377)
);

AOI21xp5_ASAP7_75t_L g1378 ( 
.A1(n_1092),
.A2(n_708),
.B(n_1036),
.Y(n_1378)
);

AOI221x1_ASAP7_75t_L g1379 ( 
.A1(n_1170),
.A2(n_1177),
.B1(n_1092),
.B2(n_1208),
.C(n_1200),
.Y(n_1379)
);

AO31x2_ASAP7_75t_L g1380 ( 
.A1(n_1092),
.A2(n_1234),
.A3(n_1252),
.B(n_1108),
.Y(n_1380)
);

AOI21xp5_ASAP7_75t_L g1381 ( 
.A1(n_1092),
.A2(n_708),
.B(n_1036),
.Y(n_1381)
);

AOI221xp5_ASAP7_75t_L g1382 ( 
.A1(n_1096),
.A2(n_970),
.B1(n_395),
.B2(n_984),
.C(n_990),
.Y(n_1382)
);

AO31x2_ASAP7_75t_L g1383 ( 
.A1(n_1092),
.A2(n_1234),
.A3(n_1252),
.B(n_1108),
.Y(n_1383)
);

OAI21xp33_ASAP7_75t_L g1384 ( 
.A1(n_1155),
.A2(n_970),
.B(n_984),
.Y(n_1384)
);

AOI21xp5_ASAP7_75t_L g1385 ( 
.A1(n_1092),
.A2(n_708),
.B(n_1036),
.Y(n_1385)
);

A2O1A1Ixp33_ASAP7_75t_L g1386 ( 
.A1(n_1095),
.A2(n_1094),
.B(n_754),
.C(n_984),
.Y(n_1386)
);

INVx5_ASAP7_75t_L g1387 ( 
.A(n_1140),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1105),
.B(n_926),
.Y(n_1388)
);

OAI21x1_ASAP7_75t_SL g1389 ( 
.A1(n_1118),
.A2(n_1122),
.B(n_1115),
.Y(n_1389)
);

NAND2x1p5_ASAP7_75t_L g1390 ( 
.A(n_1114),
.B(n_988),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1105),
.B(n_926),
.Y(n_1391)
);

O2A1O1Ixp33_ASAP7_75t_SL g1392 ( 
.A1(n_1208),
.A2(n_1118),
.B(n_1122),
.C(n_1197),
.Y(n_1392)
);

AO31x2_ASAP7_75t_L g1393 ( 
.A1(n_1092),
.A2(n_1234),
.A3(n_1252),
.B(n_1108),
.Y(n_1393)
);

HB1xp67_ASAP7_75t_L g1394 ( 
.A(n_1114),
.Y(n_1394)
);

AO21x1_ASAP7_75t_L g1395 ( 
.A1(n_1181),
.A2(n_1166),
.B(n_1171),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1093),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1093),
.Y(n_1397)
);

INVx3_ASAP7_75t_L g1398 ( 
.A(n_1167),
.Y(n_1398)
);

OR2x2_ASAP7_75t_L g1399 ( 
.A(n_1202),
.B(n_1117),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1093),
.Y(n_1400)
);

OAI22xp5_ASAP7_75t_L g1401 ( 
.A1(n_1230),
.A2(n_754),
.B1(n_926),
.B2(n_795),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1105),
.B(n_926),
.Y(n_1402)
);

AO31x2_ASAP7_75t_L g1403 ( 
.A1(n_1092),
.A2(n_1234),
.A3(n_1252),
.B(n_1108),
.Y(n_1403)
);

AOI21xp5_ASAP7_75t_L g1404 ( 
.A1(n_1092),
.A2(n_708),
.B(n_1036),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1105),
.B(n_926),
.Y(n_1405)
);

INVx2_ASAP7_75t_SL g1406 ( 
.A(n_1142),
.Y(n_1406)
);

AO21x1_ASAP7_75t_L g1407 ( 
.A1(n_1181),
.A2(n_1166),
.B(n_1171),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1093),
.Y(n_1408)
);

AOI21x1_ASAP7_75t_L g1409 ( 
.A1(n_1106),
.A2(n_1104),
.B(n_1092),
.Y(n_1409)
);

OAI22xp5_ASAP7_75t_L g1410 ( 
.A1(n_1230),
.A2(n_754),
.B1(n_926),
.B2(n_795),
.Y(n_1410)
);

AO31x2_ASAP7_75t_L g1411 ( 
.A1(n_1092),
.A2(n_1234),
.A3(n_1252),
.B(n_1108),
.Y(n_1411)
);

OAI21xp5_ASAP7_75t_L g1412 ( 
.A1(n_1244),
.A2(n_754),
.B(n_921),
.Y(n_1412)
);

AOI22xp5_ASAP7_75t_L g1413 ( 
.A1(n_1155),
.A2(n_970),
.B1(n_936),
.B2(n_933),
.Y(n_1413)
);

AOI21xp5_ASAP7_75t_L g1414 ( 
.A1(n_1092),
.A2(n_708),
.B(n_1036),
.Y(n_1414)
);

INVx3_ASAP7_75t_L g1415 ( 
.A(n_1167),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_1093),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1093),
.Y(n_1417)
);

OA21x2_ASAP7_75t_L g1418 ( 
.A1(n_1228),
.A2(n_1092),
.B(n_1108),
.Y(n_1418)
);

AOI21xp5_ASAP7_75t_L g1419 ( 
.A1(n_1092),
.A2(n_708),
.B(n_1036),
.Y(n_1419)
);

O2A1O1Ixp5_ASAP7_75t_L g1420 ( 
.A1(n_1108),
.A2(n_733),
.B(n_984),
.C(n_1092),
.Y(n_1420)
);

OAI21x1_ASAP7_75t_L g1421 ( 
.A1(n_1132),
.A2(n_1139),
.B(n_1138),
.Y(n_1421)
);

OAI21x1_ASAP7_75t_L g1422 ( 
.A1(n_1132),
.A2(n_1139),
.B(n_1138),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1202),
.B(n_1031),
.Y(n_1423)
);

BUFx4f_ASAP7_75t_L g1424 ( 
.A(n_1280),
.Y(n_1424)
);

OAI22xp5_ASAP7_75t_L g1425 ( 
.A1(n_1413),
.A2(n_1382),
.B1(n_1384),
.B2(n_1277),
.Y(n_1425)
);

INVx2_ASAP7_75t_SL g1426 ( 
.A(n_1297),
.Y(n_1426)
);

INVx4_ASAP7_75t_L g1427 ( 
.A(n_1340),
.Y(n_1427)
);

BUFx12f_ASAP7_75t_L g1428 ( 
.A(n_1297),
.Y(n_1428)
);

INVx6_ASAP7_75t_L g1429 ( 
.A(n_1340),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1287),
.Y(n_1430)
);

HB1xp67_ASAP7_75t_L g1431 ( 
.A(n_1394),
.Y(n_1431)
);

BUFx6f_ASAP7_75t_L g1432 ( 
.A(n_1254),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1296),
.Y(n_1433)
);

BUFx3_ASAP7_75t_L g1434 ( 
.A(n_1361),
.Y(n_1434)
);

OAI22xp33_ASAP7_75t_L g1435 ( 
.A1(n_1302),
.A2(n_1275),
.B1(n_1405),
.B2(n_1352),
.Y(n_1435)
);

AOI22xp33_ASAP7_75t_SL g1436 ( 
.A1(n_1273),
.A2(n_1374),
.B1(n_1410),
.B2(n_1401),
.Y(n_1436)
);

INVx1_ASAP7_75t_SL g1437 ( 
.A(n_1370),
.Y(n_1437)
);

BUFx10_ASAP7_75t_L g1438 ( 
.A(n_1359),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1276),
.Y(n_1439)
);

CKINVDCx11_ASAP7_75t_R g1440 ( 
.A(n_1268),
.Y(n_1440)
);

AOI22xp33_ASAP7_75t_L g1441 ( 
.A1(n_1342),
.A2(n_1357),
.B1(n_1372),
.B2(n_1412),
.Y(n_1441)
);

BUFx10_ASAP7_75t_L g1442 ( 
.A(n_1288),
.Y(n_1442)
);

AOI22xp5_ASAP7_75t_SL g1443 ( 
.A1(n_1329),
.A2(n_1267),
.B1(n_1388),
.B2(n_1391),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1276),
.Y(n_1444)
);

BUFx3_ASAP7_75t_L g1445 ( 
.A(n_1340),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1300),
.Y(n_1446)
);

OAI21xp5_ASAP7_75t_SL g1447 ( 
.A1(n_1328),
.A2(n_1272),
.B(n_1386),
.Y(n_1447)
);

AOI22xp33_ASAP7_75t_L g1448 ( 
.A1(n_1347),
.A2(n_1402),
.B1(n_1256),
.B2(n_1255),
.Y(n_1448)
);

BUFx12f_ASAP7_75t_L g1449 ( 
.A(n_1281),
.Y(n_1449)
);

CKINVDCx11_ASAP7_75t_R g1450 ( 
.A(n_1286),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1300),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1344),
.B(n_1346),
.Y(n_1452)
);

NOR2xp33_ASAP7_75t_L g1453 ( 
.A(n_1363),
.B(n_1399),
.Y(n_1453)
);

AOI22xp33_ASAP7_75t_L g1454 ( 
.A1(n_1293),
.A2(n_1323),
.B1(n_1395),
.B2(n_1407),
.Y(n_1454)
);

AOI22xp33_ASAP7_75t_L g1455 ( 
.A1(n_1364),
.A2(n_1375),
.B1(n_1423),
.B2(n_1265),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_1301),
.Y(n_1456)
);

AOI22xp33_ASAP7_75t_L g1457 ( 
.A1(n_1389),
.A2(n_1260),
.B1(n_1312),
.B2(n_1294),
.Y(n_1457)
);

INVx1_ASAP7_75t_SL g1458 ( 
.A(n_1406),
.Y(n_1458)
);

INVx4_ASAP7_75t_L g1459 ( 
.A(n_1387),
.Y(n_1459)
);

AOI22xp33_ASAP7_75t_L g1460 ( 
.A1(n_1333),
.A2(n_1368),
.B1(n_1408),
.B2(n_1416),
.Y(n_1460)
);

BUFx12f_ASAP7_75t_L g1461 ( 
.A(n_1254),
.Y(n_1461)
);

INVxp67_ASAP7_75t_L g1462 ( 
.A(n_1264),
.Y(n_1462)
);

NAND2x1p5_ASAP7_75t_L g1463 ( 
.A(n_1387),
.B(n_1274),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1396),
.Y(n_1464)
);

AOI22x1_ASAP7_75t_SL g1465 ( 
.A1(n_1348),
.A2(n_1417),
.B1(n_1400),
.B2(n_1396),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1397),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1319),
.B(n_1289),
.Y(n_1467)
);

INVx8_ASAP7_75t_L g1468 ( 
.A(n_1356),
.Y(n_1468)
);

BUFx3_ASAP7_75t_L g1469 ( 
.A(n_1254),
.Y(n_1469)
);

OAI22xp33_ASAP7_75t_L g1470 ( 
.A1(n_1379),
.A2(n_1350),
.B1(n_1365),
.B2(n_1354),
.Y(n_1470)
);

AOI22xp33_ASAP7_75t_SL g1471 ( 
.A1(n_1339),
.A2(n_1373),
.B1(n_1376),
.B2(n_1291),
.Y(n_1471)
);

AOI22xp33_ASAP7_75t_L g1472 ( 
.A1(n_1310),
.A2(n_1309),
.B1(n_1320),
.B2(n_1292),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1371),
.B(n_1291),
.Y(n_1473)
);

AOI22xp33_ASAP7_75t_L g1474 ( 
.A1(n_1320),
.A2(n_1339),
.B1(n_1376),
.B2(n_1373),
.Y(n_1474)
);

AOI22xp33_ASAP7_75t_L g1475 ( 
.A1(n_1303),
.A2(n_1308),
.B1(n_1324),
.B2(n_1306),
.Y(n_1475)
);

BUFx3_ASAP7_75t_L g1476 ( 
.A(n_1269),
.Y(n_1476)
);

AOI22xp33_ASAP7_75t_L g1477 ( 
.A1(n_1307),
.A2(n_1290),
.B1(n_1299),
.B2(n_1304),
.Y(n_1477)
);

BUFx2_ASAP7_75t_R g1478 ( 
.A(n_1332),
.Y(n_1478)
);

OAI22xp5_ASAP7_75t_L g1479 ( 
.A1(n_1283),
.A2(n_1298),
.B1(n_1390),
.B2(n_1278),
.Y(n_1479)
);

AOI22xp5_ASAP7_75t_L g1480 ( 
.A1(n_1290),
.A2(n_1278),
.B1(n_1392),
.B2(n_1271),
.Y(n_1480)
);

OAI22xp5_ASAP7_75t_L g1481 ( 
.A1(n_1311),
.A2(n_1321),
.B1(n_1315),
.B2(n_1348),
.Y(n_1481)
);

BUFx12f_ASAP7_75t_L g1482 ( 
.A(n_1269),
.Y(n_1482)
);

BUFx10_ASAP7_75t_L g1483 ( 
.A(n_1356),
.Y(n_1483)
);

OAI22xp5_ASAP7_75t_L g1484 ( 
.A1(n_1313),
.A2(n_1314),
.B1(n_1331),
.B2(n_1398),
.Y(n_1484)
);

BUFx2_ASAP7_75t_SL g1485 ( 
.A(n_1335),
.Y(n_1485)
);

AOI22xp5_ASAP7_75t_L g1486 ( 
.A1(n_1299),
.A2(n_1326),
.B1(n_1362),
.B2(n_1415),
.Y(n_1486)
);

INVx4_ASAP7_75t_L g1487 ( 
.A(n_1356),
.Y(n_1487)
);

AOI22xp33_ASAP7_75t_L g1488 ( 
.A1(n_1418),
.A2(n_1285),
.B1(n_1284),
.B2(n_1318),
.Y(n_1488)
);

BUFx2_ASAP7_75t_L g1489 ( 
.A(n_1338),
.Y(n_1489)
);

CKINVDCx11_ASAP7_75t_R g1490 ( 
.A(n_1337),
.Y(n_1490)
);

HB1xp67_ASAP7_75t_L g1491 ( 
.A(n_1398),
.Y(n_1491)
);

INVx8_ASAP7_75t_L g1492 ( 
.A(n_1415),
.Y(n_1492)
);

AOI22xp33_ASAP7_75t_L g1493 ( 
.A1(n_1418),
.A2(n_1285),
.B1(n_1284),
.B2(n_1279),
.Y(n_1493)
);

AOI22xp33_ASAP7_75t_L g1494 ( 
.A1(n_1330),
.A2(n_1262),
.B1(n_1419),
.B2(n_1414),
.Y(n_1494)
);

OAI22xp5_ASAP7_75t_L g1495 ( 
.A1(n_1343),
.A2(n_1353),
.B1(n_1349),
.B2(n_1345),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1334),
.Y(n_1496)
);

AOI22xp33_ASAP7_75t_SL g1497 ( 
.A1(n_1351),
.A2(n_1377),
.B1(n_1404),
.B2(n_1385),
.Y(n_1497)
);

AOI22xp33_ASAP7_75t_L g1498 ( 
.A1(n_1378),
.A2(n_1381),
.B1(n_1295),
.B2(n_1270),
.Y(n_1498)
);

BUFx3_ASAP7_75t_L g1499 ( 
.A(n_1282),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1317),
.Y(n_1500)
);

BUFx6f_ASAP7_75t_L g1501 ( 
.A(n_1317),
.Y(n_1501)
);

OAI22xp33_ASAP7_75t_L g1502 ( 
.A1(n_1327),
.A2(n_1336),
.B1(n_1263),
.B2(n_1409),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1317),
.Y(n_1503)
);

AOI22xp33_ASAP7_75t_L g1504 ( 
.A1(n_1358),
.A2(n_1360),
.B1(n_1421),
.B2(n_1369),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1282),
.B(n_1322),
.Y(n_1505)
);

CKINVDCx11_ASAP7_75t_R g1506 ( 
.A(n_1420),
.Y(n_1506)
);

AOI22xp33_ASAP7_75t_L g1507 ( 
.A1(n_1422),
.A2(n_1325),
.B1(n_1261),
.B2(n_1316),
.Y(n_1507)
);

AOI22xp33_ASAP7_75t_L g1508 ( 
.A1(n_1316),
.A2(n_1258),
.B1(n_1305),
.B2(n_1257),
.Y(n_1508)
);

AOI22xp33_ASAP7_75t_L g1509 ( 
.A1(n_1316),
.A2(n_1305),
.B1(n_1411),
.B2(n_1366),
.Y(n_1509)
);

BUFx4_ASAP7_75t_R g1510 ( 
.A(n_1266),
.Y(n_1510)
);

INVx3_ASAP7_75t_L g1511 ( 
.A(n_1341),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1322),
.B(n_1411),
.Y(n_1512)
);

OAI221xp5_ASAP7_75t_L g1513 ( 
.A1(n_1367),
.A2(n_1305),
.B1(n_1266),
.B2(n_1366),
.C(n_1380),
.Y(n_1513)
);

OAI22xp5_ASAP7_75t_L g1514 ( 
.A1(n_1266),
.A2(n_1380),
.B1(n_1403),
.B2(n_1341),
.Y(n_1514)
);

BUFx2_ASAP7_75t_L g1515 ( 
.A(n_1322),
.Y(n_1515)
);

OAI22xp33_ASAP7_75t_L g1516 ( 
.A1(n_1355),
.A2(n_1411),
.B1(n_1366),
.B2(n_1380),
.Y(n_1516)
);

BUFx2_ASAP7_75t_L g1517 ( 
.A(n_1355),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1383),
.Y(n_1518)
);

AOI22xp33_ASAP7_75t_SL g1519 ( 
.A1(n_1383),
.A2(n_1393),
.B1(n_1403),
.B2(n_1259),
.Y(n_1519)
);

CKINVDCx6p67_ASAP7_75t_R g1520 ( 
.A(n_1259),
.Y(n_1520)
);

INVx6_ASAP7_75t_L g1521 ( 
.A(n_1393),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1259),
.Y(n_1522)
);

NAND2x1p5_ASAP7_75t_L g1523 ( 
.A(n_1340),
.B(n_1387),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1287),
.Y(n_1524)
);

CKINVDCx6p67_ASAP7_75t_R g1525 ( 
.A(n_1280),
.Y(n_1525)
);

AOI22xp33_ASAP7_75t_L g1526 ( 
.A1(n_1382),
.A2(n_1384),
.B1(n_1342),
.B2(n_1374),
.Y(n_1526)
);

AOI22xp33_ASAP7_75t_SL g1527 ( 
.A1(n_1273),
.A2(n_1155),
.B1(n_1053),
.B2(n_544),
.Y(n_1527)
);

CKINVDCx14_ASAP7_75t_R g1528 ( 
.A(n_1359),
.Y(n_1528)
);

INVx1_ASAP7_75t_SL g1529 ( 
.A(n_1394),
.Y(n_1529)
);

INVx6_ASAP7_75t_L g1530 ( 
.A(n_1340),
.Y(n_1530)
);

OAI22xp5_ASAP7_75t_L g1531 ( 
.A1(n_1413),
.A2(n_1382),
.B1(n_1384),
.B2(n_970),
.Y(n_1531)
);

AOI22xp33_ASAP7_75t_SL g1532 ( 
.A1(n_1273),
.A2(n_1155),
.B1(n_1053),
.B2(n_544),
.Y(n_1532)
);

OAI22xp5_ASAP7_75t_L g1533 ( 
.A1(n_1413),
.A2(n_1382),
.B1(n_1384),
.B2(n_970),
.Y(n_1533)
);

INVx4_ASAP7_75t_L g1534 ( 
.A(n_1340),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1344),
.B(n_1346),
.Y(n_1535)
);

BUFx3_ASAP7_75t_L g1536 ( 
.A(n_1361),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1287),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1344),
.B(n_1346),
.Y(n_1538)
);

BUFx10_ASAP7_75t_L g1539 ( 
.A(n_1359),
.Y(n_1539)
);

CKINVDCx11_ASAP7_75t_R g1540 ( 
.A(n_1268),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1287),
.Y(n_1541)
);

BUFx12f_ASAP7_75t_L g1542 ( 
.A(n_1297),
.Y(n_1542)
);

INVx6_ASAP7_75t_L g1543 ( 
.A(n_1340),
.Y(n_1543)
);

BUFx10_ASAP7_75t_L g1544 ( 
.A(n_1359),
.Y(n_1544)
);

BUFx2_ASAP7_75t_L g1545 ( 
.A(n_1394),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1287),
.Y(n_1546)
);

CKINVDCx20_ASAP7_75t_R g1547 ( 
.A(n_1281),
.Y(n_1547)
);

CKINVDCx11_ASAP7_75t_R g1548 ( 
.A(n_1268),
.Y(n_1548)
);

AOI22xp33_ASAP7_75t_SL g1549 ( 
.A1(n_1273),
.A2(n_1155),
.B1(n_1053),
.B2(n_544),
.Y(n_1549)
);

AOI22xp5_ASAP7_75t_L g1550 ( 
.A1(n_1384),
.A2(n_1382),
.B1(n_970),
.B2(n_936),
.Y(n_1550)
);

AOI22xp33_ASAP7_75t_L g1551 ( 
.A1(n_1382),
.A2(n_1384),
.B1(n_1342),
.B2(n_1374),
.Y(n_1551)
);

OAI21xp5_ASAP7_75t_SL g1552 ( 
.A1(n_1382),
.A2(n_1413),
.B(n_618),
.Y(n_1552)
);

CKINVDCx11_ASAP7_75t_R g1553 ( 
.A(n_1268),
.Y(n_1553)
);

BUFx6f_ASAP7_75t_SL g1554 ( 
.A(n_1297),
.Y(n_1554)
);

BUFx2_ASAP7_75t_L g1555 ( 
.A(n_1394),
.Y(n_1555)
);

AOI22xp33_ASAP7_75t_L g1556 ( 
.A1(n_1382),
.A2(n_1384),
.B1(n_1342),
.B2(n_1374),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1287),
.Y(n_1557)
);

OAI21xp5_ASAP7_75t_L g1558 ( 
.A1(n_1342),
.A2(n_1382),
.B(n_984),
.Y(n_1558)
);

AOI22xp33_ASAP7_75t_SL g1559 ( 
.A1(n_1273),
.A2(n_1155),
.B1(n_1053),
.B2(n_544),
.Y(n_1559)
);

INVx6_ASAP7_75t_L g1560 ( 
.A(n_1340),
.Y(n_1560)
);

AOI22xp33_ASAP7_75t_SL g1561 ( 
.A1(n_1273),
.A2(n_1155),
.B1(n_1053),
.B2(n_544),
.Y(n_1561)
);

OAI22xp5_ASAP7_75t_L g1562 ( 
.A1(n_1413),
.A2(n_1382),
.B1(n_1384),
.B2(n_970),
.Y(n_1562)
);

OAI22xp33_ASAP7_75t_L g1563 ( 
.A1(n_1413),
.A2(n_1053),
.B1(n_1155),
.B2(n_544),
.Y(n_1563)
);

BUFx2_ASAP7_75t_SL g1564 ( 
.A(n_1340),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1287),
.Y(n_1565)
);

AOI21xp5_ASAP7_75t_L g1566 ( 
.A1(n_1558),
.A2(n_1457),
.B(n_1481),
.Y(n_1566)
);

AOI21x1_ASAP7_75t_L g1567 ( 
.A1(n_1495),
.A2(n_1496),
.B(n_1484),
.Y(n_1567)
);

INVxp67_ASAP7_75t_R g1568 ( 
.A(n_1452),
.Y(n_1568)
);

CKINVDCx20_ASAP7_75t_R g1569 ( 
.A(n_1440),
.Y(n_1569)
);

AND2x4_ASAP7_75t_L g1570 ( 
.A(n_1499),
.B(n_1456),
.Y(n_1570)
);

INVx3_ASAP7_75t_L g1571 ( 
.A(n_1521),
.Y(n_1571)
);

NAND2x1p5_ASAP7_75t_L g1572 ( 
.A(n_1486),
.B(n_1499),
.Y(n_1572)
);

HB1xp67_ASAP7_75t_L g1573 ( 
.A(n_1431),
.Y(n_1573)
);

BUFx2_ASAP7_75t_L g1574 ( 
.A(n_1517),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1518),
.Y(n_1575)
);

OA21x2_ASAP7_75t_L g1576 ( 
.A1(n_1507),
.A2(n_1508),
.B(n_1509),
.Y(n_1576)
);

OAI221xp5_ASAP7_75t_L g1577 ( 
.A1(n_1552),
.A2(n_1550),
.B1(n_1436),
.B2(n_1526),
.C(n_1551),
.Y(n_1577)
);

INVx1_ASAP7_75t_SL g1578 ( 
.A(n_1529),
.Y(n_1578)
);

OR2x2_ASAP7_75t_L g1579 ( 
.A(n_1501),
.B(n_1500),
.Y(n_1579)
);

NOR2xp67_ASAP7_75t_L g1580 ( 
.A(n_1480),
.B(n_1447),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1512),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1505),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1511),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1501),
.B(n_1441),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1439),
.Y(n_1585)
);

INVx1_ASAP7_75t_SL g1586 ( 
.A(n_1458),
.Y(n_1586)
);

CKINVDCx9p33_ASAP7_75t_R g1587 ( 
.A(n_1465),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1444),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1446),
.Y(n_1589)
);

INVx2_ASAP7_75t_SL g1590 ( 
.A(n_1429),
.Y(n_1590)
);

HB1xp67_ASAP7_75t_L g1591 ( 
.A(n_1489),
.Y(n_1591)
);

BUFx3_ASAP7_75t_L g1592 ( 
.A(n_1434),
.Y(n_1592)
);

INVx4_ASAP7_75t_L g1593 ( 
.A(n_1468),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1451),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1464),
.Y(n_1595)
);

OR2x2_ASAP7_75t_L g1596 ( 
.A(n_1501),
.B(n_1503),
.Y(n_1596)
);

INVx2_ASAP7_75t_L g1597 ( 
.A(n_1466),
.Y(n_1597)
);

BUFx6f_ASAP7_75t_L g1598 ( 
.A(n_1506),
.Y(n_1598)
);

OR2x6_ASAP7_75t_L g1599 ( 
.A(n_1514),
.B(n_1468),
.Y(n_1599)
);

OR2x6_ASAP7_75t_L g1600 ( 
.A(n_1468),
.B(n_1510),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1454),
.B(n_1520),
.Y(n_1601)
);

HB1xp67_ASAP7_75t_L g1602 ( 
.A(n_1545),
.Y(n_1602)
);

INVx2_ASAP7_75t_L g1603 ( 
.A(n_1522),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1515),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1510),
.Y(n_1605)
);

BUFx3_ASAP7_75t_L g1606 ( 
.A(n_1536),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1516),
.Y(n_1607)
);

AOI21x1_ASAP7_75t_L g1608 ( 
.A1(n_1531),
.A2(n_1533),
.B(n_1562),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1513),
.Y(n_1609)
);

HB1xp67_ASAP7_75t_L g1610 ( 
.A(n_1555),
.Y(n_1610)
);

O2A1O1Ixp33_ASAP7_75t_L g1611 ( 
.A1(n_1563),
.A2(n_1425),
.B(n_1526),
.C(n_1551),
.Y(n_1611)
);

AO21x2_ASAP7_75t_L g1612 ( 
.A1(n_1502),
.A2(n_1479),
.B(n_1435),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1519),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1454),
.B(n_1457),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1509),
.Y(n_1615)
);

HB1xp67_ASAP7_75t_L g1616 ( 
.A(n_1536),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1506),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1508),
.Y(n_1618)
);

OAI21x1_ASAP7_75t_L g1619 ( 
.A1(n_1498),
.A2(n_1504),
.B(n_1494),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1477),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1477),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1475),
.Y(n_1622)
);

INVx3_ASAP7_75t_L g1623 ( 
.A(n_1483),
.Y(n_1623)
);

AOI22xp33_ASAP7_75t_SL g1624 ( 
.A1(n_1443),
.A2(n_1473),
.B1(n_1467),
.B2(n_1556),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1448),
.B(n_1437),
.Y(n_1625)
);

OA21x2_ASAP7_75t_L g1626 ( 
.A1(n_1507),
.A2(n_1488),
.B(n_1493),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1475),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1430),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1433),
.Y(n_1629)
);

AOI21xp5_ASAP7_75t_L g1630 ( 
.A1(n_1493),
.A2(n_1556),
.B(n_1494),
.Y(n_1630)
);

AOI22xp33_ASAP7_75t_L g1631 ( 
.A1(n_1527),
.A2(n_1561),
.B1(n_1559),
.B2(n_1532),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1524),
.Y(n_1632)
);

CKINVDCx14_ASAP7_75t_R g1633 ( 
.A(n_1528),
.Y(n_1633)
);

NOR2xp33_ASAP7_75t_L g1634 ( 
.A(n_1462),
.B(n_1535),
.Y(n_1634)
);

AOI22xp33_ASAP7_75t_L g1635 ( 
.A1(n_1549),
.A2(n_1455),
.B1(n_1470),
.B2(n_1453),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1537),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1448),
.B(n_1541),
.Y(n_1637)
);

BUFx2_ASAP7_75t_L g1638 ( 
.A(n_1491),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1455),
.B(n_1538),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1546),
.B(n_1565),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1557),
.Y(n_1641)
);

INVx3_ASAP7_75t_L g1642 ( 
.A(n_1487),
.Y(n_1642)
);

NOR2xp33_ASAP7_75t_L g1643 ( 
.A(n_1453),
.B(n_1528),
.Y(n_1643)
);

OA21x2_ASAP7_75t_L g1644 ( 
.A1(n_1488),
.A2(n_1498),
.B(n_1504),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1460),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1460),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1497),
.Y(n_1647)
);

BUFx3_ASAP7_75t_L g1648 ( 
.A(n_1429),
.Y(n_1648)
);

BUFx10_ASAP7_75t_L g1649 ( 
.A(n_1554),
.Y(n_1649)
);

AO21x2_ASAP7_75t_L g1650 ( 
.A1(n_1490),
.A2(n_1474),
.B(n_1472),
.Y(n_1650)
);

OAI21xp5_ASAP7_75t_L g1651 ( 
.A1(n_1472),
.A2(n_1474),
.B(n_1463),
.Y(n_1651)
);

AOI22xp33_ASAP7_75t_L g1652 ( 
.A1(n_1490),
.A2(n_1471),
.B1(n_1554),
.B2(n_1428),
.Y(n_1652)
);

OR2x6_ASAP7_75t_L g1653 ( 
.A(n_1564),
.B(n_1523),
.Y(n_1653)
);

INVx8_ASAP7_75t_L g1654 ( 
.A(n_1461),
.Y(n_1654)
);

AOI21x1_ASAP7_75t_L g1655 ( 
.A1(n_1426),
.A2(n_1485),
.B(n_1463),
.Y(n_1655)
);

OAI22xp5_ASAP7_75t_L g1656 ( 
.A1(n_1478),
.A2(n_1424),
.B1(n_1560),
.B2(n_1543),
.Y(n_1656)
);

HB1xp67_ASAP7_75t_SL g1657 ( 
.A(n_1469),
.Y(n_1657)
);

OAI21x1_ASAP7_75t_L g1658 ( 
.A1(n_1492),
.A2(n_1560),
.B(n_1530),
.Y(n_1658)
);

OR2x2_ASAP7_75t_L g1659 ( 
.A(n_1445),
.B(n_1534),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1492),
.Y(n_1660)
);

HB1xp67_ASAP7_75t_L g1661 ( 
.A(n_1445),
.Y(n_1661)
);

AOI22xp33_ASAP7_75t_L g1662 ( 
.A1(n_1428),
.A2(n_1542),
.B1(n_1424),
.B2(n_1525),
.Y(n_1662)
);

OAI21xp5_ASAP7_75t_L g1663 ( 
.A1(n_1566),
.A2(n_1427),
.B(n_1459),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1637),
.B(n_1432),
.Y(n_1664)
);

OAI21x1_ASAP7_75t_SL g1665 ( 
.A1(n_1611),
.A2(n_1427),
.B(n_1534),
.Y(n_1665)
);

O2A1O1Ixp33_ASAP7_75t_SL g1666 ( 
.A1(n_1577),
.A2(n_1547),
.B(n_1560),
.C(n_1530),
.Y(n_1666)
);

AOI221xp5_ASAP7_75t_L g1667 ( 
.A1(n_1631),
.A2(n_1547),
.B1(n_1469),
.B2(n_1476),
.C(n_1459),
.Y(n_1667)
);

NOR2xp33_ASAP7_75t_SL g1668 ( 
.A(n_1569),
.B(n_1449),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1584),
.B(n_1438),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_1588),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1585),
.Y(n_1671)
);

O2A1O1Ixp33_ASAP7_75t_L g1672 ( 
.A1(n_1580),
.A2(n_1450),
.B(n_1542),
.C(n_1539),
.Y(n_1672)
);

AND2x2_ASAP7_75t_SL g1673 ( 
.A(n_1605),
.B(n_1543),
.Y(n_1673)
);

AOI21xp5_ASAP7_75t_L g1674 ( 
.A1(n_1612),
.A2(n_1543),
.B(n_1482),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_1588),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1585),
.Y(n_1676)
);

NOR2xp33_ASAP7_75t_L g1677 ( 
.A(n_1643),
.B(n_1442),
.Y(n_1677)
);

INVx2_ASAP7_75t_L g1678 ( 
.A(n_1588),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1605),
.B(n_1539),
.Y(n_1679)
);

BUFx3_ASAP7_75t_L g1680 ( 
.A(n_1648),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1581),
.B(n_1442),
.Y(n_1681)
);

AOI22x1_ASAP7_75t_SL g1682 ( 
.A1(n_1617),
.A2(n_1587),
.B1(n_1593),
.B2(n_1660),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1581),
.B(n_1544),
.Y(n_1683)
);

OR2x2_ASAP7_75t_L g1684 ( 
.A(n_1579),
.B(n_1544),
.Y(n_1684)
);

AO32x2_ASAP7_75t_L g1685 ( 
.A1(n_1579),
.A2(n_1450),
.A3(n_1449),
.B1(n_1440),
.B2(n_1540),
.Y(n_1685)
);

OAI21xp5_ASAP7_75t_L g1686 ( 
.A1(n_1608),
.A2(n_1540),
.B(n_1548),
.Y(n_1686)
);

CKINVDCx14_ASAP7_75t_R g1687 ( 
.A(n_1633),
.Y(n_1687)
);

HB1xp67_ASAP7_75t_L g1688 ( 
.A(n_1591),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1581),
.B(n_1548),
.Y(n_1689)
);

AO21x2_ASAP7_75t_L g1690 ( 
.A1(n_1630),
.A2(n_1553),
.B(n_1619),
.Y(n_1690)
);

OR2x2_ASAP7_75t_L g1691 ( 
.A(n_1596),
.B(n_1553),
.Y(n_1691)
);

OAI21xp5_ASAP7_75t_L g1692 ( 
.A1(n_1608),
.A2(n_1580),
.B(n_1635),
.Y(n_1692)
);

INVxp67_ASAP7_75t_L g1693 ( 
.A(n_1602),
.Y(n_1693)
);

CKINVDCx5p33_ASAP7_75t_R g1694 ( 
.A(n_1649),
.Y(n_1694)
);

HB1xp67_ASAP7_75t_L g1695 ( 
.A(n_1638),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1582),
.B(n_1613),
.Y(n_1696)
);

AND2x4_ASAP7_75t_L g1697 ( 
.A(n_1570),
.B(n_1571),
.Y(n_1697)
);

INVx8_ASAP7_75t_L g1698 ( 
.A(n_1654),
.Y(n_1698)
);

A2O1A1Ixp33_ASAP7_75t_L g1699 ( 
.A1(n_1624),
.A2(n_1614),
.B(n_1647),
.C(n_1651),
.Y(n_1699)
);

AOI22xp5_ASAP7_75t_L g1700 ( 
.A1(n_1612),
.A2(n_1652),
.B1(n_1617),
.B2(n_1598),
.Y(n_1700)
);

NAND2x1p5_ASAP7_75t_L g1701 ( 
.A(n_1658),
.B(n_1623),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1594),
.Y(n_1702)
);

INVxp67_ASAP7_75t_L g1703 ( 
.A(n_1610),
.Y(n_1703)
);

O2A1O1Ixp33_ASAP7_75t_L g1704 ( 
.A1(n_1625),
.A2(n_1612),
.B(n_1647),
.C(n_1617),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1582),
.B(n_1613),
.Y(n_1705)
);

OR2x6_ASAP7_75t_L g1706 ( 
.A(n_1600),
.B(n_1599),
.Y(n_1706)
);

NOR2x1_ASAP7_75t_SL g1707 ( 
.A(n_1600),
.B(n_1650),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1582),
.B(n_1615),
.Y(n_1708)
);

HB1xp67_ASAP7_75t_L g1709 ( 
.A(n_1638),
.Y(n_1709)
);

OR2x2_ASAP7_75t_L g1710 ( 
.A(n_1596),
.B(n_1639),
.Y(n_1710)
);

AOI211xp5_ASAP7_75t_L g1711 ( 
.A1(n_1598),
.A2(n_1656),
.B(n_1614),
.C(n_1609),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1573),
.B(n_1639),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1615),
.B(n_1600),
.Y(n_1713)
);

OR2x2_ASAP7_75t_L g1714 ( 
.A(n_1595),
.B(n_1597),
.Y(n_1714)
);

CKINVDCx20_ASAP7_75t_R g1715 ( 
.A(n_1592),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1600),
.B(n_1618),
.Y(n_1716)
);

NOR2xp33_ASAP7_75t_L g1717 ( 
.A(n_1634),
.B(n_1578),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1629),
.B(n_1632),
.Y(n_1718)
);

CKINVDCx20_ASAP7_75t_R g1719 ( 
.A(n_1592),
.Y(n_1719)
);

NOR2xp33_ASAP7_75t_L g1720 ( 
.A(n_1586),
.B(n_1616),
.Y(n_1720)
);

AOI21xp5_ASAP7_75t_L g1721 ( 
.A1(n_1600),
.A2(n_1572),
.B(n_1627),
.Y(n_1721)
);

CKINVDCx6p67_ASAP7_75t_R g1722 ( 
.A(n_1649),
.Y(n_1722)
);

AOI21xp5_ASAP7_75t_L g1723 ( 
.A1(n_1572),
.A2(n_1627),
.B(n_1622),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1618),
.B(n_1601),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1601),
.B(n_1570),
.Y(n_1725)
);

OAI22xp5_ASAP7_75t_L g1726 ( 
.A1(n_1598),
.A2(n_1657),
.B1(n_1568),
.B2(n_1662),
.Y(n_1726)
);

OA21x2_ASAP7_75t_L g1727 ( 
.A1(n_1609),
.A2(n_1607),
.B(n_1567),
.Y(n_1727)
);

AOI22xp5_ASAP7_75t_L g1728 ( 
.A1(n_1598),
.A2(n_1650),
.B1(n_1568),
.B2(n_1645),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1589),
.Y(n_1729)
);

NOR2xp33_ASAP7_75t_L g1730 ( 
.A(n_1677),
.B(n_1606),
.Y(n_1730)
);

OR2x2_ASAP7_75t_L g1731 ( 
.A(n_1710),
.B(n_1574),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1725),
.B(n_1576),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1725),
.B(n_1576),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1670),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1670),
.Y(n_1735)
);

INVx4_ASAP7_75t_R g1736 ( 
.A(n_1680),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1675),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1675),
.Y(n_1738)
);

INVx2_ASAP7_75t_L g1739 ( 
.A(n_1678),
.Y(n_1739)
);

OR2x2_ASAP7_75t_L g1740 ( 
.A(n_1712),
.B(n_1604),
.Y(n_1740)
);

INVxp67_ASAP7_75t_L g1741 ( 
.A(n_1688),
.Y(n_1741)
);

OR2x2_ASAP7_75t_L g1742 ( 
.A(n_1695),
.B(n_1576),
.Y(n_1742)
);

AND2x4_ASAP7_75t_L g1743 ( 
.A(n_1706),
.B(n_1599),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1716),
.B(n_1713),
.Y(n_1744)
);

AOI22xp33_ASAP7_75t_SL g1745 ( 
.A1(n_1692),
.A2(n_1598),
.B1(n_1650),
.B2(n_1572),
.Y(n_1745)
);

NOR2xp33_ASAP7_75t_L g1746 ( 
.A(n_1691),
.B(n_1598),
.Y(n_1746)
);

AND2x4_ASAP7_75t_L g1747 ( 
.A(n_1706),
.B(n_1599),
.Y(n_1747)
);

INVx3_ASAP7_75t_L g1748 ( 
.A(n_1702),
.Y(n_1748)
);

INVx1_ASAP7_75t_SL g1749 ( 
.A(n_1715),
.Y(n_1749)
);

AND2x4_ASAP7_75t_L g1750 ( 
.A(n_1706),
.B(n_1697),
.Y(n_1750)
);

AOI22xp33_ASAP7_75t_L g1751 ( 
.A1(n_1686),
.A2(n_1620),
.B1(n_1621),
.B2(n_1622),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1671),
.Y(n_1752)
);

OR2x2_ASAP7_75t_L g1753 ( 
.A(n_1709),
.B(n_1576),
.Y(n_1753)
);

OAI22xp5_ASAP7_75t_L g1754 ( 
.A1(n_1699),
.A2(n_1599),
.B1(n_1653),
.B2(n_1645),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1716),
.B(n_1599),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1676),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1729),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1714),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1724),
.B(n_1603),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1693),
.B(n_1636),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1724),
.B(n_1620),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1718),
.Y(n_1762)
);

OAI21xp5_ASAP7_75t_L g1763 ( 
.A1(n_1699),
.A2(n_1655),
.B(n_1646),
.Y(n_1763)
);

OR2x2_ASAP7_75t_L g1764 ( 
.A(n_1708),
.B(n_1696),
.Y(n_1764)
);

AND2x4_ASAP7_75t_L g1765 ( 
.A(n_1706),
.B(n_1583),
.Y(n_1765)
);

AND3x1_ASAP7_75t_L g1766 ( 
.A(n_1668),
.B(n_1640),
.C(n_1649),
.Y(n_1766)
);

OR2x2_ASAP7_75t_L g1767 ( 
.A(n_1696),
.B(n_1626),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1703),
.B(n_1636),
.Y(n_1768)
);

AND2x4_ASAP7_75t_L g1769 ( 
.A(n_1697),
.B(n_1583),
.Y(n_1769)
);

BUFx2_ASAP7_75t_L g1770 ( 
.A(n_1701),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1705),
.Y(n_1771)
);

INVx4_ASAP7_75t_L g1772 ( 
.A(n_1698),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1748),
.Y(n_1773)
);

BUFx2_ASAP7_75t_L g1774 ( 
.A(n_1770),
.Y(n_1774)
);

OR2x2_ASAP7_75t_L g1775 ( 
.A(n_1767),
.B(n_1742),
.Y(n_1775)
);

AOI221xp5_ASAP7_75t_L g1776 ( 
.A1(n_1763),
.A2(n_1704),
.B1(n_1666),
.B2(n_1667),
.C(n_1711),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1734),
.Y(n_1777)
);

OAI221xp5_ASAP7_75t_SL g1778 ( 
.A1(n_1751),
.A2(n_1700),
.B1(n_1728),
.B2(n_1672),
.C(n_1723),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1732),
.B(n_1707),
.Y(n_1779)
);

AOI222xp33_ASAP7_75t_L g1780 ( 
.A1(n_1754),
.A2(n_1646),
.B1(n_1717),
.B2(n_1726),
.C1(n_1663),
.C2(n_1689),
.Y(n_1780)
);

AND2x4_ASAP7_75t_SL g1781 ( 
.A(n_1743),
.B(n_1653),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1732),
.B(n_1690),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1734),
.Y(n_1783)
);

INVx4_ASAP7_75t_L g1784 ( 
.A(n_1772),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_SL g1785 ( 
.A(n_1766),
.B(n_1694),
.Y(n_1785)
);

NAND3xp33_ASAP7_75t_L g1786 ( 
.A(n_1745),
.B(n_1666),
.C(n_1664),
.Y(n_1786)
);

AOI31xp33_ASAP7_75t_L g1787 ( 
.A1(n_1749),
.A2(n_1687),
.A3(n_1689),
.B(n_1694),
.Y(n_1787)
);

AOI211xp5_ASAP7_75t_SL g1788 ( 
.A1(n_1746),
.A2(n_1674),
.B(n_1721),
.C(n_1642),
.Y(n_1788)
);

INVx2_ASAP7_75t_L g1789 ( 
.A(n_1767),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1762),
.B(n_1727),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1762),
.B(n_1727),
.Y(n_1791)
);

AOI33xp33_ASAP7_75t_L g1792 ( 
.A1(n_1761),
.A2(n_1752),
.A3(n_1756),
.B1(n_1757),
.B2(n_1640),
.B3(n_1683),
.Y(n_1792)
);

OAI31xp33_ASAP7_75t_L g1793 ( 
.A1(n_1741),
.A2(n_1687),
.A3(n_1679),
.B(n_1683),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1733),
.B(n_1690),
.Y(n_1794)
);

NOR2xp33_ASAP7_75t_L g1795 ( 
.A(n_1730),
.B(n_1684),
.Y(n_1795)
);

NAND2x1_ASAP7_75t_L g1796 ( 
.A(n_1736),
.B(n_1770),
.Y(n_1796)
);

INVx5_ASAP7_75t_SL g1797 ( 
.A(n_1743),
.Y(n_1797)
);

AND2x2_ASAP7_75t_L g1798 ( 
.A(n_1733),
.B(n_1690),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1735),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1735),
.Y(n_1800)
);

OAI221xp5_ASAP7_75t_SL g1801 ( 
.A1(n_1742),
.A2(n_1753),
.B1(n_1722),
.B2(n_1628),
.C(n_1641),
.Y(n_1801)
);

INVx2_ASAP7_75t_L g1802 ( 
.A(n_1739),
.Y(n_1802)
);

BUFx3_ASAP7_75t_L g1803 ( 
.A(n_1769),
.Y(n_1803)
);

AO21x2_ASAP7_75t_L g1804 ( 
.A1(n_1737),
.A2(n_1575),
.B(n_1567),
.Y(n_1804)
);

INVx3_ASAP7_75t_L g1805 ( 
.A(n_1750),
.Y(n_1805)
);

INVx4_ASAP7_75t_L g1806 ( 
.A(n_1772),
.Y(n_1806)
);

OAI31xp33_ASAP7_75t_L g1807 ( 
.A1(n_1753),
.A2(n_1679),
.A3(n_1669),
.B(n_1681),
.Y(n_1807)
);

OR2x2_ASAP7_75t_L g1808 ( 
.A(n_1731),
.B(n_1727),
.Y(n_1808)
);

NOR2xp33_ASAP7_75t_L g1809 ( 
.A(n_1760),
.B(n_1722),
.Y(n_1809)
);

AOI21xp5_ASAP7_75t_L g1810 ( 
.A1(n_1743),
.A2(n_1644),
.B(n_1626),
.Y(n_1810)
);

AND2x4_ASAP7_75t_L g1811 ( 
.A(n_1750),
.B(n_1697),
.Y(n_1811)
);

OAI22xp5_ASAP7_75t_L g1812 ( 
.A1(n_1731),
.A2(n_1673),
.B1(n_1715),
.B2(n_1719),
.Y(n_1812)
);

NOR2xp33_ASAP7_75t_L g1813 ( 
.A(n_1768),
.B(n_1649),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1738),
.Y(n_1814)
);

AOI22xp33_ASAP7_75t_L g1815 ( 
.A1(n_1776),
.A2(n_1747),
.B1(n_1673),
.B2(n_1750),
.Y(n_1815)
);

NOR2xp33_ASAP7_75t_L g1816 ( 
.A(n_1787),
.B(n_1720),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1777),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1792),
.B(n_1761),
.Y(n_1818)
);

INVx5_ASAP7_75t_SL g1819 ( 
.A(n_1804),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1777),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1783),
.Y(n_1821)
);

AND2x2_ASAP7_75t_L g1822 ( 
.A(n_1805),
.B(n_1744),
.Y(n_1822)
);

AND2x4_ASAP7_75t_L g1823 ( 
.A(n_1805),
.B(n_1750),
.Y(n_1823)
);

AND2x4_ASAP7_75t_L g1824 ( 
.A(n_1805),
.B(n_1747),
.Y(n_1824)
);

OR2x2_ASAP7_75t_L g1825 ( 
.A(n_1775),
.B(n_1764),
.Y(n_1825)
);

OR2x2_ASAP7_75t_L g1826 ( 
.A(n_1775),
.B(n_1764),
.Y(n_1826)
);

BUFx6f_ASAP7_75t_L g1827 ( 
.A(n_1796),
.Y(n_1827)
);

OR2x2_ASAP7_75t_L g1828 ( 
.A(n_1808),
.B(n_1740),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1783),
.Y(n_1829)
);

INVxp67_ASAP7_75t_L g1830 ( 
.A(n_1813),
.Y(n_1830)
);

INVxp67_ASAP7_75t_SL g1831 ( 
.A(n_1790),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1779),
.B(n_1747),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1799),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1799),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1800),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1800),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1782),
.B(n_1740),
.Y(n_1837)
);

INVx2_ASAP7_75t_SL g1838 ( 
.A(n_1796),
.Y(n_1838)
);

AND2x2_ASAP7_75t_L g1839 ( 
.A(n_1779),
.B(n_1747),
.Y(n_1839)
);

AND2x2_ASAP7_75t_L g1840 ( 
.A(n_1779),
.B(n_1755),
.Y(n_1840)
);

OR2x2_ASAP7_75t_L g1841 ( 
.A(n_1808),
.B(n_1789),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1811),
.B(n_1803),
.Y(n_1842)
);

AND2x2_ASAP7_75t_L g1843 ( 
.A(n_1811),
.B(n_1755),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1811),
.B(n_1759),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1782),
.B(n_1758),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1814),
.Y(n_1846)
);

AND2x4_ASAP7_75t_L g1847 ( 
.A(n_1811),
.B(n_1765),
.Y(n_1847)
);

AND2x2_ASAP7_75t_L g1848 ( 
.A(n_1803),
.B(n_1797),
.Y(n_1848)
);

AND2x2_ASAP7_75t_L g1849 ( 
.A(n_1803),
.B(n_1771),
.Y(n_1849)
);

INVx2_ASAP7_75t_L g1850 ( 
.A(n_1773),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1814),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1802),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1817),
.Y(n_1853)
);

INVx2_ASAP7_75t_L g1854 ( 
.A(n_1850),
.Y(n_1854)
);

INVx2_ASAP7_75t_SL g1855 ( 
.A(n_1827),
.Y(n_1855)
);

OR2x2_ASAP7_75t_L g1856 ( 
.A(n_1828),
.B(n_1790),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1817),
.Y(n_1857)
);

NOR2xp33_ASAP7_75t_L g1858 ( 
.A(n_1816),
.B(n_1787),
.Y(n_1858)
);

INVx3_ASAP7_75t_L g1859 ( 
.A(n_1827),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1827),
.B(n_1797),
.Y(n_1860)
);

AND2x2_ASAP7_75t_L g1861 ( 
.A(n_1827),
.B(n_1797),
.Y(n_1861)
);

NAND2x1p5_ASAP7_75t_L g1862 ( 
.A(n_1827),
.B(n_1784),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1820),
.Y(n_1863)
);

OR2x2_ASAP7_75t_L g1864 ( 
.A(n_1828),
.B(n_1791),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1820),
.Y(n_1865)
);

NAND3xp33_ASAP7_75t_L g1866 ( 
.A(n_1815),
.B(n_1778),
.C(n_1776),
.Y(n_1866)
);

OR2x6_ASAP7_75t_L g1867 ( 
.A(n_1838),
.B(n_1698),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1821),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1821),
.Y(n_1869)
);

INVx2_ASAP7_75t_L g1870 ( 
.A(n_1850),
.Y(n_1870)
);

INVxp67_ASAP7_75t_L g1871 ( 
.A(n_1818),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1829),
.Y(n_1872)
);

AND2x2_ASAP7_75t_L g1873 ( 
.A(n_1832),
.B(n_1797),
.Y(n_1873)
);

OR2x2_ASAP7_75t_L g1874 ( 
.A(n_1837),
.B(n_1791),
.Y(n_1874)
);

INVx2_ASAP7_75t_L g1875 ( 
.A(n_1841),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1829),
.Y(n_1876)
);

OAI21xp33_ASAP7_75t_L g1877 ( 
.A1(n_1831),
.A2(n_1778),
.B(n_1786),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1833),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1833),
.Y(n_1879)
);

AND2x2_ASAP7_75t_L g1880 ( 
.A(n_1832),
.B(n_1782),
.Y(n_1880)
);

INVx2_ASAP7_75t_L g1881 ( 
.A(n_1841),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1830),
.B(n_1794),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1844),
.B(n_1794),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1834),
.Y(n_1884)
);

AND2x4_ASAP7_75t_L g1885 ( 
.A(n_1838),
.B(n_1847),
.Y(n_1885)
);

AND2x2_ASAP7_75t_L g1886 ( 
.A(n_1839),
.B(n_1794),
.Y(n_1886)
);

AND2x2_ASAP7_75t_L g1887 ( 
.A(n_1839),
.B(n_1798),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_L g1888 ( 
.A(n_1844),
.B(n_1798),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1834),
.Y(n_1889)
);

INVx2_ASAP7_75t_L g1890 ( 
.A(n_1852),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1835),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1835),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1836),
.Y(n_1893)
);

OAI21xp5_ASAP7_75t_L g1894 ( 
.A1(n_1848),
.A2(n_1786),
.B(n_1788),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_L g1895 ( 
.A(n_1845),
.B(n_1798),
.Y(n_1895)
);

AND2x2_ASAP7_75t_L g1896 ( 
.A(n_1842),
.B(n_1774),
.Y(n_1896)
);

AND2x4_ASAP7_75t_L g1897 ( 
.A(n_1847),
.B(n_1781),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_SL g1898 ( 
.A(n_1847),
.B(n_1793),
.Y(n_1898)
);

AND2x4_ASAP7_75t_L g1899 ( 
.A(n_1885),
.B(n_1824),
.Y(n_1899)
);

AND2x2_ASAP7_75t_L g1900 ( 
.A(n_1860),
.B(n_1842),
.Y(n_1900)
);

AND2x2_ASAP7_75t_L g1901 ( 
.A(n_1860),
.B(n_1840),
.Y(n_1901)
);

INVx2_ASAP7_75t_L g1902 ( 
.A(n_1890),
.Y(n_1902)
);

AOI21xp5_ASAP7_75t_L g1903 ( 
.A1(n_1866),
.A2(n_1785),
.B(n_1788),
.Y(n_1903)
);

OR2x2_ASAP7_75t_L g1904 ( 
.A(n_1882),
.B(n_1825),
.Y(n_1904)
);

AND4x1_ASAP7_75t_L g1905 ( 
.A(n_1877),
.B(n_1780),
.C(n_1793),
.D(n_1807),
.Y(n_1905)
);

INVx1_ASAP7_75t_SL g1906 ( 
.A(n_1855),
.Y(n_1906)
);

AND3x1_ASAP7_75t_L g1907 ( 
.A(n_1858),
.B(n_1848),
.C(n_1807),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1871),
.B(n_1840),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1853),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1853),
.Y(n_1910)
);

HB1xp67_ASAP7_75t_L g1911 ( 
.A(n_1896),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1857),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1857),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1863),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1894),
.B(n_1843),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1875),
.B(n_1843),
.Y(n_1916)
);

BUFx3_ASAP7_75t_L g1917 ( 
.A(n_1859),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1863),
.Y(n_1918)
);

AND2x2_ASAP7_75t_L g1919 ( 
.A(n_1861),
.B(n_1847),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1875),
.B(n_1849),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1865),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1865),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1881),
.B(n_1849),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_SL g1924 ( 
.A(n_1861),
.B(n_1897),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1868),
.Y(n_1925)
);

AND2x2_ASAP7_75t_L g1926 ( 
.A(n_1873),
.B(n_1824),
.Y(n_1926)
);

AND2x2_ASAP7_75t_L g1927 ( 
.A(n_1873),
.B(n_1824),
.Y(n_1927)
);

OR2x2_ASAP7_75t_L g1928 ( 
.A(n_1881),
.B(n_1825),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_L g1929 ( 
.A(n_1896),
.B(n_1822),
.Y(n_1929)
);

AND2x2_ASAP7_75t_L g1930 ( 
.A(n_1885),
.B(n_1824),
.Y(n_1930)
);

NOR2xp33_ASAP7_75t_L g1931 ( 
.A(n_1898),
.B(n_1795),
.Y(n_1931)
);

AND2x2_ASAP7_75t_L g1932 ( 
.A(n_1885),
.B(n_1823),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_L g1933 ( 
.A(n_1880),
.B(n_1886),
.Y(n_1933)
);

INVx2_ASAP7_75t_L g1934 ( 
.A(n_1890),
.Y(n_1934)
);

OAI22xp5_ASAP7_75t_L g1935 ( 
.A1(n_1862),
.A2(n_1801),
.B1(n_1812),
.B2(n_1819),
.Y(n_1935)
);

OAI21xp33_ASAP7_75t_L g1936 ( 
.A1(n_1855),
.A2(n_1780),
.B(n_1801),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1909),
.Y(n_1937)
);

AOI22xp5_ASAP7_75t_L g1938 ( 
.A1(n_1907),
.A2(n_1897),
.B1(n_1867),
.B2(n_1859),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1911),
.B(n_1878),
.Y(n_1939)
);

AOI21xp5_ASAP7_75t_L g1940 ( 
.A1(n_1903),
.A2(n_1862),
.B(n_1859),
.Y(n_1940)
);

O2A1O1Ixp33_ASAP7_75t_L g1941 ( 
.A1(n_1935),
.A2(n_1862),
.B(n_1867),
.C(n_1895),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1909),
.Y(n_1942)
);

O2A1O1Ixp33_ASAP7_75t_L g1943 ( 
.A1(n_1935),
.A2(n_1867),
.B(n_1874),
.C(n_1892),
.Y(n_1943)
);

AOI22xp5_ASAP7_75t_L g1944 ( 
.A1(n_1907),
.A2(n_1897),
.B1(n_1867),
.B2(n_1812),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_L g1945 ( 
.A(n_1906),
.B(n_1868),
.Y(n_1945)
);

AOI21xp33_ASAP7_75t_SL g1946 ( 
.A1(n_1931),
.A2(n_1809),
.B(n_1654),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1910),
.Y(n_1947)
);

HB1xp67_ASAP7_75t_L g1948 ( 
.A(n_1906),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1910),
.Y(n_1949)
);

NAND2xp5_ASAP7_75t_L g1950 ( 
.A(n_1908),
.B(n_1869),
.Y(n_1950)
);

AND2x2_ASAP7_75t_L g1951 ( 
.A(n_1901),
.B(n_1880),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1912),
.Y(n_1952)
);

OR2x2_ASAP7_75t_L g1953 ( 
.A(n_1916),
.B(n_1883),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1912),
.Y(n_1954)
);

AND2x4_ASAP7_75t_L g1955 ( 
.A(n_1924),
.B(n_1823),
.Y(n_1955)
);

AOI22xp33_ASAP7_75t_L g1956 ( 
.A1(n_1936),
.A2(n_1823),
.B1(n_1819),
.B2(n_1810),
.Y(n_1956)
);

OAI221xp5_ASAP7_75t_L g1957 ( 
.A1(n_1936),
.A2(n_1874),
.B1(n_1888),
.B2(n_1856),
.C(n_1864),
.Y(n_1957)
);

OAI21xp5_ASAP7_75t_L g1958 ( 
.A1(n_1905),
.A2(n_1872),
.B(n_1869),
.Y(n_1958)
);

OAI22xp5_ASAP7_75t_SL g1959 ( 
.A1(n_1915),
.A2(n_1719),
.B1(n_1685),
.B2(n_1806),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1913),
.Y(n_1960)
);

NOR2xp33_ASAP7_75t_L g1961 ( 
.A(n_1905),
.B(n_1826),
.Y(n_1961)
);

OAI211xp5_ASAP7_75t_SL g1962 ( 
.A1(n_1920),
.A2(n_1856),
.B(n_1864),
.C(n_1891),
.Y(n_1962)
);

OR2x2_ASAP7_75t_L g1963 ( 
.A(n_1923),
.B(n_1826),
.Y(n_1963)
);

OR2x2_ASAP7_75t_L g1964 ( 
.A(n_1948),
.B(n_1945),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1945),
.Y(n_1965)
);

INVx2_ASAP7_75t_L g1966 ( 
.A(n_1955),
.Y(n_1966)
);

OAI31xp33_ASAP7_75t_L g1967 ( 
.A1(n_1961),
.A2(n_1917),
.A3(n_1900),
.B(n_1901),
.Y(n_1967)
);

NOR2xp33_ASAP7_75t_SL g1968 ( 
.A(n_1940),
.B(n_1784),
.Y(n_1968)
);

HB1xp67_ASAP7_75t_L g1969 ( 
.A(n_1955),
.Y(n_1969)
);

OAI22xp5_ASAP7_75t_L g1970 ( 
.A1(n_1959),
.A2(n_1929),
.B1(n_1933),
.B2(n_1900),
.Y(n_1970)
);

AND2x2_ASAP7_75t_L g1971 ( 
.A(n_1951),
.B(n_1919),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1937),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1942),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1947),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1949),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1952),
.Y(n_1976)
);

AOI22xp33_ASAP7_75t_L g1977 ( 
.A1(n_1956),
.A2(n_1919),
.B1(n_1927),
.B2(n_1926),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1954),
.Y(n_1978)
);

INVxp67_ASAP7_75t_SL g1979 ( 
.A(n_1938),
.Y(n_1979)
);

OAI22xp5_ASAP7_75t_L g1980 ( 
.A1(n_1944),
.A2(n_1899),
.B1(n_1904),
.B2(n_1926),
.Y(n_1980)
);

AND2x2_ASAP7_75t_L g1981 ( 
.A(n_1958),
.B(n_1927),
.Y(n_1981)
);

INVxp67_ASAP7_75t_L g1982 ( 
.A(n_1939),
.Y(n_1982)
);

INVx2_ASAP7_75t_SL g1983 ( 
.A(n_1939),
.Y(n_1983)
);

INVx2_ASAP7_75t_L g1984 ( 
.A(n_1963),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_L g1985 ( 
.A(n_1969),
.B(n_1950),
.Y(n_1985)
);

INVxp67_ASAP7_75t_SL g1986 ( 
.A(n_1964),
.Y(n_1986)
);

AOI22xp5_ASAP7_75t_L g1987 ( 
.A1(n_1979),
.A2(n_1962),
.B1(n_1957),
.B2(n_1899),
.Y(n_1987)
);

NOR3xp33_ASAP7_75t_L g1988 ( 
.A(n_1980),
.B(n_1943),
.C(n_1941),
.Y(n_1988)
);

AOI21xp5_ASAP7_75t_L g1989 ( 
.A1(n_1967),
.A2(n_1960),
.B(n_1950),
.Y(n_1989)
);

AOI322xp5_ASAP7_75t_L g1990 ( 
.A1(n_1981),
.A2(n_1930),
.A3(n_1932),
.B1(n_1899),
.B2(n_1914),
.C1(n_1925),
.C2(n_1913),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1964),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1972),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1972),
.Y(n_1993)
);

XOR2x2_ASAP7_75t_L g1994 ( 
.A(n_1981),
.B(n_1953),
.Y(n_1994)
);

OAI22xp5_ASAP7_75t_L g1995 ( 
.A1(n_1977),
.A2(n_1946),
.B1(n_1899),
.B2(n_1904),
.Y(n_1995)
);

OAI21xp5_ASAP7_75t_L g1996 ( 
.A1(n_1967),
.A2(n_1917),
.B(n_1914),
.Y(n_1996)
);

A2O1A1Ixp33_ASAP7_75t_L g1997 ( 
.A1(n_1968),
.A2(n_1917),
.B(n_1928),
.C(n_1930),
.Y(n_1997)
);

NAND3xp33_ASAP7_75t_L g1998 ( 
.A(n_1988),
.B(n_1982),
.C(n_1965),
.Y(n_1998)
);

NOR2x1_ASAP7_75t_L g1999 ( 
.A(n_1991),
.B(n_1992),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_L g2000 ( 
.A(n_1986),
.B(n_1966),
.Y(n_2000)
);

NOR2xp67_ASAP7_75t_L g2001 ( 
.A(n_1996),
.B(n_1983),
.Y(n_2001)
);

NOR2xp67_ASAP7_75t_L g2002 ( 
.A(n_1985),
.B(n_1983),
.Y(n_2002)
);

AOI211xp5_ASAP7_75t_L g2003 ( 
.A1(n_1989),
.A2(n_1970),
.B(n_1965),
.C(n_1966),
.Y(n_2003)
);

OR2x2_ASAP7_75t_L g2004 ( 
.A(n_1994),
.B(n_1984),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1993),
.Y(n_2005)
);

NAND4xp25_ASAP7_75t_L g2006 ( 
.A(n_1987),
.B(n_1984),
.C(n_1971),
.D(n_1976),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_SL g2007 ( 
.A(n_1997),
.B(n_1971),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_L g2008 ( 
.A(n_1990),
.B(n_1973),
.Y(n_2008)
);

NAND4xp25_ASAP7_75t_SL g2009 ( 
.A(n_2003),
.B(n_2008),
.C(n_1998),
.D(n_1989),
.Y(n_2009)
);

XNOR2x1_ASAP7_75t_L g2010 ( 
.A(n_2004),
.B(n_1995),
.Y(n_2010)
);

A2O1A1Ixp33_ASAP7_75t_L g2011 ( 
.A1(n_2001),
.A2(n_1978),
.B(n_1976),
.C(n_1975),
.Y(n_2011)
);

AOI211xp5_ASAP7_75t_L g2012 ( 
.A1(n_2006),
.A2(n_1975),
.B(n_1974),
.C(n_1973),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_L g2013 ( 
.A(n_2002),
.B(n_1974),
.Y(n_2013)
);

AOI22xp5_ASAP7_75t_L g2014 ( 
.A1(n_2007),
.A2(n_1978),
.B1(n_1932),
.B2(n_1922),
.Y(n_2014)
);

XNOR2xp5_ASAP7_75t_L g2015 ( 
.A(n_2010),
.B(n_2000),
.Y(n_2015)
);

INVxp67_ASAP7_75t_L g2016 ( 
.A(n_2013),
.Y(n_2016)
);

NOR2x1_ASAP7_75t_L g2017 ( 
.A(n_2009),
.B(n_1999),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_2011),
.Y(n_2018)
);

AOI22xp5_ASAP7_75t_L g2019 ( 
.A1(n_2014),
.A2(n_2005),
.B1(n_1921),
.B2(n_1918),
.Y(n_2019)
);

AOI221xp5_ASAP7_75t_L g2020 ( 
.A1(n_2012),
.A2(n_1925),
.B1(n_1922),
.B2(n_1921),
.C(n_1918),
.Y(n_2020)
);

AOI221xp5_ASAP7_75t_L g2021 ( 
.A1(n_2009),
.A2(n_1934),
.B1(n_1902),
.B2(n_1928),
.C(n_1893),
.Y(n_2021)
);

AOI22xp5_ASAP7_75t_L g2022 ( 
.A1(n_2015),
.A2(n_1934),
.B1(n_1902),
.B2(n_1893),
.Y(n_2022)
);

CKINVDCx16_ASAP7_75t_R g2023 ( 
.A(n_2017),
.Y(n_2023)
);

XOR2xp5_ASAP7_75t_L g2024 ( 
.A(n_2018),
.B(n_1682),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_2019),
.Y(n_2025)
);

NOR2x1_ASAP7_75t_L g2026 ( 
.A(n_2016),
.B(n_1902),
.Y(n_2026)
);

NOR2x1_ASAP7_75t_L g2027 ( 
.A(n_2021),
.B(n_1934),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_L g2028 ( 
.A(n_2023),
.B(n_2020),
.Y(n_2028)
);

NOR2x1_ASAP7_75t_L g2029 ( 
.A(n_2026),
.B(n_1872),
.Y(n_2029)
);

AOI221xp5_ASAP7_75t_L g2030 ( 
.A1(n_2025),
.A2(n_1892),
.B1(n_1891),
.B2(n_1889),
.C(n_1876),
.Y(n_2030)
);

NOR2x1_ASAP7_75t_L g2031 ( 
.A(n_2027),
.B(n_1876),
.Y(n_2031)
);

INVx2_ASAP7_75t_L g2032 ( 
.A(n_2029),
.Y(n_2032)
);

AOI22xp33_ASAP7_75t_L g2033 ( 
.A1(n_2032),
.A2(n_2024),
.B1(n_2028),
.B2(n_2031),
.Y(n_2033)
);

OAI22xp5_ASAP7_75t_L g2034 ( 
.A1(n_2033),
.A2(n_2022),
.B1(n_2030),
.B2(n_1889),
.Y(n_2034)
);

OAI22x1_ASAP7_75t_L g2035 ( 
.A1(n_2033),
.A2(n_1884),
.B1(n_1879),
.B2(n_1854),
.Y(n_2035)
);

OAI22xp5_ASAP7_75t_L g2036 ( 
.A1(n_2034),
.A2(n_1884),
.B1(n_1879),
.B2(n_1870),
.Y(n_2036)
);

OAI22xp5_ASAP7_75t_L g2037 ( 
.A1(n_2035),
.A2(n_1870),
.B1(n_1854),
.B2(n_1819),
.Y(n_2037)
);

AOI21xp5_ASAP7_75t_L g2038 ( 
.A1(n_2036),
.A2(n_1654),
.B(n_1886),
.Y(n_2038)
);

OAI21x1_ASAP7_75t_SL g2039 ( 
.A1(n_2037),
.A2(n_1655),
.B(n_1665),
.Y(n_2039)
);

OAI21xp5_ASAP7_75t_L g2040 ( 
.A1(n_2038),
.A2(n_1887),
.B(n_1823),
.Y(n_2040)
);

AO21x2_ASAP7_75t_L g2041 ( 
.A1(n_2040),
.A2(n_2039),
.B(n_1887),
.Y(n_2041)
);

BUFx3_ASAP7_75t_L g2042 ( 
.A(n_2041),
.Y(n_2042)
);

AOI221xp5_ASAP7_75t_L g2043 ( 
.A1(n_2042),
.A2(n_1851),
.B1(n_1846),
.B2(n_1836),
.C(n_1852),
.Y(n_2043)
);

AOI211xp5_ASAP7_75t_L g2044 ( 
.A1(n_2043),
.A2(n_1659),
.B(n_1661),
.C(n_1590),
.Y(n_2044)
);


endmodule