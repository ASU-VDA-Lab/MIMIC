module fake_jpeg_2783_n_97 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_97);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_97;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_10),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_9),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_7),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_10),
.B(n_5),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_25),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_21),
.B(n_4),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_26),
.B(n_27),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_11),
.B(n_4),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVx4_ASAP7_75t_SL g29 ( 
.A(n_20),
.Y(n_29)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

CKINVDCx12_ASAP7_75t_R g38 ( 
.A(n_31),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_0),
.Y(n_32)
);

NOR2x1_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_22),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_16),
.B(n_0),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_0),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_24),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_35),
.B(n_39),
.Y(n_56)
);

AO22x1_ASAP7_75t_L g36 ( 
.A1(n_32),
.A2(n_22),
.B1(n_19),
.B2(n_15),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_36),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_45),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_15),
.Y(n_45)
);

INVx3_ASAP7_75t_SL g46 ( 
.A(n_42),
.Y(n_46)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_41),
.A2(n_28),
.B1(n_23),
.B2(n_31),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_48),
.A2(n_36),
.B1(n_39),
.B2(n_12),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_35),
.A2(n_29),
.B1(n_14),
.B2(n_13),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_50),
.A2(n_54),
.B(n_43),
.Y(n_59)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_52),
.Y(n_62)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_40),
.A2(n_14),
.B1(n_13),
.B2(n_11),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_58),
.Y(n_66)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_57),
.B(n_36),
.Y(n_60)
);

INVx4_ASAP7_75t_SL g58 ( 
.A(n_37),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_59),
.B(n_46),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_60),
.B(n_61),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_47),
.B(n_45),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_64),
.A2(n_56),
.B1(n_58),
.B2(n_57),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g65 ( 
.A(n_53),
.B(n_44),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_65),
.B(n_68),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_44),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_64),
.A2(n_56),
.B1(n_52),
.B2(n_23),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_74),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_71),
.A2(n_66),
.B(n_65),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_72),
.A2(n_75),
.B(n_73),
.Y(n_81)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g75 ( 
.A1(n_68),
.A2(n_51),
.B(n_55),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_76),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_75),
.Y(n_77)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_77),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_80),
.A2(n_72),
.B1(n_30),
.B2(n_31),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_81),
.B(n_38),
.Y(n_86)
);

MAJx2_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_63),
.C(n_12),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_82),
.B(n_70),
.C(n_78),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_84),
.A2(n_86),
.B(n_79),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_85),
.A2(n_49),
.B1(n_25),
.B2(n_67),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_SL g91 ( 
.A(n_87),
.B(n_86),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_88),
.Y(n_92)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_83),
.Y(n_89)
);

INVxp33_ASAP7_75t_L g90 ( 
.A(n_89),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_91),
.B(n_92),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_90),
.A2(n_84),
.B(n_82),
.Y(n_93)
);

AOI322xp5_ASAP7_75t_L g95 ( 
.A1(n_93),
.A2(n_94),
.A3(n_67),
.B1(n_30),
.B2(n_17),
.C1(n_8),
.C2(n_7),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_17),
.C(n_6),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_8),
.Y(n_97)
);


endmodule