module fake_jpeg_9187_n_102 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_102);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_102;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

BUFx16f_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_18),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_15),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

CKINVDCx5p33_ASAP7_75t_R g49 ( 
.A(n_7),
.Y(n_49)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_49),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_53),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_41),
.Y(n_53)
);

BUFx12_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_0),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_0),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx4_ASAP7_75t_SL g57 ( 
.A(n_38),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_59),
.Y(n_63)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_60),
.B(n_61),
.Y(n_62)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_60),
.A2(n_44),
.B1(n_51),
.B2(n_46),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_64),
.A2(n_72),
.B1(n_73),
.B2(n_74),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_56),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_65),
.B(n_69),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_61),
.B(n_47),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_70),
.Y(n_81)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_55),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_71),
.B(n_75),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_60),
.A2(n_43),
.B1(n_38),
.B2(n_40),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_60),
.A2(n_43),
.B1(n_21),
.B2(n_24),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_60),
.A2(n_19),
.B1(n_36),
.B2(n_35),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_1),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_60),
.A2(n_17),
.B1(n_34),
.B2(n_33),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_76),
.A2(n_77),
.B1(n_4),
.B2(n_5),
.Y(n_80)
);

OA22x2_ASAP7_75t_L g77 ( 
.A1(n_53),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_57),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_78),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_82),
.Y(n_89)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_62),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_83),
.B(n_85),
.Y(n_90)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_62),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_90),
.B(n_81),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_91),
.B(n_84),
.Y(n_92)
);

OA21x2_ASAP7_75t_L g93 ( 
.A1(n_92),
.A2(n_87),
.B(n_89),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_93),
.B(n_86),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_80),
.C(n_67),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_95),
.A2(n_77),
.B(n_68),
.Y(n_96)
);

AOI21x1_ASAP7_75t_L g97 ( 
.A1(n_96),
.A2(n_88),
.B(n_79),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_88),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_98),
.A2(n_85),
.B1(n_13),
.B2(n_16),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_99),
.A2(n_12),
.B(n_20),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_100),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_31),
.Y(n_102)
);


endmodule