module real_aes_3367_n_6 (n_4, n_0, n_3, n_5, n_2, n_1, n_6);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_1;
output n_6;
wire n_17;
wire n_22;
wire n_13;
wire n_24;
wire n_12;
wire n_19;
wire n_14;
wire n_11;
wire n_16;
wire n_15;
wire n_9;
wire n_23;
wire n_20;
wire n_18;
wire n_21;
wire n_7;
wire n_8;
wire n_10;
NAND3xp33_ASAP7_75t_SL g11 ( .A(n_0), .B(n_12), .C(n_14), .Y(n_11) );
HB1xp67_ASAP7_75t_L g13 ( .A(n_1), .Y(n_13) );
INVx1_ASAP7_75t_L g8 ( .A(n_2), .Y(n_8) );
BUFx6f_ASAP7_75t_L g16 ( .A(n_3), .Y(n_16) );
INVx2_ASAP7_75t_SL g19 ( .A(n_4), .Y(n_19) );
HB1xp67_ASAP7_75t_L g21 ( .A(n_5), .Y(n_21) );
AOI22xp5_ASAP7_75t_L g6 ( .A1(n_7), .A2(n_9), .B1(n_22), .B2(n_23), .Y(n_6) );
CKINVDCx20_ASAP7_75t_R g22 ( .A(n_7), .Y(n_22) );
INVxp67_ASAP7_75t_L g7 ( .A(n_8), .Y(n_7) );
CKINVDCx20_ASAP7_75t_R g9 ( .A(n_10), .Y(n_9) );
AOI21xp5_ASAP7_75t_L g10 ( .A1(n_11), .A2(n_17), .B(n_20), .Y(n_10) );
INVx1_ASAP7_75t_L g12 ( .A(n_13), .Y(n_12) );
BUFx2_ASAP7_75t_L g14 ( .A(n_15), .Y(n_14) );
HB1xp67_ASAP7_75t_L g15 ( .A(n_16), .Y(n_15) );
NOR2xp33_ASAP7_75t_L g20 ( .A(n_17), .B(n_21), .Y(n_20) );
NOR2xp33_ASAP7_75t_L g23 ( .A(n_17), .B(n_24), .Y(n_23) );
HB1xp67_ASAP7_75t_L g17 ( .A(n_18), .Y(n_17) );
HB1xp67_ASAP7_75t_L g18 ( .A(n_19), .Y(n_18) );
CKINVDCx5p33_ASAP7_75t_R g24 ( .A(n_21), .Y(n_24) );
endmodule