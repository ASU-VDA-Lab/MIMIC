module fake_netlist_6_10_n_563 (n_52, n_16, n_1, n_91, n_119, n_46, n_18, n_21, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_125, n_77, n_106, n_92, n_42, n_96, n_8, n_90, n_24, n_105, n_54, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_100, n_13, n_121, n_11, n_17, n_23, n_20, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_41, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_563);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_125;
input n_77;
input n_106;
input n_92;
input n_42;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_54;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_100;
input n_13;
input n_121;
input n_11;
input n_17;
input n_23;
input n_20;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_41;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_563;

wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_507;
wire n_209;
wire n_367;
wire n_465;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_148;
wire n_161;
wire n_208;
wire n_462;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_144;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_524;
wire n_342;
wire n_358;
wire n_160;
wire n_449;
wire n_131;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_396;
wire n_495;
wire n_350;
wire n_392;
wire n_442;
wire n_480;
wire n_142;
wire n_143;
wire n_382;
wire n_180;
wire n_557;
wire n_349;
wire n_233;
wire n_255;
wire n_284;
wire n_400;
wire n_140;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_471;
wire n_289;
wire n_421;
wire n_424;
wire n_181;
wire n_182;
wire n_238;
wire n_202;
wire n_320;
wire n_327;
wire n_369;
wire n_280;
wire n_287;
wire n_353;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_461;
wire n_141;
wire n_383;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_222;
wire n_179;
wire n_248;
wire n_300;
wire n_517;
wire n_229;
wire n_542;
wire n_305;
wire n_532;
wire n_173;
wire n_535;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_510;
wire n_375;
wire n_338;
wire n_522;
wire n_466;
wire n_506;
wire n_360;
wire n_235;
wire n_536;
wire n_147;
wire n_191;
wire n_340;
wire n_387;
wire n_452;
wire n_344;
wire n_428;
wire n_432;
wire n_167;
wire n_174;
wire n_127;
wire n_516;
wire n_153;
wire n_525;
wire n_156;
wire n_491;
wire n_145;
wire n_133;
wire n_371;
wire n_189;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_129;
wire n_197;
wire n_137;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_155;
wire n_529;
wire n_445;
wire n_425;
wire n_454;
wire n_218;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_172;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_196;
wire n_402;
wire n_352;
wire n_478;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_374;
wire n_366;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_348;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_163;
wire n_330;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_154;
wire n_456;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_279;
wire n_252;
wire n_228;
wire n_356;
wire n_166;
wire n_184;
wire n_552;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_395;
wire n_323;
wire n_393;
wire n_411;
wire n_503;
wire n_152;
wire n_513;
wire n_321;
wire n_331;
wire n_227;
wire n_132;
wire n_406;
wire n_483;
wire n_204;
wire n_482;
wire n_527;
wire n_474;
wire n_261;
wire n_420;
wire n_312;
wire n_394;
wire n_130;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_150;
wire n_264;
wire n_263;
wire n_481;
wire n_325;
wire n_329;
wire n_464;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_505;
wire n_240;
wire n_139;
wire n_319;
wire n_134;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_311;
wire n_403;
wire n_253;
wire n_136;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_556;
wire n_159;
wire n_157;
wire n_162;
wire n_487;
wire n_550;
wire n_128;
wire n_241;
wire n_275;
wire n_553;
wire n_560;
wire n_276;
wire n_441;
wire n_221;
wire n_444;
wire n_423;
wire n_146;
wire n_318;
wire n_303;
wire n_511;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_199;
wire n_138;
wire n_266;
wire n_296;
wire n_268;
wire n_271;
wire n_404;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_453;
wire n_333;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_355;
wire n_426;
wire n_317;
wire n_149;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_257;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_401;
wire n_324;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_251;
wire n_301;
wire n_274;
wire n_151;
wire n_412;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_422;
wire n_135;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_514;
wire n_528;
wire n_391;
wire n_457;
wire n_364;
wire n_295;
wire n_385;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_554;
wire n_194;
wire n_171;
wire n_192;
wire n_169;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g127 ( 
.A(n_100),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_52),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_42),
.Y(n_129)
);

CKINVDCx5p33_ASAP7_75t_R g130 ( 
.A(n_23),
.Y(n_130)
);

CKINVDCx5p33_ASAP7_75t_R g131 ( 
.A(n_58),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_80),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_93),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_13),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_111),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_106),
.Y(n_136)
);

CKINVDCx5p33_ASAP7_75t_R g137 ( 
.A(n_27),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_76),
.Y(n_138)
);

CKINVDCx5p33_ASAP7_75t_R g139 ( 
.A(n_55),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_34),
.Y(n_140)
);

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_63),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_72),
.Y(n_142)
);

CKINVDCx5p33_ASAP7_75t_R g143 ( 
.A(n_96),
.Y(n_143)
);

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_19),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_120),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_31),
.Y(n_146)
);

CKINVDCx5p33_ASAP7_75t_R g147 ( 
.A(n_66),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_43),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_41),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_70),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_50),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_113),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_123),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_51),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_7),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_119),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_40),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_122),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_104),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_12),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_117),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_115),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_71),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_107),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_18),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_0),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_29),
.Y(n_167)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_118),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_5),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_98),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_124),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_90),
.Y(n_172)
);

BUFx2_ASAP7_75t_L g173 ( 
.A(n_9),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_26),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_36),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_87),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_57),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_68),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_44),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_67),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_17),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_69),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_14),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_28),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_62),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_125),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g187 ( 
.A(n_3),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_59),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_22),
.Y(n_189)
);

BUFx12f_ASAP7_75t_L g190 ( 
.A(n_173),
.Y(n_190)
);

INVx5_ASAP7_75t_L g191 ( 
.A(n_168),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_182),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_155),
.B(n_0),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g194 ( 
.A(n_134),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_182),
.Y(n_195)
);

AND2x6_ASAP7_75t_L g196 ( 
.A(n_168),
.B(n_15),
.Y(n_196)
);

BUFx8_ASAP7_75t_L g197 ( 
.A(n_160),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_169),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_128),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_127),
.Y(n_200)
);

BUFx12f_ASAP7_75t_L g201 ( 
.A(n_130),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_168),
.Y(n_202)
);

BUFx2_ASAP7_75t_L g203 ( 
.A(n_166),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_142),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_129),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_132),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_187),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_166),
.Y(n_208)
);

OAI22x1_ASAP7_75t_L g209 ( 
.A1(n_180),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_209)
);

BUFx12f_ASAP7_75t_L g210 ( 
.A(n_131),
.Y(n_210)
);

INVx2_ASAP7_75t_SL g211 ( 
.A(n_137),
.Y(n_211)
);

OAI21x1_ASAP7_75t_L g212 ( 
.A1(n_142),
.A2(n_64),
.B(n_121),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_128),
.B(n_4),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_177),
.B(n_5),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_164),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_177),
.B(n_6),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_139),
.Y(n_217)
);

NAND2x1p5_ASAP7_75t_L g218 ( 
.A(n_133),
.B(n_135),
.Y(n_218)
);

OAI21x1_ASAP7_75t_L g219 ( 
.A1(n_138),
.A2(n_65),
.B(n_116),
.Y(n_219)
);

NOR2x1_ASAP7_75t_L g220 ( 
.A(n_140),
.B(n_16),
.Y(n_220)
);

AND2x6_ASAP7_75t_L g221 ( 
.A(n_145),
.B(n_20),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_146),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_154),
.Y(n_223)
);

BUFx8_ASAP7_75t_SL g224 ( 
.A(n_164),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_156),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_158),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_141),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_136),
.B(n_8),
.Y(n_228)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_161),
.Y(n_229)
);

AND2x4_ASAP7_75t_L g230 ( 
.A(n_163),
.B(n_9),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_167),
.B(n_10),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_165),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_165),
.B(n_188),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_170),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_207),
.Y(n_235)
);

INVxp33_ASAP7_75t_L g236 ( 
.A(n_207),
.Y(n_236)
);

INVx2_ASAP7_75t_SL g237 ( 
.A(n_190),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_204),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_204),
.Y(n_239)
);

AND2x6_ASAP7_75t_L g240 ( 
.A(n_213),
.B(n_171),
.Y(n_240)
);

AND2x2_ASAP7_75t_SL g241 ( 
.A(n_199),
.B(n_172),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_228),
.A2(n_233),
.B1(n_193),
.B2(n_217),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_192),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_192),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g245 ( 
.A(n_192),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_211),
.B(n_179),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_195),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_225),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_225),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_225),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_230),
.B(n_188),
.Y(n_251)
);

INVx2_ASAP7_75t_SL g252 ( 
.A(n_197),
.Y(n_252)
);

BUFx2_ASAP7_75t_L g253 ( 
.A(n_224),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_230),
.B(n_175),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_200),
.B(n_227),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_195),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_195),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_206),
.Y(n_258)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_222),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_201),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_226),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_191),
.B(n_183),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_205),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_223),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_202),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_229),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_229),
.Y(n_267)
);

OR2x2_ASAP7_75t_L g268 ( 
.A(n_234),
.B(n_11),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_203),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_218),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_231),
.B(n_143),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_228),
.B(n_185),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_191),
.B(n_186),
.Y(n_273)
);

NAND3xp33_ASAP7_75t_L g274 ( 
.A(n_234),
.B(n_157),
.C(n_184),
.Y(n_274)
);

INVx5_ASAP7_75t_L g275 ( 
.A(n_196),
.Y(n_275)
);

CKINVDCx6p67_ASAP7_75t_R g276 ( 
.A(n_210),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_218),
.B(n_189),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_272),
.B(n_214),
.Y(n_278)
);

OR2x2_ASAP7_75t_L g279 ( 
.A(n_235),
.B(n_233),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_236),
.B(n_194),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_245),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_272),
.B(n_196),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_255),
.B(n_196),
.Y(n_283)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_245),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_242),
.B(n_214),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_271),
.B(n_221),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_246),
.B(n_216),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_270),
.B(n_216),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_271),
.B(n_277),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_239),
.B(n_221),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_275),
.B(n_241),
.Y(n_291)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_238),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_236),
.B(n_194),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_274),
.B(n_193),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_264),
.Y(n_295)
);

A2O1A1Ixp33_ASAP7_75t_L g296 ( 
.A1(n_235),
.A2(n_219),
.B(n_212),
.C(n_220),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_275),
.B(n_144),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_243),
.Y(n_298)
);

AND2x4_ASAP7_75t_L g299 ( 
.A(n_244),
.B(n_198),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_256),
.B(n_263),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_L g301 ( 
.A1(n_241),
.A2(n_221),
.B1(n_209),
.B2(n_198),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_247),
.B(n_147),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_238),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_251),
.B(n_148),
.Y(n_304)
);

NOR2xp67_ASAP7_75t_L g305 ( 
.A(n_237),
.B(n_149),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_257),
.B(n_150),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_251),
.B(n_151),
.Y(n_307)
);

NOR2xp67_ASAP7_75t_L g308 ( 
.A(n_252),
.B(n_152),
.Y(n_308)
);

OR2x2_ASAP7_75t_L g309 ( 
.A(n_269),
.B(n_208),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_265),
.B(n_153),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_259),
.B(n_267),
.Y(n_311)
);

HB1xp67_ASAP7_75t_L g312 ( 
.A(n_268),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_275),
.B(n_159),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_259),
.B(n_208),
.Y(n_314)
);

AOI221xp5_ASAP7_75t_L g315 ( 
.A1(n_254),
.A2(n_215),
.B1(n_232),
.B2(n_176),
.C(n_181),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_L g316 ( 
.A1(n_240),
.A2(n_215),
.B1(n_197),
.B2(n_178),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_254),
.B(n_174),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_238),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_258),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_261),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_248),
.Y(n_321)
);

NAND3xp33_ASAP7_75t_L g322 ( 
.A(n_261),
.B(n_162),
.C(n_13),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_248),
.Y(n_323)
);

NAND2xp33_ASAP7_75t_SL g324 ( 
.A(n_262),
.B(n_21),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_240),
.B(n_24),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_275),
.B(n_25),
.Y(n_326)
);

NAND3xp33_ASAP7_75t_L g327 ( 
.A(n_266),
.B(n_30),
.C(n_32),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_280),
.B(n_276),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_278),
.B(n_273),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_278),
.A2(n_266),
.B1(n_265),
.B2(n_260),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_294),
.B(n_250),
.Y(n_331)
);

OAI21x1_ASAP7_75t_L g332 ( 
.A1(n_290),
.A2(n_250),
.B(n_249),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_311),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_285),
.A2(n_250),
.B1(n_249),
.B2(n_248),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_289),
.B(n_253),
.Y(n_335)
);

AOI21xp33_ASAP7_75t_L g336 ( 
.A1(n_294),
.A2(n_249),
.B(n_248),
.Y(n_336)
);

INVx4_ASAP7_75t_L g337 ( 
.A(n_284),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_282),
.A2(n_249),
.B(n_35),
.Y(n_338)
);

INVx4_ASAP7_75t_L g339 ( 
.A(n_284),
.Y(n_339)
);

OAI21x1_ASAP7_75t_SL g340 ( 
.A1(n_301),
.A2(n_283),
.B(n_286),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_288),
.A2(n_33),
.B(n_37),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_288),
.A2(n_38),
.B(n_39),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_309),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_L g344 ( 
.A1(n_287),
.A2(n_45),
.B(n_46),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_285),
.B(n_47),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_320),
.Y(n_346)
);

BUFx2_ASAP7_75t_L g347 ( 
.A(n_293),
.Y(n_347)
);

OAI321xp33_ASAP7_75t_L g348 ( 
.A1(n_301),
.A2(n_48),
.A3(n_49),
.B1(n_53),
.B2(n_54),
.C(n_56),
.Y(n_348)
);

INVx2_ASAP7_75t_SL g349 ( 
.A(n_314),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_310),
.B(n_60),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_310),
.B(n_61),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_295),
.B(n_73),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_281),
.Y(n_353)
);

O2A1O1Ixp33_ASAP7_75t_L g354 ( 
.A1(n_291),
.A2(n_74),
.B(n_75),
.C(n_77),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_302),
.B(n_306),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_279),
.B(n_78),
.Y(n_356)
);

NAND3xp33_ASAP7_75t_L g357 ( 
.A(n_315),
.B(n_79),
.C(n_81),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_291),
.A2(n_82),
.B1(n_83),
.B2(n_84),
.Y(n_358)
);

NOR2xp67_ASAP7_75t_L g359 ( 
.A(n_305),
.B(n_126),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_302),
.B(n_85),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_304),
.B(n_307),
.Y(n_361)
);

AOI21xp5_ASAP7_75t_L g362 ( 
.A1(n_297),
.A2(n_86),
.B(n_88),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_317),
.B(n_89),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_299),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_312),
.B(n_91),
.Y(n_365)
);

HB1xp67_ASAP7_75t_L g366 ( 
.A(n_299),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_300),
.Y(n_367)
);

AND2x2_ASAP7_75t_L g368 ( 
.A(n_300),
.B(n_92),
.Y(n_368)
);

OAI21xp33_ASAP7_75t_L g369 ( 
.A1(n_316),
.A2(n_94),
.B(n_95),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_316),
.B(n_97),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_306),
.B(n_99),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_321),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_297),
.A2(n_313),
.B(n_296),
.Y(n_373)
);

INVx3_ASAP7_75t_L g374 ( 
.A(n_292),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_319),
.B(n_101),
.Y(n_375)
);

A2O1A1Ixp33_ASAP7_75t_L g376 ( 
.A1(n_325),
.A2(n_102),
.B(n_103),
.C(n_105),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_298),
.B(n_308),
.Y(n_377)
);

AOI21xp5_ASAP7_75t_L g378 ( 
.A1(n_313),
.A2(n_108),
.B(n_109),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_322),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_323),
.B(n_318),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_303),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_329),
.B(n_326),
.Y(n_382)
);

NOR2xp67_ASAP7_75t_L g383 ( 
.A(n_357),
.B(n_327),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_355),
.B(n_326),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_367),
.B(n_324),
.Y(n_385)
);

AO31x2_ASAP7_75t_L g386 ( 
.A1(n_373),
.A2(n_110),
.A3(n_112),
.B(n_114),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_346),
.Y(n_387)
);

A2O1A1Ixp33_ASAP7_75t_L g388 ( 
.A1(n_361),
.A2(n_369),
.B(n_363),
.C(n_345),
.Y(n_388)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_347),
.B(n_349),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_368),
.B(n_333),
.Y(n_390)
);

OAI21x1_ASAP7_75t_L g391 ( 
.A1(n_332),
.A2(n_334),
.B(n_374),
.Y(n_391)
);

INVx3_ASAP7_75t_L g392 ( 
.A(n_372),
.Y(n_392)
);

OAI21x1_ASAP7_75t_L g393 ( 
.A1(n_374),
.A2(n_340),
.B(n_381),
.Y(n_393)
);

BUFx2_ASAP7_75t_L g394 ( 
.A(n_364),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g395 ( 
.A1(n_331),
.A2(n_336),
.B(n_350),
.Y(n_395)
);

NOR2x1_ASAP7_75t_L g396 ( 
.A(n_344),
.B(n_371),
.Y(n_396)
);

AOI221xp5_ASAP7_75t_L g397 ( 
.A1(n_369),
.A2(n_370),
.B1(n_348),
.B2(n_335),
.C(n_365),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_379),
.A2(n_360),
.B1(n_351),
.B2(n_338),
.Y(n_398)
);

NOR2x1_ASAP7_75t_SL g399 ( 
.A(n_356),
.B(n_352),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_377),
.B(n_353),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_L g401 ( 
.A1(n_380),
.A2(n_330),
.B(n_342),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_L g402 ( 
.A1(n_341),
.A2(n_354),
.B(n_375),
.Y(n_402)
);

AO31x2_ASAP7_75t_L g403 ( 
.A1(n_376),
.A2(n_358),
.A3(n_362),
.B(n_378),
.Y(n_403)
);

BUFx6f_ASAP7_75t_SL g404 ( 
.A(n_364),
.Y(n_404)
);

BUFx2_ASAP7_75t_L g405 ( 
.A(n_364),
.Y(n_405)
);

AOI21xp5_ASAP7_75t_L g406 ( 
.A1(n_372),
.A2(n_359),
.B(n_366),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_337),
.B(n_339),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_343),
.Y(n_408)
);

BUFx8_ASAP7_75t_L g409 ( 
.A(n_328),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_329),
.B(n_278),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_355),
.A2(n_278),
.B1(n_329),
.B2(n_285),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_329),
.B(n_278),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_349),
.B(n_364),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_346),
.Y(n_414)
);

OAI21x1_ASAP7_75t_L g415 ( 
.A1(n_402),
.A2(n_395),
.B(n_401),
.Y(n_415)
);

OAI21x1_ASAP7_75t_L g416 ( 
.A1(n_398),
.A2(n_396),
.B(n_406),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_L g417 ( 
.A1(n_388),
.A2(n_411),
.B(n_410),
.Y(n_417)
);

AOI21x1_ASAP7_75t_L g418 ( 
.A1(n_396),
.A2(n_382),
.B(n_384),
.Y(n_418)
);

AOI22x1_ASAP7_75t_L g419 ( 
.A1(n_387),
.A2(n_414),
.B1(n_397),
.B2(n_392),
.Y(n_419)
);

OAI21x1_ASAP7_75t_L g420 ( 
.A1(n_392),
.A2(n_390),
.B(n_383),
.Y(n_420)
);

BUFx4f_ASAP7_75t_L g421 ( 
.A(n_408),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_386),
.Y(n_422)
);

NAND2x1p5_ASAP7_75t_L g423 ( 
.A(n_383),
.B(n_405),
.Y(n_423)
);

OAI21x1_ASAP7_75t_L g424 ( 
.A1(n_407),
.A2(n_385),
.B(n_413),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_412),
.B(n_400),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_386),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_386),
.Y(n_427)
);

OAI21x1_ASAP7_75t_L g428 ( 
.A1(n_403),
.A2(n_399),
.B(n_389),
.Y(n_428)
);

INVx1_ASAP7_75t_SL g429 ( 
.A(n_408),
.Y(n_429)
);

NAND2x1p5_ASAP7_75t_L g430 ( 
.A(n_394),
.B(n_408),
.Y(n_430)
);

AO21x2_ASAP7_75t_L g431 ( 
.A1(n_403),
.A2(n_404),
.B(n_409),
.Y(n_431)
);

O2A1O1Ixp33_ASAP7_75t_L g432 ( 
.A1(n_404),
.A2(n_411),
.B(n_388),
.C(n_410),
.Y(n_432)
);

OAI21x1_ASAP7_75t_L g433 ( 
.A1(n_409),
.A2(n_393),
.B(n_391),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_393),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_393),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_393),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_410),
.B(n_412),
.Y(n_437)
);

HB1xp67_ASAP7_75t_L g438 ( 
.A(n_408),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_425),
.B(n_437),
.Y(n_439)
);

NAND2x1p5_ASAP7_75t_L g440 ( 
.A(n_433),
.B(n_428),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_435),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_425),
.B(n_417),
.Y(n_442)
);

AO21x1_ASAP7_75t_SL g443 ( 
.A1(n_427),
.A2(n_417),
.B(n_434),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_436),
.Y(n_444)
);

BUFx2_ASAP7_75t_L g445 ( 
.A(n_438),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_419),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_423),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_423),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_434),
.Y(n_449)
);

INVx3_ASAP7_75t_L g450 ( 
.A(n_433),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_423),
.Y(n_451)
);

OR2x6_ASAP7_75t_L g452 ( 
.A(n_432),
.B(n_428),
.Y(n_452)
);

BUFx2_ASAP7_75t_L g453 ( 
.A(n_421),
.Y(n_453)
);

BUFx6f_ASAP7_75t_L g454 ( 
.A(n_421),
.Y(n_454)
);

BUFx3_ASAP7_75t_L g455 ( 
.A(n_421),
.Y(n_455)
);

BUFx2_ASAP7_75t_L g456 ( 
.A(n_430),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_431),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_424),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_419),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_442),
.B(n_431),
.Y(n_460)
);

BUFx2_ASAP7_75t_L g461 ( 
.A(n_456),
.Y(n_461)
);

BUFx3_ASAP7_75t_L g462 ( 
.A(n_455),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_449),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_439),
.B(n_429),
.Y(n_464)
);

OR2x2_ASAP7_75t_L g465 ( 
.A(n_442),
.B(n_431),
.Y(n_465)
);

HB1xp67_ASAP7_75t_L g466 ( 
.A(n_445),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_L g467 ( 
.A1(n_439),
.A2(n_429),
.B1(n_430),
.B2(n_427),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_449),
.Y(n_468)
);

INVx3_ASAP7_75t_L g469 ( 
.A(n_450),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_445),
.B(n_430),
.Y(n_470)
);

AND2x2_ASAP7_75t_L g471 ( 
.A(n_456),
.B(n_424),
.Y(n_471)
);

OR2x2_ASAP7_75t_L g472 ( 
.A(n_452),
.B(n_415),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_447),
.B(n_426),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_441),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_444),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_448),
.B(n_426),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_454),
.Y(n_477)
);

NOR2x1_ASAP7_75t_L g478 ( 
.A(n_455),
.B(n_422),
.Y(n_478)
);

INVx3_ASAP7_75t_L g479 ( 
.A(n_450),
.Y(n_479)
);

BUFx3_ASAP7_75t_L g480 ( 
.A(n_454),
.Y(n_480)
);

BUFx2_ASAP7_75t_L g481 ( 
.A(n_451),
.Y(n_481)
);

INVxp67_ASAP7_75t_SL g482 ( 
.A(n_453),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_446),
.B(n_422),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_458),
.Y(n_484)
);

INVxp67_ASAP7_75t_SL g485 ( 
.A(n_466),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_460),
.B(n_443),
.Y(n_486)
);

NOR2x1_ASAP7_75t_SL g487 ( 
.A(n_472),
.B(n_443),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_460),
.B(n_452),
.Y(n_488)
);

AOI22xp33_ASAP7_75t_SL g489 ( 
.A1(n_467),
.A2(n_415),
.B1(n_453),
.B2(n_454),
.Y(n_489)
);

INVx1_ASAP7_75t_SL g490 ( 
.A(n_464),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_465),
.B(n_452),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_468),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_468),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_484),
.Y(n_494)
);

HB1xp67_ASAP7_75t_L g495 ( 
.A(n_461),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_484),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_470),
.B(n_454),
.Y(n_497)
);

HB1xp67_ASAP7_75t_L g498 ( 
.A(n_461),
.Y(n_498)
);

AND2x2_ASAP7_75t_L g499 ( 
.A(n_465),
.B(n_452),
.Y(n_499)
);

INVx2_ASAP7_75t_SL g500 ( 
.A(n_481),
.Y(n_500)
);

INVxp67_ASAP7_75t_SL g501 ( 
.A(n_482),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g502 ( 
.A(n_471),
.B(n_457),
.Y(n_502)
);

OR2x2_ASAP7_75t_L g503 ( 
.A(n_472),
.B(n_457),
.Y(n_503)
);

NAND2x1p5_ASAP7_75t_L g504 ( 
.A(n_478),
.B(n_450),
.Y(n_504)
);

AND2x2_ASAP7_75t_L g505 ( 
.A(n_471),
.B(n_463),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_462),
.B(n_459),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_463),
.B(n_473),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_494),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_490),
.B(n_481),
.Y(n_509)
);

OAI221xp5_ASAP7_75t_L g510 ( 
.A1(n_489),
.A2(n_462),
.B1(n_454),
.B2(n_480),
.C(n_446),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_485),
.B(n_473),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_494),
.Y(n_512)
);

AND2x4_ASAP7_75t_SL g513 ( 
.A(n_495),
.B(n_477),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_496),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_486),
.B(n_457),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_507),
.B(n_476),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_496),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_486),
.B(n_476),
.Y(n_518)
);

NOR2xp67_ASAP7_75t_SL g519 ( 
.A(n_506),
.B(n_477),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_502),
.B(n_457),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_502),
.B(n_457),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_507),
.B(n_483),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_512),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_512),
.Y(n_524)
);

AND2x4_ASAP7_75t_L g525 ( 
.A(n_520),
.B(n_487),
.Y(n_525)
);

NAND4xp75_ASAP7_75t_L g526 ( 
.A(n_509),
.B(n_497),
.C(n_500),
.D(n_499),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_508),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_514),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_517),
.Y(n_529)
);

AO221x1_ASAP7_75t_L g530 ( 
.A1(n_510),
.A2(n_469),
.B1(n_479),
.B2(n_459),
.C(n_477),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_528),
.B(n_509),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_527),
.Y(n_532)
);

AND2x2_ASAP7_75t_L g533 ( 
.A(n_525),
.B(n_515),
.Y(n_533)
);

INVx3_ASAP7_75t_L g534 ( 
.A(n_525),
.Y(n_534)
);

XOR2x2_ASAP7_75t_L g535 ( 
.A(n_526),
.B(n_518),
.Y(n_535)
);

OAI22xp33_ASAP7_75t_SL g536 ( 
.A1(n_529),
.A2(n_511),
.B1(n_516),
.B2(n_522),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_527),
.B(n_498),
.Y(n_537)
);

OAI21xp5_ASAP7_75t_L g538 ( 
.A1(n_535),
.A2(n_524),
.B(n_523),
.Y(n_538)
);

NAND3xp33_ASAP7_75t_SL g539 ( 
.A(n_531),
.B(n_503),
.C(n_504),
.Y(n_539)
);

OAI21xp33_ASAP7_75t_SL g540 ( 
.A1(n_533),
.A2(n_530),
.B(n_501),
.Y(n_540)
);

OR2x2_ASAP7_75t_L g541 ( 
.A(n_537),
.B(n_503),
.Y(n_541)
);

AOI221xp5_ASAP7_75t_L g542 ( 
.A1(n_536),
.A2(n_519),
.B1(n_491),
.B2(n_499),
.C(n_488),
.Y(n_542)
);

AOI322xp5_ASAP7_75t_L g543 ( 
.A1(n_540),
.A2(n_534),
.A3(n_532),
.B1(n_515),
.B2(n_488),
.C1(n_491),
.C2(n_520),
.Y(n_543)
);

OAI221xp5_ASAP7_75t_SL g544 ( 
.A1(n_542),
.A2(n_538),
.B1(n_541),
.B2(n_534),
.C(n_539),
.Y(n_544)
);

AOI21xp5_ASAP7_75t_L g545 ( 
.A1(n_538),
.A2(n_487),
.B(n_500),
.Y(n_545)
);

AOI21xp33_ASAP7_75t_L g546 ( 
.A1(n_540),
.A2(n_492),
.B(n_493),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_542),
.B(n_521),
.Y(n_547)
);

NOR3x1_ASAP7_75t_L g548 ( 
.A(n_547),
.B(n_420),
.C(n_416),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_543),
.B(n_505),
.Y(n_549)
);

NAND5xp2_ASAP7_75t_L g550 ( 
.A(n_544),
.B(n_504),
.C(n_505),
.D(n_440),
.E(n_418),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_549),
.B(n_546),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_548),
.Y(n_552)
);

AOI21x1_ASAP7_75t_L g553 ( 
.A1(n_551),
.A2(n_545),
.B(n_550),
.Y(n_553)
);

NAND3xp33_ASAP7_75t_L g554 ( 
.A(n_553),
.B(n_552),
.C(n_477),
.Y(n_554)
);

OA22x2_ASAP7_75t_L g555 ( 
.A1(n_554),
.A2(n_513),
.B1(n_493),
.B2(n_492),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_555),
.Y(n_556)
);

XNOR2x1_ASAP7_75t_L g557 ( 
.A(n_556),
.B(n_480),
.Y(n_557)
);

AOI22xp33_ASAP7_75t_L g558 ( 
.A1(n_557),
.A2(n_477),
.B1(n_513),
.B2(n_504),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_558),
.B(n_483),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_559),
.Y(n_560)
);

XNOR2xp5_ASAP7_75t_L g561 ( 
.A(n_560),
.B(n_418),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_561),
.Y(n_562)
);

AOI22xp5_ASAP7_75t_L g563 ( 
.A1(n_562),
.A2(n_416),
.B1(n_474),
.B2(n_475),
.Y(n_563)
);


endmodule