module fake_jpeg_4335_n_334 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_334);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_334;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_11),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_SL g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx3_ASAP7_75t_SL g37 ( 
.A(n_23),
.Y(n_37)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_37),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_18),
.B(n_12),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_38),
.B(n_50),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_19),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_39),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_40),
.Y(n_83)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_41),
.B(n_48),
.Y(n_102)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_47),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_44),
.B(n_46),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_14),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_14),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_16),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_47),
.A2(n_34),
.B1(n_32),
.B2(n_30),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_52),
.A2(n_53),
.B1(n_54),
.B2(n_57),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_47),
.A2(n_32),
.B1(n_30),
.B2(n_18),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_48),
.A2(n_51),
.B1(n_50),
.B2(n_32),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_55),
.B(n_58),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_48),
.A2(n_30),
.B1(n_18),
.B2(n_24),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_42),
.A2(n_28),
.B1(n_16),
.B2(n_26),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_59),
.A2(n_79),
.B1(n_88),
.B2(n_93),
.Y(n_117)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_62),
.B(n_64),
.Y(n_128)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_65),
.B(n_73),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_51),
.Y(n_66)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_66),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_67),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_41),
.B(n_25),
.Y(n_68)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_68),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_41),
.A2(n_25),
.B1(n_24),
.B2(n_26),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_69),
.Y(n_105)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

CKINVDCx14_ASAP7_75t_R g133 ( 
.A(n_71),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_72),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_41),
.B(n_35),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_74),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_44),
.A2(n_31),
.B1(n_35),
.B2(n_29),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_75),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_44),
.B(n_29),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_77),
.B(n_81),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_39),
.B(n_28),
.C(n_21),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_78),
.B(n_8),
.C(n_1),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_L g79 ( 
.A1(n_49),
.A2(n_33),
.B1(n_20),
.B2(n_17),
.Y(n_79)
);

A2O1A1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_39),
.A2(n_19),
.B(n_23),
.C(n_21),
.Y(n_80)
);

O2A1O1Ixp33_ASAP7_75t_L g103 ( 
.A1(n_80),
.A2(n_15),
.B(n_11),
.C(n_10),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_46),
.B(n_31),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_46),
.A2(n_19),
.B1(n_23),
.B2(n_15),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_82),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_36),
.B(n_33),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_85),
.B(n_89),
.Y(n_129)
);

INVx2_ASAP7_75t_SL g87 ( 
.A(n_36),
.Y(n_87)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_87),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_40),
.A2(n_33),
.B1(n_20),
.B2(n_17),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_40),
.Y(n_89)
);

NOR2x1_ASAP7_75t_L g90 ( 
.A(n_40),
.B(n_23),
.Y(n_90)
);

NOR2x1_ASAP7_75t_L g120 ( 
.A(n_90),
.B(n_97),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_43),
.Y(n_91)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_91),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_L g93 ( 
.A1(n_43),
.A2(n_45),
.B1(n_33),
.B2(n_20),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_43),
.A2(n_23),
.B1(n_15),
.B2(n_17),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_94),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_45),
.B(n_20),
.Y(n_95)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_95),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_45),
.A2(n_15),
.B1(n_1),
.B2(n_2),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_96),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_106)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_37),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_37),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_98),
.B(n_100),
.Y(n_108)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_38),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_99),
.A2(n_15),
.B(n_9),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_38),
.B(n_12),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_38),
.B(n_11),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_101),
.B(n_8),
.Y(n_112)
);

NOR3xp33_ASAP7_75t_L g161 ( 
.A(n_103),
.B(n_4),
.C(n_5),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_106),
.A2(n_126),
.B1(n_132),
.B2(n_70),
.Y(n_147)
);

OAI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_110),
.A2(n_80),
.B1(n_58),
.B2(n_97),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_L g111 ( 
.A1(n_90),
.A2(n_79),
.B1(n_93),
.B2(n_88),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_111),
.A2(n_125),
.B1(n_56),
.B2(n_86),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_112),
.B(n_61),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_124),
.B(n_3),
.Y(n_148)
);

AO22x2_ASAP7_75t_L g125 ( 
.A1(n_92),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_55),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_99),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_128),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_134),
.B(n_136),
.Y(n_180)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_104),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_135),
.Y(n_177)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_113),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_129),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_137),
.B(n_146),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_138),
.A2(n_150),
.B1(n_161),
.B2(n_168),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_117),
.A2(n_131),
.B1(n_105),
.B2(n_111),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_139),
.A2(n_167),
.B1(n_127),
.B2(n_121),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_125),
.Y(n_140)
);

INVxp67_ASAP7_75t_SL g193 ( 
.A(n_140),
.Y(n_193)
);

O2A1O1Ixp33_ASAP7_75t_L g141 ( 
.A1(n_120),
.A2(n_96),
.B(n_63),
.C(n_92),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_141),
.A2(n_144),
.B(n_145),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_105),
.A2(n_64),
.B1(n_62),
.B2(n_71),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_142),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_120),
.B(n_59),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_143),
.B(n_149),
.C(n_158),
.Y(n_199)
);

O2A1O1Ixp33_ASAP7_75t_L g144 ( 
.A1(n_125),
.A2(n_70),
.B(n_102),
.C(n_98),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_116),
.A2(n_60),
.B(n_78),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_129),
.Y(n_146)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_147),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_148),
.B(n_152),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_110),
.B(n_89),
.C(n_76),
.Y(n_149)
);

OAI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_125),
.A2(n_84),
.B1(n_83),
.B2(n_61),
.Y(n_150)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_125),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_151),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_118),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_109),
.B(n_76),
.Y(n_153)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_153),
.Y(n_182)
);

BUFx24_ASAP7_75t_SL g154 ( 
.A(n_109),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_154),
.B(n_156),
.Y(n_206)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_104),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_155),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_123),
.Y(n_157)
);

INVx13_ASAP7_75t_L g192 ( 
.A(n_157),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_124),
.B(n_76),
.C(n_74),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_118),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_159),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_108),
.B(n_67),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_160),
.B(n_162),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_108),
.B(n_6),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_108),
.B(n_7),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_163),
.B(n_164),
.Y(n_181)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_103),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_106),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_165),
.B(n_166),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_119),
.B(n_87),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_117),
.A2(n_87),
.B1(n_83),
.B2(n_84),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_119),
.A2(n_56),
.B1(n_72),
.B2(n_91),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_169),
.A2(n_116),
.B1(n_127),
.B2(n_130),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_115),
.B(n_86),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_170),
.B(n_114),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_133),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_171),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_160),
.B(n_115),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_172),
.A2(n_187),
.B(n_178),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_173),
.A2(n_179),
.B1(n_184),
.B2(n_205),
.Y(n_236)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_166),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_183),
.B(n_186),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_139),
.A2(n_107),
.B1(n_121),
.B2(n_130),
.Y(n_184)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_144),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_143),
.B(n_107),
.Y(n_187)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_141),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_189),
.B(n_195),
.Y(n_239)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_167),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_151),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_197),
.B(n_198),
.Y(n_217)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_142),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_200),
.B(n_181),
.Y(n_234)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_162),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_201),
.B(n_202),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_137),
.B(n_112),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_146),
.B(n_112),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_204),
.B(n_208),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_165),
.A2(n_114),
.B1(n_56),
.B2(n_86),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_140),
.A2(n_122),
.B1(n_169),
.B2(n_164),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_207),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_163),
.B(n_122),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_149),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_209),
.B(n_187),
.Y(n_223)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_194),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_211),
.B(n_214),
.Y(n_257)
);

NAND2xp67_ASAP7_75t_SL g212 ( 
.A(n_193),
.B(n_170),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_212),
.A2(n_220),
.B(n_233),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_186),
.A2(n_145),
.B(n_157),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_213),
.A2(n_232),
.B(n_185),
.Y(n_248)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_194),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_177),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_215),
.Y(n_250)
);

AOI322xp5_ASAP7_75t_L g216 ( 
.A1(n_187),
.A2(n_155),
.A3(n_158),
.B1(n_196),
.B2(n_210),
.C1(n_172),
.C2(n_209),
.Y(n_216)
);

AOI221x1_ASAP7_75t_L g249 ( 
.A1(n_216),
.A2(n_202),
.B1(n_191),
.B2(n_192),
.C(n_195),
.Y(n_249)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_203),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_219),
.B(n_222),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_199),
.B(n_200),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_180),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_221),
.Y(n_242)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_208),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_223),
.B(n_230),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_175),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_224),
.B(n_229),
.Y(n_247)
);

AOI22x1_ASAP7_75t_L g226 ( 
.A1(n_188),
.A2(n_207),
.B1(n_197),
.B2(n_172),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_226),
.A2(n_188),
.B1(n_185),
.B2(n_189),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_174),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_184),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_176),
.B(n_182),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_231),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_199),
.B(n_178),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_234),
.B(n_237),
.C(n_238),
.Y(n_251)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_190),
.Y(n_235)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_235),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_183),
.B(n_196),
.C(n_210),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_179),
.B(n_201),
.C(n_198),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_232),
.B(n_181),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_240),
.B(n_245),
.C(n_254),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_234),
.B(n_204),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_243),
.B(n_225),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_244),
.A2(n_227),
.B1(n_230),
.B2(n_236),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_237),
.B(n_173),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_248),
.A2(n_252),
.B(n_261),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_249),
.B(n_244),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_226),
.A2(n_217),
.B(n_228),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_239),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_253),
.B(n_259),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_233),
.B(n_182),
.C(n_174),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_238),
.B(n_192),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_255),
.B(n_262),
.C(n_211),
.Y(n_281)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_218),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_226),
.A2(n_206),
.B(n_212),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_233),
.B(n_220),
.C(n_222),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_218),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_263),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_247),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_265),
.B(n_271),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_266),
.B(n_274),
.Y(n_296)
);

CKINVDCx14_ASAP7_75t_R g267 ( 
.A(n_257),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_267),
.B(n_277),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_270),
.B(n_272),
.Y(n_288)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_241),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_250),
.Y(n_272)
);

CKINVDCx14_ASAP7_75t_R g290 ( 
.A(n_273),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_245),
.B(n_220),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g276 ( 
.A(n_242),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_276),
.B(n_253),
.Y(n_295)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_241),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_258),
.B(n_213),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_278),
.B(n_280),
.C(n_281),
.Y(n_293)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_252),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_279),
.B(n_260),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_251),
.B(n_225),
.Y(n_280)
);

NAND3xp33_ASAP7_75t_L g282 ( 
.A(n_270),
.B(n_256),
.C(n_242),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_282),
.B(n_284),
.Y(n_299)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_283),
.Y(n_304)
);

NOR3xp33_ASAP7_75t_SL g284 ( 
.A(n_275),
.B(n_261),
.C(n_258),
.Y(n_284)
);

NOR3xp33_ASAP7_75t_SL g285 ( 
.A(n_275),
.B(n_248),
.C(n_240),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_285),
.B(n_289),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_264),
.A2(n_227),
.B1(n_236),
.B2(n_259),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_264),
.A2(n_217),
.B(n_260),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_291),
.B(n_289),
.Y(n_308)
);

XNOR2x1_ASAP7_75t_L g292 ( 
.A(n_278),
.B(n_255),
.Y(n_292)
);

MAJx2_ASAP7_75t_L g302 ( 
.A(n_292),
.B(n_294),
.C(n_280),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_SL g294 ( 
.A(n_274),
.B(n_251),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_295),
.B(n_214),
.Y(n_300)
);

BUFx2_ASAP7_75t_L g297 ( 
.A(n_295),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_297),
.B(n_306),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_293),
.B(n_269),
.C(n_281),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_298),
.B(n_301),
.Y(n_317)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_300),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_294),
.B(n_269),
.C(n_262),
.Y(n_301)
);

NAND3xp33_ASAP7_75t_L g318 ( 
.A(n_302),
.B(n_293),
.C(n_243),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_296),
.B(n_266),
.C(n_254),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_303),
.B(n_296),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_290),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_288),
.A2(n_285),
.B1(n_284),
.B2(n_263),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_307),
.Y(n_310)
);

AO21x1_ASAP7_75t_L g314 ( 
.A1(n_308),
.A2(n_268),
.B(n_292),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_309),
.B(n_301),
.C(n_303),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_297),
.B(n_219),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_311),
.A2(n_313),
.B(n_256),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_304),
.B(n_221),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_314),
.B(n_305),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_299),
.B(n_215),
.Y(n_316)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_316),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_SL g323 ( 
.A(n_318),
.B(n_302),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_319),
.B(n_324),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_320),
.A2(n_322),
.B(n_323),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_315),
.B(n_272),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_312),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_325),
.B(n_310),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_328),
.B(n_329),
.C(n_286),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_321),
.B(n_246),
.Y(n_329)
);

AOI21x1_ASAP7_75t_L g330 ( 
.A1(n_326),
.A2(n_314),
.B(n_318),
.Y(n_330)
);

OAI21xp33_ASAP7_75t_L g332 ( 
.A1(n_330),
.A2(n_331),
.B(n_327),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_317),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_287),
.Y(n_334)
);


endmodule