module fake_jpeg_2350_n_165 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_165);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_165;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_25),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_9),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_31),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_36),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_38),
.Y(n_49)
);

BUFx10_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_26),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_11),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_28),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_27),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_49),
.B(n_0),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_61),
.Y(n_66)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_59),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_39),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_57),
.A2(n_41),
.B1(n_43),
.B2(n_52),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_63),
.A2(n_73),
.B1(n_40),
.B2(n_46),
.Y(n_86)
);

HAxp5_ASAP7_75t_SL g65 ( 
.A(n_61),
.B(n_50),
.CON(n_65),
.SN(n_65)
);

OAI21xp33_ASAP7_75t_L g78 ( 
.A1(n_65),
.A2(n_50),
.B(n_55),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_62),
.B(n_41),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g79 ( 
.A(n_68),
.Y(n_79)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_72),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_60),
.A2(n_43),
.B1(n_52),
.B2(n_42),
.Y(n_73)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_71),
.Y(n_75)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

O2A1O1Ixp33_ASAP7_75t_L g76 ( 
.A1(n_65),
.A2(n_59),
.B(n_54),
.C(n_50),
.Y(n_76)
);

AOI21xp33_ASAP7_75t_L g95 ( 
.A1(n_76),
.A2(n_73),
.B(n_69),
.Y(n_95)
);

OAI32xp33_ASAP7_75t_L g77 ( 
.A1(n_66),
.A2(n_50),
.A3(n_54),
.B1(n_2),
.B2(n_3),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_78),
.Y(n_94)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_82),
.B(n_87),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_63),
.B(n_47),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_86),
.Y(n_98)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_67),
.A2(n_55),
.B(n_47),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_46),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_91),
.B(n_6),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_95),
.B(n_16),
.Y(n_108)
);

O2A1O1Ixp33_ASAP7_75t_SL g97 ( 
.A1(n_79),
.A2(n_64),
.B(n_40),
.C(n_51),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_97),
.A2(n_4),
.B(n_5),
.Y(n_111)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_99),
.Y(n_110)
);

A2O1A1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_76),
.A2(n_53),
.B(n_1),
.C(n_2),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_100),
.B(n_7),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_78),
.A2(n_42),
.B1(n_1),
.B2(n_3),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_102),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_120)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_103),
.Y(n_112)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_105),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_101),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_106),
.B(n_107),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_0),
.Y(n_107)
);

XNOR2x1_ASAP7_75t_L g126 ( 
.A(n_108),
.B(n_109),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_94),
.B(n_4),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g128 ( 
.A(n_111),
.B(n_121),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g114 ( 
.A(n_92),
.B(n_17),
.Y(n_114)
);

XNOR2x1_ASAP7_75t_L g138 ( 
.A(n_114),
.B(n_123),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_5),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_115),
.B(n_117),
.Y(n_136)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_90),
.Y(n_116)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_116),
.Y(n_133)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_104),
.Y(n_118)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_118),
.Y(n_134)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_90),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_119),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_120),
.A2(n_93),
.B1(n_97),
.B2(n_100),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_101),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_122),
.A2(n_8),
.B(n_12),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_94),
.B(n_96),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_124),
.A2(n_129),
.B1(n_131),
.B2(n_135),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_111),
.Y(n_125)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_125),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_123),
.B(n_95),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_127),
.B(n_20),
.C(n_21),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_113),
.A2(n_104),
.B1(n_10),
.B2(n_11),
.Y(n_129)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_130),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_108),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_109),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_112),
.A2(n_110),
.B1(n_118),
.B2(n_114),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_139),
.A2(n_22),
.B1(n_24),
.B2(n_30),
.Y(n_146)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_133),
.Y(n_142)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_142),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_127),
.A2(n_15),
.B(n_18),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_143),
.A2(n_128),
.B(n_137),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_144),
.B(n_148),
.C(n_143),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_146),
.B(n_147),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_132),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_132),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_149),
.A2(n_153),
.B(n_126),
.Y(n_156)
);

INVxp33_ASAP7_75t_L g154 ( 
.A(n_151),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_140),
.B(n_138),
.Y(n_153)
);

FAx1_ASAP7_75t_SL g155 ( 
.A(n_153),
.B(n_138),
.CI(n_126),
.CON(n_155),
.SN(n_155)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_155),
.B(n_144),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_156),
.A2(n_128),
.B1(n_141),
.B2(n_150),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_157),
.A2(n_158),
.B1(n_154),
.B2(n_145),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_136),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_160),
.A2(n_152),
.B(n_142),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_134),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_162),
.Y(n_163)
);

AO21x1_ASAP7_75t_L g164 ( 
.A1(n_163),
.A2(n_32),
.B(n_35),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_37),
.Y(n_165)
);


endmodule