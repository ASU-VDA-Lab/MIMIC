module fake_jpeg_26494_n_275 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_275);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_275;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_2),
.B(n_9),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_37),
.Y(n_41)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_20),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_16),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_31),
.A2(n_29),
.B1(n_24),
.B2(n_16),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_40),
.A2(n_24),
.B1(n_23),
.B2(n_27),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_37),
.A2(n_38),
.B1(n_20),
.B2(n_29),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_42),
.A2(n_15),
.B1(n_22),
.B2(n_18),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_43),
.B(n_46),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_32),
.B(n_16),
.Y(n_46)
);

A2O1A1Ixp33_ASAP7_75t_L g48 ( 
.A1(n_36),
.A2(n_14),
.B(n_26),
.C(n_27),
.Y(n_48)
);

A2O1A1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_48),
.A2(n_39),
.B(n_17),
.C(n_28),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_39),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_50),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_14),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_51),
.B(n_52),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_14),
.Y(n_52)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_57),
.B(n_59),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_35),
.B(n_26),
.Y(n_58)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_58),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_33),
.B(n_26),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_31),
.A2(n_29),
.B1(n_24),
.B2(n_27),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_60),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_63),
.A2(n_77),
.B1(n_18),
.B2(n_22),
.Y(n_85)
);

AO22x1_ASAP7_75t_SL g65 ( 
.A1(n_48),
.A2(n_60),
.B1(n_41),
.B2(n_59),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_65),
.A2(n_44),
.B1(n_19),
.B2(n_34),
.Y(n_100)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_66),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_50),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_67),
.B(n_71),
.Y(n_92)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_68),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_54),
.A2(n_15),
.B1(n_23),
.B2(n_17),
.Y(n_70)
);

CKINVDCx14_ASAP7_75t_R g101 ( 
.A(n_70),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_54),
.A2(n_23),
.B1(n_15),
.B2(n_49),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_72),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_75),
.B(n_80),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_54),
.A2(n_17),
.B1(n_21),
.B2(n_25),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_46),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_78),
.B(n_79),
.Y(n_102)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_83),
.A2(n_30),
.B(n_19),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_85),
.A2(n_104),
.B1(n_82),
.B2(n_66),
.Y(n_127)
);

OAI32xp33_ASAP7_75t_L g86 ( 
.A1(n_80),
.A2(n_41),
.A3(n_43),
.B1(n_52),
.B2(n_58),
.Y(n_86)
);

A2O1A1Ixp33_ASAP7_75t_L g112 ( 
.A1(n_86),
.A2(n_76),
.B(n_62),
.C(n_81),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_73),
.A2(n_22),
.B1(n_18),
.B2(n_49),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_87),
.A2(n_105),
.B1(n_75),
.B2(n_81),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_57),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_94),
.C(n_83),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_65),
.B(n_56),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_91),
.B(n_98),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_69),
.B(n_56),
.C(n_44),
.Y(n_94)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_61),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_96),
.B(n_99),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_65),
.B(n_44),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_64),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_100),
.B(n_45),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_65),
.B(n_47),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_103),
.B(n_47),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_73),
.A2(n_47),
.B1(n_34),
.B2(n_25),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_78),
.A2(n_25),
.B1(n_21),
.B2(n_17),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_61),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_106),
.B(n_79),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_107),
.A2(n_30),
.B(n_19),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_99),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_108),
.Y(n_137)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_102),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_109),
.B(n_119),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_110),
.A2(n_114),
.B1(n_124),
.B2(n_127),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_111),
.B(n_112),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_95),
.A2(n_64),
.B(n_67),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_115),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_95),
.A2(n_76),
.B(n_62),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_117),
.A2(n_101),
.B1(n_86),
.B2(n_85),
.Y(n_134)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_118),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_102),
.B(n_68),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_92),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_120),
.B(n_121),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_92),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_91),
.B(n_45),
.Y(n_122)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_122),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_94),
.B(n_74),
.Y(n_123)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_123),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_88),
.B(n_74),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_125),
.B(n_111),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_98),
.B(n_45),
.C(n_74),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_126),
.B(n_128),
.Y(n_152)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_103),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_129),
.B(n_131),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_107),
.A2(n_45),
.B(n_17),
.Y(n_130)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_130),
.Y(n_144)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_100),
.Y(n_131)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_108),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_132),
.B(n_138),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_134),
.A2(n_130),
.B(n_110),
.Y(n_173)
);

AOI22x1_ASAP7_75t_L g139 ( 
.A1(n_115),
.A2(n_101),
.B1(n_90),
.B2(n_104),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_139),
.A2(n_127),
.B1(n_109),
.B2(n_110),
.Y(n_170)
);

INVxp33_ASAP7_75t_L g140 ( 
.A(n_113),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_140),
.B(n_145),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_120),
.B(n_90),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_121),
.B(n_97),
.Y(n_147)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_147),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_125),
.B(n_106),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_150),
.B(n_130),
.Y(n_174)
);

INVx13_ASAP7_75t_L g151 ( 
.A(n_113),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_151),
.B(n_155),
.Y(n_177)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_118),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_153),
.B(n_154),
.Y(n_178)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_119),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_124),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_146),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_156),
.B(n_157),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_136),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_139),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_158),
.B(n_163),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_144),
.A2(n_129),
.B1(n_131),
.B2(n_148),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_159),
.A2(n_170),
.B1(n_142),
.B2(n_155),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_143),
.B(n_149),
.C(n_152),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_160),
.B(n_164),
.C(n_166),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_144),
.A2(n_122),
.B(n_116),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_161),
.A2(n_162),
.B(n_133),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_139),
.A2(n_116),
.B(n_122),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_135),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_143),
.B(n_123),
.C(n_126),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_135),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_165),
.B(n_167),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_152),
.B(n_112),
.C(n_117),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_132),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_150),
.B(n_112),
.C(n_128),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_168),
.B(n_174),
.C(n_175),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_173),
.A2(n_141),
.B(n_137),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_142),
.B(n_110),
.C(n_114),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_140),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_176),
.B(n_93),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_179),
.A2(n_187),
.B1(n_89),
.B2(n_66),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_162),
.A2(n_154),
.B(n_153),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g202 ( 
.A(n_180),
.Y(n_202)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_183),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_178),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_184),
.B(n_189),
.Y(n_200)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_167),
.Y(n_186)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_186),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_156),
.A2(n_157),
.B1(n_141),
.B2(n_172),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_158),
.A2(n_159),
.B1(n_163),
.B2(n_165),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_188),
.A2(n_191),
.B1(n_195),
.B2(n_21),
.Y(n_214)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_178),
.Y(n_189)
);

OA21x2_ASAP7_75t_SL g192 ( 
.A1(n_166),
.A2(n_151),
.B(n_133),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_192),
.B(n_198),
.Y(n_207)
);

AND2x4_ASAP7_75t_SL g193 ( 
.A(n_173),
.B(n_74),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_193),
.A2(n_199),
.B1(n_169),
.B2(n_171),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_161),
.A2(n_84),
.B(n_96),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_164),
.B(n_97),
.C(n_93),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_196),
.B(n_174),
.C(n_168),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_197),
.Y(n_206)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_177),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_175),
.A2(n_89),
.B1(n_84),
.B2(n_82),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_194),
.B(n_160),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_203),
.B(n_212),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_205),
.B(n_216),
.C(n_189),
.Y(n_224)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_182),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_208),
.B(n_211),
.Y(n_221)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_209),
.Y(n_217)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_210),
.Y(n_225)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_185),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_194),
.B(n_17),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_190),
.B(n_25),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_213),
.B(n_191),
.Y(n_222)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_214),
.Y(n_227)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_185),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_215),
.B(n_180),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_196),
.B(n_21),
.C(n_7),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_203),
.B(n_190),
.C(n_198),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_218),
.B(n_219),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_213),
.B(n_183),
.C(n_199),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_222),
.B(n_226),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_207),
.A2(n_179),
.B1(n_184),
.B2(n_181),
.Y(n_223)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_223),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_224),
.B(n_216),
.C(n_204),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_205),
.B(n_188),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_212),
.B(n_186),
.C(n_195),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_228),
.B(n_229),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_209),
.B(n_193),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_230),
.B(n_231),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_204),
.B(n_193),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_232),
.B(n_243),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_224),
.Y(n_234)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_234),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_226),
.B(n_206),
.C(n_208),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_236),
.B(n_239),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_225),
.A2(n_201),
.B1(n_214),
.B2(n_202),
.Y(n_237)
);

O2A1O1Ixp33_ASAP7_75t_SL g244 ( 
.A1(n_237),
.A2(n_217),
.B(n_227),
.C(n_230),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_220),
.B(n_200),
.C(n_7),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_221),
.A2(n_6),
.B(n_12),
.Y(n_242)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_242),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_220),
.B(n_6),
.C(n_12),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_244),
.A2(n_11),
.B(n_9),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_238),
.A2(n_240),
.B(n_241),
.Y(n_245)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_245),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_233),
.B(n_222),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_246),
.B(n_249),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_233),
.B(n_231),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_235),
.B(n_13),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_251),
.B(n_0),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_239),
.A2(n_11),
.B(n_10),
.Y(n_253)
);

AOI21xp33_ASAP7_75t_L g259 ( 
.A1(n_253),
.A2(n_0),
.B(n_1),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_248),
.B(n_243),
.C(n_237),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_254),
.B(n_249),
.C(n_246),
.Y(n_264)
);

AO21x1_ASAP7_75t_L g255 ( 
.A1(n_247),
.A2(n_244),
.B(n_252),
.Y(n_255)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_255),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_256),
.A2(n_259),
.B(n_0),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_250),
.A2(n_11),
.B1(n_9),
.B2(n_2),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_257),
.A2(n_260),
.B1(n_251),
.B2(n_1),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_263),
.B(n_265),
.Y(n_270)
);

MAJx2_ASAP7_75t_L g267 ( 
.A(n_264),
.B(n_266),
.C(n_258),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_261),
.B(n_1),
.C(n_2),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_267),
.A2(n_268),
.B(n_269),
.Y(n_271)
);

OAI21x1_ASAP7_75t_L g268 ( 
.A1(n_262),
.A2(n_255),
.B(n_258),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_262),
.A2(n_1),
.B(n_3),
.Y(n_269)
);

AOI321xp33_ASAP7_75t_L g272 ( 
.A1(n_270),
.A2(n_3),
.A3(n_4),
.B1(n_5),
.B2(n_261),
.C(n_262),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_272),
.B(n_4),
.Y(n_273)
);

BUFx24_ASAP7_75t_SL g274 ( 
.A(n_273),
.Y(n_274)
);

OR2x2_ASAP7_75t_L g275 ( 
.A(n_274),
.B(n_271),
.Y(n_275)
);


endmodule