module real_jpeg_30141_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_300;
wire n_215;
wire n_286;
wire n_288;
wire n_292;
wire n_194;
wire n_153;
wire n_104;
wire n_161;
wire n_207;
wire n_301;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_255;
wire n_243;
wire n_115;
wire n_299;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_164;
wire n_48;
wire n_184;
wire n_275;
wire n_293;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_290;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_302;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_298;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_134;
wire n_270;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_289;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_150;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_70;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_297;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_240;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_167;
wire n_128;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_295;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_283;
wire n_181;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_0),
.A2(n_32),
.B1(n_33),
.B2(n_147),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_0),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_0),
.A2(n_76),
.B1(n_77),
.B2(n_147),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_0),
.A2(n_29),
.B1(n_30),
.B2(n_147),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_0),
.A2(n_47),
.B1(n_50),
.B2(n_147),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_1),
.Y(n_90)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_1),
.Y(n_91)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_1),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_2),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_2),
.B(n_72),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_2),
.B(n_32),
.Y(n_193)
);

AOI21xp33_ASAP7_75t_L g197 ( 
.A1(n_2),
.A2(n_32),
.B(n_193),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_2),
.A2(n_29),
.B1(n_30),
.B2(n_151),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_2),
.A2(n_47),
.B(n_51),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_2),
.B(n_119),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_2),
.A2(n_88),
.B1(n_170),
.B2(n_241),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_3),
.A2(n_76),
.B1(n_77),
.B2(n_153),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_3),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_3),
.A2(n_32),
.B1(n_33),
.B2(n_153),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_3),
.A2(n_29),
.B1(n_30),
.B2(n_153),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_3),
.A2(n_47),
.B1(n_50),
.B2(n_153),
.Y(n_241)
);

BUFx12_ASAP7_75t_L g74 ( 
.A(n_4),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_5),
.A2(n_29),
.B1(n_30),
.B2(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_5),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_5),
.A2(n_32),
.B1(n_33),
.B2(n_57),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_5),
.A2(n_57),
.B1(n_76),
.B2(n_77),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_5),
.A2(n_47),
.B1(n_50),
.B2(n_57),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx13_ASAP7_75t_L g76 ( 
.A(n_7),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_8),
.A2(n_32),
.B1(n_33),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_8),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_8),
.A2(n_38),
.B1(n_76),
.B2(n_77),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_8),
.A2(n_29),
.B1(n_30),
.B2(n_38),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_8),
.A2(n_38),
.B1(n_47),
.B2(n_50),
.Y(n_169)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_10),
.A2(n_76),
.B1(n_77),
.B2(n_125),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_10),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_10),
.A2(n_32),
.B1(n_33),
.B2(n_125),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_10),
.A2(n_29),
.B1(n_30),
.B2(n_125),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_10),
.A2(n_47),
.B1(n_50),
.B2(n_125),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_11),
.A2(n_32),
.B1(n_33),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_11),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_11),
.A2(n_29),
.B1(n_30),
.B2(n_40),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_11),
.A2(n_40),
.B1(n_47),
.B2(n_50),
.Y(n_138)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_13),
.A2(n_32),
.B1(n_33),
.B2(n_35),
.Y(n_31)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_14),
.A2(n_29),
.B1(n_30),
.B2(n_44),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_14),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_14),
.A2(n_44),
.B1(n_47),
.B2(n_50),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_14),
.A2(n_44),
.B1(n_76),
.B2(n_77),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_14),
.A2(n_32),
.B1(n_33),
.B2(n_44),
.Y(n_164)
);

INVx11_ASAP7_75t_SL g48 ( 
.A(n_15),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_129),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_127),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_101),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_19),
.B(n_101),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_85),
.B2(n_86),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_58),
.B2(n_59),
.Y(n_21)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_23),
.A2(n_24),
.B(n_41),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_41),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_36),
.B2(n_39),
.Y(n_24)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_25),
.B(n_69),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_25),
.A2(n_26),
.B1(n_146),
.B2(n_148),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_25),
.A2(n_26),
.B1(n_146),
.B2(n_179),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_25),
.A2(n_26),
.B1(n_179),
.B2(n_197),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_31),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_26),
.B(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_26),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_26),
.B(n_164),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_26)
);

INVx6_ASAP7_75t_L g192 ( 
.A(n_27),
.Y(n_192)
);

NAND2xp33_ASAP7_75t_SL g194 ( 
.A(n_27),
.B(n_30),
.Y(n_194)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp33_ASAP7_75t_L g55 ( 
.A1(n_29),
.A2(n_30),
.B1(n_49),
.B2(n_51),
.Y(n_55)
);

AOI32xp33_ASAP7_75t_L g191 ( 
.A1(n_29),
.A2(n_33),
.A3(n_192),
.B1(n_193),
.B2(n_194),
.Y(n_191)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

A2O1A1Ixp33_ASAP7_75t_L g219 ( 
.A1(n_30),
.A2(n_49),
.B(n_151),
.C(n_220),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_32),
.A2(n_33),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_32),
.B(n_73),
.Y(n_167)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_33),
.A2(n_80),
.B1(n_150),
.B2(n_167),
.Y(n_166)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_37),
.A2(n_119),
.B(n_120),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_39),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_52),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_42),
.A2(n_54),
.B(n_201),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_43),
.B(n_45),
.Y(n_42)
);

CKINVDCx14_ASAP7_75t_R g63 ( 
.A(n_43),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_45),
.B(n_56),
.Y(n_97)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_55),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_46),
.A2(n_54),
.B(n_63),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_46),
.A2(n_54),
.B1(n_96),
.B2(n_117),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_46),
.A2(n_52),
.B(n_117),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_46),
.A2(n_54),
.B1(n_200),
.B2(n_201),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_46),
.A2(n_54),
.B1(n_217),
.B2(n_218),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_46),
.A2(n_54),
.B1(n_200),
.B2(n_218),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_46),
.B(n_151),
.Y(n_239)
);

OA22x2_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_49),
.B1(n_50),
.B2(n_51),
.Y(n_46)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_47),
.Y(n_50)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_49),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_50),
.B(n_90),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_50),
.B(n_246),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_56),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_54),
.A2(n_96),
.B(n_97),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_54),
.A2(n_63),
.B(n_97),
.Y(n_143)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_60),
.A2(n_70),
.B1(n_83),
.B2(n_84),
.Y(n_59)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_62),
.B1(n_64),
.B2(n_65),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_67),
.B(n_68),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_66),
.A2(n_162),
.B(n_163),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_66),
.A2(n_68),
.B(n_280),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_70),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_75),
.B(n_78),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_71),
.B(n_82),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_71),
.A2(n_123),
.B1(n_158),
.B2(n_159),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_71),
.A2(n_123),
.B1(n_124),
.B2(n_159),
.Y(n_277)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

O2A1O1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_72),
.A2(n_73),
.B(n_77),
.C(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_72),
.B(n_99),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_72),
.A2(n_79),
.B1(n_150),
.B2(n_152),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_73),
.B(n_77),
.Y(n_80)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_76),
.Y(n_77)
);

HAxp5_ASAP7_75t_SL g150 ( 
.A(n_77),
.B(n_151),
.CON(n_150),
.SN(n_150)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_79),
.B(n_81),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_79),
.A2(n_99),
.B(n_100),
.Y(n_98)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_79),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

AOI21xp33_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_94),
.B(n_98),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_87),
.B(n_95),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_87),
.A2(n_98),
.B1(n_104),
.B2(n_105),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_87),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_87),
.A2(n_95),
.B1(n_105),
.B2(n_294),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_91),
.B(n_92),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_88),
.A2(n_138),
.B(n_139),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_88),
.A2(n_138),
.B1(n_169),
.B2(n_170),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_88),
.A2(n_114),
.B(n_228),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_88),
.A2(n_233),
.B1(n_241),
.B2(n_242),
.Y(n_240)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_112),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_89),
.A2(n_93),
.B(n_140),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_89),
.A2(n_115),
.B1(n_232),
.B2(n_234),
.Y(n_231)
);

INVx11_ASAP7_75t_L g115 ( 
.A(n_91),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_91),
.B(n_113),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_91),
.B(n_151),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_115),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_94),
.B(n_103),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_95),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_98),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_106),
.C(n_107),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_102),
.B(n_106),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_SL g299 ( 
.A1(n_107),
.A2(n_108),
.B1(n_300),
.B2(n_301),
.Y(n_299)
);

CKINVDCx14_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_118),
.C(n_121),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_109),
.B(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_116),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_110),
.B(n_116),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_114),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_111),
.A2(n_169),
.B(n_170),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx11_ASAP7_75t_L g242 ( 
.A(n_115),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_118),
.A2(n_121),
.B1(n_122),
.B2(n_291),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_118),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_123),
.A2(n_124),
.B(n_126),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_297),
.B(n_302),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_284),
.B(n_296),
.Y(n_130)
);

O2A1O1Ixp33_ASAP7_75t_SL g131 ( 
.A1(n_132),
.A2(n_183),
.B(n_265),
.C(n_283),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_171),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_133),
.B(n_171),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_154),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_141),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_135),
.B(n_141),
.C(n_154),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_137),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_136),
.B(n_137),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_144),
.C(n_149),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_142),
.A2(n_143),
.B1(n_144),
.B2(n_145),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_148),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_149),
.B(n_174),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_152),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_155),
.B(n_165),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_156),
.A2(n_157),
.B1(n_160),
.B2(n_161),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_156),
.B(n_161),
.C(n_165),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_164),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_168),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_166),
.B(n_168),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_175),
.C(n_177),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_172),
.A2(n_173),
.B1(n_260),
.B2(n_262),
.Y(n_259)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_175),
.A2(n_176),
.B1(n_177),
.B2(n_261),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_177),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_180),
.C(n_182),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_178),
.B(n_205),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_180),
.A2(n_181),
.B1(n_182),
.B2(n_206),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_182),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_184),
.B(n_264),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_257),
.B(n_263),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_211),
.B(n_256),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_202),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_187),
.B(n_202),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_195),
.C(n_198),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_188),
.A2(n_189),
.B1(n_253),
.B2(n_254),
.Y(n_252)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_191),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_190),
.B(n_191),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_195),
.A2(n_196),
.B1(n_198),
.B2(n_199),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_196),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_199),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_203),
.A2(n_204),
.B1(n_207),
.B2(n_208),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_203),
.B(n_209),
.C(n_210),
.Y(n_258)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_250),
.B(n_255),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_229),
.B(n_249),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_221),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_214),
.B(n_221),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_215),
.B(n_219),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_215),
.A2(n_216),
.B1(n_219),
.B2(n_236),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_219),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_227),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_224),
.B1(n_225),
.B2(n_226),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_223),
.B(n_226),
.C(n_227),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_224),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_226),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_228),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_237),
.B(n_248),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_235),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_231),
.B(n_235),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_238),
.A2(n_243),
.B(n_247),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_239),
.B(n_240),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_251),
.B(n_252),
.Y(n_255)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_258),
.B(n_259),
.Y(n_263)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_260),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_266),
.B(n_267),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_268),
.A2(n_269),
.B1(n_281),
.B2(n_282),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_271),
.B1(n_272),
.B2(n_273),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_270),
.B(n_273),
.C(n_282),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_274),
.B(n_276),
.C(n_279),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_276),
.A2(n_277),
.B1(n_278),
.B2(n_279),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_277),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_281),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_285),
.B(n_286),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_295),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_288),
.A2(n_289),
.B1(n_292),
.B2(n_293),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_288),
.B(n_293),
.C(n_295),
.Y(n_298)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_298),
.B(n_299),
.Y(n_302)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);


endmodule