module real_aes_7744_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_555;
wire n_364;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_545;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_537;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_453;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_288;
wire n_147;
wire n_150;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g241 ( .A1(n_0), .A2(n_242), .B(n_243), .C(n_247), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_1), .B(n_183), .Y(n_248) );
NAND3xp33_ASAP7_75t_SL g109 ( .A(n_2), .B(n_110), .C(n_111), .Y(n_109) );
INVx1_ASAP7_75t_L g465 ( .A(n_2), .Y(n_465) );
AOI22xp5_ASAP7_75t_L g104 ( .A1(n_3), .A2(n_105), .B1(n_114), .B2(n_757), .Y(n_104) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_4), .B(n_155), .Y(n_231) );
A2O1A1Ixp33_ASAP7_75t_L g512 ( .A1(n_5), .A2(n_141), .B(n_146), .C(n_513), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g550 ( .A1(n_6), .A2(n_136), .B(n_551), .Y(n_550) );
AOI21xp5_ASAP7_75t_L g173 ( .A1(n_7), .A2(n_136), .B(n_174), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_8), .B(n_183), .Y(n_557) );
AO21x2_ASAP7_75t_L g186 ( .A1(n_9), .A2(n_171), .B(n_187), .Y(n_186) );
AND2x6_ASAP7_75t_L g141 ( .A(n_10), .B(n_142), .Y(n_141) );
A2O1A1Ixp33_ASAP7_75t_L g256 ( .A1(n_11), .A2(n_141), .B(n_146), .C(n_257), .Y(n_256) );
INVx1_ASAP7_75t_L g495 ( .A(n_12), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_13), .B(n_108), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g466 ( .A(n_13), .B(n_42), .Y(n_466) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_14), .B(n_246), .Y(n_515) );
INVx1_ASAP7_75t_L g165 ( .A(n_15), .Y(n_165) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_16), .B(n_155), .Y(n_193) );
A2O1A1Ixp33_ASAP7_75t_L g502 ( .A1(n_17), .A2(n_156), .B(n_503), .C(n_505), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_18), .B(n_183), .Y(n_506) );
AOI22xp5_ASAP7_75t_SL g470 ( .A1(n_19), .A2(n_463), .B1(n_471), .B2(n_752), .Y(n_470) );
AOI22xp5_ASAP7_75t_L g122 ( .A1(n_20), .A2(n_48), .B1(n_123), .B2(n_124), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_20), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_20), .B(n_220), .Y(n_594) );
A2O1A1Ixp33_ASAP7_75t_L g215 ( .A1(n_21), .A2(n_146), .B(n_197), .C(n_216), .Y(n_215) );
A2O1A1Ixp33_ASAP7_75t_L g524 ( .A1(n_22), .A2(n_195), .B(n_245), .C(n_525), .Y(n_524) );
NAND2xp5_ASAP7_75t_SL g546 ( .A(n_23), .B(n_246), .Y(n_546) );
NAND2xp5_ASAP7_75t_SL g535 ( .A(n_24), .B(n_246), .Y(n_535) );
CKINVDCx16_ASAP7_75t_R g542 ( .A(n_25), .Y(n_542) );
INVx1_ASAP7_75t_L g534 ( .A(n_26), .Y(n_534) );
A2O1A1Ixp33_ASAP7_75t_L g189 ( .A1(n_27), .A2(n_146), .B(n_190), .C(n_197), .Y(n_189) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_28), .Y(n_140) );
CKINVDCx20_ASAP7_75t_R g511 ( .A(n_29), .Y(n_511) );
INVx1_ASAP7_75t_L g591 ( .A(n_30), .Y(n_591) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_31), .A2(n_136), .B(n_239), .Y(n_238) );
INVx2_ASAP7_75t_L g139 ( .A(n_32), .Y(n_139) );
A2O1A1Ixp33_ASAP7_75t_L g204 ( .A1(n_33), .A2(n_144), .B(n_159), .C(n_205), .Y(n_204) );
CKINVDCx20_ASAP7_75t_R g518 ( .A(n_34), .Y(n_518) );
A2O1A1Ixp33_ASAP7_75t_L g553 ( .A1(n_35), .A2(n_245), .B(n_554), .C(n_556), .Y(n_553) );
INVxp67_ASAP7_75t_L g592 ( .A(n_36), .Y(n_592) );
OAI22xp5_ASAP7_75t_SL g126 ( .A1(n_37), .A2(n_47), .B1(n_127), .B2(n_128), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_37), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_38), .B(n_192), .Y(n_191) );
A2O1A1Ixp33_ASAP7_75t_L g532 ( .A1(n_39), .A2(n_146), .B(n_197), .C(n_533), .Y(n_532) );
CKINVDCx14_ASAP7_75t_R g552 ( .A(n_40), .Y(n_552) );
OAI22xp5_ASAP7_75t_L g477 ( .A1(n_41), .A2(n_46), .B1(n_478), .B2(n_479), .Y(n_477) );
INVx1_ASAP7_75t_L g479 ( .A(n_41), .Y(n_479) );
INVx1_ASAP7_75t_L g108 ( .A(n_42), .Y(n_108) );
A2O1A1Ixp33_ASAP7_75t_L g492 ( .A1(n_43), .A2(n_247), .B(n_493), .C(n_494), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_44), .B(n_214), .Y(n_213) );
CKINVDCx20_ASAP7_75t_R g261 ( .A(n_45), .Y(n_261) );
CKINVDCx20_ASAP7_75t_R g478 ( .A(n_46), .Y(n_478) );
INVx1_ASAP7_75t_L g128 ( .A(n_47), .Y(n_128) );
INVx1_ASAP7_75t_L g124 ( .A(n_48), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_49), .B(n_155), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_50), .B(n_136), .Y(n_188) );
CKINVDCx20_ASAP7_75t_R g537 ( .A(n_51), .Y(n_537) );
CKINVDCx20_ASAP7_75t_R g588 ( .A(n_52), .Y(n_588) );
A2O1A1Ixp33_ASAP7_75t_L g143 ( .A1(n_53), .A2(n_144), .B(n_149), .C(n_159), .Y(n_143) );
INVx1_ASAP7_75t_L g244 ( .A(n_54), .Y(n_244) );
INVx1_ASAP7_75t_L g150 ( .A(n_55), .Y(n_150) );
INVx1_ASAP7_75t_L g523 ( .A(n_56), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_57), .B(n_136), .Y(n_135) );
CKINVDCx20_ASAP7_75t_R g223 ( .A(n_58), .Y(n_223) );
CKINVDCx14_ASAP7_75t_R g491 ( .A(n_59), .Y(n_491) );
INVx1_ASAP7_75t_L g142 ( .A(n_60), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_61), .B(n_136), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_62), .B(n_183), .Y(n_182) );
A2O1A1Ixp33_ASAP7_75t_L g176 ( .A1(n_63), .A2(n_177), .B(n_179), .C(n_181), .Y(n_176) );
INVx1_ASAP7_75t_L g164 ( .A(n_64), .Y(n_164) );
INVx1_ASAP7_75t_SL g555 ( .A(n_65), .Y(n_555) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_66), .Y(n_119) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_67), .B(n_155), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_68), .B(n_183), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_69), .B(n_156), .Y(n_258) );
INVx1_ASAP7_75t_L g545 ( .A(n_70), .Y(n_545) );
CKINVDCx16_ASAP7_75t_R g240 ( .A(n_71), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_72), .B(n_152), .Y(n_217) );
A2O1A1Ixp33_ASAP7_75t_L g228 ( .A1(n_73), .A2(n_146), .B(n_159), .C(n_229), .Y(n_228) );
CKINVDCx16_ASAP7_75t_R g175 ( .A(n_74), .Y(n_175) );
INVx1_ASAP7_75t_L g113 ( .A(n_75), .Y(n_113) );
AOI21xp5_ASAP7_75t_L g489 ( .A1(n_76), .A2(n_136), .B(n_490), .Y(n_489) );
CKINVDCx20_ASAP7_75t_R g548 ( .A(n_77), .Y(n_548) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_78), .A2(n_136), .B(n_500), .Y(n_499) );
OAI22xp5_ASAP7_75t_SL g472 ( .A1(n_79), .A2(n_473), .B1(n_474), .B2(n_480), .Y(n_472) );
CKINVDCx20_ASAP7_75t_R g480 ( .A(n_79), .Y(n_480) );
AOI21xp5_ASAP7_75t_L g586 ( .A1(n_80), .A2(n_214), .B(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g501 ( .A(n_81), .Y(n_501) );
CKINVDCx16_ASAP7_75t_R g531 ( .A(n_82), .Y(n_531) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_83), .B(n_151), .Y(n_218) );
AOI22xp5_ASAP7_75t_L g474 ( .A1(n_84), .A2(n_475), .B1(n_476), .B2(n_477), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_84), .Y(n_475) );
CKINVDCx20_ASAP7_75t_R g209 ( .A(n_85), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_86), .A2(n_136), .B(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g504 ( .A(n_87), .Y(n_504) );
INVx2_ASAP7_75t_L g162 ( .A(n_88), .Y(n_162) );
INVx1_ASAP7_75t_L g514 ( .A(n_89), .Y(n_514) );
CKINVDCx20_ASAP7_75t_R g236 ( .A(n_90), .Y(n_236) );
NAND2xp5_ASAP7_75t_SL g259 ( .A(n_91), .B(n_246), .Y(n_259) );
INVx2_ASAP7_75t_L g110 ( .A(n_92), .Y(n_110) );
OR2x2_ASAP7_75t_L g462 ( .A(n_92), .B(n_463), .Y(n_462) );
A2O1A1Ixp33_ASAP7_75t_L g543 ( .A1(n_93), .A2(n_146), .B(n_159), .C(n_544), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_94), .B(n_136), .Y(n_203) );
NAND2xp5_ASAP7_75t_SL g467 ( .A(n_95), .B(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g206 ( .A(n_96), .Y(n_206) );
INVxp67_ASAP7_75t_L g180 ( .A(n_97), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_98), .B(n_171), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_99), .B(n_113), .Y(n_112) );
INVx1_ASAP7_75t_L g230 ( .A(n_100), .Y(n_230) );
INVx1_ASAP7_75t_L g254 ( .A(n_101), .Y(n_254) );
INVx2_ASAP7_75t_L g526 ( .A(n_102), .Y(n_526) );
AND2x2_ASAP7_75t_L g166 ( .A(n_103), .B(n_161), .Y(n_166) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_SL g758 ( .A(n_106), .Y(n_758) );
OR2x2_ASAP7_75t_L g106 ( .A(n_107), .B(n_109), .Y(n_106) );
INVx2_ASAP7_75t_L g482 ( .A(n_110), .Y(n_482) );
INVx1_ASAP7_75t_L g751 ( .A(n_110), .Y(n_751) );
NOR2x2_ASAP7_75t_L g754 ( .A(n_110), .B(n_463), .Y(n_754) );
INVx1_ASAP7_75t_SL g111 ( .A(n_112), .Y(n_111) );
OA21x2_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_120), .B(n_469), .Y(n_114) );
INVx1_ASAP7_75t_SL g115 ( .A(n_116), .Y(n_115) );
INVx1_ASAP7_75t_SL g116 ( .A(n_117), .Y(n_116) );
BUFx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx2_ASAP7_75t_SL g756 ( .A(n_118), .Y(n_756) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
OAI21xp5_ASAP7_75t_SL g120 ( .A1(n_121), .A2(n_459), .B(n_467), .Y(n_120) );
XNOR2xp5_ASAP7_75t_L g121 ( .A(n_122), .B(n_125), .Y(n_121) );
XOR2xp5_ASAP7_75t_L g125 ( .A(n_126), .B(n_129), .Y(n_125) );
AOI22xp5_ASAP7_75t_L g481 ( .A1(n_129), .A2(n_482), .B1(n_483), .B2(n_750), .Y(n_481) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
OR5x1_ASAP7_75t_L g130 ( .A(n_131), .B(n_332), .C(n_410), .D(n_434), .E(n_451), .Y(n_130) );
OAI211xp5_ASAP7_75t_SL g131 ( .A1(n_132), .A2(n_198), .B(n_249), .C(n_309), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_133), .B(n_167), .Y(n_132) );
AND2x2_ASAP7_75t_L g263 ( .A(n_133), .B(n_169), .Y(n_263) );
INVx5_ASAP7_75t_SL g291 ( .A(n_133), .Y(n_291) );
AND2x2_ASAP7_75t_L g327 ( .A(n_133), .B(n_312), .Y(n_327) );
OR2x2_ASAP7_75t_L g366 ( .A(n_133), .B(n_168), .Y(n_366) );
OR2x2_ASAP7_75t_L g397 ( .A(n_133), .B(n_288), .Y(n_397) );
NOR2xp33_ASAP7_75t_L g433 ( .A(n_133), .B(n_301), .Y(n_433) );
AND2x2_ASAP7_75t_L g445 ( .A(n_133), .B(n_288), .Y(n_445) );
OR2x6_ASAP7_75t_L g133 ( .A(n_134), .B(n_166), .Y(n_133) );
AOI21xp5_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_143), .B(n_161), .Y(n_134) );
BUFx2_ASAP7_75t_L g214 ( .A(n_136), .Y(n_214) );
AND2x4_ASAP7_75t_L g136 ( .A(n_137), .B(n_141), .Y(n_136) );
NAND2x1p5_ASAP7_75t_L g255 ( .A(n_137), .B(n_141), .Y(n_255) );
AND2x2_ASAP7_75t_L g137 ( .A(n_138), .B(n_140), .Y(n_137) );
INVx1_ASAP7_75t_L g181 ( .A(n_138), .Y(n_181) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx2_ASAP7_75t_L g147 ( .A(n_139), .Y(n_147) );
INVx1_ASAP7_75t_L g196 ( .A(n_139), .Y(n_196) );
INVx1_ASAP7_75t_L g148 ( .A(n_140), .Y(n_148) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_140), .Y(n_153) );
INVx3_ASAP7_75t_L g156 ( .A(n_140), .Y(n_156) );
INVx1_ASAP7_75t_L g192 ( .A(n_140), .Y(n_192) );
BUFx6f_ASAP7_75t_L g246 ( .A(n_140), .Y(n_246) );
INVx4_ASAP7_75t_SL g160 ( .A(n_141), .Y(n_160) );
BUFx3_ASAP7_75t_L g197 ( .A(n_141), .Y(n_197) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
O2A1O1Ixp33_ASAP7_75t_L g174 ( .A1(n_145), .A2(n_160), .B(n_175), .C(n_176), .Y(n_174) );
O2A1O1Ixp33_ASAP7_75t_SL g239 ( .A1(n_145), .A2(n_160), .B(n_240), .C(n_241), .Y(n_239) );
O2A1O1Ixp33_ASAP7_75t_SL g490 ( .A1(n_145), .A2(n_160), .B(n_491), .C(n_492), .Y(n_490) );
O2A1O1Ixp33_ASAP7_75t_SL g500 ( .A1(n_145), .A2(n_160), .B(n_501), .C(n_502), .Y(n_500) );
O2A1O1Ixp33_ASAP7_75t_SL g522 ( .A1(n_145), .A2(n_160), .B(n_523), .C(n_524), .Y(n_522) );
O2A1O1Ixp33_ASAP7_75t_L g551 ( .A1(n_145), .A2(n_160), .B(n_552), .C(n_553), .Y(n_551) );
O2A1O1Ixp33_ASAP7_75t_SL g587 ( .A1(n_145), .A2(n_160), .B(n_588), .C(n_589), .Y(n_587) );
INVx5_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
AND2x6_ASAP7_75t_L g146 ( .A(n_147), .B(n_148), .Y(n_146) );
BUFx3_ASAP7_75t_L g158 ( .A(n_147), .Y(n_158) );
BUFx6f_ASAP7_75t_L g233 ( .A(n_147), .Y(n_233) );
O2A1O1Ixp33_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_151), .B(n_154), .C(n_157), .Y(n_149) );
O2A1O1Ixp33_ASAP7_75t_L g205 ( .A1(n_151), .A2(n_157), .B(n_206), .C(n_207), .Y(n_205) );
O2A1O1Ixp5_ASAP7_75t_L g513 ( .A1(n_151), .A2(n_514), .B(n_515), .C(n_516), .Y(n_513) );
O2A1O1Ixp33_ASAP7_75t_L g544 ( .A1(n_151), .A2(n_516), .B(n_545), .C(n_546), .Y(n_544) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx4_ASAP7_75t_L g178 ( .A(n_153), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g179 ( .A(n_155), .B(n_180), .Y(n_179) );
INVx2_ASAP7_75t_L g242 ( .A(n_155), .Y(n_242) );
O2A1O1Ixp33_ASAP7_75t_L g533 ( .A1(n_155), .A2(n_219), .B(n_534), .C(n_535), .Y(n_533) );
OAI22xp33_ASAP7_75t_L g590 ( .A1(n_155), .A2(n_178), .B1(n_591), .B2(n_592), .Y(n_590) );
INVx5_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_156), .B(n_495), .Y(n_494) );
HB1xp67_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx2_ASAP7_75t_L g247 ( .A(n_158), .Y(n_247) );
INVx1_ASAP7_75t_L g505 ( .A(n_158), .Y(n_505) );
INVx1_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
AOI21xp5_ASAP7_75t_L g202 ( .A1(n_161), .A2(n_203), .B(n_204), .Y(n_202) );
INVx2_ASAP7_75t_L g221 ( .A(n_161), .Y(n_221) );
INVx1_ASAP7_75t_L g224 ( .A(n_161), .Y(n_224) );
OA21x2_ASAP7_75t_L g488 ( .A1(n_161), .A2(n_489), .B(n_496), .Y(n_488) );
O2A1O1Ixp33_ASAP7_75t_L g530 ( .A1(n_161), .A2(n_255), .B(n_531), .C(n_532), .Y(n_530) );
AND2x2_ASAP7_75t_SL g161 ( .A(n_162), .B(n_163), .Y(n_161) );
AND2x2_ASAP7_75t_L g172 ( .A(n_162), .B(n_163), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_164), .B(n_165), .Y(n_163) );
AND2x2_ASAP7_75t_L g444 ( .A(n_167), .B(n_445), .Y(n_444) );
INVx1_ASAP7_75t_SL g167 ( .A(n_168), .Y(n_167) );
OR2x2_ASAP7_75t_L g307 ( .A(n_168), .B(n_308), .Y(n_307) );
OR2x2_ASAP7_75t_L g168 ( .A(n_169), .B(n_185), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_169), .B(n_288), .Y(n_287) );
HB1xp67_ASAP7_75t_L g300 ( .A(n_169), .Y(n_300) );
INVx3_ASAP7_75t_L g315 ( .A(n_169), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_169), .B(n_185), .Y(n_339) );
OR2x2_ASAP7_75t_L g348 ( .A(n_169), .B(n_291), .Y(n_348) );
AND2x2_ASAP7_75t_L g352 ( .A(n_169), .B(n_312), .Y(n_352) );
AND2x2_ASAP7_75t_L g358 ( .A(n_169), .B(n_359), .Y(n_358) );
INVxp67_ASAP7_75t_L g395 ( .A(n_169), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_169), .B(n_252), .Y(n_409) );
OA21x2_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_173), .B(n_182), .Y(n_169) );
OA21x2_ASAP7_75t_L g498 ( .A1(n_170), .A2(n_499), .B(n_506), .Y(n_498) );
OA21x2_ASAP7_75t_L g520 ( .A1(n_170), .A2(n_521), .B(n_527), .Y(n_520) );
OA21x2_ASAP7_75t_L g549 ( .A1(n_170), .A2(n_550), .B(n_557), .Y(n_549) );
HB1xp67_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx4_ASAP7_75t_L g184 ( .A(n_171), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g187 ( .A1(n_171), .A2(n_188), .B(n_189), .Y(n_187) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx1_ASAP7_75t_L g262 ( .A(n_172), .Y(n_262) );
O2A1O1Ixp33_ASAP7_75t_L g229 ( .A1(n_177), .A2(n_230), .B(n_231), .C(n_232), .Y(n_229) );
INVx1_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g503 ( .A(n_178), .B(n_504), .Y(n_503) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_178), .B(n_526), .Y(n_525) );
INVx2_ASAP7_75t_L g219 ( .A(n_181), .Y(n_219) );
NAND2xp5_ASAP7_75t_SL g589 ( .A(n_181), .B(n_590), .Y(n_589) );
OA21x2_ASAP7_75t_L g237 ( .A1(n_183), .A2(n_238), .B(n_248), .Y(n_237) );
INVx3_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
NOR2xp33_ASAP7_75t_L g208 ( .A(n_184), .B(n_209), .Y(n_208) );
AO21x2_ASAP7_75t_L g226 ( .A1(n_184), .A2(n_227), .B(n_235), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_184), .B(n_236), .Y(n_235) );
AO21x2_ASAP7_75t_L g252 ( .A1(n_184), .A2(n_253), .B(n_260), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g517 ( .A(n_184), .B(n_518), .Y(n_517) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_184), .B(n_537), .Y(n_536) );
AO21x2_ASAP7_75t_L g540 ( .A1(n_184), .A2(n_541), .B(n_547), .Y(n_540) );
OR2x2_ASAP7_75t_L g301 ( .A(n_185), .B(n_252), .Y(n_301) );
AND2x2_ASAP7_75t_L g312 ( .A(n_185), .B(n_288), .Y(n_312) );
AND2x2_ASAP7_75t_L g324 ( .A(n_185), .B(n_315), .Y(n_324) );
NAND2xp5_ASAP7_75t_SL g347 ( .A(n_185), .B(n_252), .Y(n_347) );
INVx1_ASAP7_75t_SL g359 ( .A(n_185), .Y(n_359) );
INVx2_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
AND2x2_ASAP7_75t_L g251 ( .A(n_186), .B(n_252), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_186), .B(n_291), .Y(n_290) );
AOI21xp5_ASAP7_75t_L g190 ( .A1(n_191), .A2(n_193), .B(n_194), .Y(n_190) );
AOI21xp5_ASAP7_75t_L g257 ( .A1(n_194), .A2(n_258), .B(n_259), .Y(n_257) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
INVx3_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
INVx1_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
AND2x2_ASAP7_75t_L g199 ( .A(n_200), .B(n_210), .Y(n_199) );
AND2x2_ASAP7_75t_L g272 ( .A(n_200), .B(n_273), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_200), .B(n_225), .Y(n_276) );
AND2x2_ASAP7_75t_L g279 ( .A(n_200), .B(n_280), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_200), .B(n_282), .Y(n_281) );
OR2x2_ASAP7_75t_L g304 ( .A(n_200), .B(n_295), .Y(n_304) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_200), .Y(n_323) );
AND2x2_ASAP7_75t_L g344 ( .A(n_200), .B(n_345), .Y(n_344) );
OR2x2_ASAP7_75t_L g354 ( .A(n_200), .B(n_355), .Y(n_354) );
AND2x2_ASAP7_75t_L g400 ( .A(n_200), .B(n_283), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_200), .B(n_306), .Y(n_427) );
INVx5_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
BUFx2_ASAP7_75t_L g297 ( .A(n_201), .Y(n_297) );
AND2x2_ASAP7_75t_L g363 ( .A(n_201), .B(n_295), .Y(n_363) );
AND2x2_ASAP7_75t_L g447 ( .A(n_201), .B(n_315), .Y(n_447) );
OR2x6_ASAP7_75t_L g201 ( .A(n_202), .B(n_208), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_210), .B(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g436 ( .A(n_210), .Y(n_436) );
AND2x2_ASAP7_75t_L g210 ( .A(n_211), .B(n_225), .Y(n_210) );
AND2x2_ASAP7_75t_L g266 ( .A(n_211), .B(n_267), .Y(n_266) );
AND2x4_ASAP7_75t_L g275 ( .A(n_211), .B(n_273), .Y(n_275) );
INVx5_ASAP7_75t_L g283 ( .A(n_211), .Y(n_283) );
AND2x2_ASAP7_75t_L g306 ( .A(n_211), .B(n_237), .Y(n_306) );
HB1xp67_ASAP7_75t_L g343 ( .A(n_211), .Y(n_343) );
OR2x6_ASAP7_75t_L g211 ( .A(n_212), .B(n_222), .Y(n_211) );
AOI21xp5_ASAP7_75t_SL g212 ( .A1(n_213), .A2(n_215), .B(n_220), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_217), .A2(n_218), .B(n_219), .Y(n_216) );
INVx1_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g547 ( .A(n_221), .B(n_548), .Y(n_547) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_223), .B(n_224), .Y(n_222) );
AO21x2_ASAP7_75t_L g509 ( .A1(n_224), .A2(n_510), .B(n_517), .Y(n_509) );
INVx1_ASAP7_75t_L g384 ( .A(n_225), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_225), .B(n_400), .Y(n_399) );
AND2x2_ASAP7_75t_L g417 ( .A(n_225), .B(n_283), .Y(n_417) );
A2O1A1Ixp33_ASAP7_75t_L g446 ( .A1(n_225), .A2(n_340), .B(n_447), .C(n_448), .Y(n_446) );
AND2x2_ASAP7_75t_L g225 ( .A(n_226), .B(n_237), .Y(n_225) );
BUFx2_ASAP7_75t_L g267 ( .A(n_226), .Y(n_267) );
INVx2_ASAP7_75t_L g271 ( .A(n_226), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_228), .B(n_234), .Y(n_227) );
HB1xp67_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
INVx3_ASAP7_75t_L g556 ( .A(n_233), .Y(n_556) );
INVx2_ASAP7_75t_L g273 ( .A(n_237), .Y(n_273) );
AND2x2_ASAP7_75t_L g280 ( .A(n_237), .B(n_271), .Y(n_280) );
AND2x2_ASAP7_75t_L g371 ( .A(n_237), .B(n_283), .Y(n_371) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_244), .B(n_245), .Y(n_243) );
NOR2xp33_ASAP7_75t_L g554 ( .A(n_245), .B(n_555), .Y(n_554) );
INVx4_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
INVx2_ASAP7_75t_L g493 ( .A(n_246), .Y(n_493) );
INVx2_ASAP7_75t_L g516 ( .A(n_247), .Y(n_516) );
AOI211x1_ASAP7_75t_SL g249 ( .A1(n_250), .A2(n_264), .B(n_277), .C(n_302), .Y(n_249) );
INVx1_ASAP7_75t_L g368 ( .A(n_250), .Y(n_368) );
AND2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_263), .Y(n_250) );
INVx5_ASAP7_75t_SL g288 ( .A(n_252), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_252), .B(n_358), .Y(n_357) );
AOI311xp33_ASAP7_75t_L g376 ( .A1(n_252), .A2(n_377), .A3(n_379), .B(n_380), .C(n_386), .Y(n_376) );
A2O1A1Ixp33_ASAP7_75t_L g411 ( .A1(n_252), .A2(n_324), .B(n_412), .C(n_415), .Y(n_411) );
OAI21xp5_ASAP7_75t_L g253 ( .A1(n_254), .A2(n_255), .B(n_256), .Y(n_253) );
OAI21xp5_ASAP7_75t_L g510 ( .A1(n_255), .A2(n_511), .B(n_512), .Y(n_510) );
OAI21xp5_ASAP7_75t_L g541 ( .A1(n_255), .A2(n_542), .B(n_543), .Y(n_541) );
NOR2xp33_ASAP7_75t_L g260 ( .A(n_261), .B(n_262), .Y(n_260) );
INVx2_ASAP7_75t_L g584 ( .A(n_262), .Y(n_584) );
INVxp67_ASAP7_75t_L g331 ( .A(n_263), .Y(n_331) );
NAND4xp25_ASAP7_75t_SL g264 ( .A(n_265), .B(n_268), .C(n_274), .D(n_276), .Y(n_264) );
NOR2xp33_ASAP7_75t_L g329 ( .A(n_265), .B(n_330), .Y(n_329) );
INVx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g322 ( .A(n_266), .B(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_269), .B(n_272), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_269), .B(n_275), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_269), .B(n_282), .Y(n_402) );
BUFx2_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_270), .B(n_283), .Y(n_420) );
HB1xp67_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
INVx2_ASAP7_75t_L g295 ( .A(n_271), .Y(n_295) );
INVxp67_ASAP7_75t_L g330 ( .A(n_272), .Y(n_330) );
AND2x4_ASAP7_75t_L g282 ( .A(n_273), .B(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g356 ( .A(n_273), .B(n_295), .Y(n_356) );
INVx1_ASAP7_75t_L g383 ( .A(n_273), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_273), .B(n_370), .Y(n_430) );
NOR2xp33_ASAP7_75t_L g364 ( .A(n_274), .B(n_344), .Y(n_364) );
INVx1_ASAP7_75t_SL g274 ( .A(n_275), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_275), .B(n_297), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_275), .B(n_344), .Y(n_443) );
INVx1_ASAP7_75t_L g454 ( .A(n_276), .Y(n_454) );
A2O1A1Ixp33_ASAP7_75t_L g277 ( .A1(n_278), .A2(n_281), .B(n_284), .C(n_292), .Y(n_277) );
INVx1_ASAP7_75t_SL g278 ( .A(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g296 ( .A(n_280), .B(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g334 ( .A(n_280), .B(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g316 ( .A(n_281), .Y(n_316) );
AND2x2_ASAP7_75t_L g293 ( .A(n_282), .B(n_294), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_282), .B(n_344), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_282), .B(n_363), .Y(n_387) );
OR2x2_ASAP7_75t_L g303 ( .A(n_283), .B(n_304), .Y(n_303) );
INVx2_ASAP7_75t_L g335 ( .A(n_283), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_283), .B(n_295), .Y(n_350) );
AND2x2_ASAP7_75t_L g407 ( .A(n_283), .B(n_363), .Y(n_407) );
HB1xp67_ASAP7_75t_L g414 ( .A(n_283), .Y(n_414) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AOI221xp5_ASAP7_75t_L g418 ( .A1(n_285), .A2(n_297), .B1(n_419), .B2(n_421), .C(n_424), .Y(n_418) );
AND2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_289), .Y(n_285) );
INVx1_ASAP7_75t_SL g286 ( .A(n_287), .Y(n_286) );
OR2x2_ASAP7_75t_L g308 ( .A(n_288), .B(n_291), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_288), .B(n_358), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_288), .B(n_315), .Y(n_423) );
INVx1_ASAP7_75t_SL g289 ( .A(n_290), .Y(n_289) );
OR2x2_ASAP7_75t_L g408 ( .A(n_290), .B(n_409), .Y(n_408) );
OR2x2_ASAP7_75t_L g422 ( .A(n_290), .B(n_423), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_291), .B(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g319 ( .A(n_291), .B(n_312), .Y(n_319) );
AND2x2_ASAP7_75t_L g389 ( .A(n_291), .B(n_390), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_291), .B(n_338), .Y(n_435) );
NOR2xp33_ASAP7_75t_L g438 ( .A(n_291), .B(n_439), .Y(n_438) );
OAI21xp5_ASAP7_75t_SL g292 ( .A1(n_293), .A2(n_296), .B(n_298), .Y(n_292) );
INVx2_ASAP7_75t_L g325 ( .A(n_293), .Y(n_325) );
HB1xp67_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
INVx1_ASAP7_75t_L g345 ( .A(n_295), .Y(n_345) );
OR2x2_ASAP7_75t_L g349 ( .A(n_297), .B(n_350), .Y(n_349) );
OR2x2_ASAP7_75t_L g452 ( .A(n_297), .B(n_420), .Y(n_452) );
INVx1_ASAP7_75t_SL g298 ( .A(n_299), .Y(n_298) );
OR2x2_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
AOI21xp33_ASAP7_75t_SL g302 ( .A1(n_303), .A2(n_305), .B(n_307), .Y(n_302) );
INVx1_ASAP7_75t_L g456 ( .A(n_303), .Y(n_456) );
INVx2_ASAP7_75t_SL g370 ( .A(n_304), .Y(n_370) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
A2O1A1Ixp33_ASAP7_75t_L g451 ( .A1(n_307), .A2(n_388), .B(n_452), .C(n_453), .Y(n_451) );
OAI322xp33_ASAP7_75t_SL g320 ( .A1(n_308), .A2(n_321), .A3(n_324), .B1(n_325), .B2(n_326), .C1(n_328), .C2(n_331), .Y(n_320) );
INVx2_ASAP7_75t_L g340 ( .A(n_308), .Y(n_340) );
AOI221xp5_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_316), .B1(n_317), .B2(n_319), .C(n_320), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
OAI22xp33_ASAP7_75t_SL g386 ( .A1(n_311), .A2(n_387), .B1(n_388), .B2(n_391), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_312), .B(n_315), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_312), .B(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
OR2x2_ASAP7_75t_L g385 ( .A(n_314), .B(n_347), .Y(n_385) );
INVx1_ASAP7_75t_L g375 ( .A(n_315), .Y(n_375) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
AOI21xp5_ASAP7_75t_L g428 ( .A1(n_319), .A2(n_429), .B(n_431), .Y(n_428) );
AOI21xp33_ASAP7_75t_L g353 ( .A1(n_321), .A2(n_354), .B(n_357), .Y(n_353) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
NOR2xp67_ASAP7_75t_SL g382 ( .A(n_323), .B(n_383), .Y(n_382) );
NOR2xp33_ASAP7_75t_L g415 ( .A(n_323), .B(n_416), .Y(n_415) );
INVx1_ASAP7_75t_SL g439 ( .A(n_324), .Y(n_439) );
INVx1_ASAP7_75t_SL g326 ( .A(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
NAND4xp25_ASAP7_75t_L g332 ( .A(n_333), .B(n_360), .C(n_376), .D(n_392), .Y(n_332) );
AOI211xp5_ASAP7_75t_L g333 ( .A1(n_334), .A2(n_336), .B(n_341), .C(n_353), .Y(n_333) );
INVx1_ASAP7_75t_L g425 ( .A(n_334), .Y(n_425) );
AND2x2_ASAP7_75t_L g373 ( .A(n_335), .B(n_356), .Y(n_373) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_338), .B(n_340), .Y(n_337) );
INVx1_ASAP7_75t_SL g338 ( .A(n_339), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_340), .B(n_375), .Y(n_374) );
OAI22xp33_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_346), .B1(n_349), .B2(n_351), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_343), .B(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g391 ( .A(n_344), .Y(n_391) );
O2A1O1Ixp33_ASAP7_75t_L g405 ( .A1(n_344), .A2(n_383), .B(n_406), .C(n_408), .Y(n_405) );
OR2x2_ASAP7_75t_L g346 ( .A(n_347), .B(n_348), .Y(n_346) );
INVx1_ASAP7_75t_L g390 ( .A(n_347), .Y(n_390) );
INVx1_ASAP7_75t_L g450 ( .A(n_348), .Y(n_450) );
NAND2xp33_ASAP7_75t_SL g440 ( .A(n_349), .B(n_441), .Y(n_440) );
INVx1_ASAP7_75t_SL g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx2_ASAP7_75t_L g379 ( .A(n_358), .Y(n_379) );
O2A1O1Ixp33_ASAP7_75t_L g360 ( .A1(n_361), .A2(n_364), .B(n_365), .C(n_367), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
OAI22xp5_ASAP7_75t_L g367 ( .A1(n_368), .A2(n_369), .B1(n_372), .B2(n_374), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_370), .B(n_371), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_370), .B(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_375), .B(n_396), .Y(n_458) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
AOI21xp33_ASAP7_75t_SL g380 ( .A1(n_381), .A2(n_384), .B(n_385), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_SL g388 ( .A(n_389), .Y(n_388) );
AOI221xp5_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_398), .B1(n_401), .B2(n_403), .C(n_405), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_395), .B(n_396), .Y(n_394) );
INVx1_ASAP7_75t_SL g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVxp67_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
OAI22xp5_ASAP7_75t_L g424 ( .A1(n_408), .A2(n_425), .B1(n_426), .B2(n_427), .Y(n_424) );
NAND3xp33_ASAP7_75t_SL g410 ( .A(n_411), .B(n_418), .C(n_428), .Y(n_410) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_SL g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
CKINVDCx16_ASAP7_75t_R g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVxp67_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
OAI211xp5_ASAP7_75t_L g434 ( .A1(n_435), .A2(n_436), .B(n_437), .C(n_446), .Y(n_434) );
INVx1_ASAP7_75t_L g455 ( .A(n_435), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g437 ( .A1(n_438), .A2(n_440), .B1(n_442), .B2(n_444), .Y(n_437) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
AOI22xp5_ASAP7_75t_L g453 ( .A1(n_454), .A2(n_455), .B1(n_456), .B2(n_457), .Y(n_453) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_SL g460 ( .A(n_461), .Y(n_460) );
INVx1_ASAP7_75t_SL g461 ( .A(n_462), .Y(n_461) );
INVx2_ASAP7_75t_L g468 ( .A(n_462), .Y(n_468) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_465), .B(n_466), .Y(n_464) );
NAND3xp33_ASAP7_75t_L g469 ( .A(n_467), .B(n_470), .C(n_755), .Y(n_469) );
XNOR2xp5_ASAP7_75t_L g471 ( .A(n_472), .B(n_481), .Y(n_471) );
CKINVDCx20_ASAP7_75t_R g473 ( .A(n_474), .Y(n_473) );
CKINVDCx16_ASAP7_75t_R g476 ( .A(n_477), .Y(n_476) );
OR2x2_ASAP7_75t_L g483 ( .A(n_484), .B(n_680), .Y(n_483) );
NAND5xp2_ASAP7_75t_L g484 ( .A(n_485), .B(n_595), .C(n_627), .D(n_644), .E(n_667), .Y(n_484) );
AOI221xp5_ASAP7_75t_L g485 ( .A1(n_486), .A2(n_528), .B1(n_558), .B2(n_562), .C(n_566), .Y(n_485) );
INVx1_ASAP7_75t_L g707 ( .A(n_486), .Y(n_707) );
AND2x2_ASAP7_75t_L g486 ( .A(n_487), .B(n_507), .Y(n_486) );
AND3x2_ASAP7_75t_L g682 ( .A(n_487), .B(n_509), .C(n_683), .Y(n_682) );
AND2x2_ASAP7_75t_L g487 ( .A(n_488), .B(n_497), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_488), .B(n_564), .Y(n_563) );
BUFx3_ASAP7_75t_L g573 ( .A(n_488), .Y(n_573) );
AND2x2_ASAP7_75t_L g577 ( .A(n_488), .B(n_519), .Y(n_577) );
INVx2_ASAP7_75t_L g604 ( .A(n_488), .Y(n_604) );
OR2x2_ASAP7_75t_L g615 ( .A(n_488), .B(n_520), .Y(n_615) );
NOR2xp33_ASAP7_75t_L g634 ( .A(n_488), .B(n_508), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_488), .B(n_653), .Y(n_652) );
AND2x2_ASAP7_75t_L g694 ( .A(n_488), .B(n_520), .Y(n_694) );
HB1xp67_ASAP7_75t_L g576 ( .A(n_497), .Y(n_576) );
AND2x2_ASAP7_75t_L g635 ( .A(n_497), .B(n_636), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_497), .B(n_508), .Y(n_654) );
INVx1_ASAP7_75t_SL g497 ( .A(n_498), .Y(n_497) );
OR2x2_ASAP7_75t_L g565 ( .A(n_498), .B(n_508), .Y(n_565) );
HB1xp67_ASAP7_75t_L g572 ( .A(n_498), .Y(n_572) );
AND2x2_ASAP7_75t_L g621 ( .A(n_498), .B(n_520), .Y(n_621) );
NAND3xp33_ASAP7_75t_L g646 ( .A(n_498), .B(n_507), .C(n_604), .Y(n_646) );
AND2x2_ASAP7_75t_L g711 ( .A(n_498), .B(n_509), .Y(n_711) );
AND2x2_ASAP7_75t_L g745 ( .A(n_498), .B(n_508), .Y(n_745) );
INVxp67_ASAP7_75t_L g574 ( .A(n_507), .Y(n_574) );
AND2x2_ASAP7_75t_L g507 ( .A(n_508), .B(n_519), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_508), .B(n_604), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_508), .B(n_635), .Y(n_643) );
AND2x2_ASAP7_75t_L g693 ( .A(n_508), .B(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g721 ( .A(n_508), .Y(n_721) );
INVx4_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
AND2x2_ASAP7_75t_L g628 ( .A(n_509), .B(n_621), .Y(n_628) );
BUFx3_ASAP7_75t_L g660 ( .A(n_509), .Y(n_660) );
INVx2_ASAP7_75t_L g636 ( .A(n_519), .Y(n_636) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
HB1xp67_ASAP7_75t_L g605 ( .A(n_520), .Y(n_605) );
AOI22xp33_ASAP7_75t_L g695 ( .A1(n_528), .A2(n_696), .B1(n_698), .B2(n_699), .Y(n_695) );
AND2x2_ASAP7_75t_L g528 ( .A(n_529), .B(n_538), .Y(n_528) );
AND2x2_ASAP7_75t_L g558 ( .A(n_529), .B(n_559), .Y(n_558) );
INVx3_ASAP7_75t_SL g569 ( .A(n_529), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_529), .B(n_599), .Y(n_631) );
OR2x2_ASAP7_75t_L g650 ( .A(n_529), .B(n_539), .Y(n_650) );
AND2x2_ASAP7_75t_L g655 ( .A(n_529), .B(n_607), .Y(n_655) );
AND2x2_ASAP7_75t_L g658 ( .A(n_529), .B(n_600), .Y(n_658) );
AND2x2_ASAP7_75t_L g670 ( .A(n_529), .B(n_549), .Y(n_670) );
AND2x2_ASAP7_75t_L g686 ( .A(n_529), .B(n_540), .Y(n_686) );
AND2x4_ASAP7_75t_L g689 ( .A(n_529), .B(n_560), .Y(n_689) );
OR2x2_ASAP7_75t_L g706 ( .A(n_529), .B(n_642), .Y(n_706) );
OR2x2_ASAP7_75t_L g737 ( .A(n_529), .B(n_582), .Y(n_737) );
NAND2xp5_ASAP7_75t_SL g739 ( .A(n_529), .B(n_665), .Y(n_739) );
OR2x6_ASAP7_75t_L g529 ( .A(n_530), .B(n_536), .Y(n_529) );
AND2x2_ASAP7_75t_L g613 ( .A(n_538), .B(n_580), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_538), .B(n_600), .Y(n_732) );
AND2x2_ASAP7_75t_L g538 ( .A(n_539), .B(n_549), .Y(n_538) );
AND2x2_ASAP7_75t_L g568 ( .A(n_539), .B(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g599 ( .A(n_539), .B(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g607 ( .A(n_539), .B(n_582), .Y(n_607) );
AND2x2_ASAP7_75t_L g625 ( .A(n_539), .B(n_560), .Y(n_625) );
OR2x2_ASAP7_75t_L g642 ( .A(n_539), .B(n_600), .Y(n_642) );
INVx2_ASAP7_75t_SL g539 ( .A(n_540), .Y(n_539) );
BUFx2_ASAP7_75t_L g561 ( .A(n_540), .Y(n_561) );
AND2x2_ASAP7_75t_L g665 ( .A(n_540), .B(n_549), .Y(n_665) );
INVx2_ASAP7_75t_L g560 ( .A(n_549), .Y(n_560) );
INVx1_ASAP7_75t_L g677 ( .A(n_549), .Y(n_677) );
AND2x2_ASAP7_75t_L g727 ( .A(n_549), .B(n_569), .Y(n_727) );
AND2x2_ASAP7_75t_L g579 ( .A(n_559), .B(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g611 ( .A(n_559), .B(n_569), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_559), .B(n_658), .Y(n_657) );
AND2x2_ASAP7_75t_L g559 ( .A(n_560), .B(n_561), .Y(n_559) );
AND2x2_ASAP7_75t_L g598 ( .A(n_560), .B(n_569), .Y(n_598) );
OR2x2_ASAP7_75t_L g714 ( .A(n_561), .B(n_688), .Y(n_714) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_564), .B(n_694), .Y(n_700) );
INVx2_ASAP7_75t_SL g564 ( .A(n_565), .Y(n_564) );
OAI32xp33_ASAP7_75t_L g656 ( .A1(n_565), .A2(n_657), .A3(n_659), .B1(n_661), .B2(n_662), .Y(n_656) );
OR2x2_ASAP7_75t_L g673 ( .A(n_565), .B(n_615), .Y(n_673) );
OAI21xp33_ASAP7_75t_SL g698 ( .A1(n_565), .A2(n_575), .B(n_603), .Y(n_698) );
OAI22xp33_ASAP7_75t_L g566 ( .A1(n_567), .A2(n_570), .B1(n_575), .B2(n_578), .Y(n_566) );
INVxp33_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_568), .B(n_639), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_569), .B(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g624 ( .A(n_569), .B(n_625), .Y(n_624) );
AND2x2_ASAP7_75t_L g724 ( .A(n_569), .B(n_665), .Y(n_724) );
OR2x2_ASAP7_75t_L g748 ( .A(n_569), .B(n_642), .Y(n_748) );
AOI21xp33_ASAP7_75t_L g731 ( .A1(n_570), .A2(n_630), .B(n_732), .Y(n_731) );
OR2x2_ASAP7_75t_L g570 ( .A(n_571), .B(n_574), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_572), .B(n_573), .Y(n_571) );
INVx1_ASAP7_75t_L g608 ( .A(n_572), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_572), .B(n_577), .Y(n_626) );
AND2x2_ASAP7_75t_L g648 ( .A(n_573), .B(n_621), .Y(n_648) );
INVx1_ASAP7_75t_L g661 ( .A(n_573), .Y(n_661) );
OR2x2_ASAP7_75t_L g666 ( .A(n_573), .B(n_600), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
NOR2xp33_ASAP7_75t_L g614 ( .A(n_576), .B(n_615), .Y(n_614) );
OAI22xp33_ASAP7_75t_L g596 ( .A1(n_577), .A2(n_597), .B1(n_602), .B2(n_606), .Y(n_596) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
OAI22xp5_ASAP7_75t_L g645 ( .A1(n_580), .A2(n_639), .B1(n_646), .B2(n_647), .Y(n_645) );
AND2x2_ASAP7_75t_L g723 ( .A(n_580), .B(n_724), .Y(n_723) );
INVx2_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx1_ASAP7_75t_SL g581 ( .A(n_582), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_582), .B(n_677), .Y(n_676) );
AND2x2_ASAP7_75t_L g742 ( .A(n_582), .B(n_625), .Y(n_742) );
AO21x2_ASAP7_75t_L g582 ( .A1(n_583), .A2(n_585), .B(n_593), .Y(n_582) );
INVx1_ASAP7_75t_L g601 ( .A(n_583), .Y(n_601) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
OA21x2_ASAP7_75t_L g600 ( .A1(n_586), .A2(n_594), .B(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
AOI221xp5_ASAP7_75t_L g595 ( .A1(n_596), .A2(n_608), .B1(n_609), .B2(n_614), .C(n_616), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_598), .B(n_599), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_598), .B(n_600), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_598), .B(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g617 ( .A(n_599), .Y(n_617) );
O2A1O1Ixp33_ASAP7_75t_L g704 ( .A1(n_599), .A2(n_705), .B(n_706), .C(n_707), .Y(n_704) );
AND2x2_ASAP7_75t_L g709 ( .A(n_599), .B(n_689), .Y(n_709) );
O2A1O1Ixp33_ASAP7_75t_SL g747 ( .A1(n_599), .A2(n_688), .B(n_748), .C(n_749), .Y(n_747) );
BUFx3_ASAP7_75t_L g639 ( .A(n_600), .Y(n_639) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_603), .B(n_660), .Y(n_703) );
AOI211xp5_ASAP7_75t_L g722 ( .A1(n_603), .A2(n_723), .B(n_725), .C(n_731), .Y(n_722) );
AND2x2_ASAP7_75t_L g603 ( .A(n_604), .B(n_605), .Y(n_603) );
INVxp67_ASAP7_75t_L g683 ( .A(n_605), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_607), .B(n_727), .Y(n_726) );
NAND2xp5_ASAP7_75t_SL g609 ( .A(n_610), .B(n_612), .Y(n_609) );
INVx1_ASAP7_75t_SL g610 ( .A(n_611), .Y(n_610) );
AOI211xp5_ASAP7_75t_L g627 ( .A1(n_611), .A2(n_628), .B(n_629), .C(n_637), .Y(n_627) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g712 ( .A(n_615), .Y(n_712) );
OR2x2_ASAP7_75t_L g729 ( .A(n_615), .B(n_659), .Y(n_729) );
OAI22xp5_ASAP7_75t_L g616 ( .A1(n_617), .A2(n_618), .B1(n_623), .B2(n_626), .Y(n_616) );
OAI22xp33_ASAP7_75t_L g629 ( .A1(n_618), .A2(n_630), .B1(n_631), .B2(n_632), .Y(n_629) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
NOR2xp33_ASAP7_75t_L g619 ( .A(n_620), .B(n_622), .Y(n_619) );
OR2x2_ASAP7_75t_L g716 ( .A(n_620), .B(n_660), .Y(n_716) );
INVx1_ASAP7_75t_SL g620 ( .A(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g671 ( .A(n_621), .B(n_661), .Y(n_671) );
INVx1_ASAP7_75t_L g679 ( .A(n_622), .Y(n_679) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_625), .B(n_639), .Y(n_687) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
AND2x2_ASAP7_75t_L g633 ( .A(n_634), .B(n_635), .Y(n_633) );
NAND2xp5_ASAP7_75t_SL g678 ( .A(n_635), .B(n_679), .Y(n_678) );
INVx2_ASAP7_75t_L g744 ( .A(n_636), .Y(n_744) );
AOI21xp33_ASAP7_75t_L g637 ( .A1(n_638), .A2(n_640), .B(n_643), .Y(n_637) );
INVx1_ASAP7_75t_L g674 ( .A(n_638), .Y(n_674) );
NAND2xp5_ASAP7_75t_SL g649 ( .A(n_639), .B(n_650), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_639), .B(n_670), .Y(n_669) );
NAND2x1p5_ASAP7_75t_L g690 ( .A(n_639), .B(n_665), .Y(n_690) );
NAND2xp5_ASAP7_75t_SL g697 ( .A(n_639), .B(n_686), .Y(n_697) );
OAI211xp5_ASAP7_75t_L g701 ( .A1(n_639), .A2(n_649), .B(n_689), .C(n_702), .Y(n_701) );
INVx1_ASAP7_75t_SL g641 ( .A(n_642), .Y(n_641) );
AOI221xp5_ASAP7_75t_SL g644 ( .A1(n_645), .A2(n_649), .B1(n_651), .B2(n_655), .C(n_656), .Y(n_644) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVxp67_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_653), .B(n_661), .Y(n_735) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
O2A1O1Ixp33_ASAP7_75t_L g746 ( .A1(n_655), .A2(n_670), .B(n_672), .C(n_747), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_658), .B(n_665), .Y(n_730) );
NAND2xp5_ASAP7_75t_SL g749 ( .A(n_659), .B(n_712), .Y(n_749) );
CKINVDCx16_ASAP7_75t_R g659 ( .A(n_660), .Y(n_659) );
INVxp33_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
NOR2xp33_ASAP7_75t_L g663 ( .A(n_664), .B(n_666), .Y(n_663) );
AOI21xp33_ASAP7_75t_SL g675 ( .A1(n_664), .A2(n_676), .B(n_678), .Y(n_675) );
NOR2xp33_ASAP7_75t_L g736 ( .A(n_664), .B(n_737), .Y(n_736) );
INVx2_ASAP7_75t_SL g664 ( .A(n_665), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_665), .B(n_719), .Y(n_718) );
AOI221xp5_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_671), .B1(n_672), .B2(n_674), .C(n_675), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_671), .B(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g705 ( .A(n_677), .Y(n_705) );
NAND5xp2_ASAP7_75t_L g680 ( .A(n_681), .B(n_708), .C(n_722), .D(n_733), .E(n_746), .Y(n_680) );
AOI211xp5_ASAP7_75t_L g681 ( .A1(n_682), .A2(n_684), .B(n_691), .C(n_704), .Y(n_681) );
INVx2_ASAP7_75t_SL g728 ( .A(n_682), .Y(n_728) );
NAND4xp25_ASAP7_75t_SL g684 ( .A(n_685), .B(n_687), .C(n_688), .D(n_690), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx3_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
OAI211xp5_ASAP7_75t_SL g691 ( .A1(n_690), .A2(n_692), .B(n_695), .C(n_701), .Y(n_691) );
CKINVDCx20_ASAP7_75t_R g692 ( .A(n_693), .Y(n_692) );
AOI221xp5_ASAP7_75t_L g733 ( .A1(n_693), .A2(n_734), .B1(n_736), .B2(n_738), .C(n_740), .Y(n_733) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
AOI221xp5_ASAP7_75t_SL g708 ( .A1(n_709), .A2(n_710), .B1(n_713), .B2(n_715), .C(n_717), .Y(n_708) );
AND2x2_ASAP7_75t_L g710 ( .A(n_711), .B(n_712), .Y(n_710) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
OAI22xp5_ASAP7_75t_L g740 ( .A1(n_716), .A2(n_739), .B1(n_741), .B2(n_743), .Y(n_740) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_SL g719 ( .A(n_720), .Y(n_719) );
OAI22xp5_ASAP7_75t_L g725 ( .A1(n_726), .A2(n_728), .B1(n_729), .B2(n_730), .Y(n_725) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_SL g741 ( .A(n_742), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_744), .B(n_745), .Y(n_743) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx2_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx2_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
endmodule