module real_aes_7311_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_754;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_602;
wire n_552;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_741;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g499 ( .A1(n_0), .A2(n_163), .B(n_500), .C(n_503), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_1), .B(n_495), .Y(n_504) );
AOI22xp33_ASAP7_75t_L g100 ( .A1(n_2), .A2(n_101), .B1(n_112), .B2(n_754), .Y(n_100) );
INVx1_ASAP7_75t_L g110 ( .A(n_3), .Y(n_110) );
INVx1_ASAP7_75t_L g161 ( .A(n_4), .Y(n_161) );
NAND2xp5_ASAP7_75t_SL g568 ( .A(n_5), .B(n_164), .Y(n_568) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_6), .A2(n_463), .B(n_539), .Y(n_538) );
AO21x2_ASAP7_75t_L g517 ( .A1(n_7), .A2(n_171), .B(n_518), .Y(n_517) );
AOI22xp33_ASAP7_75t_L g217 ( .A1(n_8), .A2(n_36), .B1(n_151), .B2(n_199), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_9), .B(n_171), .Y(n_179) );
AND2x6_ASAP7_75t_L g166 ( .A(n_10), .B(n_167), .Y(n_166) );
A2O1A1Ixp33_ASAP7_75t_L g511 ( .A1(n_11), .A2(n_166), .B(n_468), .C(n_512), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g111 ( .A(n_12), .B(n_37), .Y(n_111) );
INVx1_ASAP7_75t_L g145 ( .A(n_13), .Y(n_145) );
INVx1_ASAP7_75t_L g142 ( .A(n_14), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_15), .B(n_147), .Y(n_208) );
NAND2xp5_ASAP7_75t_SL g523 ( .A(n_16), .B(n_164), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_17), .B(n_138), .Y(n_245) );
AO32x2_ASAP7_75t_L g215 ( .A1(n_18), .A2(n_137), .A3(n_171), .B1(n_190), .B2(n_216), .Y(n_215) );
AOI222xp33_ASAP7_75t_SL g121 ( .A1(n_19), .A2(n_40), .B1(n_122), .B2(n_741), .C1(n_742), .C2(n_744), .Y(n_121) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_20), .B(n_151), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_21), .B(n_138), .Y(n_168) );
AOI22xp33_ASAP7_75t_L g218 ( .A1(n_22), .A2(n_54), .B1(n_151), .B2(n_199), .Y(n_218) );
AOI22xp33_ASAP7_75t_SL g201 ( .A1(n_23), .A2(n_80), .B1(n_147), .B2(n_151), .Y(n_201) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_24), .B(n_151), .Y(n_231) );
A2O1A1Ixp33_ASAP7_75t_L g485 ( .A1(n_25), .A2(n_190), .B(n_468), .C(n_486), .Y(n_485) );
A2O1A1Ixp33_ASAP7_75t_L g520 ( .A1(n_26), .A2(n_190), .B(n_468), .C(n_521), .Y(n_520) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_27), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_28), .B(n_192), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g496 ( .A1(n_29), .A2(n_463), .B(n_497), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_30), .B(n_192), .Y(n_233) );
INVx2_ASAP7_75t_L g149 ( .A(n_31), .Y(n_149) );
A2O1A1Ixp33_ASAP7_75t_L g465 ( .A1(n_32), .A2(n_466), .B(n_470), .C(n_476), .Y(n_465) );
NAND2xp5_ASAP7_75t_SL g183 ( .A(n_33), .B(n_151), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_34), .B(n_192), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_35), .B(n_210), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_38), .B(n_484), .Y(n_483) );
CKINVDCx20_ASAP7_75t_R g516 ( .A(n_39), .Y(n_516) );
INVx1_ASAP7_75t_L g741 ( .A(n_40), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_41), .B(n_164), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_42), .B(n_463), .Y(n_519) );
OAI22xp5_ASAP7_75t_SL g124 ( .A1(n_43), .A2(n_125), .B1(n_126), .B2(n_447), .Y(n_124) );
INVx1_ASAP7_75t_L g447 ( .A(n_43), .Y(n_447) );
OAI22xp5_ASAP7_75t_SL g752 ( .A1(n_43), .A2(n_45), .B1(n_447), .B2(n_753), .Y(n_752) );
A2O1A1Ixp33_ASAP7_75t_L g530 ( .A1(n_44), .A2(n_466), .B(n_476), .C(n_531), .Y(n_530) );
CKINVDCx20_ASAP7_75t_R g753 ( .A(n_45), .Y(n_753) );
NAND2xp5_ASAP7_75t_SL g174 ( .A(n_46), .B(n_151), .Y(n_174) );
INVx1_ASAP7_75t_L g501 ( .A(n_47), .Y(n_501) );
AOI22xp33_ASAP7_75t_L g198 ( .A1(n_48), .A2(n_89), .B1(n_199), .B2(n_200), .Y(n_198) );
INVx1_ASAP7_75t_L g532 ( .A(n_49), .Y(n_532) );
NAND2xp5_ASAP7_75t_SL g177 ( .A(n_50), .B(n_151), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_51), .B(n_151), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_52), .B(n_463), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_53), .B(n_159), .Y(n_178) );
AOI22xp33_ASAP7_75t_SL g243 ( .A1(n_55), .A2(n_59), .B1(n_147), .B2(n_151), .Y(n_243) );
CKINVDCx20_ASAP7_75t_R g491 ( .A(n_56), .Y(n_491) );
NAND2xp5_ASAP7_75t_SL g187 ( .A(n_57), .B(n_151), .Y(n_187) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_58), .B(n_151), .Y(n_207) );
INVx1_ASAP7_75t_L g167 ( .A(n_60), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_61), .B(n_463), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_62), .B(n_495), .Y(n_544) );
A2O1A1Ixp33_ASAP7_75t_L g541 ( .A1(n_63), .A2(n_153), .B(n_159), .C(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_64), .B(n_151), .Y(n_162) );
INVx1_ASAP7_75t_L g141 ( .A(n_65), .Y(n_141) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_66), .Y(n_117) );
NAND2xp5_ASAP7_75t_SL g474 ( .A(n_67), .B(n_164), .Y(n_474) );
AO32x2_ASAP7_75t_L g196 ( .A1(n_68), .A2(n_171), .A3(n_190), .B1(n_197), .B2(n_202), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_69), .B(n_165), .Y(n_513) );
INVx1_ASAP7_75t_L g186 ( .A(n_70), .Y(n_186) );
INVx1_ASAP7_75t_L g228 ( .A(n_71), .Y(n_228) );
CKINVDCx16_ASAP7_75t_R g498 ( .A(n_72), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_73), .B(n_473), .Y(n_487) );
A2O1A1Ixp33_ASAP7_75t_L g565 ( .A1(n_74), .A2(n_468), .B(n_476), .C(n_566), .Y(n_565) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_75), .B(n_147), .Y(n_229) );
CKINVDCx16_ASAP7_75t_R g540 ( .A(n_76), .Y(n_540) );
INVx1_ASAP7_75t_L g105 ( .A(n_77), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_78), .Y(n_120) );
NAND2xp5_ASAP7_75t_SL g488 ( .A(n_79), .B(n_472), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_81), .B(n_199), .Y(n_213) );
CKINVDCx20_ASAP7_75t_R g479 ( .A(n_82), .Y(n_479) );
NAND2xp5_ASAP7_75t_SL g232 ( .A(n_83), .B(n_147), .Y(n_232) );
INVx2_ASAP7_75t_L g139 ( .A(n_84), .Y(n_139) );
CKINVDCx20_ASAP7_75t_R g572 ( .A(n_85), .Y(n_572) );
NAND2xp5_ASAP7_75t_SL g514 ( .A(n_86), .B(n_189), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_87), .B(n_147), .Y(n_175) );
OR2x2_ASAP7_75t_L g107 ( .A(n_88), .B(n_108), .Y(n_107) );
OR2x2_ASAP7_75t_L g450 ( .A(n_88), .B(n_109), .Y(n_450) );
INVx2_ASAP7_75t_L g454 ( .A(n_88), .Y(n_454) );
AOI22xp33_ASAP7_75t_L g242 ( .A1(n_90), .A2(n_99), .B1(n_147), .B2(n_148), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_91), .B(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g471 ( .A(n_92), .Y(n_471) );
INVxp67_ASAP7_75t_L g543 ( .A(n_93), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_94), .B(n_147), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g104 ( .A(n_95), .B(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g509 ( .A(n_96), .Y(n_509) );
INVx1_ASAP7_75t_L g567 ( .A(n_97), .Y(n_567) );
AND2x2_ASAP7_75t_L g534 ( .A(n_98), .B(n_192), .Y(n_534) );
INVx1_ASAP7_75t_SL g101 ( .A(n_102), .Y(n_101) );
INVx1_ASAP7_75t_L g755 ( .A(n_102), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g102 ( .A(n_103), .B(n_106), .Y(n_102) );
INVx1_ASAP7_75t_SL g103 ( .A(n_104), .Y(n_103) );
INVx1_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
HB1xp67_ASAP7_75t_L g119 ( .A(n_107), .Y(n_119) );
AOI21xp5_ASAP7_75t_L g749 ( .A1(n_107), .A2(n_118), .B(n_750), .Y(n_749) );
NOR2x2_ASAP7_75t_L g746 ( .A(n_108), .B(n_454), .Y(n_746) );
INVx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
OR2x2_ASAP7_75t_L g453 ( .A(n_109), .B(n_454), .Y(n_453) );
AND2x2_ASAP7_75t_L g109 ( .A(n_110), .B(n_111), .Y(n_109) );
BUFx3_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
AOI22xp5_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_121), .B1(n_747), .B2(n_749), .Y(n_113) );
NOR2xp33_ASAP7_75t_L g114 ( .A(n_115), .B(n_118), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx2_ASAP7_75t_L g748 ( .A(n_117), .Y(n_748) );
NOR2xp33_ASAP7_75t_SL g118 ( .A(n_119), .B(n_120), .Y(n_118) );
OAI22x1_ASAP7_75t_SL g122 ( .A1(n_123), .A2(n_448), .B1(n_451), .B2(n_455), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
OAI22xp5_ASAP7_75t_SL g742 ( .A1(n_124), .A2(n_448), .B1(n_453), .B2(n_743), .Y(n_742) );
OAI22xp5_ASAP7_75t_SL g750 ( .A1(n_125), .A2(n_126), .B1(n_751), .B2(n_752), .Y(n_750) );
INVx1_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
AND2x2_ASAP7_75t_SL g126 ( .A(n_127), .B(n_413), .Y(n_126) );
NOR3xp33_ASAP7_75t_L g127 ( .A(n_128), .B(n_317), .C(n_401), .Y(n_127) );
NAND4xp25_ASAP7_75t_L g128 ( .A(n_129), .B(n_260), .C(n_282), .D(n_298), .Y(n_128) );
AOI221xp5_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_193), .B1(n_219), .B2(n_238), .C(n_246), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_132), .B(n_169), .Y(n_131) );
NAND2xp5_ASAP7_75t_SL g272 ( .A(n_132), .B(n_238), .Y(n_272) );
NAND4xp25_ASAP7_75t_L g312 ( .A(n_132), .B(n_300), .C(n_313), .D(n_315), .Y(n_312) );
INVxp67_ASAP7_75t_L g429 ( .A(n_132), .Y(n_429) );
INVx3_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
OR2x2_ASAP7_75t_L g311 ( .A(n_133), .B(n_249), .Y(n_311) );
AND2x2_ASAP7_75t_L g335 ( .A(n_133), .B(n_169), .Y(n_335) );
INVx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
AND2x2_ASAP7_75t_L g302 ( .A(n_134), .B(n_237), .Y(n_302) );
AND2x2_ASAP7_75t_L g342 ( .A(n_134), .B(n_323), .Y(n_342) );
AND2x2_ASAP7_75t_L g359 ( .A(n_134), .B(n_360), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_134), .B(n_170), .Y(n_383) );
INVx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
AND2x2_ASAP7_75t_L g236 ( .A(n_135), .B(n_237), .Y(n_236) );
AND2x2_ASAP7_75t_L g254 ( .A(n_135), .B(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g266 ( .A(n_135), .B(n_170), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_135), .B(n_180), .Y(n_288) );
OA21x2_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_143), .B(n_168), .Y(n_135) );
OA21x2_ASAP7_75t_L g180 ( .A1(n_136), .A2(n_181), .B(n_191), .Y(n_180) );
INVx2_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
NOR2xp33_ASAP7_75t_L g515 ( .A(n_137), .B(n_516), .Y(n_515) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_138), .Y(n_171) );
AND2x2_ASAP7_75t_L g138 ( .A(n_139), .B(n_140), .Y(n_138) );
AND2x2_ASAP7_75t_SL g192 ( .A(n_139), .B(n_140), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_141), .B(n_142), .Y(n_140) );
OAI21xp5_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_157), .B(n_166), .Y(n_143) );
O2A1O1Ixp33_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_146), .B(n_150), .C(n_153), .Y(n_144) );
AOI21xp5_ASAP7_75t_L g512 ( .A1(n_146), .A2(n_513), .B(n_514), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_146), .A2(n_522), .B(n_523), .Y(n_521) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx3_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx2_ASAP7_75t_L g152 ( .A(n_149), .Y(n_152) );
INVx1_ASAP7_75t_L g160 ( .A(n_149), .Y(n_160) );
INVx3_ASAP7_75t_L g227 ( .A(n_151), .Y(n_227) );
HB1xp67_ASAP7_75t_L g569 ( .A(n_151), .Y(n_569) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g199 ( .A(n_152), .Y(n_199) );
BUFx3_ASAP7_75t_L g200 ( .A(n_152), .Y(n_200) );
AND2x6_ASAP7_75t_L g468 ( .A(n_152), .B(n_469), .Y(n_468) );
O2A1O1Ixp33_ASAP7_75t_L g566 ( .A1(n_153), .A2(n_567), .B(n_568), .C(n_569), .Y(n_566) );
INVx1_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_154), .A2(n_231), .B(n_232), .Y(n_230) );
INVx4_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx2_ASAP7_75t_L g473 ( .A(n_155), .Y(n_473) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx3_ASAP7_75t_L g165 ( .A(n_156), .Y(n_165) );
BUFx6f_ASAP7_75t_L g189 ( .A(n_156), .Y(n_189) );
INVx1_ASAP7_75t_L g210 ( .A(n_156), .Y(n_210) );
AND2x2_ASAP7_75t_L g464 ( .A(n_156), .B(n_160), .Y(n_464) );
INVx1_ASAP7_75t_L g469 ( .A(n_156), .Y(n_469) );
O2A1O1Ixp33_ASAP7_75t_L g157 ( .A1(n_158), .A2(n_161), .B(n_162), .C(n_163), .Y(n_157) );
O2A1O1Ixp5_ASAP7_75t_L g185 ( .A1(n_158), .A2(n_186), .B(n_187), .C(n_188), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g486 ( .A1(n_158), .A2(n_487), .B(n_488), .Y(n_486) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
AOI21xp5_ASAP7_75t_L g176 ( .A1(n_163), .A2(n_177), .B(n_178), .Y(n_176) );
OAI22xp5_ASAP7_75t_L g216 ( .A1(n_163), .A2(n_189), .B1(n_217), .B2(n_218), .Y(n_216) );
OAI22xp5_ASAP7_75t_L g241 ( .A1(n_163), .A2(n_189), .B1(n_242), .B2(n_243), .Y(n_241) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
AOI21xp5_ASAP7_75t_L g173 ( .A1(n_164), .A2(n_174), .B(n_175), .Y(n_173) );
AOI21xp5_ASAP7_75t_L g182 ( .A1(n_164), .A2(n_183), .B(n_184), .Y(n_182) );
O2A1O1Ixp5_ASAP7_75t_SL g226 ( .A1(n_164), .A2(n_227), .B(n_228), .C(n_229), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g542 ( .A(n_164), .B(n_543), .Y(n_542) );
INVx5_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
OAI22xp5_ASAP7_75t_SL g197 ( .A1(n_165), .A2(n_189), .B1(n_198), .B2(n_201), .Y(n_197) );
OAI21xp5_ASAP7_75t_L g172 ( .A1(n_166), .A2(n_173), .B(n_176), .Y(n_172) );
BUFx3_ASAP7_75t_L g190 ( .A(n_166), .Y(n_190) );
OAI21xp5_ASAP7_75t_L g205 ( .A1(n_166), .A2(n_206), .B(n_211), .Y(n_205) );
OAI21xp5_ASAP7_75t_L g225 ( .A1(n_166), .A2(n_226), .B(n_230), .Y(n_225) );
AND2x4_ASAP7_75t_L g463 ( .A(n_166), .B(n_464), .Y(n_463) );
INVx4_ASAP7_75t_SL g477 ( .A(n_166), .Y(n_477) );
NAND2x1p5_ASAP7_75t_L g510 ( .A(n_166), .B(n_464), .Y(n_510) );
AND2x2_ASAP7_75t_L g269 ( .A(n_169), .B(n_270), .Y(n_269) );
AOI221xp5_ASAP7_75t_L g318 ( .A1(n_169), .A2(n_319), .B1(n_322), .B2(n_324), .C(n_328), .Y(n_318) );
AND2x2_ASAP7_75t_L g377 ( .A(n_169), .B(n_342), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_169), .B(n_359), .Y(n_411) );
AND2x2_ASAP7_75t_L g169 ( .A(n_170), .B(n_180), .Y(n_169) );
INVx3_ASAP7_75t_L g237 ( .A(n_170), .Y(n_237) );
AND2x2_ASAP7_75t_L g286 ( .A(n_170), .B(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g340 ( .A(n_170), .B(n_255), .Y(n_340) );
AND2x2_ASAP7_75t_L g398 ( .A(n_170), .B(n_399), .Y(n_398) );
OA21x2_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_172), .B(n_179), .Y(n_170) );
INVx4_ASAP7_75t_L g240 ( .A(n_171), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_171), .A2(n_519), .B(n_520), .Y(n_518) );
HB1xp67_ASAP7_75t_L g537 ( .A(n_171), .Y(n_537) );
AND2x2_ASAP7_75t_L g238 ( .A(n_180), .B(n_239), .Y(n_238) );
INVx2_ASAP7_75t_L g255 ( .A(n_180), .Y(n_255) );
INVx1_ASAP7_75t_L g310 ( .A(n_180), .Y(n_310) );
HB1xp67_ASAP7_75t_L g316 ( .A(n_180), .Y(n_316) );
AND2x2_ASAP7_75t_L g361 ( .A(n_180), .B(n_237), .Y(n_361) );
OR2x2_ASAP7_75t_L g400 ( .A(n_180), .B(n_239), .Y(n_400) );
OAI21xp5_ASAP7_75t_L g181 ( .A1(n_182), .A2(n_185), .B(n_190), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_188), .A2(n_212), .B(n_213), .Y(n_211) );
INVx2_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
INVx4_ASAP7_75t_L g502 ( .A(n_189), .Y(n_502) );
NAND3xp33_ASAP7_75t_L g259 ( .A(n_190), .B(n_240), .C(n_241), .Y(n_259) );
INVx2_ASAP7_75t_L g202 ( .A(n_192), .Y(n_202) );
OA21x2_ASAP7_75t_L g204 ( .A1(n_192), .A2(n_205), .B(n_214), .Y(n_204) );
OA21x2_ASAP7_75t_L g224 ( .A1(n_192), .A2(n_225), .B(n_233), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g461 ( .A1(n_192), .A2(n_462), .B(n_465), .Y(n_461) );
INVx1_ASAP7_75t_L g492 ( .A(n_192), .Y(n_492) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_192), .A2(n_529), .B(n_530), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_193), .B(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g193 ( .A(n_194), .B(n_203), .Y(n_193) );
AND2x2_ASAP7_75t_L g396 ( .A(n_194), .B(n_393), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_194), .B(n_378), .Y(n_428) );
BUFx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
AND2x2_ASAP7_75t_L g327 ( .A(n_195), .B(n_251), .Y(n_327) );
AND2x2_ASAP7_75t_L g376 ( .A(n_195), .B(n_222), .Y(n_376) );
INVx1_ASAP7_75t_L g422 ( .A(n_195), .Y(n_422) );
INVx1_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
BUFx6f_ASAP7_75t_L g235 ( .A(n_196), .Y(n_235) );
AND2x2_ASAP7_75t_L g277 ( .A(n_196), .B(n_251), .Y(n_277) );
INVx1_ASAP7_75t_L g294 ( .A(n_196), .Y(n_294) );
AND2x2_ASAP7_75t_L g300 ( .A(n_196), .B(n_215), .Y(n_300) );
HB1xp67_ASAP7_75t_L g475 ( .A(n_200), .Y(n_475) );
INVx2_ASAP7_75t_L g503 ( .A(n_200), .Y(n_503) );
INVx1_ASAP7_75t_L g489 ( .A(n_202), .Y(n_489) );
AND2x2_ASAP7_75t_L g368 ( .A(n_203), .B(n_276), .Y(n_368) );
INVx2_ASAP7_75t_L g433 ( .A(n_203), .Y(n_433) );
AND2x2_ASAP7_75t_L g203 ( .A(n_204), .B(n_215), .Y(n_203) );
AND2x2_ASAP7_75t_L g250 ( .A(n_204), .B(n_251), .Y(n_250) );
OR2x2_ASAP7_75t_L g263 ( .A(n_204), .B(n_223), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_204), .B(n_222), .Y(n_291) );
INVx1_ASAP7_75t_L g297 ( .A(n_204), .Y(n_297) );
INVx1_ASAP7_75t_L g314 ( .A(n_204), .Y(n_314) );
HB1xp67_ASAP7_75t_L g326 ( .A(n_204), .Y(n_326) );
INVx2_ASAP7_75t_L g394 ( .A(n_204), .Y(n_394) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_207), .A2(n_208), .B(n_209), .Y(n_206) );
INVx1_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
INVx2_ASAP7_75t_L g251 ( .A(n_215), .Y(n_251) );
BUFx2_ASAP7_75t_L g348 ( .A(n_215), .Y(n_348) );
AND2x2_ASAP7_75t_L g393 ( .A(n_215), .B(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_221), .B(n_234), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_221), .B(n_330), .Y(n_329) );
AOI21xp5_ASAP7_75t_L g416 ( .A1(n_221), .A2(n_392), .B(n_406), .Y(n_416) );
AND2x2_ASAP7_75t_L g441 ( .A(n_221), .B(n_327), .Y(n_441) );
BUFx2_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVx1_ASAP7_75t_L g363 ( .A(n_223), .Y(n_363) );
AND2x2_ASAP7_75t_L g392 ( .A(n_223), .B(n_393), .Y(n_392) );
INVx2_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
HB1xp67_ASAP7_75t_L g276 ( .A(n_224), .Y(n_276) );
INVx2_ASAP7_75t_L g295 ( .A(n_224), .Y(n_295) );
OR2x2_ASAP7_75t_L g296 ( .A(n_224), .B(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g234 ( .A(n_235), .B(n_236), .Y(n_234) );
INVx2_ASAP7_75t_L g249 ( .A(n_235), .Y(n_249) );
OR2x2_ASAP7_75t_L g262 ( .A(n_235), .B(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g330 ( .A(n_235), .B(n_326), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_235), .B(n_426), .Y(n_425) );
OR2x2_ASAP7_75t_L g431 ( .A(n_235), .B(n_432), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_235), .B(n_368), .Y(n_443) );
AND2x2_ASAP7_75t_L g322 ( .A(n_236), .B(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g345 ( .A(n_236), .B(n_238), .Y(n_345) );
INVx2_ASAP7_75t_L g257 ( .A(n_237), .Y(n_257) );
AND2x2_ASAP7_75t_L g285 ( .A(n_237), .B(n_258), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_237), .B(n_310), .Y(n_366) );
AND2x2_ASAP7_75t_L g280 ( .A(n_238), .B(n_281), .Y(n_280) );
INVx1_ASAP7_75t_L g427 ( .A(n_238), .Y(n_427) );
AND2x2_ASAP7_75t_L g439 ( .A(n_238), .B(n_302), .Y(n_439) );
AND2x2_ASAP7_75t_L g265 ( .A(n_239), .B(n_255), .Y(n_265) );
INVx1_ASAP7_75t_L g360 ( .A(n_239), .Y(n_360) );
AO21x1_ASAP7_75t_L g239 ( .A1(n_240), .A2(n_241), .B(n_244), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g478 ( .A(n_240), .B(n_479), .Y(n_478) );
INVx3_ASAP7_75t_L g495 ( .A(n_240), .Y(n_495) );
AO21x2_ASAP7_75t_L g507 ( .A1(n_240), .A2(n_508), .B(n_515), .Y(n_507) );
AO21x2_ASAP7_75t_L g563 ( .A1(n_240), .A2(n_564), .B(n_571), .Y(n_563) );
NOR2xp33_ASAP7_75t_L g571 ( .A(n_240), .B(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
AND2x4_ASAP7_75t_L g258 ( .A(n_245), .B(n_259), .Y(n_258) );
INVxp67_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_248), .B(n_252), .Y(n_247) );
AND2x2_ASAP7_75t_L g248 ( .A(n_249), .B(n_250), .Y(n_248) );
NOR2xp33_ASAP7_75t_L g305 ( .A(n_249), .B(n_296), .Y(n_305) );
OR2x2_ASAP7_75t_L g437 ( .A(n_249), .B(n_438), .Y(n_437) );
AND2x2_ASAP7_75t_L g354 ( .A(n_250), .B(n_295), .Y(n_354) );
AND2x2_ASAP7_75t_L g362 ( .A(n_250), .B(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_L g421 ( .A(n_250), .B(n_422), .Y(n_421) );
AND2x2_ASAP7_75t_L g445 ( .A(n_250), .B(n_292), .Y(n_445) );
NOR2xp67_ASAP7_75t_L g403 ( .A(n_251), .B(n_404), .Y(n_403) );
OR2x2_ASAP7_75t_L g432 ( .A(n_251), .B(n_295), .Y(n_432) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
NAND2x1p5_ASAP7_75t_L g253 ( .A(n_254), .B(n_256), .Y(n_253) );
AND2x2_ASAP7_75t_L g284 ( .A(n_254), .B(n_285), .Y(n_284) );
INVxp67_ASAP7_75t_L g446 ( .A(n_254), .Y(n_446) );
NOR2x1_ASAP7_75t_L g256 ( .A(n_257), .B(n_258), .Y(n_256) );
INVx1_ASAP7_75t_L g281 ( .A(n_257), .Y(n_281) );
AND2x2_ASAP7_75t_L g332 ( .A(n_257), .B(n_265), .Y(n_332) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_257), .B(n_400), .Y(n_426) );
INVx2_ASAP7_75t_L g271 ( .A(n_258), .Y(n_271) );
INVx3_ASAP7_75t_L g323 ( .A(n_258), .Y(n_323) );
OR2x2_ASAP7_75t_L g351 ( .A(n_258), .B(n_352), .Y(n_351) );
AOI311xp33_ASAP7_75t_L g260 ( .A1(n_261), .A2(n_264), .A3(n_266), .B(n_267), .C(n_278), .Y(n_260) );
O2A1O1Ixp33_ASAP7_75t_L g298 ( .A1(n_261), .A2(n_299), .B(n_301), .C(n_303), .Y(n_298) );
INVx2_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
INVx2_ASAP7_75t_SL g283 ( .A(n_263), .Y(n_283) );
INVx2_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
AND2x2_ASAP7_75t_L g301 ( .A(n_265), .B(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_265), .B(n_281), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_265), .B(n_266), .Y(n_434) );
AND2x2_ASAP7_75t_L g356 ( .A(n_266), .B(n_270), .Y(n_356) );
AOI21xp33_ASAP7_75t_L g267 ( .A1(n_268), .A2(n_272), .B(n_273), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g414 ( .A(n_270), .B(n_302), .Y(n_414) );
INVx2_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
NOR2xp33_ASAP7_75t_L g287 ( .A(n_271), .B(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g308 ( .A(n_271), .Y(n_308) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_277), .Y(n_274) );
AND2x2_ASAP7_75t_L g299 ( .A(n_275), .B(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
INVx1_ASAP7_75t_L g344 ( .A(n_277), .Y(n_344) );
AND2x4_ASAP7_75t_L g406 ( .A(n_277), .B(n_375), .Y(n_406) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AOI222xp33_ASAP7_75t_L g357 ( .A1(n_280), .A2(n_346), .B1(n_358), .B2(n_362), .C1(n_364), .C2(n_368), .Y(n_357) );
A2O1A1Ixp33_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_284), .B(n_286), .C(n_289), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_283), .B(n_327), .Y(n_350) );
INVx1_ASAP7_75t_L g372 ( .A(n_285), .Y(n_372) );
INVx1_ASAP7_75t_L g306 ( .A(n_287), .Y(n_306) );
OR2x2_ASAP7_75t_L g371 ( .A(n_288), .B(n_372), .Y(n_371) );
OAI21xp33_ASAP7_75t_SL g289 ( .A1(n_290), .A2(n_292), .B(n_296), .Y(n_289) );
NAND3xp33_ASAP7_75t_L g307 ( .A(n_290), .B(n_308), .C(n_309), .Y(n_307) );
AOI21xp5_ASAP7_75t_L g405 ( .A1(n_290), .A2(n_327), .B(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx1_ASAP7_75t_SL g292 ( .A(n_293), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_294), .B(n_295), .Y(n_293) );
HB1xp67_ASAP7_75t_L g347 ( .A(n_294), .Y(n_347) );
AND2x2_ASAP7_75t_SL g313 ( .A(n_295), .B(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g404 ( .A(n_295), .Y(n_404) );
HB1xp67_ASAP7_75t_L g420 ( .A(n_295), .Y(n_420) );
INVx2_ASAP7_75t_L g378 ( .A(n_296), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_300), .B(n_321), .Y(n_320) );
INVx2_ASAP7_75t_L g352 ( .A(n_302), .Y(n_352) );
OAI221xp5_ASAP7_75t_L g303 ( .A1(n_304), .A2(n_306), .B1(n_307), .B2(n_311), .C(n_312), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_SL g385 ( .A(n_306), .B(n_386), .Y(n_385) );
INVx1_ASAP7_75t_SL g440 ( .A(n_306), .Y(n_440) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx2_ASAP7_75t_L g321 ( .A(n_313), .Y(n_321) );
NOR2xp33_ASAP7_75t_L g343 ( .A(n_313), .B(n_344), .Y(n_343) );
AND2x2_ASAP7_75t_L g379 ( .A(n_313), .B(n_327), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_313), .B(n_389), .Y(n_388) );
AND2x2_ASAP7_75t_L g412 ( .A(n_313), .B(n_347), .Y(n_412) );
BUFx3_ASAP7_75t_L g375 ( .A(n_314), .Y(n_375) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
NAND5xp2_ASAP7_75t_L g317 ( .A(n_318), .B(n_336), .C(n_357), .D(n_369), .E(n_384), .Y(n_317) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
AOI32xp33_ASAP7_75t_L g409 ( .A1(n_321), .A2(n_348), .A3(n_364), .B1(n_410), .B2(n_412), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_323), .B(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_L g324 ( .A(n_325), .B(n_327), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx1_ASAP7_75t_SL g333 ( .A(n_327), .Y(n_333) );
OAI22xp5_ASAP7_75t_L g328 ( .A1(n_329), .A2(n_331), .B1(n_333), .B2(n_334), .Y(n_328) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx1_ASAP7_75t_SL g334 ( .A(n_335), .Y(n_334) );
AOI221xp5_ASAP7_75t_L g336 ( .A1(n_337), .A2(n_343), .B1(n_345), .B2(n_346), .C(n_349), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
OR2x2_ASAP7_75t_L g338 ( .A(n_339), .B(n_341), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g408 ( .A(n_340), .B(n_359), .Y(n_408) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
AOI221xp5_ASAP7_75t_L g423 ( .A1(n_345), .A2(n_406), .B1(n_424), .B2(n_429), .C(n_430), .Y(n_423) );
AND2x2_ASAP7_75t_L g346 ( .A(n_347), .B(n_348), .Y(n_346) );
INVx2_ASAP7_75t_L g389 ( .A(n_348), .Y(n_389) );
OAI22xp5_ASAP7_75t_L g349 ( .A1(n_350), .A2(n_351), .B1(n_353), .B2(n_355), .Y(n_349) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx1_ASAP7_75t_SL g355 ( .A(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g358 ( .A(n_359), .B(n_361), .Y(n_358) );
INVx1_ASAP7_75t_L g367 ( .A(n_359), .Y(n_367) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
OR2x2_ASAP7_75t_L g365 ( .A(n_366), .B(n_367), .Y(n_365) );
AOI222xp33_ASAP7_75t_L g369 ( .A1(n_370), .A2(n_373), .B1(n_377), .B2(n_378), .C1(n_379), .C2(n_380), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g373 ( .A(n_374), .B(n_376), .Y(n_373) );
INVxp67_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
OAI22xp33_ASAP7_75t_L g424 ( .A1(n_378), .A2(n_425), .B1(n_427), .B2(n_428), .Y(n_424) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_SL g382 ( .A(n_383), .Y(n_382) );
AOI21xp5_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_387), .B(n_390), .Y(n_384) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
AOI21xp33_ASAP7_75t_L g390 ( .A1(n_391), .A2(n_395), .B(n_397), .Y(n_390) );
INVx2_ASAP7_75t_SL g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g438 ( .A(n_393), .Y(n_438) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_SL g399 ( .A(n_400), .Y(n_399) );
A2O1A1Ixp33_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_405), .B(n_407), .C(n_409), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
AOI211xp5_ASAP7_75t_L g413 ( .A1(n_414), .A2(n_415), .B(n_417), .C(n_442), .Y(n_413) );
CKINVDCx16_ASAP7_75t_R g418 ( .A(n_414), .Y(n_418) );
INVxp67_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
OAI211xp5_ASAP7_75t_L g417 ( .A1(n_418), .A2(n_419), .B(n_423), .C(n_435), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_420), .B(n_421), .Y(n_419) );
AOI21xp33_ASAP7_75t_L g430 ( .A1(n_431), .A2(n_433), .B(n_434), .Y(n_430) );
AOI22xp5_ASAP7_75t_L g435 ( .A1(n_436), .A2(n_439), .B1(n_440), .B2(n_441), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
AOI21xp33_ASAP7_75t_L g442 ( .A1(n_443), .A2(n_444), .B(n_446), .Y(n_442) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx2_ASAP7_75t_L g743 ( .A(n_455), .Y(n_743) );
OR3x2_ASAP7_75t_L g455 ( .A(n_456), .B(n_655), .C(n_698), .Y(n_455) );
NAND5xp2_ASAP7_75t_L g456 ( .A(n_457), .B(n_582), .C(n_612), .D(n_629), .E(n_644), .Y(n_456) );
AOI221xp5_ASAP7_75t_SL g457 ( .A1(n_458), .A2(n_505), .B1(n_545), .B2(n_551), .C(n_555), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_459), .B(n_480), .Y(n_458) );
OR2x2_ASAP7_75t_L g560 ( .A(n_459), .B(n_561), .Y(n_560) );
AND2x2_ASAP7_75t_L g599 ( .A(n_459), .B(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g617 ( .A(n_459), .B(n_618), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_459), .B(n_553), .Y(n_634) );
OR2x2_ASAP7_75t_L g646 ( .A(n_459), .B(n_647), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_459), .B(n_605), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_459), .B(n_679), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_459), .B(n_583), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_459), .B(n_591), .Y(n_697) );
AND2x2_ASAP7_75t_L g729 ( .A(n_459), .B(n_493), .Y(n_729) );
HB1xp67_ASAP7_75t_L g737 ( .A(n_459), .Y(n_737) );
INVx5_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_460), .B(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g557 ( .A(n_460), .B(n_535), .Y(n_557) );
BUFx2_ASAP7_75t_L g579 ( .A(n_460), .Y(n_579) );
AND2x2_ASAP7_75t_L g608 ( .A(n_460), .B(n_481), .Y(n_608) );
AND2x2_ASAP7_75t_L g663 ( .A(n_460), .B(n_561), .Y(n_663) );
OR2x6_ASAP7_75t_L g460 ( .A(n_461), .B(n_478), .Y(n_460) );
BUFx2_ASAP7_75t_L g484 ( .A(n_463), .Y(n_484) );
INVx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
O2A1O1Ixp33_ASAP7_75t_SL g497 ( .A1(n_467), .A2(n_477), .B(n_498), .C(n_499), .Y(n_497) );
O2A1O1Ixp33_ASAP7_75t_L g539 ( .A1(n_467), .A2(n_477), .B(n_540), .C(n_541), .Y(n_539) );
INVx5_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
O2A1O1Ixp33_ASAP7_75t_L g470 ( .A1(n_471), .A2(n_472), .B(n_474), .C(n_475), .Y(n_470) );
O2A1O1Ixp33_ASAP7_75t_L g531 ( .A1(n_472), .A2(n_475), .B(n_532), .C(n_533), .Y(n_531) );
INVx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_480), .B(n_617), .Y(n_626) );
OAI32xp33_ASAP7_75t_L g640 ( .A1(n_480), .A2(n_576), .A3(n_641), .B1(n_642), .B2(n_643), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_480), .B(n_642), .Y(n_672) );
NOR2xp33_ASAP7_75t_L g683 ( .A(n_480), .B(n_560), .Y(n_683) );
INVx1_ASAP7_75t_SL g712 ( .A(n_480), .Y(n_712) );
NAND4xp25_ASAP7_75t_L g721 ( .A(n_480), .B(n_507), .C(n_663), .D(n_722), .Y(n_721) );
AND2x4_ASAP7_75t_L g480 ( .A(n_481), .B(n_493), .Y(n_480) );
INVx5_ASAP7_75t_L g554 ( .A(n_481), .Y(n_554) );
AND2x2_ASAP7_75t_L g583 ( .A(n_481), .B(n_494), .Y(n_583) );
HB1xp67_ASAP7_75t_L g662 ( .A(n_481), .Y(n_662) );
AND2x2_ASAP7_75t_L g732 ( .A(n_481), .B(n_679), .Y(n_732) );
OR2x6_ASAP7_75t_L g481 ( .A(n_482), .B(n_490), .Y(n_481) );
AOI21xp5_ASAP7_75t_SL g482 ( .A1(n_483), .A2(n_485), .B(n_489), .Y(n_482) );
NOR2xp33_ASAP7_75t_L g490 ( .A(n_491), .B(n_492), .Y(n_490) );
AND2x4_ASAP7_75t_L g605 ( .A(n_493), .B(n_554), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_493), .B(n_615), .Y(n_614) );
AND2x2_ASAP7_75t_L g639 ( .A(n_493), .B(n_561), .Y(n_639) );
INVx2_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
AND2x2_ASAP7_75t_L g553 ( .A(n_494), .B(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g591 ( .A(n_494), .B(n_563), .Y(n_591) );
AND2x2_ASAP7_75t_L g600 ( .A(n_494), .B(n_562), .Y(n_600) );
OA21x2_ASAP7_75t_L g494 ( .A1(n_495), .A2(n_496), .B(n_504), .Y(n_494) );
NOR2xp33_ASAP7_75t_L g500 ( .A(n_501), .B(n_502), .Y(n_500) );
AOI222xp33_ASAP7_75t_L g668 ( .A1(n_505), .A2(n_669), .B1(n_671), .B2(n_673), .C1(n_676), .C2(n_677), .Y(n_668) );
AND2x4_ASAP7_75t_L g505 ( .A(n_506), .B(n_524), .Y(n_505) );
AND2x2_ASAP7_75t_L g601 ( .A(n_506), .B(n_602), .Y(n_601) );
NAND3xp33_ASAP7_75t_L g718 ( .A(n_506), .B(n_579), .C(n_719), .Y(n_718) );
AND2x2_ASAP7_75t_L g506 ( .A(n_507), .B(n_517), .Y(n_506) );
INVx5_ASAP7_75t_SL g550 ( .A(n_507), .Y(n_550) );
OAI322xp33_ASAP7_75t_L g555 ( .A1(n_507), .A2(n_556), .A3(n_558), .B1(n_559), .B2(n_573), .C1(n_576), .C2(n_578), .Y(n_555) );
NAND2xp5_ASAP7_75t_SL g621 ( .A(n_507), .B(n_548), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_507), .B(n_536), .Y(n_727) );
OAI21xp5_ASAP7_75t_L g508 ( .A1(n_509), .A2(n_510), .B(n_511), .Y(n_508) );
INVx2_ASAP7_75t_L g548 ( .A(n_517), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_517), .B(n_526), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_524), .B(n_586), .Y(n_641) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
OR2x2_ASAP7_75t_L g620 ( .A(n_525), .B(n_621), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_526), .B(n_535), .Y(n_525) );
OR2x2_ASAP7_75t_L g549 ( .A(n_526), .B(n_550), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_526), .B(n_557), .Y(n_556) );
OR2x2_ASAP7_75t_L g588 ( .A(n_526), .B(n_536), .Y(n_588) );
AND2x2_ASAP7_75t_L g611 ( .A(n_526), .B(n_548), .Y(n_611) );
NOR2xp33_ASAP7_75t_L g622 ( .A(n_526), .B(n_623), .Y(n_622) );
AND2x2_ASAP7_75t_L g627 ( .A(n_526), .B(n_586), .Y(n_627) );
AND2x2_ASAP7_75t_L g635 ( .A(n_526), .B(n_636), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_526), .B(n_595), .Y(n_685) );
INVx5_ASAP7_75t_SL g526 ( .A(n_527), .Y(n_526) );
AND2x2_ASAP7_75t_L g575 ( .A(n_527), .B(n_550), .Y(n_575) );
OR2x2_ASAP7_75t_L g576 ( .A(n_527), .B(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g602 ( .A(n_527), .B(n_536), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_527), .B(n_649), .Y(n_690) );
OR2x2_ASAP7_75t_L g706 ( .A(n_527), .B(n_650), .Y(n_706) );
AND2x2_ASAP7_75t_SL g713 ( .A(n_527), .B(n_667), .Y(n_713) );
HB1xp67_ASAP7_75t_L g720 ( .A(n_527), .Y(n_720) );
OR2x6_ASAP7_75t_L g527 ( .A(n_528), .B(n_534), .Y(n_527) );
AND2x2_ASAP7_75t_L g574 ( .A(n_535), .B(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g624 ( .A(n_535), .B(n_548), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_535), .B(n_550), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_535), .B(n_586), .Y(n_708) );
INVx3_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_536), .B(n_550), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_536), .B(n_548), .Y(n_596) );
OR2x2_ASAP7_75t_L g650 ( .A(n_536), .B(n_548), .Y(n_650) );
AND2x2_ASAP7_75t_L g667 ( .A(n_536), .B(n_547), .Y(n_667) );
INVxp67_ASAP7_75t_L g689 ( .A(n_536), .Y(n_689) );
AND2x2_ASAP7_75t_L g716 ( .A(n_536), .B(n_586), .Y(n_716) );
HB1xp67_ASAP7_75t_L g723 ( .A(n_536), .Y(n_723) );
OA21x2_ASAP7_75t_L g536 ( .A1(n_537), .A2(n_538), .B(n_544), .Y(n_536) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
OR2x2_ASAP7_75t_L g546 ( .A(n_547), .B(n_549), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_547), .B(n_597), .Y(n_670) );
INVx1_ASAP7_75t_SL g547 ( .A(n_548), .Y(n_547) );
AND2x2_ASAP7_75t_L g586 ( .A(n_548), .B(n_550), .Y(n_586) );
OR2x2_ASAP7_75t_L g653 ( .A(n_548), .B(n_654), .Y(n_653) );
INVx2_ASAP7_75t_L g597 ( .A(n_549), .Y(n_597) );
OR2x2_ASAP7_75t_L g658 ( .A(n_549), .B(n_650), .Y(n_658) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx1_ASAP7_75t_L g558 ( .A(n_553), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_553), .B(n_617), .Y(n_616) );
OR2x2_ASAP7_75t_L g559 ( .A(n_554), .B(n_560), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_554), .B(n_581), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_554), .B(n_561), .Y(n_593) );
INVx2_ASAP7_75t_L g638 ( .A(n_554), .Y(n_638) );
AND2x2_ASAP7_75t_L g651 ( .A(n_554), .B(n_591), .Y(n_651) );
AND2x2_ASAP7_75t_L g676 ( .A(n_554), .B(n_600), .Y(n_676) );
INVx1_ASAP7_75t_L g628 ( .A(n_559), .Y(n_628) );
INVx2_ASAP7_75t_SL g615 ( .A(n_560), .Y(n_615) );
INVx1_ASAP7_75t_L g618 ( .A(n_561), .Y(n_618) );
INVx2_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
HB1xp67_ASAP7_75t_L g581 ( .A(n_562), .Y(n_581) );
INVx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
BUFx2_ASAP7_75t_L g679 ( .A(n_563), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_565), .B(n_570), .Y(n_564) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g648 ( .A(n_575), .B(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g654 ( .A(n_575), .Y(n_654) );
AOI22xp5_ASAP7_75t_L g656 ( .A1(n_575), .A2(n_657), .B1(n_659), .B2(n_664), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_575), .B(n_667), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_576), .B(n_670), .Y(n_669) );
INVx1_ASAP7_75t_SL g610 ( .A(n_577), .Y(n_610) );
OR2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_580), .Y(n_578) );
OR2x2_ASAP7_75t_L g592 ( .A(n_579), .B(n_593), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_579), .B(n_583), .Y(n_643) );
AND2x2_ASAP7_75t_L g666 ( .A(n_579), .B(n_667), .Y(n_666) );
BUFx2_ASAP7_75t_L g642 ( .A(n_581), .Y(n_642) );
AOI211xp5_ASAP7_75t_L g582 ( .A1(n_583), .A2(n_584), .B(n_589), .C(n_603), .Y(n_582) );
INVx1_ASAP7_75t_L g606 ( .A(n_583), .Y(n_606) );
OAI221xp5_ASAP7_75t_SL g714 ( .A1(n_583), .A2(n_715), .B1(n_717), .B2(n_718), .C(n_721), .Y(n_714) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_586), .B(n_587), .Y(n_585) );
INVx1_ASAP7_75t_L g733 ( .A(n_586), .Y(n_733) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
OR2x2_ASAP7_75t_L g682 ( .A(n_588), .B(n_621), .Y(n_682) );
A2O1A1Ixp33_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_592), .B(n_594), .C(n_598), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_595), .B(n_597), .Y(n_594) );
INVx1_ASAP7_75t_SL g595 ( .A(n_596), .Y(n_595) );
OAI32xp33_ASAP7_75t_L g707 ( .A1(n_596), .A2(n_597), .A3(n_660), .B1(n_697), .B2(n_708), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_599), .B(n_601), .Y(n_598) );
AND2x2_ASAP7_75t_L g739 ( .A(n_599), .B(n_638), .Y(n_739) );
AND2x2_ASAP7_75t_L g686 ( .A(n_600), .B(n_638), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_600), .B(n_608), .Y(n_704) );
AOI31xp33_ASAP7_75t_SL g603 ( .A1(n_604), .A2(n_606), .A3(n_607), .B(n_609), .Y(n_603) );
INVxp67_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_605), .B(n_617), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_605), .B(n_615), .Y(n_702) );
AOI221xp5_ASAP7_75t_L g724 ( .A1(n_605), .A2(n_635), .B1(n_725), .B2(n_728), .C(n_730), .Y(n_724) );
CKINVDCx16_ASAP7_75t_R g607 ( .A(n_608), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_610), .B(n_611), .Y(n_609) );
AND2x2_ASAP7_75t_L g630 ( .A(n_610), .B(n_631), .Y(n_630) );
AOI222xp33_ASAP7_75t_L g612 ( .A1(n_613), .A2(n_619), .B1(n_622), .B2(n_625), .C1(n_627), .C2(n_628), .Y(n_612) );
NAND2xp5_ASAP7_75t_SL g613 ( .A(n_614), .B(n_616), .Y(n_613) );
INVx1_ASAP7_75t_L g695 ( .A(n_614), .Y(n_695) );
INVx1_ASAP7_75t_L g717 ( .A(n_617), .Y(n_717) );
INVx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
OAI22xp5_ASAP7_75t_L g730 ( .A1(n_620), .A2(n_731), .B1(n_733), .B2(n_734), .Y(n_730) );
INVx1_ASAP7_75t_L g636 ( .A(n_621), .Y(n_636) );
INVx1_ASAP7_75t_SL g623 ( .A(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
AOI221xp5_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_633), .B1(n_635), .B2(n_637), .C(n_640), .Y(n_629) );
INVx1_ASAP7_75t_SL g631 ( .A(n_632), .Y(n_631) );
OR2x2_ASAP7_75t_L g674 ( .A(n_632), .B(n_675), .Y(n_674) );
OR2x2_ASAP7_75t_L g726 ( .A(n_632), .B(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g701 ( .A(n_637), .Y(n_701) );
AND2x2_ASAP7_75t_L g637 ( .A(n_638), .B(n_639), .Y(n_637) );
INVx1_ASAP7_75t_L g665 ( .A(n_638), .Y(n_665) );
INVx1_ASAP7_75t_L g647 ( .A(n_639), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_642), .B(n_729), .Y(n_734) );
AOI22xp33_ASAP7_75t_L g644 ( .A1(n_645), .A2(n_648), .B1(n_651), .B2(n_652), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx1_ASAP7_75t_SL g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_SL g738 ( .A(n_651), .Y(n_738) );
INVxp33_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
NOR2xp33_ASAP7_75t_L g696 ( .A(n_653), .B(n_697), .Y(n_696) );
OAI32xp33_ASAP7_75t_L g687 ( .A1(n_654), .A2(n_688), .A3(n_689), .B1(n_690), .B2(n_691), .Y(n_687) );
NAND4xp25_ASAP7_75t_L g655 ( .A(n_656), .B(n_668), .C(n_680), .D(n_692), .Y(n_655) );
INVx1_ASAP7_75t_SL g657 ( .A(n_658), .Y(n_657) );
NAND2xp33_ASAP7_75t_SL g659 ( .A(n_660), .B(n_661), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_662), .B(n_663), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_663), .B(n_712), .Y(n_711) );
AND2x2_ASAP7_75t_L g664 ( .A(n_665), .B(n_666), .Y(n_664) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
CKINVDCx16_ASAP7_75t_R g673 ( .A(n_674), .Y(n_673) );
AOI221xp5_ASAP7_75t_L g709 ( .A1(n_677), .A2(n_693), .B1(n_710), .B2(n_713), .C(n_714), .Y(n_709) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
AND2x2_ASAP7_75t_L g728 ( .A(n_679), .B(n_729), .Y(n_728) );
AOI221xp5_ASAP7_75t_L g680 ( .A1(n_681), .A2(n_683), .B1(n_684), .B2(n_686), .C(n_687), .Y(n_680) );
INVx1_ASAP7_75t_SL g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
NOR2xp33_ASAP7_75t_L g719 ( .A(n_689), .B(n_720), .Y(n_719) );
AOI21xp5_ASAP7_75t_L g692 ( .A1(n_693), .A2(n_695), .B(n_696), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
NAND4xp25_ASAP7_75t_L g698 ( .A(n_699), .B(n_709), .C(n_724), .D(n_735), .Y(n_698) );
O2A1O1Ixp33_ASAP7_75t_L g699 ( .A1(n_700), .A2(n_703), .B(n_705), .C(n_707), .Y(n_699) );
NAND2xp5_ASAP7_75t_SL g700 ( .A(n_701), .B(n_702), .Y(n_700) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVxp67_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_SL g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g740 ( .A(n_727), .Y(n_740) );
INVx2_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
OAI21xp5_ASAP7_75t_L g735 ( .A1(n_736), .A2(n_739), .B(n_740), .Y(n_735) );
NOR2xp33_ASAP7_75t_L g736 ( .A(n_737), .B(n_738), .Y(n_736) );
INVx1_ASAP7_75t_SL g744 ( .A(n_745), .Y(n_744) );
INVx2_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx2_ASAP7_75t_SL g747 ( .A(n_748), .Y(n_747) );
CKINVDCx20_ASAP7_75t_R g751 ( .A(n_752), .Y(n_751) );
INVx1_ASAP7_75t_SL g754 ( .A(n_755), .Y(n_754) );
endmodule