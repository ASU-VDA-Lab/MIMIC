module fake_jpeg_8016_n_143 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_143);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_143;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx8_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_2),
.B(n_5),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_6),
.B(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_1),
.B(n_12),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_34),
.Y(n_43)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_20),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_20),
.B(n_1),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_36),
.Y(n_44)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

BUFx2_ASAP7_75t_SL g38 ( 
.A(n_16),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_40),
.B(n_52),
.Y(n_72)
);

BUFx16f_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

INVxp33_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_51),
.A2(n_33),
.B1(n_32),
.B2(n_22),
.Y(n_66)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_34),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_55),
.B(n_68),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_48),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_56),
.B(n_57),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_48),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_58),
.B(n_59),
.Y(n_79)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_50),
.B(n_36),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_60),
.B(n_64),
.Y(n_82)
);

AND2x6_ASAP7_75t_L g61 ( 
.A(n_49),
.B(n_3),
.Y(n_61)
);

AOI21xp33_ASAP7_75t_L g77 ( 
.A1(n_61),
.A2(n_63),
.B(n_67),
.Y(n_77)
);

AND2x6_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_3),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_35),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_51),
.A2(n_21),
.B1(n_14),
.B2(n_25),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_65),
.A2(n_70),
.B1(n_71),
.B2(n_24),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g74 ( 
.A(n_66),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_53),
.B(n_22),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_53),
.A2(n_25),
.B(n_14),
.Y(n_68)
);

OA22x2_ASAP7_75t_SL g70 ( 
.A1(n_47),
.A2(n_19),
.B1(n_16),
.B2(n_28),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_41),
.A2(n_15),
.B1(n_17),
.B2(n_29),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_55),
.B(n_29),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_76),
.Y(n_90)
);

INVx13_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_88),
.Y(n_96)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_72),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_46),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_84),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_83),
.A2(n_70),
.B1(n_41),
.B2(n_63),
.Y(n_92)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_59),
.B(n_24),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_85),
.B(n_86),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_68),
.B(n_15),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_3),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_62),
.B(n_17),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_SL g89 ( 
.A(n_81),
.B(n_67),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_SL g103 ( 
.A(n_89),
.B(n_91),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_92),
.B(n_99),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_70),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_93),
.B(n_83),
.C(n_82),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_77),
.A2(n_61),
.B1(n_40),
.B2(n_45),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_94),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_84),
.A2(n_45),
.B1(n_69),
.B2(n_54),
.Y(n_95)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_95),
.Y(n_106)
);

OAI22x1_ASAP7_75t_L g97 ( 
.A1(n_74),
.A2(n_27),
.B1(n_28),
.B2(n_18),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_97),
.A2(n_98),
.B(n_88),
.Y(n_104)
);

A2O1A1Ixp33_ASAP7_75t_SL g98 ( 
.A1(n_87),
.A2(n_58),
.B(n_27),
.C(n_28),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_78),
.A2(n_54),
.B1(n_26),
.B2(n_28),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_80),
.B(n_8),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_100),
.B(n_102),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_103),
.B(n_108),
.C(n_111),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_104),
.A2(n_105),
.B(n_113),
.Y(n_115)
);

NOR4xp25_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_82),
.C(n_86),
.D(n_79),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_96),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_107),
.B(n_85),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_73),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_94),
.A2(n_79),
.B(n_76),
.Y(n_113)
);

A2O1A1Ixp33_ASAP7_75t_L g114 ( 
.A1(n_112),
.A2(n_92),
.B(n_108),
.C(n_110),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_114),
.B(n_118),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_109),
.B(n_101),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_116),
.Y(n_125)
);

INVxp33_ASAP7_75t_L g118 ( 
.A(n_106),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_103),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_119),
.B(n_120),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_112),
.A2(n_98),
.B(n_93),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_121),
.A2(n_97),
.B1(n_98),
.B2(n_75),
.Y(n_123)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_123),
.Y(n_130)
);

HB1xp67_ASAP7_75t_L g126 ( 
.A(n_118),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_126),
.B(n_4),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_117),
.B(n_111),
.C(n_98),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_127),
.B(n_121),
.C(n_75),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_125),
.B(n_115),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_128),
.B(n_131),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_129),
.B(n_127),
.C(n_123),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_122),
.A2(n_4),
.B(n_6),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_132),
.A2(n_124),
.B1(n_9),
.B2(n_11),
.Y(n_133)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_133),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_135),
.B(n_136),
.C(n_18),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_129),
.B(n_130),
.Y(n_136)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_137),
.Y(n_140)
);

O2A1O1Ixp33_ASAP7_75t_L g138 ( 
.A1(n_134),
.A2(n_7),
.B(n_13),
.C(n_18),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_138),
.A2(n_7),
.B(n_18),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_141),
.A2(n_139),
.B(n_136),
.Y(n_142)
);

HAxp5_ASAP7_75t_SL g143 ( 
.A(n_142),
.B(n_140),
.CON(n_143),
.SN(n_143)
);


endmodule