module fake_jpeg_4528_n_89 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_89);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_89;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

BUFx4f_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

INVx6_ASAP7_75t_SL g12 ( 
.A(n_7),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

INVx6_ASAP7_75t_SL g19 ( 
.A(n_12),
.Y(n_19)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_21),
.B(n_23),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_SL g23 ( 
.A1(n_18),
.A2(n_2),
.B(n_3),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_24),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_21),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_26),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_19),
.B(n_13),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_13),
.Y(n_36)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_32),
.B(n_15),
.Y(n_35)
);

OAI22xp33_ASAP7_75t_L g33 ( 
.A1(n_27),
.A2(n_22),
.B1(n_20),
.B2(n_10),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_33),
.A2(n_29),
.B1(n_28),
.B2(n_32),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_35),
.B(n_36),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_15),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_39),
.Y(n_41)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_31),
.B(n_17),
.Y(n_40)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_31),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_16),
.Y(n_56)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_33),
.Y(n_45)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_46),
.Y(n_50)
);

O2A1O1Ixp33_ASAP7_75t_L g48 ( 
.A1(n_34),
.A2(n_29),
.B(n_28),
.C(n_16),
.Y(n_48)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

BUFx24_ASAP7_75t_SL g52 ( 
.A(n_47),
.Y(n_52)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_29),
.C(n_28),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_54),
.B(n_55),
.Y(n_64)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_56),
.B(n_57),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_25),
.C(n_15),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_58),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_59),
.B(n_61),
.Y(n_68)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_50),
.A2(n_45),
.B1(n_44),
.B2(n_46),
.Y(n_62)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

NAND3xp33_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_44),
.C(n_45),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_63),
.A2(n_14),
.B(n_11),
.Y(n_72)
);

AO221x1_ASAP7_75t_L g65 ( 
.A1(n_58),
.A2(n_43),
.B1(n_49),
.B2(n_48),
.C(n_14),
.Y(n_65)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_64),
.B(n_51),
.Y(n_70)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_66),
.B(n_62),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_71),
.B(n_73),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_72),
.A2(n_14),
.B(n_11),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_49),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_67),
.A2(n_69),
.B1(n_73),
.B2(n_71),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_74),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_68),
.B(n_60),
.Y(n_76)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_76),
.Y(n_82)
);

AOI31xp67_ASAP7_75t_SL g79 ( 
.A1(n_78),
.A2(n_11),
.A3(n_1),
.B(n_0),
.Y(n_79)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_79),
.Y(n_83)
);

NAND3xp33_ASAP7_75t_L g84 ( 
.A(n_80),
.B(n_8),
.C(n_9),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_75),
.B(n_5),
.Y(n_81)
);

BUFx24_ASAP7_75t_SL g85 ( 
.A(n_81),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_84),
.B(n_8),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_83),
.A2(n_77),
.B1(n_82),
.B2(n_1),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_86),
.A2(n_87),
.B(n_85),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_88),
.B(n_1),
.Y(n_89)
);


endmodule