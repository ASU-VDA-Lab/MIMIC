module fake_jpeg_3373_n_126 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_126);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_126;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g33 ( 
.A(n_32),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_21),
.B(n_6),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_27),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_30),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_23),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

BUFx4f_ASAP7_75t_SL g44 ( 
.A(n_33),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_44),
.Y(n_56)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_34),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_43),
.Y(n_53)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_50),
.B(n_41),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_44),
.B(n_34),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_43),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_53),
.B(n_54),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_41),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_55),
.B(n_38),
.Y(n_62)
);

NOR2x1_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_33),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_59),
.B(n_38),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_61),
.B(n_65),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_62),
.B(n_67),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_52),
.B(n_46),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_64),
.B(n_70),
.Y(n_73)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_56),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_56),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_68),
.B(n_69),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_59),
.B(n_39),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_57),
.A2(n_56),
.B(n_51),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_39),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_71),
.B(n_42),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_64),
.A2(n_58),
.B1(n_45),
.B2(n_51),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_72),
.A2(n_81),
.B1(n_19),
.B2(n_18),
.Y(n_92)
);

AO22x2_ASAP7_75t_L g75 ( 
.A1(n_70),
.A2(n_60),
.B1(n_48),
.B2(n_42),
.Y(n_75)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_75),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_80),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_35),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_65),
.A2(n_60),
.B1(n_43),
.B2(n_40),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_62),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_82),
.B(n_83),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_36),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_73),
.A2(n_36),
.B1(n_31),
.B2(n_28),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_84),
.A2(n_88),
.B1(n_15),
.B2(n_2),
.Y(n_98)
);

NOR2xp67_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_0),
.Y(n_85)
);

NAND3xp33_ASAP7_75t_L g99 ( 
.A(n_85),
.B(n_0),
.C(n_2),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_75),
.A2(n_26),
.B1(n_25),
.B2(n_24),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_22),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_89),
.B(n_91),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_72),
.B(n_20),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_93),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_79),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_75),
.B(n_16),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_94),
.B(n_8),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_75),
.A2(n_78),
.B(n_1),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_95),
.A2(n_78),
.B(n_1),
.Y(n_97)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_90),
.Y(n_96)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_96),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_97),
.A2(n_100),
.B1(n_103),
.B2(n_84),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_98),
.B(n_99),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_87),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_100)
);

CKINVDCx12_ASAP7_75t_R g101 ( 
.A(n_86),
.Y(n_101)
);

BUFx12_ASAP7_75t_L g111 ( 
.A(n_101),
.Y(n_111)
);

A2O1A1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_94),
.A2(n_3),
.B(n_4),
.C(n_5),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_102),
.B(n_91),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_88),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_106),
.B(n_89),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_107),
.B(n_112),
.Y(n_116)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_104),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_110),
.B(n_100),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_113),
.B(n_9),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_114),
.A2(n_115),
.B1(n_108),
.B2(n_116),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_109),
.A2(n_105),
.B1(n_99),
.B2(n_102),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_117),
.A2(n_113),
.B(n_111),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_118),
.B(n_119),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_116),
.B(n_10),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_120),
.B(n_111),
.Y(n_122)
);

AOI321xp33_ASAP7_75t_L g123 ( 
.A1(n_122),
.A2(n_11),
.A3(n_12),
.B1(n_13),
.B2(n_14),
.C(n_121),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_123),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_122),
.C(n_13),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_125),
.B(n_11),
.Y(n_126)
);


endmodule