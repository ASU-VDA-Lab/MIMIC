module fake_jpeg_2659_n_527 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_527);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_527;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx2_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_17),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_16),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx2_ASAP7_75t_SL g39 ( 
.A(n_11),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_0),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_14),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_8),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_18),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

BUFx12_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

BUFx4f_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_9),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_8),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_10),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_2),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_6),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g153 ( 
.A(n_57),
.Y(n_153)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_58),
.Y(n_131)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_59),
.Y(n_129)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_60),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_23),
.B(n_7),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_61),
.B(n_67),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g192 ( 
.A(n_62),
.Y(n_192)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g178 ( 
.A(n_63),
.Y(n_178)
);

BUFx12_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g140 ( 
.A(n_64),
.Y(n_140)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_65),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_31),
.B(n_0),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_66),
.B(n_71),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_23),
.B(n_7),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_31),
.B(n_36),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_68),
.B(n_103),
.Y(n_172)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_69),
.Y(n_201)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_70),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_36),
.B(n_0),
.Y(n_71)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_72),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_73),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_74),
.Y(n_144)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_32),
.Y(n_75)
);

INVx11_ASAP7_75t_L g150 ( 
.A(n_75),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_24),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_76),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_24),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_77),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_78),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_39),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_79),
.B(n_117),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_41),
.Y(n_80)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_80),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_51),
.B(n_21),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_81),
.B(n_104),
.Y(n_162)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

INVx5_ASAP7_75t_L g197 ( 
.A(n_82),
.Y(n_197)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_19),
.Y(n_83)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_83),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_41),
.Y(n_84)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_84),
.Y(n_147)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

INVx8_ASAP7_75t_L g170 ( 
.A(n_85),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

INVx6_ASAP7_75t_L g188 ( 
.A(n_86),
.Y(n_188)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_87),
.Y(n_135)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_21),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g205 ( 
.A(n_88),
.Y(n_205)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_32),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g155 ( 
.A(n_89),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_32),
.Y(n_90)
);

INVx8_ASAP7_75t_L g204 ( 
.A(n_90),
.Y(n_204)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_26),
.Y(n_91)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_91),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_28),
.B(n_10),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_92),
.B(n_95),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_35),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_93),
.Y(n_196)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_35),
.Y(n_94)
);

INVx11_ASAP7_75t_L g171 ( 
.A(n_94),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_28),
.B(n_10),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_27),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_96),
.B(n_99),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_35),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g199 ( 
.A(n_97),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_35),
.Y(n_98)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_98),
.Y(n_191)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_19),
.B(n_11),
.Y(n_99)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_27),
.Y(n_100)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_100),
.Y(n_137)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_56),
.Y(n_101)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_101),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_33),
.Y(n_102)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_102),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_42),
.B(n_5),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_42),
.B(n_5),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_51),
.B(n_1),
.Y(n_105)
);

AND2x2_ASAP7_75t_SL g200 ( 
.A(n_105),
.B(n_1),
.Y(n_200)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_25),
.Y(n_106)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_106),
.Y(n_143)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_33),
.Y(n_107)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_107),
.Y(n_182)
);

BUFx12f_ASAP7_75t_L g108 ( 
.A(n_44),
.Y(n_108)
);

INVx11_ASAP7_75t_L g179 ( 
.A(n_108),
.Y(n_179)
);

BUFx5_ASAP7_75t_L g109 ( 
.A(n_30),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g149 ( 
.A(n_109),
.Y(n_149)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_44),
.Y(n_110)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_110),
.Y(n_206)
);

BUFx12f_ASAP7_75t_L g111 ( 
.A(n_56),
.Y(n_111)
);

BUFx24_ASAP7_75t_L g202 ( 
.A(n_111),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_21),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_112),
.B(n_119),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_46),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_113),
.Y(n_151)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_25),
.Y(n_114)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_114),
.Y(n_146)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_46),
.Y(n_115)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_115),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_34),
.Y(n_116)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_116),
.Y(n_165)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_30),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g118 ( 
.A(n_30),
.Y(n_118)
);

BUFx5_ASAP7_75t_L g163 ( 
.A(n_118),
.Y(n_163)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_34),
.B(n_12),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_43),
.B(n_12),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_120),
.B(n_121),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_43),
.Y(n_121)
);

INVx2_ASAP7_75t_SL g122 ( 
.A(n_37),
.Y(n_122)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_122),
.Y(n_166)
);

BUFx12f_ASAP7_75t_L g123 ( 
.A(n_20),
.Y(n_123)
);

BUFx12_ASAP7_75t_L g133 ( 
.A(n_123),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_108),
.A2(n_53),
.B1(n_52),
.B2(n_47),
.Y(n_128)
);

OA22x2_ASAP7_75t_L g251 ( 
.A1(n_128),
.A2(n_152),
.B1(n_161),
.B2(n_187),
.Y(n_251)
);

OAI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_73),
.A2(n_74),
.B1(n_80),
.B2(n_78),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_130),
.A2(n_189),
.B1(n_151),
.B2(n_175),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_66),
.A2(n_53),
.B1(n_52),
.B2(n_47),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_134),
.A2(n_175),
.B1(n_194),
.B2(n_180),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_116),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_136),
.B(n_138),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_113),
.Y(n_138)
);

INVx6_ASAP7_75t_SL g142 ( 
.A(n_64),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g235 ( 
.A(n_142),
.Y(n_235)
);

INVx13_ASAP7_75t_L g145 ( 
.A(n_59),
.Y(n_145)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_145),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_111),
.A2(n_54),
.B1(n_49),
.B2(n_45),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_88),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_157),
.B(n_176),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_118),
.A2(n_54),
.B1(n_49),
.B2(n_45),
.Y(n_161)
);

BUFx12_ASAP7_75t_L g169 ( 
.A(n_70),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_169),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_76),
.A2(n_40),
.B1(n_29),
.B2(n_20),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_61),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_67),
.B(n_38),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_177),
.B(n_183),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_92),
.B(n_104),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_95),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_184),
.B(n_198),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_103),
.B(n_38),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_185),
.B(n_190),
.Y(n_243)
);

BUFx12_ASAP7_75t_L g186 ( 
.A(n_82),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_186),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_122),
.A2(n_37),
.B1(n_40),
.B2(n_29),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_71),
.A2(n_13),
.B1(n_15),
.B2(n_18),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_120),
.B(n_15),
.Y(n_190)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_81),
.Y(n_193)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_193),
.Y(n_217)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_90),
.Y(n_195)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_195),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_77),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_200),
.B(n_3),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_105),
.B(n_2),
.Y(n_203)
);

AOI21xp33_ASAP7_75t_L g223 ( 
.A1(n_203),
.A2(n_159),
.B(n_162),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_123),
.B(n_2),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_207),
.B(n_140),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_168),
.Y(n_208)
);

INVxp33_ASAP7_75t_L g298 ( 
.A(n_208),
.Y(n_298)
);

INVx6_ASAP7_75t_L g209 ( 
.A(n_141),
.Y(n_209)
);

INVx3_ASAP7_75t_L g305 ( 
.A(n_209),
.Y(n_305)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_205),
.Y(n_213)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_213),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_172),
.B(n_102),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g328 ( 
.A(n_214),
.B(n_223),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_215),
.B(n_218),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_168),
.B(n_98),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g314 ( 
.A(n_216),
.Y(n_314)
);

AO22x1_ASAP7_75t_L g218 ( 
.A1(n_203),
.A2(n_86),
.B1(n_93),
.B2(n_97),
.Y(n_218)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_139),
.Y(n_221)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_221),
.Y(n_278)
);

INVx2_ASAP7_75t_SL g222 ( 
.A(n_205),
.Y(n_222)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_222),
.Y(n_287)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_143),
.Y(n_224)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_224),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_187),
.A2(n_85),
.B(n_4),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_225),
.A2(n_241),
.B(n_274),
.Y(n_284)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_145),
.Y(n_226)
);

INVx5_ASAP7_75t_SL g303 ( 
.A(n_226),
.Y(n_303)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_165),
.Y(n_228)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_228),
.Y(n_320)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_191),
.Y(n_229)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_229),
.Y(n_308)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_166),
.Y(n_230)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_230),
.Y(n_323)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_135),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_231),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_200),
.A2(n_84),
.B1(n_3),
.B2(n_4),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_232),
.A2(n_215),
.B1(n_218),
.B2(n_208),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_156),
.B(n_4),
.C(n_146),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_233),
.B(n_252),
.C(n_275),
.Y(n_301)
);

NAND2x1_ASAP7_75t_SL g234 ( 
.A(n_201),
.B(n_158),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_234),
.A2(n_163),
.B(n_186),
.Y(n_293)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_153),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_236),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_125),
.B(n_160),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_237),
.B(n_240),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_238),
.A2(n_254),
.B1(n_271),
.B2(n_209),
.Y(n_319)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_153),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_239),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_178),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_161),
.A2(n_152),
.B(n_128),
.Y(n_241)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_191),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_242),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_127),
.A2(n_132),
.B1(n_192),
.B2(n_131),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g296 ( 
.A1(n_244),
.A2(n_276),
.B1(n_226),
.B2(n_220),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_167),
.B(n_182),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_245),
.B(n_257),
.Y(n_285)
);

INVx4_ASAP7_75t_L g246 ( 
.A(n_179),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_246),
.B(n_250),
.Y(n_300)
);

INVx11_ASAP7_75t_L g247 ( 
.A(n_155),
.Y(n_247)
);

BUFx24_ASAP7_75t_L g288 ( 
.A(n_247),
.Y(n_288)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_137),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_248),
.B(n_256),
.Y(n_280)
);

INVx6_ASAP7_75t_L g249 ( 
.A(n_141),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_249),
.Y(n_315)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_173),
.Y(n_250)
);

MAJx2_ASAP7_75t_L g252 ( 
.A(n_148),
.B(n_206),
.C(n_178),
.Y(n_252)
);

A2O1A1Ixp33_ASAP7_75t_L g253 ( 
.A1(n_130),
.A2(n_133),
.B(n_154),
.C(n_164),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_253),
.B(n_273),
.Y(n_329)
);

OAI22xp33_ASAP7_75t_L g254 ( 
.A1(n_188),
.A2(n_126),
.B1(n_147),
.B2(n_144),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_154),
.B(n_140),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_124),
.B(n_188),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_124),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_258),
.B(n_259),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_202),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_126),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_260),
.B(n_261),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_147),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_202),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_262),
.B(n_264),
.Y(n_295)
);

AO22x1_ASAP7_75t_L g263 ( 
.A1(n_179),
.A2(n_192),
.B1(n_171),
.B2(n_150),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_263),
.B(n_265),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_202),
.Y(n_264)
);

INVx2_ASAP7_75t_SL g265 ( 
.A(n_155),
.Y(n_265)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_144),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_267),
.B(n_268),
.Y(n_306)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_204),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_174),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_269),
.B(n_222),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_169),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_270),
.B(n_272),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_140),
.B(n_129),
.Y(n_272)
);

O2A1O1Ixp33_ASAP7_75t_L g274 ( 
.A1(n_196),
.A2(n_133),
.B(n_149),
.C(n_150),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_196),
.B(n_180),
.C(n_174),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_181),
.A2(n_197),
.B1(n_155),
.B2(n_199),
.Y(n_276)
);

NAND2x1_ASAP7_75t_L g277 ( 
.A(n_194),
.B(n_199),
.Y(n_277)
);

OR2x2_ASAP7_75t_L g313 ( 
.A(n_277),
.B(n_220),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_215),
.B(n_199),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_279),
.B(n_289),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_238),
.A2(n_204),
.B1(n_170),
.B2(n_171),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_281),
.A2(n_294),
.B1(n_302),
.B2(n_312),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_283),
.A2(n_235),
.B1(n_277),
.B2(n_265),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_252),
.B(n_133),
.Y(n_289)
);

NAND3xp33_ASAP7_75t_SL g292 ( 
.A(n_210),
.B(n_169),
.C(n_186),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_292),
.B(n_311),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_293),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_241),
.A2(n_170),
.B1(n_225),
.B2(n_217),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_296),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_251),
.A2(n_227),
.B1(n_253),
.B2(n_255),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_232),
.B(n_233),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_304),
.B(n_316),
.Y(n_341)
);

MAJx3_ASAP7_75t_L g307 ( 
.A(n_251),
.B(n_234),
.C(n_216),
.Y(n_307)
);

NOR2x1_ASAP7_75t_L g352 ( 
.A(n_307),
.B(n_311),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_216),
.B(n_231),
.C(n_251),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_251),
.A2(n_254),
.B1(n_267),
.B2(n_250),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_313),
.B(n_325),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_266),
.B(n_275),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_243),
.B(n_219),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_318),
.B(n_320),
.Y(n_354)
);

AOI22xp33_ASAP7_75t_L g366 ( 
.A1(n_319),
.A2(n_315),
.B1(n_279),
.B2(n_309),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_249),
.A2(n_268),
.B1(n_242),
.B2(n_229),
.Y(n_321)
);

AO22x1_ASAP7_75t_L g355 ( 
.A1(n_321),
.A2(n_312),
.B1(n_281),
.B2(n_327),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_212),
.B(n_270),
.C(n_213),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_326),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_SL g330 ( 
.A1(n_307),
.A2(n_247),
.B1(n_265),
.B2(n_274),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g385 ( 
.A(n_330),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_332),
.B(n_355),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_307),
.A2(n_222),
.B1(n_263),
.B2(n_246),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_334),
.A2(n_360),
.B1(n_321),
.B2(n_323),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_282),
.B(n_211),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_335),
.B(n_337),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_285),
.B(n_211),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_287),
.Y(n_338)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_338),
.Y(n_370)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_287),
.Y(n_339)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_339),
.Y(n_377)
);

OR2x2_ASAP7_75t_L g340 ( 
.A(n_329),
.B(n_259),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_340),
.B(n_354),
.Y(n_371)
);

INVx3_ASAP7_75t_L g342 ( 
.A(n_305),
.Y(n_342)
);

INVx3_ASAP7_75t_L g372 ( 
.A(n_342),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_SL g343 ( 
.A(n_328),
.B(n_318),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_343),
.B(n_347),
.Y(n_378)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_306),
.Y(n_344)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_344),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_L g346 ( 
.A1(n_289),
.A2(n_262),
.B(n_264),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_SL g387 ( 
.A1(n_346),
.A2(n_352),
.B(n_361),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_328),
.B(n_280),
.Y(n_347)
);

INVx6_ASAP7_75t_SL g349 ( 
.A(n_303),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_349),
.Y(n_379)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_305),
.Y(n_350)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_350),
.Y(n_388)
);

INVx2_ASAP7_75t_SL g351 ( 
.A(n_288),
.Y(n_351)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_351),
.Y(n_390)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_322),
.Y(n_353)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_353),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_283),
.A2(n_291),
.B1(n_304),
.B2(n_316),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_356),
.A2(n_365),
.B1(n_366),
.B2(n_308),
.Y(n_392)
);

A2O1A1Ixp33_ASAP7_75t_L g357 ( 
.A1(n_291),
.A2(n_301),
.B(n_302),
.C(n_284),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_357),
.B(n_359),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_SL g358 ( 
.A(n_298),
.B(n_317),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_358),
.B(n_363),
.Y(n_384)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_278),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_291),
.A2(n_284),
.B1(n_314),
.B2(n_294),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_SL g361 ( 
.A1(n_313),
.A2(n_314),
.B(n_293),
.Y(n_361)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_278),
.Y(n_363)
);

INVx3_ASAP7_75t_L g364 ( 
.A(n_308),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_364),
.B(n_369),
.Y(n_394)
);

OAI22xp33_ASAP7_75t_L g365 ( 
.A1(n_315),
.A2(n_327),
.B1(n_301),
.B2(n_309),
.Y(n_365)
);

O2A1O1Ixp33_ASAP7_75t_L g368 ( 
.A1(n_327),
.A2(n_303),
.B(n_325),
.C(n_299),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_368),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_299),
.B(n_310),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_341),
.B(n_320),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_SL g428 ( 
.A(n_375),
.B(n_381),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_341),
.B(n_310),
.C(n_323),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_376),
.B(n_396),
.C(n_399),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_333),
.B(n_295),
.Y(n_381)
);

AND2x6_ASAP7_75t_L g382 ( 
.A(n_357),
.B(n_290),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_382),
.B(n_331),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_349),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_386),
.B(n_393),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_SL g418 ( 
.A1(n_391),
.A2(n_397),
.B(n_348),
.Y(n_418)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_392),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_358),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_362),
.A2(n_286),
.B1(n_300),
.B2(n_324),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_395),
.A2(n_334),
.B1(n_355),
.B2(n_360),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_333),
.B(n_365),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_SL g397 ( 
.A1(n_361),
.A2(n_324),
.B(n_300),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_352),
.B(n_286),
.C(n_297),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_336),
.B(n_300),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_400),
.B(n_348),
.C(n_344),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_343),
.B(n_297),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_SL g417 ( 
.A(n_401),
.B(n_345),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g402 ( 
.A1(n_398),
.A2(n_353),
.B1(n_362),
.B2(n_345),
.Y(n_402)
);

AOI22xp33_ASAP7_75t_L g439 ( 
.A1(n_402),
.A2(n_376),
.B1(n_377),
.B2(n_368),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_384),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_403),
.B(n_405),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_381),
.B(n_336),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_404),
.B(n_411),
.C(n_415),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_407),
.A2(n_408),
.B1(n_410),
.B2(n_422),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_389),
.A2(n_355),
.B1(n_331),
.B2(n_340),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_389),
.A2(n_331),
.B1(n_340),
.B2(n_354),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_396),
.B(n_336),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_394),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_412),
.B(n_414),
.Y(n_432)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_370),
.Y(n_413)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_413),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_374),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_375),
.B(n_346),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_417),
.B(n_359),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_SL g437 ( 
.A1(n_418),
.A2(n_387),
.B(n_367),
.Y(n_437)
);

BUFx2_ASAP7_75t_L g419 ( 
.A(n_372),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_419),
.Y(n_436)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_370),
.Y(n_420)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_420),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_421),
.B(n_424),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_389),
.A2(n_395),
.B1(n_383),
.B2(n_373),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_380),
.B(n_363),
.Y(n_423)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_423),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_400),
.B(n_399),
.C(n_387),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_371),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_425),
.B(n_377),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_380),
.B(n_398),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_426),
.B(n_427),
.Y(n_444)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_397),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_427),
.A2(n_385),
.B1(n_367),
.B2(n_373),
.Y(n_429)
);

HB1xp67_ASAP7_75t_L g457 ( 
.A(n_429),
.Y(n_457)
);

A2O1A1Ixp33_ASAP7_75t_SL g430 ( 
.A1(n_405),
.A2(n_371),
.B(n_391),
.C(n_385),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_430),
.B(n_433),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_406),
.B(n_379),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_SL g435 ( 
.A(n_426),
.B(n_378),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_435),
.B(n_438),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_437),
.B(n_447),
.Y(n_459)
);

INVxp67_ASAP7_75t_L g438 ( 
.A(n_419),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_439),
.B(n_441),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_442),
.A2(n_446),
.B1(n_448),
.B2(n_420),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_422),
.B(n_338),
.Y(n_445)
);

CKINVDCx16_ASAP7_75t_R g471 ( 
.A(n_445),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_423),
.B(n_388),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_428),
.B(n_404),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_409),
.A2(n_382),
.B1(n_390),
.B2(n_388),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_428),
.B(n_372),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_451),
.B(n_415),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_L g482 ( 
.A1(n_453),
.A2(n_456),
.B1(n_467),
.B2(n_468),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_434),
.B(n_416),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_455),
.B(n_464),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_435),
.A2(n_409),
.B1(n_407),
.B2(n_413),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_440),
.B(n_424),
.C(n_416),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_460),
.B(n_465),
.C(n_429),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_461),
.B(n_432),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_433),
.B(n_421),
.Y(n_462)
);

CKINVDCx16_ASAP7_75t_R g480 ( 
.A(n_462),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_SL g463 ( 
.A(n_434),
.B(n_411),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_SL g479 ( 
.A(n_463),
.B(n_470),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_440),
.B(n_410),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_443),
.B(n_418),
.C(n_408),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_431),
.A2(n_390),
.B1(n_339),
.B2(n_351),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_445),
.A2(n_444),
.B1(n_437),
.B2(n_452),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_444),
.B(n_350),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_469),
.B(n_446),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_SL g470 ( 
.A(n_443),
.B(n_342),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_473),
.B(n_477),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_458),
.Y(n_474)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_474),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_475),
.B(n_478),
.Y(n_492)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_469),
.Y(n_476)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_476),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_455),
.B(n_448),
.C(n_452),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_460),
.B(n_441),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_481),
.B(n_485),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_464),
.B(n_463),
.C(n_465),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_483),
.B(n_457),
.C(n_466),
.Y(n_487)
);

INVx1_ASAP7_75t_SL g484 ( 
.A(n_468),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_484),
.B(n_436),
.Y(n_497)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_471),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g503 ( 
.A(n_487),
.B(n_483),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_484),
.A2(n_454),
.B1(n_459),
.B2(n_430),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_488),
.B(n_438),
.Y(n_507)
);

OAI21xp5_ASAP7_75t_SL g489 ( 
.A1(n_482),
.A2(n_430),
.B(n_470),
.Y(n_489)
);

AOI21xp5_ASAP7_75t_SL g502 ( 
.A1(n_489),
.A2(n_475),
.B(n_479),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_480),
.A2(n_430),
.B1(n_450),
.B2(n_449),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_491),
.A2(n_495),
.B1(n_497),
.B2(n_496),
.Y(n_500)
);

INVxp67_ASAP7_75t_L g494 ( 
.A(n_473),
.Y(n_494)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_494),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_474),
.A2(n_430),
.B1(n_450),
.B2(n_449),
.Y(n_495)
);

OR2x2_ASAP7_75t_L g499 ( 
.A(n_497),
.B(n_491),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_490),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_498),
.B(n_505),
.Y(n_514)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_499),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_500),
.A2(n_507),
.B1(n_486),
.B2(n_472),
.Y(n_510)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_489),
.B(n_478),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_501),
.B(n_503),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_L g508 ( 
.A1(n_502),
.A2(n_488),
.B(n_487),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_492),
.B(n_472),
.C(n_479),
.Y(n_505)
);

OR2x2_ASAP7_75t_L g506 ( 
.A(n_495),
.B(n_436),
.Y(n_506)
);

OAI21x1_ASAP7_75t_L g509 ( 
.A1(n_506),
.A2(n_493),
.B(n_494),
.Y(n_509)
);

AOI21xp5_ASAP7_75t_L g518 ( 
.A1(n_508),
.A2(n_511),
.B(n_499),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_509),
.B(n_510),
.Y(n_516)
);

NOR2xp67_ASAP7_75t_SL g511 ( 
.A(n_502),
.B(n_364),
.Y(n_511)
);

INVx5_ASAP7_75t_L g515 ( 
.A(n_514),
.Y(n_515)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_515),
.Y(n_522)
);

XOR2xp5_ASAP7_75t_L g517 ( 
.A(n_513),
.B(n_501),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_517),
.B(n_518),
.C(n_351),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_512),
.B(n_504),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_SL g520 ( 
.A(n_519),
.B(n_506),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_520),
.B(n_521),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_522),
.B(n_516),
.C(n_517),
.Y(n_524)
);

OAI21xp5_ASAP7_75t_L g525 ( 
.A1(n_524),
.A2(n_515),
.B(n_288),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_525),
.B(n_523),
.C(n_288),
.Y(n_526)
);

OR2x2_ASAP7_75t_L g527 ( 
.A(n_526),
.B(n_288),
.Y(n_527)
);


endmodule