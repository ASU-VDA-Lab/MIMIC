module fake_jpeg_976_n_207 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_207);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_207;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx12_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_51),
.Y(n_53)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_21),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_13),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_10),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_8),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_2),
.Y(n_62)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_45),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_9),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_6),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_10),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_8),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_24),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_7),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_19),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_77),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_67),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_81),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_80),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_67),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_83),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_84),
.Y(n_93)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_77),
.Y(n_85)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_78),
.B(n_61),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_64),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_83),
.B(n_74),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_89),
.B(n_97),
.Y(n_112)
);

CKINVDCx12_ASAP7_75t_R g92 ( 
.A(n_77),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_92),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_81),
.A2(n_66),
.B1(n_68),
.B2(n_56),
.Y(n_94)
);

BUFx5_ASAP7_75t_L g105 ( 
.A(n_94),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_79),
.B(n_57),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_93),
.Y(n_98)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_88),
.Y(n_99)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_99),
.Y(n_130)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_101),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_103),
.B(n_104),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_87),
.B(n_62),
.Y(n_104)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

BUFx4f_ASAP7_75t_SL g119 ( 
.A(n_106),
.Y(n_119)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_91),
.Y(n_107)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_107),
.Y(n_137)
);

A2O1A1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_94),
.A2(n_68),
.B(n_75),
.C(n_55),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_108),
.B(n_111),
.Y(n_125)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_109),
.Y(n_128)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_95),
.Y(n_110)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_110),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_60),
.Y(n_111)
);

INVx3_ASAP7_75t_SL g113 ( 
.A(n_96),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_113),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_71),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_114),
.B(n_0),
.Y(n_135)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_96),
.B(n_80),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_115),
.Y(n_126)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_96),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_116),
.A2(n_72),
.B1(n_63),
.B2(n_59),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_105),
.A2(n_84),
.B1(n_82),
.B2(n_79),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_117),
.A2(n_31),
.B1(n_49),
.B2(n_15),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_108),
.A2(n_76),
.B(n_73),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_121),
.A2(n_52),
.B(n_4),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_112),
.B(n_69),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_122),
.B(n_133),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_100),
.B(n_63),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_124),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_115),
.A2(n_53),
.B1(n_65),
.B2(n_54),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_127),
.A2(n_131),
.B1(n_5),
.B2(n_6),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_106),
.A2(n_53),
.B1(n_65),
.B2(n_54),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_102),
.B(n_0),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_134),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_135),
.B(n_3),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_99),
.B(n_1),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_136),
.B(n_138),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_116),
.B(n_1),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_113),
.B(n_2),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_139),
.B(n_33),
.Y(n_144)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_128),
.Y(n_140)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_140),
.Y(n_169)
);

OA22x2_ASAP7_75t_L g142 ( 
.A1(n_117),
.A2(n_107),
.B1(n_110),
.B2(n_72),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_142),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_125),
.A2(n_59),
.B(n_52),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_143),
.A2(n_148),
.B(n_151),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_144),
.B(n_156),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_119),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_145),
.B(n_150),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_126),
.A2(n_52),
.B(n_4),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_149),
.B(n_153),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_132),
.Y(n_150)
);

INVx13_ASAP7_75t_L g152 ( 
.A(n_132),
.Y(n_152)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_152),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_120),
.B(n_3),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_123),
.B(n_5),
.Y(n_154)
);

NOR4xp25_ASAP7_75t_L g177 ( 
.A(n_154),
.B(n_14),
.C(n_16),
.D(n_18),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_155),
.A2(n_157),
.B1(n_161),
.B2(n_20),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_118),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_134),
.A2(n_7),
.B1(n_9),
.B2(n_11),
.Y(n_157)
);

BUFx12_ASAP7_75t_L g158 ( 
.A(n_119),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_158),
.B(n_159),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_130),
.B(n_11),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_130),
.A2(n_12),
.B(n_13),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_160),
.A2(n_129),
.B(n_137),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_164),
.A2(n_177),
.B(n_160),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_146),
.B(n_137),
.C(n_119),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_165),
.B(n_168),
.C(n_147),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_146),
.B(n_32),
.C(n_47),
.Y(n_168)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_156),
.Y(n_173)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_173),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_162),
.B(n_12),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_174),
.B(n_176),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_141),
.B(n_14),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_178),
.A2(n_155),
.B1(n_147),
.B2(n_157),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_179),
.B(n_181),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_180),
.B(n_186),
.C(n_38),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_167),
.Y(n_181)
);

CKINVDCx14_ASAP7_75t_R g191 ( 
.A(n_182),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_165),
.A2(n_158),
.B(n_152),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_183),
.A2(n_185),
.B1(n_188),
.B2(n_25),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_172),
.A2(n_166),
.B1(n_164),
.B2(n_169),
.Y(n_185)
);

AOI322xp5_ASAP7_75t_L g186 ( 
.A1(n_172),
.A2(n_158),
.A3(n_142),
.B1(n_28),
.B2(n_29),
.C1(n_30),
.C2(n_34),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_175),
.A2(n_142),
.B(n_26),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_180),
.B(n_168),
.C(n_170),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_189),
.B(n_194),
.C(n_195),
.Y(n_197)
);

FAx1_ASAP7_75t_SL g190 ( 
.A(n_181),
.B(n_171),
.CI(n_163),
.CON(n_190),
.SN(n_190)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_190),
.B(n_192),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_184),
.B(n_35),
.C(n_37),
.Y(n_194)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_193),
.Y(n_196)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_196),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_194),
.B(n_187),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_199),
.B(n_189),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_201),
.B(n_197),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_202),
.B(n_200),
.Y(n_203)
);

OR2x2_ASAP7_75t_L g204 ( 
.A(n_203),
.B(n_190),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_204),
.B(n_198),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_205),
.A2(n_191),
.B1(n_40),
.B2(n_44),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_206),
.B(n_39),
.Y(n_207)
);


endmodule