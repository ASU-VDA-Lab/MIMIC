module real_aes_17819_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_357;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_549;
wire n_376;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_666;
wire n_320;
wire n_537;
wire n_551;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_746;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_527;
wire n_434;
wire n_502;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_554;
wire n_475;
wire n_855;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
AND2x4_ASAP7_75t_L g106 ( .A(n_0), .B(n_107), .Y(n_106) );
AOI22xp5_ASAP7_75t_L g529 ( .A1(n_1), .A2(n_4), .B1(n_252), .B2(n_530), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g146 ( .A1(n_2), .A2(n_40), .B1(n_147), .B2(n_149), .Y(n_146) );
AOI22xp33_ASAP7_75t_L g504 ( .A1(n_3), .A2(n_22), .B1(n_149), .B2(n_192), .Y(n_504) );
AOI22xp5_ASAP7_75t_L g242 ( .A1(n_5), .A2(n_15), .B1(n_174), .B2(n_243), .Y(n_242) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_6), .A2(n_57), .B1(n_194), .B2(n_219), .Y(n_555) );
AOI22xp5_ASAP7_75t_L g608 ( .A1(n_7), .A2(n_16), .B1(n_147), .B2(n_178), .Y(n_608) );
INVx1_ASAP7_75t_L g107 ( .A(n_8), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g591 ( .A(n_9), .Y(n_591) );
CKINVDCx5p33_ASAP7_75t_R g206 ( .A(n_10), .Y(n_206) );
AOI22xp5_ASAP7_75t_L g217 ( .A1(n_11), .A2(n_17), .B1(n_176), .B2(n_218), .Y(n_217) );
OR2x2_ASAP7_75t_L g114 ( .A(n_12), .B(n_36), .Y(n_114) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_13), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g246 ( .A(n_14), .Y(n_246) );
AOI22xp5_ASAP7_75t_L g251 ( .A1(n_18), .A2(n_97), .B1(n_174), .B2(n_252), .Y(n_251) );
AOI22xp33_ASAP7_75t_L g239 ( .A1(n_19), .A2(n_37), .B1(n_210), .B2(n_240), .Y(n_239) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_20), .B(n_175), .Y(n_207) );
OAI21x1_ASAP7_75t_L g163 ( .A1(n_21), .A2(n_54), .B(n_164), .Y(n_163) );
CKINVDCx5p33_ASAP7_75t_R g256 ( .A(n_23), .Y(n_256) );
CKINVDCx5p33_ASAP7_75t_R g509 ( .A(n_24), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_25), .B(n_153), .Y(n_516) );
INVx4_ASAP7_75t_R g571 ( .A(n_26), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g154 ( .A1(n_27), .A2(n_44), .B1(n_155), .B2(n_157), .Y(n_154) );
AOI22xp33_ASAP7_75t_L g230 ( .A1(n_28), .A2(n_50), .B1(n_157), .B2(n_174), .Y(n_230) );
CKINVDCx5p33_ASAP7_75t_R g200 ( .A(n_29), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_30), .B(n_210), .Y(n_209) );
CKINVDCx5p33_ASAP7_75t_R g184 ( .A(n_31), .Y(n_184) );
NAND2xp5_ASAP7_75t_SL g523 ( .A(n_32), .B(n_149), .Y(n_523) );
INVx1_ASAP7_75t_L g532 ( .A(n_33), .Y(n_532) );
A2O1A1Ixp33_ASAP7_75t_SL g589 ( .A1(n_34), .A2(n_147), .B(n_159), .C(n_590), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g505 ( .A1(n_35), .A2(n_51), .B1(n_147), .B2(n_157), .Y(n_505) );
AOI22xp5_ASAP7_75t_L g190 ( .A1(n_38), .A2(n_83), .B1(n_147), .B2(n_191), .Y(n_190) );
AOI22xp33_ASAP7_75t_L g221 ( .A1(n_39), .A2(n_43), .B1(n_147), .B2(n_178), .Y(n_221) );
CKINVDCx5p33_ASAP7_75t_R g587 ( .A(n_41), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g254 ( .A1(n_42), .A2(n_56), .B1(n_174), .B2(n_229), .Y(n_254) );
INVx1_ASAP7_75t_L g520 ( .A(n_45), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_46), .B(n_147), .Y(n_522) );
CKINVDCx5p33_ASAP7_75t_R g541 ( .A(n_47), .Y(n_541) );
INVx2_ASAP7_75t_L g126 ( .A(n_48), .Y(n_126) );
INVx1_ASAP7_75t_L g109 ( .A(n_49), .Y(n_109) );
BUFx3_ASAP7_75t_L g129 ( .A(n_49), .Y(n_129) );
AOI22xp33_ASAP7_75t_L g130 ( .A1(n_52), .A2(n_131), .B1(n_837), .B2(n_838), .Y(n_130) );
INVx1_ASAP7_75t_L g837 ( .A(n_52), .Y(n_837) );
CKINVDCx5p33_ASAP7_75t_R g572 ( .A(n_53), .Y(n_572) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_55), .A2(n_85), .B1(n_147), .B2(n_157), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g228 ( .A1(n_58), .A2(n_71), .B1(n_155), .B2(n_229), .Y(n_228) );
CKINVDCx5p33_ASAP7_75t_R g611 ( .A(n_59), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g177 ( .A1(n_60), .A2(n_73), .B1(n_147), .B2(n_178), .Y(n_177) );
AOI22xp5_ASAP7_75t_L g173 ( .A1(n_61), .A2(n_95), .B1(n_174), .B2(n_176), .Y(n_173) );
AND2x4_ASAP7_75t_L g143 ( .A(n_62), .B(n_144), .Y(n_143) );
INVx1_ASAP7_75t_L g164 ( .A(n_63), .Y(n_164) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_64), .Y(n_117) );
AOI22xp33_ASAP7_75t_L g528 ( .A1(n_65), .A2(n_88), .B1(n_155), .B2(n_157), .Y(n_528) );
AO22x1_ASAP7_75t_L g558 ( .A1(n_66), .A2(n_72), .B1(n_240), .B2(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g144 ( .A(n_67), .Y(n_144) );
AND2x2_ASAP7_75t_L g592 ( .A(n_68), .B(n_161), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_69), .B(n_194), .Y(n_547) );
CKINVDCx5p33_ASAP7_75t_R g585 ( .A(n_70), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_74), .B(n_149), .Y(n_542) );
INVx2_ASAP7_75t_L g153 ( .A(n_75), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_76), .B(n_161), .Y(n_513) );
CKINVDCx5p33_ASAP7_75t_R g568 ( .A(n_77), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g193 ( .A1(n_78), .A2(n_96), .B1(n_157), .B2(n_194), .Y(n_193) );
CKINVDCx5p33_ASAP7_75t_R g232 ( .A(n_79), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_80), .B(n_171), .Y(n_556) );
AOI22xp33_ASAP7_75t_L g99 ( .A1(n_81), .A2(n_100), .B1(n_115), .B2(n_858), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g166 ( .A(n_82), .Y(n_166) );
CKINVDCx5p33_ASAP7_75t_R g851 ( .A(n_84), .Y(n_851) );
AOI22xp5_ASAP7_75t_L g844 ( .A1(n_86), .A2(n_132), .B1(n_845), .B2(n_846), .Y(n_844) );
INVx1_ASAP7_75t_L g845 ( .A(n_86), .Y(n_845) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_87), .B(n_161), .Y(n_213) );
CKINVDCx5p33_ASAP7_75t_R g223 ( .A(n_89), .Y(n_223) );
NAND2xp5_ASAP7_75t_SL g538 ( .A(n_90), .B(n_161), .Y(n_538) );
INVx1_ASAP7_75t_L g111 ( .A(n_91), .Y(n_111) );
NAND2xp33_ASAP7_75t_L g211 ( .A(n_92), .B(n_175), .Y(n_211) );
A2O1A1Ixp33_ASAP7_75t_L g566 ( .A1(n_93), .A2(n_180), .B(n_194), .C(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g573 ( .A(n_94), .B(n_574), .Y(n_573) );
NAND2xp33_ASAP7_75t_L g546 ( .A(n_98), .B(n_156), .Y(n_546) );
INVx2_ASAP7_75t_SL g100 ( .A(n_101), .Y(n_100) );
INVx3_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
BUFx6f_ASAP7_75t_SL g102 ( .A(n_103), .Y(n_102) );
BUFx6f_ASAP7_75t_SL g859 ( .A(n_103), .Y(n_859) );
AND2x2_ASAP7_75t_SL g103 ( .A(n_104), .B(n_112), .Y(n_103) );
NOR3xp33_ASAP7_75t_L g104 ( .A(n_105), .B(n_108), .C(n_110), .Y(n_104) );
INVx2_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
AND3x2_ASAP7_75t_L g119 ( .A(n_108), .B(n_110), .C(n_120), .Y(n_119) );
HB1xp67_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
BUFx2_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
INVx2_ASAP7_75t_L g491 ( .A(n_111), .Y(n_491) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_113), .Y(n_112) );
BUFx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
INVx1_ASAP7_75t_L g120 ( .A(n_114), .Y(n_120) );
NOR2x1_ASAP7_75t_L g857 ( .A(n_114), .B(n_129), .Y(n_857) );
OR2x6_ASAP7_75t_L g115 ( .A(n_116), .B(n_121), .Y(n_115) );
INVxp67_ASAP7_75t_SL g847 ( .A(n_116), .Y(n_847) );
NOR2x1_ASAP7_75t_R g116 ( .A(n_117), .B(n_118), .Y(n_116) );
INVx3_ASAP7_75t_L g843 ( .A(n_118), .Y(n_843) );
INVx4_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_120), .B(n_128), .Y(n_127) );
OAI21xp5_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_130), .B(n_839), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_123), .Y(n_122) );
BUFx12f_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
AND2x6_ASAP7_75t_SL g124 ( .A(n_125), .B(n_127), .Y(n_124) );
BUFx3_ASAP7_75t_L g849 ( .A(n_125), .Y(n_849) );
INVx1_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
NOR2xp33_ASAP7_75t_L g854 ( .A(n_126), .B(n_855), .Y(n_854) );
INVx1_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx2_ASAP7_75t_L g838 ( .A(n_131), .Y(n_838) );
OA22x2_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_488), .B1(n_492), .B2(n_494), .Y(n_131) );
INVx2_ASAP7_75t_L g846 ( .A(n_132), .Y(n_846) );
AND2x4_ASAP7_75t_L g132 ( .A(n_133), .B(n_384), .Y(n_132) );
NOR2x1_ASAP7_75t_L g133 ( .A(n_134), .B(n_336), .Y(n_133) );
NAND3xp33_ASAP7_75t_L g134 ( .A(n_135), .B(n_283), .C(n_321), .Y(n_134) );
AOI221xp5_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_214), .B1(n_234), .B2(n_262), .C(n_268), .Y(n_135) );
AOI22xp5_ASAP7_75t_L g460 ( .A1(n_136), .A2(n_461), .B1(n_464), .B2(n_465), .Y(n_460) );
INVx2_ASAP7_75t_SL g136 ( .A(n_137), .Y(n_136) );
OR2x2_ASAP7_75t_L g137 ( .A(n_138), .B(n_185), .Y(n_137) );
INVx1_ASAP7_75t_L g375 ( .A(n_138), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_139), .B(n_167), .Y(n_138) );
INVx1_ASAP7_75t_L g327 ( .A(n_139), .Y(n_327) );
AND2x4_ASAP7_75t_L g370 ( .A(n_139), .B(n_291), .Y(n_370) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
AND2x2_ASAP7_75t_L g298 ( .A(n_140), .B(n_201), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_140), .B(n_267), .Y(n_358) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
AND2x2_ASAP7_75t_L g266 ( .A(n_141), .B(n_267), .Y(n_266) );
OR2x2_ASAP7_75t_L g282 ( .A(n_141), .B(n_187), .Y(n_282) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_141), .Y(n_289) );
INVx1_ASAP7_75t_L g345 ( .A(n_141), .Y(n_345) );
AO31x2_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_145), .A3(n_160), .B(n_165), .Y(n_141) );
INVx2_ASAP7_75t_L g182 ( .A(n_142), .Y(n_182) );
AO31x2_ASAP7_75t_L g215 ( .A1(n_142), .A2(n_169), .A3(n_216), .B(n_222), .Y(n_215) );
AO31x2_ASAP7_75t_L g237 ( .A1(n_142), .A2(n_188), .A3(n_238), .B(n_245), .Y(n_237) );
AO31x2_ASAP7_75t_L g606 ( .A1(n_142), .A2(n_233), .A3(n_607), .B(n_610), .Y(n_606) );
BUFx10_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx1_ASAP7_75t_L g197 ( .A(n_143), .Y(n_197) );
BUFx10_ASAP7_75t_L g507 ( .A(n_143), .Y(n_507) );
INVx1_ASAP7_75t_L g562 ( .A(n_143), .Y(n_562) );
OAI22xp5_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_150), .B1(n_154), .B2(n_158), .Y(n_145) );
INVx1_ASAP7_75t_L g176 ( .A(n_147), .Y(n_176) );
INVx4_ASAP7_75t_L g178 ( .A(n_147), .Y(n_178) );
INVx1_ASAP7_75t_L g229 ( .A(n_147), .Y(n_229) );
INVx3_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_148), .Y(n_149) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_148), .Y(n_156) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_148), .Y(n_157) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_148), .Y(n_175) );
INVx2_ASAP7_75t_L g192 ( .A(n_148), .Y(n_192) );
INVx1_ASAP7_75t_L g194 ( .A(n_148), .Y(n_194) );
INVx1_ASAP7_75t_L g220 ( .A(n_148), .Y(n_220) );
INVx1_ASAP7_75t_L g241 ( .A(n_148), .Y(n_241) );
INVx1_ASAP7_75t_L g244 ( .A(n_148), .Y(n_244) );
INVx1_ASAP7_75t_L g253 ( .A(n_148), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g584 ( .A(n_149), .B(n_585), .Y(n_584) );
OAI22xp5_ASAP7_75t_L g227 ( .A1(n_150), .A2(n_158), .B1(n_228), .B2(n_230), .Y(n_227) );
OAI22xp5_ASAP7_75t_L g238 ( .A1(n_150), .A2(n_158), .B1(n_239), .B2(n_242), .Y(n_238) );
OAI22xp5_ASAP7_75t_L g250 ( .A1(n_150), .A2(n_158), .B1(n_251), .B2(n_254), .Y(n_250) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g506 ( .A(n_151), .Y(n_506) );
BUFx3_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g544 ( .A(n_152), .Y(n_544) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
BUFx8_ASAP7_75t_L g159 ( .A(n_153), .Y(n_159) );
INVx1_ASAP7_75t_L g180 ( .A(n_153), .Y(n_180) );
INVx1_ASAP7_75t_L g519 ( .A(n_153), .Y(n_519) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx1_ASAP7_75t_L g210 ( .A(n_156), .Y(n_210) );
OAI22xp33_ASAP7_75t_L g570 ( .A1(n_156), .A2(n_244), .B1(n_571), .B2(n_572), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_157), .B(n_518), .Y(n_517) );
INVx2_ASAP7_75t_L g530 ( .A(n_157), .Y(n_530) );
OAI22xp5_ASAP7_75t_L g172 ( .A1(n_158), .A2(n_173), .B1(n_177), .B2(n_179), .Y(n_172) );
OAI22xp5_ASAP7_75t_L g189 ( .A1(n_158), .A2(n_190), .B1(n_193), .B2(n_195), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_158), .A2(n_209), .B(n_211), .Y(n_208) );
OAI22xp5_ASAP7_75t_L g216 ( .A1(n_158), .A2(n_179), .B1(n_217), .B2(n_221), .Y(n_216) );
OAI22xp5_ASAP7_75t_L g503 ( .A1(n_158), .A2(n_504), .B1(n_505), .B2(n_506), .Y(n_503) );
OAI22xp5_ASAP7_75t_L g527 ( .A1(n_158), .A2(n_195), .B1(n_528), .B2(n_529), .Y(n_527) );
OAI22x1_ASAP7_75t_L g607 ( .A1(n_158), .A2(n_195), .B1(n_608), .B2(n_609), .Y(n_607) );
INVx6_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
O2A1O1Ixp5_ASAP7_75t_L g205 ( .A1(n_159), .A2(n_178), .B(n_206), .C(n_207), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g545 ( .A1(n_159), .A2(n_546), .B(n_547), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_159), .B(n_558), .Y(n_557) );
A2O1A1Ixp33_ASAP7_75t_L g620 ( .A1(n_159), .A2(n_554), .B(n_558), .C(n_561), .Y(n_620) );
AO31x2_ASAP7_75t_L g502 ( .A1(n_160), .A2(n_503), .A3(n_507), .B(n_508), .Y(n_502) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
NOR2x1_ASAP7_75t_L g548 ( .A(n_161), .B(n_549), .Y(n_548) );
INVx4_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
NOR2xp33_ASAP7_75t_L g165 ( .A(n_162), .B(n_166), .Y(n_165) );
NOR2xp33_ASAP7_75t_L g183 ( .A(n_162), .B(n_184), .Y(n_183) );
BUFx3_ASAP7_75t_L g188 ( .A(n_162), .Y(n_188) );
INVx2_ASAP7_75t_SL g203 ( .A(n_162), .Y(n_203) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_162), .B(n_246), .Y(n_245) );
AND2x2_ASAP7_75t_L g524 ( .A(n_162), .B(n_507), .Y(n_524) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx2_ASAP7_75t_L g171 ( .A(n_163), .Y(n_171) );
INVx3_ASAP7_75t_L g265 ( .A(n_167), .Y(n_265) );
AND2x2_ASAP7_75t_L g280 ( .A(n_167), .B(n_201), .Y(n_280) );
INVx2_ASAP7_75t_L g286 ( .A(n_167), .Y(n_286) );
AND2x4_ASAP7_75t_L g348 ( .A(n_167), .B(n_187), .Y(n_348) );
HB1xp67_ASAP7_75t_L g426 ( .A(n_167), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_167), .B(n_481), .Y(n_480) );
INVx3_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
AND2x2_ASAP7_75t_L g297 ( .A(n_168), .B(n_187), .Y(n_297) );
AND2x2_ASAP7_75t_L g325 ( .A(n_168), .B(n_326), .Y(n_325) );
BUFx2_ASAP7_75t_L g404 ( .A(n_168), .Y(n_404) );
AO31x2_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_172), .A3(n_181), .B(n_183), .Y(n_168) );
AO31x2_ASAP7_75t_L g526 ( .A1(n_169), .A2(n_196), .A3(n_527), .B(n_531), .Y(n_526) );
AOI21x1_ASAP7_75t_L g581 ( .A1(n_169), .A2(n_582), .B(n_592), .Y(n_581) );
BUFx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g508 ( .A(n_170), .B(n_509), .Y(n_508) );
NOR2xp33_ASAP7_75t_L g531 ( .A(n_170), .B(n_532), .Y(n_531) );
INVx2_ASAP7_75t_L g574 ( .A(n_170), .Y(n_574) );
NOR2xp33_ASAP7_75t_L g610 ( .A(n_170), .B(n_611), .Y(n_610) );
INVx2_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx2_ASAP7_75t_L g199 ( .A(n_171), .Y(n_199) );
INVx2_ASAP7_75t_L g233 ( .A(n_171), .Y(n_233) );
OAI21xp33_ASAP7_75t_L g561 ( .A1(n_171), .A2(n_556), .B(n_562), .Y(n_561) );
INVx3_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVxp67_ASAP7_75t_SL g559 ( .A(n_175), .Y(n_559) );
O2A1O1Ixp33_ASAP7_75t_L g540 ( .A1(n_178), .A2(n_541), .B(n_542), .C(n_543), .Y(n_540) );
INVx1_ASAP7_75t_SL g179 ( .A(n_180), .Y(n_179) );
INVx1_ASAP7_75t_L g195 ( .A(n_180), .Y(n_195) );
AO31x2_ASAP7_75t_L g249 ( .A1(n_181), .A2(n_225), .A3(n_250), .B(n_255), .Y(n_249) );
INVx1_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g565 ( .A1(n_182), .A2(n_566), .B(n_569), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_186), .B(n_201), .Y(n_185) );
INVx1_ASAP7_75t_L g360 ( .A(n_186), .Y(n_360) );
NAND2x1_ASAP7_75t_L g388 ( .A(n_186), .B(n_280), .Y(n_388) );
BUFx2_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
OR2x2_ASAP7_75t_L g290 ( .A(n_187), .B(n_291), .Y(n_290) );
INVx2_ASAP7_75t_L g326 ( .A(n_187), .Y(n_326) );
INVx1_ASAP7_75t_L g402 ( .A(n_187), .Y(n_402) );
AO31x2_ASAP7_75t_L g187 ( .A1(n_188), .A2(n_189), .A3(n_196), .B(n_198), .Y(n_187) );
INVx2_ASAP7_75t_SL g191 ( .A(n_192), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g590 ( .A(n_192), .B(n_591), .Y(n_590) );
NAND2xp5_ASAP7_75t_SL g569 ( .A(n_195), .B(n_570), .Y(n_569) );
AO31x2_ASAP7_75t_L g224 ( .A1(n_196), .A2(n_225), .A3(n_227), .B(n_231), .Y(n_224) );
INVx2_ASAP7_75t_SL g196 ( .A(n_197), .Y(n_196) );
INVx2_ASAP7_75t_SL g212 ( .A(n_197), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g198 ( .A(n_199), .B(n_200), .Y(n_198) );
NOR2xp33_ASAP7_75t_SL g222 ( .A(n_199), .B(n_223), .Y(n_222) );
INVx2_ASAP7_75t_L g226 ( .A(n_199), .Y(n_226) );
AND2x4_ASAP7_75t_L g341 ( .A(n_201), .B(n_326), .Y(n_341) );
INVx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
BUFx2_ASAP7_75t_L g363 ( .A(n_202), .Y(n_363) );
OAI21x1_ASAP7_75t_L g202 ( .A1(n_203), .A2(n_204), .B(n_213), .Y(n_202) );
OAI21x1_ASAP7_75t_L g267 ( .A1(n_203), .A2(n_204), .B(n_213), .Y(n_267) );
OAI21x1_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_208), .B(n_212), .Y(n_204) );
AND2x4_ASAP7_75t_L g235 ( .A(n_214), .B(n_236), .Y(n_235) );
AND2x2_ASAP7_75t_L g214 ( .A(n_215), .B(n_224), .Y(n_214) );
INVx4_ASAP7_75t_SL g259 ( .A(n_215), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_215), .B(n_261), .Y(n_271) );
BUFx2_ASAP7_75t_L g335 ( .A(n_215), .Y(n_335) );
AND2x2_ASAP7_75t_L g379 ( .A(n_215), .B(n_237), .Y(n_379) );
INVx1_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g567 ( .A(n_220), .B(n_568), .Y(n_567) );
INVx2_ASAP7_75t_L g257 ( .A(n_224), .Y(n_257) );
OR2x2_ASAP7_75t_L g295 ( .A(n_224), .B(n_237), .Y(n_295) );
INVx2_ASAP7_75t_L g306 ( .A(n_224), .Y(n_306) );
AND2x4_ASAP7_75t_L g309 ( .A(n_224), .B(n_310), .Y(n_309) );
HB1xp67_ASAP7_75t_L g350 ( .A(n_224), .Y(n_350) );
INVx1_ASAP7_75t_L g391 ( .A(n_224), .Y(n_391) );
AO21x2_ASAP7_75t_L g564 ( .A1(n_225), .A2(n_565), .B(n_573), .Y(n_564) );
INVx2_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_232), .B(n_233), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g255 ( .A(n_233), .B(n_256), .Y(n_255) );
OR2x2_ASAP7_75t_L g234 ( .A(n_235), .B(n_247), .Y(n_234) );
INVx2_ASAP7_75t_L g484 ( .A(n_235), .Y(n_484) );
AND2x4_ASAP7_75t_L g445 ( .A(n_236), .B(n_248), .Y(n_445) );
HB1xp67_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
INVx1_ASAP7_75t_L g261 ( .A(n_237), .Y(n_261) );
INVx2_ASAP7_75t_L g310 ( .A(n_237), .Y(n_310) );
INVx1_ASAP7_75t_L g366 ( .A(n_237), .Y(n_366) );
AND2x2_ASAP7_75t_L g392 ( .A(n_237), .B(n_317), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_237), .B(n_305), .Y(n_396) );
OAI21xp33_ASAP7_75t_SL g515 ( .A1(n_240), .A2(n_516), .B(n_517), .Y(n_515) );
INVx1_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
AND2x2_ASAP7_75t_L g247 ( .A(n_248), .B(n_258), .Y(n_247) );
INVx3_ASAP7_75t_L g373 ( .A(n_248), .Y(n_373) );
AND2x4_ASAP7_75t_L g248 ( .A(n_249), .B(n_257), .Y(n_248) );
INVx2_ASAP7_75t_L g277 ( .A(n_249), .Y(n_277) );
INVx2_ASAP7_75t_L g317 ( .A(n_249), .Y(n_317) );
INVx2_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g586 ( .A(n_253), .B(n_587), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_257), .B(n_259), .Y(n_318) );
AND2x2_ASAP7_75t_L g346 ( .A(n_257), .B(n_317), .Y(n_346) );
INVx1_ASAP7_75t_L g272 ( .A(n_258), .Y(n_272) );
NAND2x1_ASAP7_75t_L g408 ( .A(n_258), .B(n_382), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_258), .B(n_346), .Y(n_457) );
AND2x4_ASAP7_75t_L g258 ( .A(n_259), .B(n_260), .Y(n_258) );
INVx2_ASAP7_75t_L g275 ( .A(n_259), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_259), .B(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g365 ( .A(n_259), .B(n_366), .Y(n_365) );
HB1xp67_ASAP7_75t_L g442 ( .A(n_259), .Y(n_442) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
AOI22xp5_ASAP7_75t_L g454 ( .A1(n_262), .A2(n_455), .B1(n_456), .B2(n_458), .Y(n_454) );
INVx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_264), .B(n_266), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_264), .B(n_298), .Y(n_333) );
INVx2_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
AND2x4_ASAP7_75t_L g356 ( .A(n_265), .B(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g455 ( .A(n_265), .B(n_266), .Y(n_455) );
AND2x2_ASAP7_75t_L g328 ( .A(n_266), .B(n_297), .Y(n_328) );
AND2x4_ASAP7_75t_L g347 ( .A(n_266), .B(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g398 ( .A(n_266), .B(n_325), .Y(n_398) );
INVx1_ASAP7_75t_L g291 ( .A(n_267), .Y(n_291) );
AOI31xp33_ASAP7_75t_L g268 ( .A1(n_269), .A2(n_272), .A3(n_273), .B(n_278), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_270), .B(n_313), .Y(n_312) );
HB1xp67_ASAP7_75t_L g464 ( .A(n_270), .Y(n_464) );
OAI21xp33_ASAP7_75t_L g482 ( .A1(n_270), .A2(n_272), .B(n_302), .Y(n_482) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
INVx1_ASAP7_75t_L g324 ( .A(n_271), .Y(n_324) );
HB1xp67_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
OR2x2_ASAP7_75t_L g459 ( .A(n_274), .B(n_295), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
INVx2_ASAP7_75t_L g293 ( .A(n_275), .Y(n_293) );
INVx1_ASAP7_75t_L g314 ( .A(n_276), .Y(n_314) );
HB1xp67_ASAP7_75t_L g421 ( .A(n_276), .Y(n_421) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
INVx2_ASAP7_75t_L g303 ( .A(n_277), .Y(n_303) );
OR2x2_ASAP7_75t_L g331 ( .A(n_277), .B(n_306), .Y(n_331) );
INVx2_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
NOR2x1p5_ASAP7_75t_L g320 ( .A(n_282), .B(n_286), .Y(n_320) );
AOI221xp5_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_292), .B1(n_296), .B2(n_299), .C(n_311), .Y(n_283) );
AND2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_287), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
NOR2x1_ASAP7_75t_L g287 ( .A(n_288), .B(n_290), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g400 ( .A(n_289), .B(n_303), .Y(n_400) );
AND2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
OR2x2_ASAP7_75t_L g330 ( .A(n_293), .B(n_331), .Y(n_330) );
AND2x4_ASAP7_75t_L g417 ( .A(n_293), .B(n_309), .Y(n_417) );
AND2x4_ASAP7_75t_L g334 ( .A(n_294), .B(n_335), .Y(n_334) );
INVx2_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
OR2x2_ASAP7_75t_L g353 ( .A(n_295), .B(n_316), .Y(n_353) );
AND2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
AND2x4_ASAP7_75t_SL g369 ( .A(n_297), .B(n_370), .Y(n_369) );
INVx1_ASAP7_75t_SL g410 ( .A(n_297), .Y(n_410) );
INVx2_ASAP7_75t_L g419 ( .A(n_297), .Y(n_419) );
AND2x2_ASAP7_75t_L g433 ( .A(n_297), .B(n_363), .Y(n_433) );
INVx1_ASAP7_75t_L g411 ( .A(n_298), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_300), .B(n_307), .Y(n_299) );
OR2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_304), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_301), .B(n_395), .Y(n_394) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
NAND2x1p5_ASAP7_75t_L g343 ( .A(n_302), .B(n_309), .Y(n_343) );
AND2x2_ASAP7_75t_L g364 ( .A(n_302), .B(n_365), .Y(n_364) );
NAND2x1_ASAP7_75t_L g472 ( .A(n_302), .B(n_334), .Y(n_472) );
INVx3_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
HB1xp67_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
AOI21xp5_ASAP7_75t_L g311 ( .A1(n_312), .A2(n_315), .B(n_319), .Y(n_311) );
NAND2x1_ASAP7_75t_L g473 ( .A(n_313), .B(n_417), .Y(n_473) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_314), .B(n_324), .Y(n_323) );
OR2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_318), .Y(n_315) );
INVx4_ASAP7_75t_L g382 ( .A(n_316), .Y(n_382) );
AND2x2_ASAP7_75t_L g452 ( .A(n_316), .B(n_357), .Y(n_452) );
INVx3_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g349 ( .A(n_317), .B(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g362 ( .A(n_320), .B(n_363), .Y(n_362) );
NOR2x1_ASAP7_75t_L g432 ( .A(n_320), .B(n_433), .Y(n_432) );
AOI322xp5_ASAP7_75t_L g321 ( .A1(n_322), .A2(n_325), .A3(n_327), .B1(n_328), .B2(n_329), .C1(n_332), .C2(n_334), .Y(n_321) );
INVxp67_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g415 ( .A(n_325), .B(n_363), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_325), .B(n_429), .Y(n_428) );
AND2x2_ASAP7_75t_L g439 ( .A(n_325), .B(n_440), .Y(n_439) );
AND2x2_ASAP7_75t_L g444 ( .A(n_325), .B(n_429), .Y(n_444) );
INVx1_ASAP7_75t_L g453 ( .A(n_325), .Y(n_453) );
OR2x2_ASAP7_75t_L g339 ( .A(n_327), .B(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g466 ( .A(n_327), .Y(n_466) );
AND2x2_ASAP7_75t_L g469 ( .A(n_328), .B(n_470), .Y(n_469) );
INVx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
NOR3xp33_ASAP7_75t_L g405 ( .A(n_331), .B(n_345), .C(n_406), .Y(n_405) );
INVx2_ASAP7_75t_L g447 ( .A(n_331), .Y(n_447) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
NAND3xp33_ASAP7_75t_SL g336 ( .A(n_337), .B(n_351), .C(n_361), .Y(n_336) );
AOI222xp33_ASAP7_75t_L g337 ( .A1(n_338), .A2(n_342), .B1(n_344), .B2(n_346), .C1(n_347), .C2(n_349), .Y(n_337) );
INVxp67_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
OAI22x1_ASAP7_75t_L g483 ( .A1(n_340), .A2(n_484), .B1(n_485), .B2(n_486), .Y(n_483) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
AND2x4_ASAP7_75t_L g344 ( .A(n_341), .B(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_341), .B(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g437 ( .A(n_341), .B(n_403), .Y(n_437) );
AND2x4_ASAP7_75t_L g467 ( .A(n_341), .B(n_404), .Y(n_467) );
AND2x2_ASAP7_75t_L g448 ( .A(n_342), .B(n_415), .Y(n_448) );
INVx2_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx2_ASAP7_75t_L g440 ( .A(n_345), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_346), .B(n_379), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_346), .B(n_365), .Y(n_463) );
INVx1_ASAP7_75t_L g383 ( .A(n_347), .Y(n_383) );
INVx2_ASAP7_75t_L g427 ( .A(n_349), .Y(n_427) );
INVx1_ASAP7_75t_L g377 ( .A(n_350), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_352), .B(n_354), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
NAND2x1p5_ASAP7_75t_L g355 ( .A(n_356), .B(n_359), .Y(n_355) );
AOI221xp5_ASAP7_75t_SL g443 ( .A1(n_356), .A2(n_444), .B1(n_445), .B2(n_446), .C(n_448), .Y(n_443) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g429 ( .A(n_358), .Y(n_429) );
INVxp67_ASAP7_75t_SL g481 ( .A(n_358), .Y(n_481) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
NOR2xp33_ASAP7_75t_L g475 ( .A(n_360), .B(n_466), .Y(n_475) );
AOI221xp5_ASAP7_75t_L g361 ( .A1(n_362), .A2(n_364), .B1(n_367), .B2(n_378), .C(n_380), .Y(n_361) );
OR2x2_ASAP7_75t_L g418 ( .A(n_363), .B(n_419), .Y(n_418) );
AOI32xp33_ASAP7_75t_L g399 ( .A1(n_365), .A2(n_379), .A3(n_400), .B1(n_401), .B2(n_405), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_365), .B(n_421), .Y(n_420) );
OAI22xp5_ASAP7_75t_L g367 ( .A1(n_368), .A2(n_371), .B1(n_374), .B2(n_376), .Y(n_367) );
INVx3_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_370), .B(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
OR2x2_ASAP7_75t_L g441 ( .A(n_373), .B(n_442), .Y(n_441) );
HB1xp67_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
AND2x2_ASAP7_75t_L g434 ( .A(n_377), .B(n_379), .Y(n_434) );
AND2x2_ASAP7_75t_L g487 ( .A(n_377), .B(n_392), .Y(n_487) );
AND2x2_ASAP7_75t_L g446 ( .A(n_378), .B(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_379), .B(n_382), .Y(n_381) );
NOR2xp33_ASAP7_75t_L g380 ( .A(n_381), .B(n_383), .Y(n_380) );
NOR2x1_ASAP7_75t_L g384 ( .A(n_385), .B(n_449), .Y(n_384) );
NAND4xp75_ASAP7_75t_L g385 ( .A(n_386), .B(n_412), .C(n_430), .D(n_443), .Y(n_385) );
AOI211x1_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_389), .B(n_393), .C(n_407), .Y(n_386) );
INVxp67_ASAP7_75t_L g485 ( .A(n_387), .Y(n_485) );
INVx2_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
AND2x2_ASAP7_75t_L g389 ( .A(n_390), .B(n_392), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
OAI21xp33_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_397), .B(n_399), .Y(n_393) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVxp67_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
AND2x2_ASAP7_75t_L g401 ( .A(n_402), .B(n_403), .Y(n_401) );
BUFx2_ASAP7_75t_L g406 ( .A(n_402), .Y(n_406) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g478 ( .A(n_406), .Y(n_478) );
NOR3xp33_ASAP7_75t_L g407 ( .A(n_408), .B(n_409), .C(n_411), .Y(n_407) );
INVx2_ASAP7_75t_L g470 ( .A(n_408), .Y(n_470) );
INVx2_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
NOR2x1_ASAP7_75t_L g412 ( .A(n_413), .B(n_422), .Y(n_412) );
OAI22xp5_ASAP7_75t_L g413 ( .A1(n_414), .A2(n_416), .B1(n_418), .B2(n_420), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx2_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
OAI22xp5_ASAP7_75t_L g422 ( .A1(n_423), .A2(n_424), .B1(n_427), .B2(n_428), .Y(n_422) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
AOI21xp5_ASAP7_75t_L g430 ( .A1(n_431), .A2(n_434), .B(n_435), .Y(n_430) );
INVxp67_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
AOI21xp33_ASAP7_75t_L g435 ( .A1(n_436), .A2(n_438), .B(n_441), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_442), .B(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g462 ( .A(n_445), .Y(n_462) );
NAND4xp75_ASAP7_75t_SL g449 ( .A(n_450), .B(n_460), .C(n_468), .D(n_476), .Y(n_449) );
OA21x2_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_453), .B(n_454), .Y(n_450) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_462), .B(n_463), .Y(n_461) );
AND2x2_ASAP7_75t_L g465 ( .A(n_466), .B(n_467), .Y(n_465) );
NOR2xp67_ASAP7_75t_SL g468 ( .A(n_469), .B(n_471), .Y(n_468) );
AOI21xp5_ASAP7_75t_L g471 ( .A1(n_472), .A2(n_473), .B(n_474), .Y(n_471) );
INVxp67_ASAP7_75t_SL g474 ( .A(n_475), .Y(n_474) );
AOI21x1_ASAP7_75t_L g476 ( .A1(n_477), .A2(n_482), .B(n_483), .Y(n_476) );
AND2x4_ASAP7_75t_L g477 ( .A(n_478), .B(n_479), .Y(n_477) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx8_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
BUFx12f_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
CKINVDCx5p33_ASAP7_75t_R g490 ( .A(n_491), .Y(n_490) );
BUFx8_ASAP7_75t_SL g493 ( .A(n_491), .Y(n_493) );
AND2x2_ASAP7_75t_L g856 ( .A(n_491), .B(n_857), .Y(n_856) );
INVx3_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
AND2x4_ASAP7_75t_L g494 ( .A(n_495), .B(n_727), .Y(n_494) );
NOR4xp25_ASAP7_75t_L g495 ( .A(n_496), .B(n_627), .C(n_669), .D(n_701), .Y(n_495) );
OAI211xp5_ASAP7_75t_L g496 ( .A1(n_497), .A2(n_533), .B(n_575), .C(n_612), .Y(n_496) );
HB1xp67_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
AND2x4_ASAP7_75t_L g499 ( .A(n_500), .B(n_510), .Y(n_499) );
INVx2_ASAP7_75t_L g640 ( .A(n_500), .Y(n_640) );
INVx2_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
AND2x2_ASAP7_75t_L g719 ( .A(n_501), .B(n_512), .Y(n_719) );
BUFx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_502), .B(n_526), .Y(n_578) );
AND2x2_ASAP7_75t_L g601 ( .A(n_502), .B(n_602), .Y(n_601) );
INVx2_ASAP7_75t_SL g626 ( .A(n_502), .Y(n_626) );
OR2x2_ASAP7_75t_L g689 ( .A(n_502), .B(n_526), .Y(n_689) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_506), .A2(n_522), .B(n_523), .Y(n_521) );
OAI21x1_ASAP7_75t_L g554 ( .A1(n_506), .A2(n_555), .B(n_556), .Y(n_554) );
INVx1_ASAP7_75t_L g549 ( .A(n_507), .Y(n_549) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
OR2x2_ASAP7_75t_L g623 ( .A(n_511), .B(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g635 ( .A(n_511), .Y(n_635) );
INVxp67_ASAP7_75t_SL g813 ( .A(n_511), .Y(n_813) );
OR2x2_ASAP7_75t_L g826 ( .A(n_511), .B(n_827), .Y(n_826) );
OR2x2_ASAP7_75t_L g511 ( .A(n_512), .B(n_525), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_512), .B(n_580), .Y(n_579) );
INVx3_ASAP7_75t_L g599 ( .A(n_512), .Y(n_599) );
AND2x2_ASAP7_75t_L g646 ( .A(n_512), .B(n_647), .Y(n_646) );
NAND2x1p5_ASAP7_75t_SL g665 ( .A(n_512), .B(n_666), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_512), .B(n_600), .Y(n_715) );
INVx1_ASAP7_75t_L g804 ( .A(n_512), .Y(n_804) );
AND2x2_ASAP7_75t_L g833 ( .A(n_512), .B(n_526), .Y(n_833) );
AND2x4_ASAP7_75t_L g512 ( .A(n_513), .B(n_514), .Y(n_512) );
OAI21xp5_ASAP7_75t_L g514 ( .A1(n_515), .A2(n_521), .B(n_524), .Y(n_514) );
NOR2xp33_ASAP7_75t_L g518 ( .A(n_519), .B(n_520), .Y(n_518) );
BUFx4f_ASAP7_75t_L g588 ( .A(n_519), .Y(n_588) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g600 ( .A(n_526), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_526), .B(n_626), .Y(n_648) );
INVx1_ASAP7_75t_L g668 ( .A(n_526), .Y(n_668) );
NOR2xp33_ASAP7_75t_L g720 ( .A(n_526), .B(n_602), .Y(n_720) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_535), .B(n_550), .Y(n_534) );
OR2x2_ASAP7_75t_L g617 ( .A(n_535), .B(n_618), .Y(n_617) );
OR2x2_ASAP7_75t_L g724 ( .A(n_535), .B(n_673), .Y(n_724) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx1_ASAP7_75t_L g633 ( .A(n_536), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_536), .B(n_653), .Y(n_652) );
NOR2x1_ASAP7_75t_L g738 ( .A(n_536), .B(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx2_ASAP7_75t_L g596 ( .A(n_537), .Y(n_596) );
BUFx3_ASAP7_75t_L g644 ( .A(n_537), .Y(n_644) );
AND2x2_ASAP7_75t_L g680 ( .A(n_537), .B(n_661), .Y(n_680) );
AND2x2_ASAP7_75t_L g760 ( .A(n_537), .B(n_606), .Y(n_760) );
AND2x2_ASAP7_75t_L g773 ( .A(n_537), .B(n_564), .Y(n_773) );
NAND2x1p5_ASAP7_75t_L g537 ( .A(n_538), .B(n_539), .Y(n_537) );
OAI21x1_ASAP7_75t_L g539 ( .A1(n_540), .A2(n_545), .B(n_548), .Y(n_539) );
INVx2_ASAP7_75t_SL g543 ( .A(n_544), .Y(n_543) );
INVx2_ASAP7_75t_L g713 ( .A(n_550), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_550), .B(n_643), .Y(n_721) );
AND2x2_ASAP7_75t_L g550 ( .A(n_551), .B(n_563), .Y(n_550) );
AND2x2_ASAP7_75t_L g632 ( .A(n_551), .B(n_564), .Y(n_632) );
INVx1_ASAP7_75t_L g740 ( .A(n_551), .Y(n_740) );
INVx2_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
AND2x4_ASAP7_75t_L g594 ( .A(n_552), .B(n_564), .Y(n_594) );
AND2x2_ASAP7_75t_L g657 ( .A(n_552), .B(n_563), .Y(n_657) );
AOI21x1_ASAP7_75t_L g552 ( .A1(n_553), .A2(n_557), .B(n_560), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
AOI21xp5_ASAP7_75t_L g582 ( .A1(n_562), .A2(n_583), .B(n_589), .Y(n_582) );
AND2x2_ASAP7_75t_L g615 ( .A(n_563), .B(n_606), .Y(n_615) );
INVx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g605 ( .A(n_564), .B(n_606), .Y(n_605) );
OR2x2_ASAP7_75t_L g673 ( .A(n_564), .B(n_606), .Y(n_673) );
INVx1_ASAP7_75t_L g684 ( .A(n_564), .Y(n_684) );
AND2x2_ASAP7_75t_L g747 ( .A(n_564), .B(n_596), .Y(n_747) );
AOI22xp33_ASAP7_75t_L g575 ( .A1(n_576), .A2(n_593), .B1(n_597), .B2(n_603), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g645 ( .A1(n_576), .A2(n_646), .B1(n_649), .B2(n_651), .Y(n_645) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
OR2x2_ASAP7_75t_L g577 ( .A(n_578), .B(n_579), .Y(n_577) );
OR2x2_ASAP7_75t_L g725 ( .A(n_578), .B(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g831 ( .A(n_578), .Y(n_831) );
INVx1_ASAP7_75t_L g690 ( .A(n_579), .Y(n_690) );
OR2x2_ASAP7_75t_L g753 ( .A(n_579), .B(n_648), .Y(n_753) );
OR2x2_ASAP7_75t_L g624 ( .A(n_580), .B(n_625), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_580), .B(n_599), .Y(n_700) );
AND2x2_ASAP7_75t_L g717 ( .A(n_580), .B(n_644), .Y(n_717) );
HB1xp67_ASAP7_75t_L g734 ( .A(n_580), .Y(n_734) );
INVxp67_ASAP7_75t_L g782 ( .A(n_580), .Y(n_782) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx2_ASAP7_75t_L g602 ( .A(n_581), .Y(n_602) );
OAI21xp5_ASAP7_75t_L g583 ( .A1(n_584), .A2(n_586), .B(n_588), .Y(n_583) );
AND2x2_ASAP7_75t_L g593 ( .A(n_594), .B(n_595), .Y(n_593) );
HB1xp67_ASAP7_75t_L g692 ( .A(n_594), .Y(n_692) );
INVx3_ASAP7_75t_L g697 ( .A(n_594), .Y(n_697) );
AND2x2_ASAP7_75t_L g710 ( .A(n_594), .B(n_711), .Y(n_710) );
AND2x2_ASAP7_75t_L g810 ( .A(n_594), .B(n_772), .Y(n_810) );
INVx1_ASAP7_75t_L g604 ( .A(n_595), .Y(n_604) );
OR2x2_ASAP7_75t_L g787 ( .A(n_595), .B(n_762), .Y(n_787) );
BUFx2_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
AND2x2_ASAP7_75t_L g711 ( .A(n_596), .B(n_621), .Y(n_711) );
AND2x2_ASAP7_75t_L g732 ( .A(n_596), .B(n_657), .Y(n_732) );
AND2x2_ASAP7_75t_L g597 ( .A(n_598), .B(n_601), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_598), .B(n_640), .Y(n_639) );
INVx2_ASAP7_75t_L g733 ( .A(n_598), .Y(n_733) );
AND2x2_ASAP7_75t_L g775 ( .A(n_598), .B(n_776), .Y(n_775) );
AND2x4_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
INVx2_ASAP7_75t_L g676 ( .A(n_599), .Y(n_676) );
AND2x2_ASAP7_75t_L g707 ( .A(n_599), .B(n_708), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_599), .B(n_666), .Y(n_726) );
AND2x2_ASAP7_75t_L g675 ( .A(n_601), .B(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g791 ( .A(n_601), .Y(n_791) );
AND2x2_ASAP7_75t_L g814 ( .A(n_601), .B(n_804), .Y(n_814) );
INVx1_ASAP7_75t_L g827 ( .A(n_601), .Y(n_827) );
INVx2_ASAP7_75t_L g666 ( .A(n_602), .Y(n_666) );
OR2x2_ASAP7_75t_L g762 ( .A(n_602), .B(n_626), .Y(n_762) );
AND2x2_ASAP7_75t_L g603 ( .A(n_604), .B(n_605), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_605), .B(n_643), .Y(n_650) );
INVx2_ASAP7_75t_L g621 ( .A(n_606), .Y(n_621) );
INVx2_ASAP7_75t_L g661 ( .A(n_606), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_606), .B(n_619), .Y(n_683) );
OAI21xp33_ASAP7_75t_L g612 ( .A1(n_613), .A2(n_616), .B(n_622), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx2_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_615), .B(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
OR2x2_ASAP7_75t_L g756 ( .A(n_618), .B(n_757), .Y(n_756) );
OR2x2_ASAP7_75t_L g618 ( .A(n_619), .B(n_621), .Y(n_618) );
INVx2_ASAP7_75t_L g662 ( .A(n_619), .Y(n_662) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g653 ( .A(n_621), .Y(n_653) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g636 ( .A(n_624), .Y(n_636) );
INVxp67_ASAP7_75t_L g807 ( .A(n_624), .Y(n_807) );
OR2x2_ASAP7_75t_L g709 ( .A(n_625), .B(n_666), .Y(n_709) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
NAND4xp25_ASAP7_75t_L g627 ( .A(n_628), .B(n_637), .C(n_645), .D(n_654), .Y(n_627) );
NAND3xp33_ASAP7_75t_L g628 ( .A(n_629), .B(n_634), .C(n_636), .Y(n_628) );
INVx3_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
A2O1A1Ixp33_ASAP7_75t_L g823 ( .A1(n_630), .A2(n_824), .B(n_826), .C(n_828), .Y(n_823) );
OR2x6_ASAP7_75t_L g630 ( .A(n_631), .B(n_633), .Y(n_630) );
INVx2_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_632), .B(n_680), .Y(n_679) );
NOR3xp33_ASAP7_75t_L g735 ( .A(n_632), .B(n_736), .C(n_738), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g816 ( .A(n_632), .B(n_711), .Y(n_816) );
AOI221xp5_ASAP7_75t_L g828 ( .A1(n_632), .A2(n_737), .B1(n_829), .B2(n_832), .C(n_834), .Y(n_828) );
INVx1_ASAP7_75t_L g819 ( .A(n_633), .Y(n_819) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_638), .B(n_641), .Y(n_637) );
AOI221xp5_ASAP7_75t_L g754 ( .A1(n_638), .A2(n_646), .B1(n_681), .B2(n_755), .C(n_758), .Y(n_754) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g812 ( .A(n_640), .B(n_813), .Y(n_812) );
INVx1_ASAP7_75t_L g705 ( .A(n_641), .Y(n_705) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
NAND2x1p5_ASAP7_75t_L g659 ( .A(n_643), .B(n_660), .Y(n_659) );
AND2x2_ASAP7_75t_L g820 ( .A(n_643), .B(n_671), .Y(n_820) );
INVx3_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
BUFx2_ASAP7_75t_L g656 ( .A(n_644), .Y(n_656) );
AND3x1_ASAP7_75t_L g829 ( .A(n_644), .B(n_830), .C(n_831), .Y(n_829) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
OR2x2_ASAP7_75t_L g699 ( .A(n_648), .B(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g769 ( .A(n_651), .Y(n_769) );
INVx2_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
OR2x2_ASAP7_75t_L g745 ( .A(n_653), .B(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g772 ( .A(n_653), .Y(n_772) );
OAI21xp5_ASAP7_75t_L g654 ( .A1(n_655), .A2(n_658), .B(n_663), .Y(n_654) );
AND2x2_ASAP7_75t_L g655 ( .A(n_656), .B(n_657), .Y(n_655) );
NAND2x1_ASAP7_75t_L g670 ( .A(n_656), .B(n_671), .Y(n_670) );
INVx2_ASAP7_75t_L g737 ( .A(n_657), .Y(n_737) );
INVxp67_ASAP7_75t_SL g658 ( .A(n_659), .Y(n_658) );
AND2x2_ASAP7_75t_L g660 ( .A(n_661), .B(n_662), .Y(n_660) );
INVx1_ASAP7_75t_L g693 ( .A(n_661), .Y(n_693) );
OR2x2_ASAP7_75t_L g672 ( .A(n_662), .B(n_673), .Y(n_672) );
INVx2_ASAP7_75t_L g785 ( .A(n_662), .Y(n_785) );
INVx2_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g811 ( .A(n_664), .B(n_812), .Y(n_811) );
OR2x2_ASAP7_75t_L g664 ( .A(n_665), .B(n_667), .Y(n_664) );
OR2x2_ASAP7_75t_L g741 ( .A(n_665), .B(n_689), .Y(n_741) );
INVx2_ASAP7_75t_L g830 ( .A(n_665), .Y(n_830) );
INVx1_ASAP7_75t_L g704 ( .A(n_666), .Y(n_704) );
NOR4xp25_ASAP7_75t_L g834 ( .A(n_666), .B(n_697), .C(n_835), .D(n_836), .Y(n_834) );
INVx1_ASAP7_75t_L g836 ( .A(n_667), .Y(n_836) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
BUFx3_ASAP7_75t_L g822 ( .A(n_668), .Y(n_822) );
OAI211xp5_ASAP7_75t_SL g669 ( .A1(n_670), .A2(n_674), .B(n_677), .C(n_685), .Y(n_669) );
INVx2_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g809 ( .A(n_672), .Y(n_809) );
INVx2_ASAP7_75t_L g794 ( .A(n_673), .Y(n_794) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
OAI21xp5_ASAP7_75t_L g677 ( .A1(n_675), .A2(n_678), .B(n_681), .Y(n_677) );
OR2x2_ASAP7_75t_L g761 ( .A(n_676), .B(n_762), .Y(n_761) );
AND2x2_ASAP7_75t_L g779 ( .A(n_676), .B(n_780), .Y(n_779) );
INVxp67_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g695 ( .A(n_680), .Y(n_695) );
AND2x4_ASAP7_75t_SL g784 ( .A(n_680), .B(n_785), .Y(n_784) );
INVx3_ASAP7_75t_R g681 ( .A(n_682), .Y(n_681) );
OR2x2_ASAP7_75t_L g682 ( .A(n_683), .B(n_684), .Y(n_682) );
HB1xp67_ASAP7_75t_L g750 ( .A(n_683), .Y(n_750) );
INVx1_ASAP7_75t_L g757 ( .A(n_684), .Y(n_757) );
AOI32xp33_ASAP7_75t_L g685 ( .A1(n_686), .A2(n_691), .A3(n_693), .B1(n_694), .B2(n_698), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_688), .B(n_690), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_688), .B(n_704), .Y(n_703) );
HB1xp67_ASAP7_75t_L g749 ( .A(n_688), .Y(n_749) );
INVx2_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
OR2x2_ASAP7_75t_L g766 ( .A(n_689), .B(n_704), .Y(n_766) );
INVx2_ASAP7_75t_L g780 ( .A(n_689), .Y(n_780) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
NOR2xp33_ASAP7_75t_L g694 ( .A(n_695), .B(n_696), .Y(n_694) );
INVx2_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
NAND2xp5_ASAP7_75t_SL g759 ( .A(n_697), .B(n_760), .Y(n_759) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
OAI211xp5_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_705), .B(n_706), .C(n_722), .Y(n_701) );
HB1xp67_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
AOI21xp5_ASAP7_75t_L g706 ( .A1(n_707), .A2(n_710), .B(n_712), .Y(n_706) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g763 ( .A(n_711), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g797 ( .A(n_711), .B(n_798), .Y(n_797) );
OAI32xp33_ASAP7_75t_L g712 ( .A1(n_713), .A2(n_714), .A3(n_716), .B1(n_718), .B2(n_721), .Y(n_712) );
INVx1_ASAP7_75t_L g798 ( .A(n_713), .Y(n_798) );
HB1xp67_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
OR2x2_ASAP7_75t_L g790 ( .A(n_715), .B(n_791), .Y(n_790) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_719), .B(n_720), .Y(n_718) );
INVxp67_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
NOR2xp33_ASAP7_75t_L g723 ( .A(n_724), .B(n_725), .Y(n_723) );
NOR2x1_ASAP7_75t_L g727 ( .A(n_728), .B(n_799), .Y(n_727) );
NAND4xp25_ASAP7_75t_L g728 ( .A(n_729), .B(n_754), .C(n_767), .D(n_795), .Y(n_728) );
NOR2xp67_ASAP7_75t_L g729 ( .A(n_730), .B(n_742), .Y(n_729) );
OAI32xp33_ASAP7_75t_L g730 ( .A1(n_731), .A2(n_733), .A3(n_734), .B1(n_735), .B2(n_741), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
OR2x2_ASAP7_75t_L g781 ( .A(n_733), .B(n_782), .Y(n_781) );
OAI32xp33_ASAP7_75t_L g786 ( .A1(n_733), .A2(n_787), .A3(n_788), .B1(n_790), .B2(n_792), .Y(n_786) );
NOR2xp33_ASAP7_75t_L g821 ( .A(n_734), .B(n_822), .Y(n_821) );
NAND2xp5_ASAP7_75t_SL g800 ( .A(n_736), .B(n_801), .Y(n_800) );
INVx3_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
AND2x2_ASAP7_75t_L g793 ( .A(n_739), .B(n_794), .Y(n_793) );
INVx1_ASAP7_75t_L g825 ( .A(n_739), .Y(n_825) );
INVx2_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g789 ( .A(n_740), .Y(n_789) );
OAI22x1_ASAP7_75t_L g742 ( .A1(n_743), .A2(n_748), .B1(n_750), .B2(n_751), .Y(n_742) );
INVx2_ASAP7_75t_SL g743 ( .A(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx2_ASAP7_75t_SL g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g795 ( .A(n_752), .B(n_796), .Y(n_795) );
INVx2_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx3_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
NOR2x1_ASAP7_75t_L g818 ( .A(n_756), .B(n_819), .Y(n_818) );
OAI22xp5_ASAP7_75t_L g758 ( .A1(n_759), .A2(n_761), .B1(n_763), .B2(n_764), .Y(n_758) );
NAND2x1_ASAP7_75t_L g824 ( .A(n_760), .B(n_825), .Y(n_824) );
INVx2_ASAP7_75t_L g835 ( .A(n_760), .Y(n_835) );
INVx2_ASAP7_75t_L g776 ( .A(n_762), .Y(n_776) );
INVx2_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
INVx2_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
NOR3xp33_ASAP7_75t_SL g767 ( .A(n_768), .B(n_777), .C(n_786), .Y(n_767) );
AOI21xp5_ASAP7_75t_L g768 ( .A1(n_769), .A2(n_770), .B(n_774), .Y(n_768) );
NAND2xp33_ASAP7_75t_L g796 ( .A(n_770), .B(n_797), .Y(n_796) );
INVx2_ASAP7_75t_SL g770 ( .A(n_771), .Y(n_770) );
AND2x2_ASAP7_75t_L g771 ( .A(n_772), .B(n_773), .Y(n_771) );
INVx1_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
AND2x4_ASAP7_75t_L g832 ( .A(n_776), .B(n_833), .Y(n_832) );
AOI21xp5_ASAP7_75t_L g777 ( .A1(n_778), .A2(n_781), .B(n_783), .Y(n_777) );
INVx1_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
AND2x4_ASAP7_75t_L g803 ( .A(n_780), .B(n_804), .Y(n_803) );
INVxp67_ASAP7_75t_SL g802 ( .A(n_782), .Y(n_802) );
INVx1_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
INVxp67_ASAP7_75t_SL g788 ( .A(n_789), .Y(n_788) );
INVx2_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
NAND3xp33_ASAP7_75t_SL g799 ( .A(n_800), .B(n_805), .C(n_817), .Y(n_799) );
AND2x2_ASAP7_75t_L g801 ( .A(n_802), .B(n_803), .Y(n_801) );
INVx1_ASAP7_75t_L g808 ( .A(n_804), .Y(n_808) );
AOI222xp33_ASAP7_75t_L g805 ( .A1(n_806), .A2(n_809), .B1(n_810), .B2(n_811), .C1(n_814), .C2(n_815), .Y(n_805) );
AND2x2_ASAP7_75t_L g806 ( .A(n_807), .B(n_808), .Y(n_806) );
INVx1_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
O2A1O1Ixp5_ASAP7_75t_L g817 ( .A1(n_818), .A2(n_820), .B(n_821), .C(n_823), .Y(n_817) );
AOI21xp5_ASAP7_75t_L g839 ( .A1(n_840), .A2(n_848), .B(n_850), .Y(n_839) );
OAI21xp5_ASAP7_75t_L g840 ( .A1(n_841), .A2(n_844), .B(n_847), .Y(n_840) );
INVx1_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
INVx2_ASAP7_75t_L g842 ( .A(n_843), .Y(n_842) );
INVx1_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
NOR2xp33_ASAP7_75t_L g850 ( .A(n_851), .B(n_852), .Y(n_850) );
INVx6_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
BUFx10_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
INVx1_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
INVx4_ASAP7_75t_SL g858 ( .A(n_859), .Y(n_858) );
endmodule