module fake_netlist_1_7619_n_725 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_725);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_725;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_560;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_695;
wire n_625;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVxp67_ASAP7_75t_L g80 ( .A(n_16), .Y(n_80) );
CKINVDCx16_ASAP7_75t_R g81 ( .A(n_44), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_20), .Y(n_82) );
HB1xp67_ASAP7_75t_L g83 ( .A(n_3), .Y(n_83) );
INVxp67_ASAP7_75t_SL g84 ( .A(n_77), .Y(n_84) );
HB1xp67_ASAP7_75t_L g85 ( .A(n_3), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_6), .Y(n_86) );
INVx1_ASAP7_75t_SL g87 ( .A(n_19), .Y(n_87) );
INVx2_ASAP7_75t_L g88 ( .A(n_72), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_59), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_65), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_41), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_53), .Y(n_92) );
CKINVDCx20_ASAP7_75t_R g93 ( .A(n_55), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_35), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_6), .Y(n_95) );
CKINVDCx14_ASAP7_75t_R g96 ( .A(n_18), .Y(n_96) );
CKINVDCx5p33_ASAP7_75t_R g97 ( .A(n_30), .Y(n_97) );
INVxp67_ASAP7_75t_SL g98 ( .A(n_9), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_26), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_75), .Y(n_100) );
INVxp67_ASAP7_75t_SL g101 ( .A(n_27), .Y(n_101) );
HB1xp67_ASAP7_75t_L g102 ( .A(n_36), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_73), .Y(n_103) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_13), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_79), .Y(n_105) );
INVxp67_ASAP7_75t_SL g106 ( .A(n_49), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_42), .Y(n_107) );
INVxp33_ASAP7_75t_SL g108 ( .A(n_10), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_74), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_69), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g111 ( .A(n_37), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_28), .Y(n_112) );
INVx2_ASAP7_75t_L g113 ( .A(n_17), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_8), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_5), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_12), .Y(n_116) );
INVxp67_ASAP7_75t_L g117 ( .A(n_56), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_40), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_58), .Y(n_119) );
INVxp67_ASAP7_75t_SL g120 ( .A(n_38), .Y(n_120) );
INVxp67_ASAP7_75t_L g121 ( .A(n_25), .Y(n_121) );
BUFx3_ASAP7_75t_L g122 ( .A(n_2), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_29), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_46), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_52), .Y(n_125) );
INVxp67_ASAP7_75t_SL g126 ( .A(n_76), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_23), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_10), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_122), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_102), .B(n_0), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_88), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_88), .Y(n_132) );
AND2x2_ASAP7_75t_L g133 ( .A(n_81), .B(n_0), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_122), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_122), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_86), .B(n_1), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_113), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_86), .B(n_1), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_88), .Y(n_139) );
AND2x2_ASAP7_75t_L g140 ( .A(n_81), .B(n_2), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_95), .B(n_4), .Y(n_141) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_123), .Y(n_142) );
BUFx3_ASAP7_75t_L g143 ( .A(n_123), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_123), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_113), .Y(n_145) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_125), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_113), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_95), .B(n_4), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_82), .Y(n_149) );
INVx2_ASAP7_75t_SL g150 ( .A(n_125), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_125), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_127), .Y(n_152) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_127), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_82), .Y(n_154) );
HB1xp67_ASAP7_75t_L g155 ( .A(n_83), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_89), .Y(n_156) );
INVx3_ASAP7_75t_L g157 ( .A(n_127), .Y(n_157) );
CKINVDCx5p33_ASAP7_75t_R g158 ( .A(n_93), .Y(n_158) );
INVx3_ASAP7_75t_L g159 ( .A(n_89), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_90), .Y(n_160) );
NAND2x1p5_ASAP7_75t_L g161 ( .A(n_90), .B(n_91), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_91), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_92), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_92), .Y(n_164) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_94), .Y(n_165) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_94), .Y(n_166) );
OA21x2_ASAP7_75t_L g167 ( .A1(n_99), .A2(n_39), .B(n_71), .Y(n_167) );
HB1xp67_ASAP7_75t_L g168 ( .A(n_85), .Y(n_168) );
OA21x2_ASAP7_75t_L g169 ( .A1(n_99), .A2(n_34), .B(n_70), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_100), .Y(n_170) );
AND2x2_ASAP7_75t_L g171 ( .A(n_96), .B(n_5), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_100), .Y(n_172) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_142), .Y(n_173) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_142), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_149), .B(n_97), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_142), .Y(n_176) );
AND2x2_ASAP7_75t_SL g177 ( .A(n_171), .B(n_105), .Y(n_177) );
HB1xp67_ASAP7_75t_L g178 ( .A(n_155), .Y(n_178) );
OAI22xp5_ASAP7_75t_L g179 ( .A1(n_168), .A2(n_114), .B1(n_115), .B2(n_116), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_149), .B(n_117), .Y(n_180) );
INVx3_ASAP7_75t_L g181 ( .A(n_165), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_161), .Y(n_182) );
INVx4_ASAP7_75t_L g183 ( .A(n_159), .Y(n_183) );
AND2x6_ASAP7_75t_L g184 ( .A(n_133), .B(n_109), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g185 ( .A(n_154), .B(n_121), .Y(n_185) );
BUFx3_ASAP7_75t_L g186 ( .A(n_129), .Y(n_186) );
INVx5_ASAP7_75t_L g187 ( .A(n_165), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_142), .Y(n_188) );
OR2x6_ASAP7_75t_L g189 ( .A(n_133), .B(n_114), .Y(n_189) );
INVx4_ASAP7_75t_L g190 ( .A(n_159), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_154), .B(n_107), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_156), .B(n_108), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_142), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_161), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_161), .Y(n_195) );
INVx3_ASAP7_75t_L g196 ( .A(n_165), .Y(n_196) );
INVxp67_ASAP7_75t_SL g197 ( .A(n_171), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_161), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_142), .Y(n_199) );
BUFx2_ASAP7_75t_L g200 ( .A(n_171), .Y(n_200) );
INVx8_ASAP7_75t_L g201 ( .A(n_133), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_150), .Y(n_202) );
OAI22xp33_ASAP7_75t_L g203 ( .A1(n_130), .A2(n_115), .B1(n_116), .B2(n_98), .Y(n_203) );
AO22x2_ASAP7_75t_L g204 ( .A1(n_140), .A2(n_109), .B1(n_103), .B2(n_124), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_165), .Y(n_205) );
AND2x2_ASAP7_75t_SL g206 ( .A(n_140), .B(n_110), .Y(n_206) );
INVx3_ASAP7_75t_L g207 ( .A(n_165), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_156), .B(n_80), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_150), .Y(n_209) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_159), .B(n_110), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_160), .B(n_112), .Y(n_211) );
INVx6_ASAP7_75t_L g212 ( .A(n_165), .Y(n_212) );
AND2x4_ASAP7_75t_L g213 ( .A(n_160), .B(n_124), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_165), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_150), .Y(n_215) );
AOI22xp33_ASAP7_75t_L g216 ( .A1(n_162), .A2(n_103), .B1(n_105), .B2(n_119), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_142), .Y(n_217) );
BUFx3_ASAP7_75t_L g218 ( .A(n_129), .Y(n_218) );
AND2x4_ASAP7_75t_L g219 ( .A(n_162), .B(n_112), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g220 ( .A(n_163), .B(n_118), .Y(n_220) );
AOI22xp33_ASAP7_75t_L g221 ( .A1(n_163), .A2(n_118), .B1(n_119), .B2(n_111), .Y(n_221) );
AND2x4_ASAP7_75t_L g222 ( .A(n_164), .B(n_84), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_159), .Y(n_223) );
INVx8_ASAP7_75t_L g224 ( .A(n_157), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_146), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_172), .Y(n_226) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_164), .B(n_87), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_170), .B(n_126), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_172), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_166), .Y(n_230) );
BUFx6f_ASAP7_75t_L g231 ( .A(n_146), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_166), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_146), .Y(n_233) );
BUFx3_ASAP7_75t_L g234 ( .A(n_134), .Y(n_234) );
INVx4_ASAP7_75t_L g235 ( .A(n_167), .Y(n_235) );
AND2x2_ASAP7_75t_L g236 ( .A(n_170), .B(n_120), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_172), .Y(n_237) );
INVx2_ASAP7_75t_L g238 ( .A(n_183), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_224), .Y(n_239) );
INVx2_ASAP7_75t_L g240 ( .A(n_183), .Y(n_240) );
BUFx6f_ASAP7_75t_L g241 ( .A(n_224), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_192), .B(n_130), .Y(n_242) );
BUFx3_ASAP7_75t_L g243 ( .A(n_224), .Y(n_243) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_222), .B(n_158), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_224), .Y(n_245) );
INVx2_ASAP7_75t_L g246 ( .A(n_183), .Y(n_246) );
AO22x1_ASAP7_75t_L g247 ( .A1(n_184), .A2(n_101), .B1(n_106), .B2(n_141), .Y(n_247) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_222), .B(n_136), .Y(n_248) );
INVx2_ASAP7_75t_L g249 ( .A(n_190), .Y(n_249) );
AND2x4_ASAP7_75t_L g250 ( .A(n_189), .B(n_148), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_190), .Y(n_251) );
HB1xp67_ASAP7_75t_L g252 ( .A(n_178), .Y(n_252) );
OAI22xp5_ASAP7_75t_L g253 ( .A1(n_206), .A2(n_136), .B1(n_138), .B2(n_141), .Y(n_253) );
INVx1_ASAP7_75t_SL g254 ( .A(n_200), .Y(n_254) );
BUFx2_ASAP7_75t_L g255 ( .A(n_201), .Y(n_255) );
AND2x4_ASAP7_75t_L g256 ( .A(n_189), .B(n_148), .Y(n_256) );
INVx1_ASAP7_75t_SL g257 ( .A(n_200), .Y(n_257) );
NAND2xp5_ASAP7_75t_SL g258 ( .A(n_182), .B(n_166), .Y(n_258) );
HB1xp67_ASAP7_75t_L g259 ( .A(n_189), .Y(n_259) );
INVx3_ASAP7_75t_L g260 ( .A(n_190), .Y(n_260) );
NAND2x1p5_ASAP7_75t_L g261 ( .A(n_194), .B(n_169), .Y(n_261) );
INVx2_ASAP7_75t_SL g262 ( .A(n_201), .Y(n_262) );
BUFx3_ASAP7_75t_L g263 ( .A(n_195), .Y(n_263) );
INVx2_ASAP7_75t_L g264 ( .A(n_223), .Y(n_264) );
OR2x6_ASAP7_75t_L g265 ( .A(n_201), .B(n_138), .Y(n_265) );
AND3x2_ASAP7_75t_SL g266 ( .A(n_201), .B(n_104), .C(n_128), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_202), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_226), .Y(n_268) );
INVx1_ASAP7_75t_SL g269 ( .A(n_189), .Y(n_269) );
AND2x2_ASAP7_75t_L g270 ( .A(n_197), .B(n_143), .Y(n_270) );
OR2x6_ASAP7_75t_L g271 ( .A(n_204), .B(n_143), .Y(n_271) );
HB1xp67_ASAP7_75t_L g272 ( .A(n_184), .Y(n_272) );
INVx5_ASAP7_75t_L g273 ( .A(n_212), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_222), .B(n_143), .Y(n_274) );
AOI21xp5_ASAP7_75t_L g275 ( .A1(n_198), .A2(n_169), .B(n_167), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_236), .B(n_213), .Y(n_276) );
AND2x4_ASAP7_75t_L g277 ( .A(n_236), .B(n_147), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_229), .Y(n_278) );
NOR2xp33_ASAP7_75t_L g279 ( .A(n_208), .B(n_135), .Y(n_279) );
NOR2xp33_ASAP7_75t_L g280 ( .A(n_227), .B(n_135), .Y(n_280) );
INVx2_ASAP7_75t_SL g281 ( .A(n_213), .Y(n_281) );
BUFx3_ASAP7_75t_L g282 ( .A(n_186), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_237), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_176), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_209), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_176), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_188), .Y(n_287) );
OR2x6_ASAP7_75t_L g288 ( .A(n_204), .B(n_169), .Y(n_288) );
NOR2xp33_ASAP7_75t_L g289 ( .A(n_227), .B(n_134), .Y(n_289) );
OAI22xp5_ASAP7_75t_L g290 ( .A1(n_206), .A2(n_157), .B1(n_132), .B2(n_139), .Y(n_290) );
AOI22xp33_ASAP7_75t_L g291 ( .A1(n_184), .A2(n_166), .B1(n_157), .B2(n_146), .Y(n_291) );
AND2x4_ASAP7_75t_SL g292 ( .A(n_221), .B(n_157), .Y(n_292) );
NAND3xp33_ASAP7_75t_L g293 ( .A(n_216), .B(n_169), .C(n_167), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_215), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_213), .Y(n_295) );
O2A1O1Ixp5_ASAP7_75t_L g296 ( .A1(n_235), .A2(n_131), .B(n_132), .C(n_144), .Y(n_296) );
AOI22xp33_ASAP7_75t_L g297 ( .A1(n_184), .A2(n_166), .B1(n_146), .B2(n_153), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_219), .Y(n_298) );
BUFx4f_ASAP7_75t_L g299 ( .A(n_184), .Y(n_299) );
OR2x4_ASAP7_75t_L g300 ( .A(n_180), .B(n_147), .Y(n_300) );
AND2x2_ASAP7_75t_L g301 ( .A(n_177), .B(n_145), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_219), .Y(n_302) );
BUFx6f_ASAP7_75t_L g303 ( .A(n_173), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_219), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_204), .Y(n_305) );
AND2x4_ASAP7_75t_L g306 ( .A(n_184), .B(n_145), .Y(n_306) );
BUFx6f_ASAP7_75t_L g307 ( .A(n_173), .Y(n_307) );
AND2x2_ASAP7_75t_L g308 ( .A(n_301), .B(n_177), .Y(n_308) );
BUFx12f_ASAP7_75t_L g309 ( .A(n_271), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_268), .Y(n_310) );
INVx4_ASAP7_75t_L g311 ( .A(n_241), .Y(n_311) );
INVxp67_ASAP7_75t_L g312 ( .A(n_252), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_268), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_278), .Y(n_314) );
CKINVDCx8_ASAP7_75t_R g315 ( .A(n_271), .Y(n_315) );
INVxp67_ASAP7_75t_SL g316 ( .A(n_263), .Y(n_316) );
INVxp67_ASAP7_75t_L g317 ( .A(n_254), .Y(n_317) );
AND2x2_ASAP7_75t_L g318 ( .A(n_301), .B(n_204), .Y(n_318) );
BUFx6f_ASAP7_75t_L g319 ( .A(n_241), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_278), .Y(n_320) );
INVx3_ASAP7_75t_L g321 ( .A(n_260), .Y(n_321) );
HB1xp67_ASAP7_75t_L g322 ( .A(n_271), .Y(n_322) );
AND2x6_ASAP7_75t_L g323 ( .A(n_269), .B(n_186), .Y(n_323) );
AND2x4_ASAP7_75t_L g324 ( .A(n_255), .B(n_228), .Y(n_324) );
OR2x2_ASAP7_75t_L g325 ( .A(n_257), .B(n_179), .Y(n_325) );
INVx4_ASAP7_75t_L g326 ( .A(n_241), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_283), .Y(n_327) );
BUFx3_ASAP7_75t_L g328 ( .A(n_241), .Y(n_328) );
BUFx6f_ASAP7_75t_L g329 ( .A(n_263), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_283), .Y(n_330) );
AOI21xp33_ASAP7_75t_L g331 ( .A1(n_262), .A2(n_244), .B(n_253), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_264), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_264), .Y(n_333) );
OR2x6_ASAP7_75t_L g334 ( .A(n_271), .B(n_211), .Y(n_334) );
OAI22xp5_ASAP7_75t_L g335 ( .A1(n_299), .A2(n_175), .B1(n_191), .B2(n_185), .Y(n_335) );
NOR3xp33_ASAP7_75t_L g336 ( .A(n_259), .B(n_203), .C(n_220), .Y(n_336) );
HB1xp67_ASAP7_75t_L g337 ( .A(n_255), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_260), .Y(n_338) );
BUFx2_ASAP7_75t_L g339 ( .A(n_243), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_250), .B(n_210), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_260), .Y(n_341) );
OAI21xp5_ASAP7_75t_L g342 ( .A1(n_296), .A2(n_235), .B(n_210), .Y(n_342) );
AOI221xp5_ASAP7_75t_L g343 ( .A1(n_242), .A2(n_248), .B1(n_276), .B2(n_277), .C(n_256), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_238), .Y(n_344) );
INVxp67_ASAP7_75t_SL g345 ( .A(n_243), .Y(n_345) );
BUFx3_ASAP7_75t_L g346 ( .A(n_299), .Y(n_346) );
BUFx6f_ASAP7_75t_L g347 ( .A(n_299), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_250), .B(n_218), .Y(n_348) );
BUFx12f_ASAP7_75t_L g349 ( .A(n_265), .Y(n_349) );
OR2x2_ASAP7_75t_L g350 ( .A(n_250), .B(n_218), .Y(n_350) );
AND2x2_ASAP7_75t_L g351 ( .A(n_256), .B(n_234), .Y(n_351) );
AND2x2_ASAP7_75t_SL g352 ( .A(n_305), .B(n_235), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_256), .B(n_234), .Y(n_353) );
CKINVDCx6p67_ASAP7_75t_R g354 ( .A(n_265), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_238), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_240), .Y(n_356) );
BUFx3_ASAP7_75t_L g357 ( .A(n_282), .Y(n_357) );
BUFx3_ASAP7_75t_L g358 ( .A(n_282), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_240), .Y(n_359) );
BUFx6f_ASAP7_75t_L g360 ( .A(n_246), .Y(n_360) );
O2A1O1Ixp33_ASAP7_75t_SL g361 ( .A1(n_258), .A2(n_232), .B(n_230), .C(n_205), .Y(n_361) );
OAI22xp5_ASAP7_75t_L g362 ( .A1(n_315), .A2(n_288), .B1(n_265), .B2(n_281), .Y(n_362) );
OAI22xp33_ASAP7_75t_SL g363 ( .A1(n_315), .A2(n_288), .B1(n_265), .B2(n_290), .Y(n_363) );
AOI221xp5_ASAP7_75t_L g364 ( .A1(n_343), .A2(n_277), .B1(n_279), .B2(n_292), .C(n_270), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_310), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_308), .B(n_270), .Y(n_366) );
OAI22xp5_ASAP7_75t_L g367 ( .A1(n_334), .A2(n_281), .B1(n_302), .B2(n_304), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_313), .Y(n_368) );
CKINVDCx20_ASAP7_75t_R g369 ( .A(n_317), .Y(n_369) );
INVx2_ASAP7_75t_SL g370 ( .A(n_309), .Y(n_370) );
BUFx2_ASAP7_75t_L g371 ( .A(n_309), .Y(n_371) );
INVx3_ASAP7_75t_L g372 ( .A(n_329), .Y(n_372) );
OA21x2_ASAP7_75t_L g373 ( .A1(n_342), .A2(n_275), .B(n_293), .Y(n_373) );
BUFx3_ASAP7_75t_L g374 ( .A(n_319), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_324), .B(n_277), .Y(n_375) );
AND2x2_ASAP7_75t_L g376 ( .A(n_308), .B(n_306), .Y(n_376) );
OR2x2_ASAP7_75t_L g377 ( .A(n_325), .B(n_274), .Y(n_377) );
BUFx6f_ASAP7_75t_L g378 ( .A(n_319), .Y(n_378) );
AOI22xp33_ASAP7_75t_L g379 ( .A1(n_318), .A2(n_306), .B1(n_292), .B2(n_272), .Y(n_379) );
A2O1A1Ixp33_ASAP7_75t_L g380 ( .A1(n_331), .A2(n_280), .B(n_289), .C(n_267), .Y(n_380) );
AOI22xp33_ASAP7_75t_L g381 ( .A1(n_318), .A2(n_306), .B1(n_262), .B2(n_298), .Y(n_381) );
OAI22xp5_ASAP7_75t_L g382 ( .A1(n_334), .A2(n_295), .B1(n_300), .B2(n_288), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_313), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_310), .Y(n_384) );
OAI22xp5_ASAP7_75t_L g385 ( .A1(n_334), .A2(n_288), .B1(n_300), .B2(n_261), .Y(n_385) );
INVx4_ASAP7_75t_L g386 ( .A(n_329), .Y(n_386) );
AOI22xp33_ASAP7_75t_L g387 ( .A1(n_325), .A2(n_245), .B1(n_239), .B2(n_251), .Y(n_387) );
INVx4_ASAP7_75t_L g388 ( .A(n_329), .Y(n_388) );
CKINVDCx20_ASAP7_75t_R g389 ( .A(n_312), .Y(n_389) );
OAI22x1_ASAP7_75t_L g390 ( .A1(n_322), .A2(n_266), .B1(n_261), .B2(n_167), .Y(n_390) );
OAI21x1_ASAP7_75t_L g391 ( .A1(n_313), .A2(n_261), .B(n_167), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_324), .B(n_246), .Y(n_392) );
AOI22xp33_ASAP7_75t_L g393 ( .A1(n_336), .A2(n_249), .B1(n_251), .B2(n_285), .Y(n_393) );
OAI22xp33_ASAP7_75t_L g394 ( .A1(n_334), .A2(n_300), .B1(n_266), .B2(n_294), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_314), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_365), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_365), .Y(n_397) );
NAND2x1_ASAP7_75t_L g398 ( .A(n_368), .B(n_330), .Y(n_398) );
AND2x4_ASAP7_75t_L g399 ( .A(n_376), .B(n_334), .Y(n_399) );
BUFx6f_ASAP7_75t_L g400 ( .A(n_378), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_366), .B(n_324), .Y(n_401) );
AOI21xp5_ASAP7_75t_L g402 ( .A1(n_380), .A2(n_316), .B(n_361), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_384), .Y(n_403) );
BUFx2_ASAP7_75t_L g404 ( .A(n_369), .Y(n_404) );
OAI221xp5_ASAP7_75t_L g405 ( .A1(n_364), .A2(n_337), .B1(n_335), .B2(n_350), .C(n_353), .Y(n_405) );
OAI211xp5_ASAP7_75t_L g406 ( .A1(n_387), .A2(n_137), .B(n_291), .C(n_297), .Y(n_406) );
AOI221xp5_ASAP7_75t_L g407 ( .A1(n_394), .A2(n_375), .B1(n_366), .B2(n_377), .C(n_363), .Y(n_407) );
AOI221xp5_ASAP7_75t_L g408 ( .A1(n_377), .A2(n_324), .B1(n_137), .B2(n_340), .C(n_247), .Y(n_408) );
OAI221xp5_ASAP7_75t_L g409 ( .A1(n_381), .A2(n_350), .B1(n_314), .B2(n_320), .C(n_327), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_384), .Y(n_410) );
AOI22xp33_ASAP7_75t_L g411 ( .A1(n_362), .A2(n_349), .B1(n_354), .B2(n_352), .Y(n_411) );
AOI22xp33_ASAP7_75t_L g412 ( .A1(n_362), .A2(n_349), .B1(n_354), .B2(n_352), .Y(n_412) );
INVx5_ASAP7_75t_L g413 ( .A(n_378), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_395), .Y(n_414) );
AOI22xp5_ASAP7_75t_L g415 ( .A1(n_389), .A2(n_348), .B1(n_351), .B2(n_340), .Y(n_415) );
AND2x4_ASAP7_75t_L g416 ( .A(n_376), .B(n_348), .Y(n_416) );
OAI22xp5_ASAP7_75t_L g417 ( .A1(n_379), .A2(n_327), .B1(n_320), .B2(n_333), .Y(n_417) );
AOI22xp33_ASAP7_75t_L g418 ( .A1(n_363), .A2(n_352), .B1(n_351), .B2(n_323), .Y(n_418) );
AO21x2_ASAP7_75t_L g419 ( .A1(n_391), .A2(n_332), .B(n_333), .Y(n_419) );
OAI22xp5_ASAP7_75t_L g420 ( .A1(n_385), .A2(n_332), .B1(n_330), .B2(n_329), .Y(n_420) );
OAI22xp33_ASAP7_75t_L g421 ( .A1(n_371), .A2(n_385), .B1(n_370), .B2(n_382), .Y(n_421) );
AOI22xp33_ASAP7_75t_SL g422 ( .A1(n_371), .A2(n_323), .B1(n_339), .B2(n_329), .Y(n_422) );
OAI221xp5_ASAP7_75t_L g423 ( .A1(n_393), .A2(n_330), .B1(n_339), .B2(n_345), .C(n_131), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_392), .B(n_359), .Y(n_424) );
OAI21x1_ASAP7_75t_L g425 ( .A1(n_402), .A2(n_391), .B(n_373), .Y(n_425) );
NAND3xp33_ASAP7_75t_L g426 ( .A(n_407), .B(n_368), .C(n_383), .Y(n_426) );
OAI221xp5_ASAP7_75t_L g427 ( .A1(n_415), .A2(n_370), .B1(n_367), .B2(n_395), .C(n_132), .Y(n_427) );
OAI31xp33_ASAP7_75t_L g428 ( .A1(n_409), .A2(n_392), .A3(n_383), .B(n_368), .Y(n_428) );
OAI222xp33_ASAP7_75t_L g429 ( .A1(n_421), .A2(n_383), .B1(n_388), .B2(n_386), .C1(n_390), .C2(n_372), .Y(n_429) );
OAI21xp33_ASAP7_75t_L g430 ( .A1(n_409), .A2(n_390), .B(n_131), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_424), .B(n_386), .Y(n_431) );
NAND4xp25_ASAP7_75t_SL g432 ( .A(n_411), .B(n_139), .C(n_144), .D(n_151), .Y(n_432) );
OA21x2_ASAP7_75t_L g433 ( .A1(n_420), .A2(n_152), .B(n_151), .Y(n_433) );
BUFx2_ASAP7_75t_SL g434 ( .A(n_413), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_396), .B(n_386), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_397), .B(n_373), .Y(n_436) );
NOR2xp33_ASAP7_75t_L g437 ( .A(n_404), .B(n_311), .Y(n_437) );
NAND3xp33_ASAP7_75t_L g438 ( .A(n_418), .B(n_373), .C(n_146), .Y(n_438) );
INVxp67_ASAP7_75t_L g439 ( .A(n_401), .Y(n_439) );
OAI21xp5_ASAP7_75t_L g440 ( .A1(n_405), .A2(n_373), .B(n_344), .Y(n_440) );
A2O1A1Ixp33_ASAP7_75t_L g441 ( .A1(n_412), .A2(n_328), .B(n_357), .C(n_358), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_403), .B(n_386), .Y(n_442) );
AOI22xp33_ASAP7_75t_L g443 ( .A1(n_405), .A2(n_323), .B1(n_357), .B2(n_358), .Y(n_443) );
AOI221x1_ASAP7_75t_SL g444 ( .A1(n_410), .A2(n_139), .B1(n_144), .B2(n_151), .C(n_152), .Y(n_444) );
OAI22xp5_ASAP7_75t_L g445 ( .A1(n_423), .A2(n_388), .B1(n_374), .B2(n_357), .Y(n_445) );
AOI22xp33_ASAP7_75t_L g446 ( .A1(n_399), .A2(n_323), .B1(n_358), .B2(n_388), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_419), .Y(n_447) );
OAI211xp5_ASAP7_75t_SL g448 ( .A1(n_408), .A2(n_152), .B(n_258), .C(n_230), .Y(n_448) );
OAI33xp33_ASAP7_75t_L g449 ( .A1(n_417), .A2(n_232), .A3(n_214), .B1(n_205), .B2(n_338), .B3(n_341), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_414), .B(n_388), .Y(n_450) );
OAI211xp5_ASAP7_75t_L g451 ( .A1(n_408), .A2(n_169), .B(n_166), .C(n_153), .Y(n_451) );
OAI221xp5_ASAP7_75t_L g452 ( .A1(n_423), .A2(n_341), .B1(n_338), .B2(n_166), .C(n_321), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_399), .B(n_372), .Y(n_453) );
HB1xp67_ASAP7_75t_L g454 ( .A(n_416), .Y(n_454) );
AOI22xp33_ASAP7_75t_L g455 ( .A1(n_416), .A2(n_323), .B1(n_321), .B2(n_311), .Y(n_455) );
AOI221xp5_ASAP7_75t_L g456 ( .A1(n_422), .A2(n_146), .B1(n_153), .B2(n_344), .C(n_359), .Y(n_456) );
INVx1_ASAP7_75t_SL g457 ( .A(n_413), .Y(n_457) );
AOI22xp33_ASAP7_75t_L g458 ( .A1(n_398), .A2(n_323), .B1(n_321), .B2(n_326), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_413), .B(n_372), .Y(n_459) );
NOR3xp33_ASAP7_75t_L g460 ( .A(n_406), .B(n_326), .C(n_311), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_436), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_447), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_436), .Y(n_463) );
INVx4_ASAP7_75t_L g464 ( .A(n_459), .Y(n_464) );
OR2x2_ASAP7_75t_L g465 ( .A(n_431), .B(n_419), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_431), .B(n_413), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_447), .Y(n_467) );
AO21x2_ASAP7_75t_L g468 ( .A1(n_430), .A2(n_233), .B(n_225), .Y(n_468) );
NOR3xp33_ASAP7_75t_L g469 ( .A(n_437), .B(n_311), .C(n_326), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_447), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_435), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_425), .Y(n_472) );
INVx2_ASAP7_75t_SL g473 ( .A(n_457), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_439), .B(n_372), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_435), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_454), .B(n_442), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_442), .Y(n_477) );
HB1xp67_ASAP7_75t_L g478 ( .A(n_450), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_450), .B(n_323), .Y(n_479) );
INVx5_ASAP7_75t_SL g480 ( .A(n_434), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_425), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_453), .B(n_153), .Y(n_482) );
NAND3xp33_ASAP7_75t_L g483 ( .A(n_438), .B(n_153), .C(n_231), .Y(n_483) );
BUFx8_ASAP7_75t_L g484 ( .A(n_459), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_433), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_440), .Y(n_486) );
AND2x4_ASAP7_75t_L g487 ( .A(n_457), .B(n_400), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_440), .B(n_374), .Y(n_488) );
OAI33xp33_ASAP7_75t_L g489 ( .A1(n_430), .A2(n_214), .A3(n_8), .B1(n_9), .B2(n_11), .B3(n_12), .Y(n_489) );
INVx1_ASAP7_75t_SL g490 ( .A(n_434), .Y(n_490) );
AND2x4_ASAP7_75t_SL g491 ( .A(n_453), .B(n_326), .Y(n_491) );
OAI221xp5_ASAP7_75t_L g492 ( .A1(n_444), .A2(n_153), .B1(n_374), .B2(n_321), .C(n_328), .Y(n_492) );
OR2x2_ASAP7_75t_L g493 ( .A(n_428), .B(n_400), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_433), .Y(n_494) );
OAI31xp33_ASAP7_75t_L g495 ( .A1(n_428), .A2(n_328), .A3(n_359), .B(n_355), .Y(n_495) );
OR2x2_ASAP7_75t_L g496 ( .A(n_426), .B(n_438), .Y(n_496) );
INVx2_ASAP7_75t_L g497 ( .A(n_433), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_426), .Y(n_498) );
AOI211xp5_ASAP7_75t_L g499 ( .A1(n_432), .A2(n_153), .B(n_319), .C(n_378), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_433), .B(n_400), .Y(n_500) );
OAI33xp33_ASAP7_75t_L g501 ( .A1(n_445), .A2(n_7), .A3(n_11), .B1(n_13), .B2(n_14), .B3(n_15), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_444), .Y(n_502) );
OAI31xp33_ASAP7_75t_L g503 ( .A1(n_427), .A2(n_355), .A3(n_356), .B(n_346), .Y(n_503) );
INVxp67_ASAP7_75t_SL g504 ( .A(n_445), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_443), .B(n_378), .Y(n_505) );
INVx2_ASAP7_75t_L g506 ( .A(n_452), .Y(n_506) );
INVx1_ASAP7_75t_SL g507 ( .A(n_432), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_451), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_460), .Y(n_509) );
INVx2_ASAP7_75t_L g510 ( .A(n_429), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_458), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_446), .B(n_378), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_466), .B(n_7), .Y(n_513) );
NAND2xp5_ASAP7_75t_SL g514 ( .A(n_499), .B(n_456), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_462), .Y(n_515) );
NAND2xp33_ASAP7_75t_L g516 ( .A(n_490), .B(n_455), .Y(n_516) );
OR2x2_ASAP7_75t_SL g517 ( .A(n_478), .B(n_378), .Y(n_517) );
OR2x2_ASAP7_75t_L g518 ( .A(n_471), .B(n_14), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_462), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_466), .B(n_15), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_471), .Y(n_521) );
NAND2xp5_ASAP7_75t_SL g522 ( .A(n_499), .B(n_441), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_475), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_475), .B(n_16), .Y(n_524) );
AND2x4_ASAP7_75t_L g525 ( .A(n_464), .B(n_17), .Y(n_525) );
A2O1A1Ixp33_ASAP7_75t_L g526 ( .A1(n_495), .A2(n_448), .B(n_449), .C(n_346), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_477), .B(n_18), .Y(n_527) );
OR2x2_ASAP7_75t_L g528 ( .A(n_477), .B(n_356), .Y(n_528) );
NAND4xp25_ASAP7_75t_L g529 ( .A(n_476), .B(n_199), .C(n_233), .D(n_193), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_502), .B(n_360), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_464), .B(n_319), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_465), .Y(n_532) );
OR2x2_ASAP7_75t_L g533 ( .A(n_465), .B(n_319), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_502), .B(n_360), .Y(n_534) );
NOR3xp33_ASAP7_75t_L g535 ( .A(n_501), .B(n_193), .C(n_225), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_461), .Y(n_536) );
AOI221xp5_ASAP7_75t_L g537 ( .A1(n_489), .A2(n_181), .B1(n_196), .B2(n_207), .C(n_173), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_461), .Y(n_538) );
INVx2_ASAP7_75t_L g539 ( .A(n_467), .Y(n_539) );
OAI221xp5_ASAP7_75t_L g540 ( .A1(n_507), .A2(n_188), .B1(n_199), .B2(n_217), .C(n_173), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_463), .Y(n_541) );
INVx1_ASAP7_75t_SL g542 ( .A(n_491), .Y(n_542) );
OR2x6_ASAP7_75t_SL g543 ( .A(n_480), .B(n_217), .Y(n_543) );
NAND3xp33_ASAP7_75t_SL g544 ( .A(n_503), .B(n_21), .C(n_22), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_464), .B(n_24), .Y(n_545) );
INVx2_ASAP7_75t_L g546 ( .A(n_467), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_463), .B(n_360), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_474), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_473), .Y(n_549) );
NAND2xp5_ASAP7_75t_SL g550 ( .A(n_495), .B(n_347), .Y(n_550) );
AOI221xp5_ASAP7_75t_L g551 ( .A1(n_482), .A2(n_511), .B1(n_498), .B2(n_486), .C(n_508), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_473), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_470), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_470), .Y(n_554) );
AND2x4_ASAP7_75t_L g555 ( .A(n_488), .B(n_31), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_491), .B(n_32), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_479), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_511), .B(n_360), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_509), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_509), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_493), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_493), .Y(n_562) );
INVx1_ASAP7_75t_SL g563 ( .A(n_487), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_510), .B(n_33), .Y(n_564) );
NAND4xp25_ASAP7_75t_L g565 ( .A(n_503), .B(n_196), .C(n_181), .D(n_207), .Y(n_565) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_510), .B(n_43), .Y(n_566) );
NAND2xp33_ASAP7_75t_SL g567 ( .A(n_480), .B(n_347), .Y(n_567) );
INVx3_ASAP7_75t_L g568 ( .A(n_480), .Y(n_568) );
INVx2_ASAP7_75t_L g569 ( .A(n_485), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_484), .Y(n_570) );
NOR3xp33_ASAP7_75t_L g571 ( .A(n_492), .B(n_181), .C(n_207), .Y(n_571) );
INVx1_ASAP7_75t_SL g572 ( .A(n_487), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_536), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_548), .B(n_486), .Y(n_574) );
NAND2x1p5_ASAP7_75t_L g575 ( .A(n_525), .B(n_480), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_559), .B(n_498), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_532), .B(n_504), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_538), .Y(n_578) );
NAND3xp33_ASAP7_75t_L g579 ( .A(n_560), .B(n_508), .C(n_469), .Y(n_579) );
INVx2_ASAP7_75t_L g580 ( .A(n_569), .Y(n_580) );
AND2x4_ASAP7_75t_L g581 ( .A(n_561), .B(n_488), .Y(n_581) );
INVx2_ASAP7_75t_L g582 ( .A(n_569), .Y(n_582) );
OAI21xp33_ASAP7_75t_L g583 ( .A1(n_566), .A2(n_496), .B(n_506), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_562), .B(n_485), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_521), .B(n_506), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_523), .B(n_541), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_515), .B(n_494), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_557), .B(n_496), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_551), .B(n_484), .Y(n_589) );
INVxp33_ASAP7_75t_L g590 ( .A(n_525), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_549), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_552), .B(n_484), .Y(n_592) );
INVxp67_ASAP7_75t_L g593 ( .A(n_543), .Y(n_593) );
OAI31xp33_ASAP7_75t_L g594 ( .A1(n_522), .A2(n_483), .A3(n_500), .B(n_487), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_530), .B(n_484), .Y(n_595) );
OR2x2_ASAP7_75t_L g596 ( .A(n_517), .B(n_497), .Y(n_596) );
INVxp67_ASAP7_75t_L g597 ( .A(n_566), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_534), .Y(n_598) );
AND2x2_ASAP7_75t_L g599 ( .A(n_515), .B(n_497), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_513), .B(n_487), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_553), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_554), .Y(n_602) );
AOI21xp5_ASAP7_75t_L g603 ( .A1(n_522), .A2(n_483), .B(n_494), .Y(n_603) );
OR2x2_ASAP7_75t_L g604 ( .A(n_533), .B(n_472), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_519), .Y(n_605) );
OAI322xp33_ASAP7_75t_L g606 ( .A1(n_518), .A2(n_472), .A3(n_481), .B1(n_505), .B2(n_500), .C1(n_512), .C2(n_231), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_519), .Y(n_607) );
AND2x2_ASAP7_75t_L g608 ( .A(n_539), .B(n_481), .Y(n_608) );
NOR3xp33_ASAP7_75t_L g609 ( .A(n_544), .B(n_512), .C(n_505), .Y(n_609) );
AND2x2_ASAP7_75t_L g610 ( .A(n_539), .B(n_546), .Y(n_610) );
HB1xp67_ASAP7_75t_L g611 ( .A(n_542), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_546), .B(n_468), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_520), .B(n_468), .Y(n_613) );
NOR2x1p5_ASAP7_75t_L g614 ( .A(n_568), .B(n_346), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_528), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_558), .Y(n_616) );
OAI21x1_ASAP7_75t_SL g617 ( .A1(n_570), .A2(n_468), .B(n_47), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_524), .Y(n_618) );
OAI222xp33_ASAP7_75t_L g619 ( .A1(n_514), .A2(n_187), .B1(n_48), .B2(n_50), .C1(n_51), .C2(n_54), .Y(n_619) );
INVx2_ASAP7_75t_L g620 ( .A(n_547), .Y(n_620) );
NOR2x1_ASAP7_75t_SL g621 ( .A(n_545), .B(n_347), .Y(n_621) );
INVxp67_ASAP7_75t_L g622 ( .A(n_564), .Y(n_622) );
AND2x2_ASAP7_75t_L g623 ( .A(n_563), .B(n_231), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_527), .B(n_231), .Y(n_624) );
AND2x2_ASAP7_75t_L g625 ( .A(n_572), .B(n_231), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_555), .B(n_174), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_598), .B(n_577), .Y(n_627) );
NAND4xp25_ASAP7_75t_L g628 ( .A(n_589), .B(n_544), .C(n_555), .D(n_571), .Y(n_628) );
OR2x2_ASAP7_75t_L g629 ( .A(n_588), .B(n_577), .Y(n_629) );
XNOR2x1_ASAP7_75t_L g630 ( .A(n_575), .B(n_556), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_586), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_586), .B(n_516), .Y(n_632) );
INVx2_ASAP7_75t_L g633 ( .A(n_580), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_618), .B(n_531), .Y(n_634) );
NAND2xp5_ASAP7_75t_SL g635 ( .A(n_596), .B(n_567), .Y(n_635) );
AOI21xp33_ASAP7_75t_SL g636 ( .A1(n_593), .A2(n_514), .B(n_568), .Y(n_636) );
NOR2xp33_ASAP7_75t_L g637 ( .A(n_597), .B(n_529), .Y(n_637) );
NAND3xp33_ASAP7_75t_L g638 ( .A(n_594), .B(n_537), .C(n_571), .Y(n_638) );
AND2x2_ASAP7_75t_L g639 ( .A(n_581), .B(n_550), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_622), .B(n_526), .Y(n_640) );
AND2x2_ASAP7_75t_L g641 ( .A(n_584), .B(n_550), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_573), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_615), .B(n_526), .Y(n_643) );
NOR2xp33_ASAP7_75t_L g644 ( .A(n_611), .B(n_540), .Y(n_644) );
OR2x2_ASAP7_75t_L g645 ( .A(n_581), .B(n_567), .Y(n_645) );
NOR2xp33_ASAP7_75t_L g646 ( .A(n_590), .B(n_565), .Y(n_646) );
INVx2_ASAP7_75t_L g647 ( .A(n_580), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_591), .B(n_535), .Y(n_648) );
AOI21xp33_ASAP7_75t_L g649 ( .A1(n_590), .A2(n_174), .B(n_173), .Y(n_649) );
AND2x2_ASAP7_75t_L g650 ( .A(n_581), .B(n_535), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_578), .Y(n_651) );
AND2x4_ASAP7_75t_SL g652 ( .A(n_584), .B(n_360), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_601), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_602), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_576), .Y(n_655) );
NAND4xp75_ASAP7_75t_L g656 ( .A(n_595), .B(n_45), .C(n_57), .D(n_60), .Y(n_656) );
INVx2_ASAP7_75t_L g657 ( .A(n_582), .Y(n_657) );
NAND2xp5_ASAP7_75t_SL g658 ( .A(n_596), .B(n_174), .Y(n_658) );
AOI22xp33_ASAP7_75t_L g659 ( .A1(n_609), .A2(n_174), .B1(n_212), .B2(n_347), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_574), .B(n_174), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_585), .Y(n_661) );
OAI21xp5_ASAP7_75t_L g662 ( .A1(n_579), .A2(n_187), .B(n_196), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_616), .B(n_61), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_620), .B(n_62), .Y(n_664) );
OAI22xp5_ASAP7_75t_SL g665 ( .A1(n_575), .A2(n_592), .B1(n_600), .B2(n_621), .Y(n_665) );
INVx2_ASAP7_75t_L g666 ( .A(n_582), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_620), .B(n_63), .Y(n_667) );
INVx3_ASAP7_75t_L g668 ( .A(n_575), .Y(n_668) );
OAI21xp5_ASAP7_75t_SL g669 ( .A1(n_619), .A2(n_347), .B(n_66), .Y(n_669) );
XOR2xp5_ASAP7_75t_L g670 ( .A(n_621), .B(n_64), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_610), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_610), .Y(n_672) );
AOI22xp5_ASAP7_75t_L g673 ( .A1(n_583), .A2(n_212), .B1(n_187), .B2(n_307), .Y(n_673) );
NAND4xp25_ASAP7_75t_L g674 ( .A(n_603), .B(n_286), .C(n_284), .D(n_287), .Y(n_674) );
OAI21xp5_ASAP7_75t_L g675 ( .A1(n_626), .A2(n_187), .B(n_249), .Y(n_675) );
AOI22xp5_ASAP7_75t_L g676 ( .A1(n_613), .A2(n_212), .B1(n_187), .B2(n_307), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_587), .B(n_599), .Y(n_677) );
OAI21xp33_ASAP7_75t_L g678 ( .A1(n_604), .A2(n_67), .B(n_68), .Y(n_678) );
OAI211xp5_ASAP7_75t_L g679 ( .A1(n_626), .A2(n_78), .B(n_273), .C(n_284), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_605), .Y(n_680) );
AND2x2_ASAP7_75t_L g681 ( .A(n_587), .B(n_273), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_599), .B(n_286), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_607), .B(n_287), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_608), .B(n_273), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_608), .Y(n_685) );
NOR3xp33_ASAP7_75t_L g686 ( .A(n_624), .B(n_273), .C(n_303), .Y(n_686) );
AOI22xp5_ASAP7_75t_L g687 ( .A1(n_614), .A2(n_303), .B1(n_307), .B2(n_273), .Y(n_687) );
XOR2xp5_ASAP7_75t_L g688 ( .A(n_604), .B(n_623), .Y(n_688) );
AOI22xp5_ASAP7_75t_L g689 ( .A1(n_646), .A2(n_637), .B1(n_628), .B2(n_640), .Y(n_689) );
AOI22xp5_ASAP7_75t_L g690 ( .A1(n_646), .A2(n_637), .B1(n_669), .B2(n_650), .Y(n_690) );
INVx2_ASAP7_75t_L g691 ( .A(n_633), .Y(n_691) );
OAI22xp5_ASAP7_75t_L g692 ( .A1(n_630), .A2(n_665), .B1(n_668), .B2(n_669), .Y(n_692) );
AOI22xp5_ASAP7_75t_L g693 ( .A1(n_639), .A2(n_630), .B1(n_644), .B2(n_632), .Y(n_693) );
AOI222xp33_ASAP7_75t_L g694 ( .A1(n_638), .A2(n_643), .B1(n_661), .B2(n_655), .C1(n_634), .C2(n_635), .Y(n_694) );
AOI221xp5_ASAP7_75t_L g695 ( .A1(n_636), .A2(n_642), .B1(n_651), .B2(n_631), .C(n_627), .Y(n_695) );
NOR2x1_ASAP7_75t_L g696 ( .A(n_635), .B(n_668), .Y(n_696) );
OAI211xp5_ASAP7_75t_L g697 ( .A1(n_659), .A2(n_644), .B(n_658), .C(n_670), .Y(n_697) );
AOI22xp5_ASAP7_75t_L g698 ( .A1(n_641), .A2(n_688), .B1(n_648), .B2(n_671), .Y(n_698) );
AOI222xp33_ASAP7_75t_L g699 ( .A1(n_641), .A2(n_653), .B1(n_654), .B2(n_672), .C1(n_685), .C2(n_680), .Y(n_699) );
AOI21xp5_ASAP7_75t_L g700 ( .A1(n_658), .A2(n_662), .B(n_679), .Y(n_700) );
NAND2xp33_ASAP7_75t_SL g701 ( .A(n_645), .B(n_659), .Y(n_701) );
AOI22xp5_ASAP7_75t_L g702 ( .A1(n_629), .A2(n_677), .B1(n_652), .B2(n_681), .Y(n_702) );
NAND2x1_ASAP7_75t_L g703 ( .A(n_696), .B(n_617), .Y(n_703) );
NAND4xp25_ASAP7_75t_L g704 ( .A(n_692), .B(n_673), .C(n_678), .D(n_687), .Y(n_704) );
HB1xp67_ASAP7_75t_L g705 ( .A(n_691), .Y(n_705) );
NOR4xp25_ASAP7_75t_L g706 ( .A(n_695), .B(n_663), .C(n_674), .D(n_684), .Y(n_706) );
AOI221xp5_ASAP7_75t_L g707 ( .A1(n_701), .A2(n_606), .B1(n_649), .B2(n_657), .C(n_647), .Y(n_707) );
NAND3xp33_ASAP7_75t_SL g708 ( .A(n_690), .B(n_686), .C(n_675), .Y(n_708) );
OAI221xp5_ASAP7_75t_L g709 ( .A1(n_689), .A2(n_674), .B1(n_676), .B2(n_647), .C(n_657), .Y(n_709) );
OAI221xp5_ASAP7_75t_L g710 ( .A1(n_693), .A2(n_633), .B1(n_666), .B2(n_667), .C(n_664), .Y(n_710) );
OAI22xp5_ASAP7_75t_L g711 ( .A1(n_703), .A2(n_698), .B1(n_702), .B2(n_697), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_705), .Y(n_712) );
NOR3xp33_ASAP7_75t_L g713 ( .A(n_708), .B(n_656), .C(n_700), .Y(n_713) );
AOI22xp5_ASAP7_75t_L g714 ( .A1(n_704), .A2(n_694), .B1(n_699), .B2(n_652), .Y(n_714) );
CKINVDCx20_ASAP7_75t_R g715 ( .A(n_706), .Y(n_715) );
NOR3xp33_ASAP7_75t_L g716 ( .A(n_713), .B(n_709), .C(n_710), .Y(n_716) );
OA22x2_ASAP7_75t_L g717 ( .A1(n_714), .A2(n_617), .B1(n_707), .B2(n_682), .Y(n_717) );
NAND3xp33_ASAP7_75t_L g718 ( .A(n_715), .B(n_660), .C(n_683), .Y(n_718) );
NAND3xp33_ASAP7_75t_SL g719 ( .A(n_716), .B(n_711), .C(n_712), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_718), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_720), .B(n_717), .Y(n_721) );
OAI22x1_ASAP7_75t_L g722 ( .A1(n_719), .A2(n_625), .B1(n_623), .B2(n_612), .Y(n_722) );
OR2x6_ASAP7_75t_L g723 ( .A(n_721), .B(n_625), .Y(n_723) );
AOI22xp5_ASAP7_75t_SL g724 ( .A1(n_723), .A2(n_722), .B1(n_612), .B2(n_307), .Y(n_724) );
AOI221xp5_ASAP7_75t_L g725 ( .A1(n_724), .A2(n_303), .B1(n_307), .B2(n_719), .C(n_721), .Y(n_725) );
endmodule