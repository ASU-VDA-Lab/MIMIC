module fake_ariane_683_n_1690 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_1690);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1690;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_1654;
wire n_1560;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_155;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_727;
wire n_590;
wire n_699;
wire n_301;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_211;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_640;
wire n_197;
wire n_463;
wire n_1476;
wire n_1524;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_154;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_571;
wire n_414;
wire n_1521;
wire n_284;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_443;
wire n_1412;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1323;
wire n_1235;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_153;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1670;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_156;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_121),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_115),
.Y(n_154)
);

BUFx10_ASAP7_75t_L g155 ( 
.A(n_64),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_86),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_40),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_23),
.Y(n_158)
);

BUFx2_ASAP7_75t_L g159 ( 
.A(n_96),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_39),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_53),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_132),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_81),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_57),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_83),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_54),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_44),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_26),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_16),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_133),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_88),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_5),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_143),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_106),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_140),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_144),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_53),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_32),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_55),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_39),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_142),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_79),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_120),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_21),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_6),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_119),
.Y(n_186)
);

BUFx5_ASAP7_75t_L g187 ( 
.A(n_73),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_23),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_55),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_8),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_18),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_12),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_90),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_68),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_59),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_125),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_93),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_74),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_148),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_110),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_10),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_139),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_114),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_40),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_138),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_62),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_50),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_63),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_99),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_17),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_60),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_108),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_152),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_145),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_147),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_7),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_35),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_80),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_28),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_67),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_75),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_17),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_12),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_92),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_109),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_137),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_19),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_102),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_48),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_127),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_58),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_2),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_18),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_4),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_69),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_6),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g237 ( 
.A(n_76),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_130),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_59),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_26),
.Y(n_240)
);

INVx2_ASAP7_75t_SL g241 ( 
.A(n_27),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_89),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_103),
.Y(n_243)
);

BUFx10_ASAP7_75t_L g244 ( 
.A(n_111),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_0),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_151),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_27),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_33),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_126),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_129),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_49),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_113),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_77),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_51),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_134),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_112),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_131),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_29),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_85),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_149),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_50),
.Y(n_261)
);

BUFx10_ASAP7_75t_L g262 ( 
.A(n_14),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_48),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_3),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_38),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_100),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_118),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_37),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_46),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_14),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_28),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_38),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_34),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_32),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_34),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_54),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_42),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_49),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_47),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_33),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_52),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_71),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_56),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_136),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_31),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_51),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_122),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_41),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_21),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_95),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_41),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_56),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_47),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_7),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_36),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_61),
.Y(n_296)
);

INVx1_ASAP7_75t_SL g297 ( 
.A(n_37),
.Y(n_297)
);

BUFx3_ASAP7_75t_L g298 ( 
.A(n_25),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_1),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_87),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_52),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_19),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_185),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_194),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_169),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_185),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_178),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_159),
.B(n_0),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_185),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_185),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_185),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_202),
.Y(n_312)
);

INVxp67_ASAP7_75t_SL g313 ( 
.A(n_233),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_218),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_273),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_273),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_273),
.Y(n_317)
);

INVxp33_ASAP7_75t_L g318 ( 
.A(n_158),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_273),
.Y(n_319)
);

BUFx2_ASAP7_75t_L g320 ( 
.A(n_233),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_273),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_246),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_277),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_267),
.Y(n_324)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_193),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_241),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_287),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_277),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_300),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_219),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_184),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_270),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_188),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_189),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_277),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_277),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_277),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_190),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_241),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_157),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_295),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_271),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_154),
.B(n_1),
.Y(n_343)
);

INVx1_ASAP7_75t_SL g344 ( 
.A(n_289),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_295),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_191),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_295),
.Y(n_347)
);

INVxp67_ASAP7_75t_SL g348 ( 
.A(n_298),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_295),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_291),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_298),
.B(n_2),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_295),
.Y(n_352)
);

BUFx2_ASAP7_75t_L g353 ( 
.A(n_157),
.Y(n_353)
);

CKINVDCx16_ASAP7_75t_R g354 ( 
.A(n_282),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_192),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_187),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_299),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_294),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_207),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_262),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_155),
.Y(n_361)
);

CKINVDCx16_ASAP7_75t_R g362 ( 
.A(n_155),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_217),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_155),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_294),
.Y(n_365)
);

NOR2xp67_ASAP7_75t_L g366 ( 
.A(n_166),
.B(n_3),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_213),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_227),
.Y(n_368)
);

INVxp67_ASAP7_75t_SL g369 ( 
.A(n_172),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_213),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_244),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_259),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_231),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_232),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_244),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_187),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_162),
.B(n_4),
.Y(n_377)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_320),
.B(n_244),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_356),
.Y(n_379)
);

AND2x4_ASAP7_75t_L g380 ( 
.A(n_367),
.B(n_214),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_356),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_356),
.Y(n_382)
);

AND2x4_ASAP7_75t_L g383 ( 
.A(n_367),
.B(n_214),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_376),
.Y(n_384)
);

AND2x2_ASAP7_75t_SL g385 ( 
.A(n_308),
.B(n_259),
.Y(n_385)
);

AND2x4_ASAP7_75t_L g386 ( 
.A(n_370),
.B(n_237),
.Y(n_386)
);

AND3x2_ASAP7_75t_L g387 ( 
.A(n_360),
.B(n_236),
.C(n_170),
.Y(n_387)
);

AND2x4_ASAP7_75t_L g388 ( 
.A(n_370),
.B(n_237),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_376),
.Y(n_389)
);

BUFx2_ASAP7_75t_L g390 ( 
.A(n_305),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_320),
.B(n_180),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_376),
.Y(n_392)
);

CKINVDCx11_ASAP7_75t_R g393 ( 
.A(n_330),
.Y(n_393)
);

HB1xp67_ASAP7_75t_L g394 ( 
.A(n_353),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_372),
.B(n_165),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_317),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_317),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_317),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_303),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_303),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_306),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_306),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_309),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_309),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_313),
.B(n_195),
.Y(n_405)
);

XNOR2x2_ASAP7_75t_R g406 ( 
.A(n_304),
.B(n_5),
.Y(n_406)
);

HB1xp67_ASAP7_75t_L g407 ( 
.A(n_353),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_310),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_310),
.Y(n_409)
);

OA21x2_ASAP7_75t_L g410 ( 
.A1(n_311),
.A2(n_316),
.B(n_315),
.Y(n_410)
);

AND2x4_ASAP7_75t_L g411 ( 
.A(n_372),
.B(n_348),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_307),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_311),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_315),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_340),
.Y(n_415)
);

INVx2_ASAP7_75t_SL g416 ( 
.A(n_316),
.Y(n_416)
);

AND2x4_ASAP7_75t_L g417 ( 
.A(n_369),
.B(n_201),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_319),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_319),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_321),
.Y(n_420)
);

HB1xp67_ASAP7_75t_L g421 ( 
.A(n_331),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_321),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_323),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_323),
.Y(n_424)
);

HB1xp67_ASAP7_75t_L g425 ( 
.A(n_333),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_318),
.B(n_204),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_328),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_328),
.Y(n_428)
);

OAI21x1_ASAP7_75t_L g429 ( 
.A1(n_343),
.A2(n_182),
.B(n_175),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_335),
.Y(n_430)
);

AND2x4_ASAP7_75t_L g431 ( 
.A(n_326),
.B(n_339),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_335),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_336),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_336),
.Y(n_434)
);

INVx3_ASAP7_75t_L g435 ( 
.A(n_337),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_337),
.Y(n_436)
);

HB1xp67_ASAP7_75t_L g437 ( 
.A(n_334),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_341),
.B(n_196),
.Y(n_438)
);

AND2x4_ASAP7_75t_L g439 ( 
.A(n_358),
.B(n_210),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_358),
.B(n_216),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_341),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_345),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_345),
.Y(n_443)
);

OR2x6_ASAP7_75t_L g444 ( 
.A(n_366),
.B(n_222),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_347),
.B(n_198),
.Y(n_445)
);

HB1xp67_ASAP7_75t_L g446 ( 
.A(n_338),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_384),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_385),
.B(n_325),
.Y(n_448)
);

AND2x2_ASAP7_75t_SL g449 ( 
.A(n_385),
.B(n_362),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_384),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_385),
.A2(n_354),
.B1(n_325),
.B2(n_362),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_410),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_384),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_410),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_385),
.B(n_354),
.Y(n_455)
);

NAND3xp33_ASAP7_75t_L g456 ( 
.A(n_385),
.B(n_355),
.C(n_346),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_389),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_440),
.Y(n_458)
);

NAND3xp33_ASAP7_75t_L g459 ( 
.A(n_378),
.B(n_363),
.C(n_359),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_389),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_378),
.B(n_368),
.Y(n_461)
);

AND2x6_ASAP7_75t_L g462 ( 
.A(n_378),
.B(n_255),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_389),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_410),
.Y(n_464)
);

INVxp67_ASAP7_75t_L g465 ( 
.A(n_390),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_410),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_410),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_410),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_379),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_401),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_401),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_379),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_379),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_411),
.B(n_373),
.Y(n_474)
);

AND2x4_ASAP7_75t_L g475 ( 
.A(n_444),
.B(n_411),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_401),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_379),
.Y(n_477)
);

AND2x6_ASAP7_75t_L g478 ( 
.A(n_378),
.B(n_255),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_411),
.B(n_374),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_381),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_408),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_381),
.Y(n_482)
);

INVxp67_ASAP7_75t_SL g483 ( 
.A(n_381),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_431),
.B(n_421),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_408),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_411),
.B(n_377),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_440),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_381),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_411),
.B(n_417),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_440),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_440),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_431),
.B(n_312),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_408),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_382),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_382),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_418),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_382),
.Y(n_497)
);

INVx2_ASAP7_75t_SL g498 ( 
.A(n_431),
.Y(n_498)
);

INVx2_ASAP7_75t_SL g499 ( 
.A(n_431),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_417),
.B(n_361),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_418),
.Y(n_501)
);

INVx2_ASAP7_75t_SL g502 ( 
.A(n_431),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_382),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_418),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_431),
.B(n_322),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_392),
.Y(n_506)
);

AND2x4_ASAP7_75t_L g507 ( 
.A(n_444),
.B(n_366),
.Y(n_507)
);

NAND3xp33_ASAP7_75t_L g508 ( 
.A(n_394),
.B(n_351),
.C(n_161),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_421),
.B(n_329),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_420),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_426),
.B(n_439),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_425),
.B(n_153),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_417),
.B(n_347),
.Y(n_513)
);

BUFx3_ASAP7_75t_L g514 ( 
.A(n_392),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_420),
.Y(n_515)
);

AND2x6_ASAP7_75t_L g516 ( 
.A(n_392),
.B(n_255),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_392),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_420),
.Y(n_518)
);

BUFx3_ASAP7_75t_L g519 ( 
.A(n_380),
.Y(n_519)
);

INVx3_ASAP7_75t_L g520 ( 
.A(n_435),
.Y(n_520)
);

BUFx8_ASAP7_75t_SL g521 ( 
.A(n_390),
.Y(n_521)
);

INVx2_ASAP7_75t_SL g522 ( 
.A(n_444),
.Y(n_522)
);

AND2x6_ASAP7_75t_L g523 ( 
.A(n_380),
.B(n_255),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_SL g524 ( 
.A(n_412),
.B(n_364),
.Y(n_524)
);

NAND2xp33_ASAP7_75t_L g525 ( 
.A(n_425),
.B(n_187),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_435),
.Y(n_526)
);

AND2x6_ASAP7_75t_L g527 ( 
.A(n_380),
.B(n_255),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_426),
.B(n_365),
.Y(n_528)
);

INVx2_ASAP7_75t_SL g529 ( 
.A(n_444),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_422),
.Y(n_530)
);

INVx5_ASAP7_75t_L g531 ( 
.A(n_396),
.Y(n_531)
);

OR2x6_ASAP7_75t_L g532 ( 
.A(n_444),
.B(n_365),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_417),
.B(n_349),
.Y(n_533)
);

INVx3_ASAP7_75t_L g534 ( 
.A(n_435),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_417),
.B(n_349),
.Y(n_535)
);

BUFx3_ASAP7_75t_L g536 ( 
.A(n_380),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_417),
.B(n_371),
.Y(n_537)
);

AND2x4_ASAP7_75t_L g538 ( 
.A(n_444),
.B(n_405),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_422),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_422),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_380),
.B(n_352),
.Y(n_541)
);

INVx4_ASAP7_75t_L g542 ( 
.A(n_444),
.Y(n_542)
);

AND2x6_ASAP7_75t_L g543 ( 
.A(n_380),
.B(n_205),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_423),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_423),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_383),
.B(n_352),
.Y(n_546)
);

AND2x6_ASAP7_75t_L g547 ( 
.A(n_383),
.B(n_209),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_383),
.B(n_183),
.Y(n_548)
);

OR2x6_ASAP7_75t_L g549 ( 
.A(n_444),
.B(n_223),
.Y(n_549)
);

AOI22xp33_ASAP7_75t_L g550 ( 
.A1(n_383),
.A2(n_229),
.B1(n_263),
.B2(n_302),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_423),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_435),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_437),
.B(n_153),
.Y(n_553)
);

HB1xp67_ASAP7_75t_L g554 ( 
.A(n_394),
.Y(n_554)
);

INVx4_ASAP7_75t_L g555 ( 
.A(n_383),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_435),
.Y(n_556)
);

OR2x2_ASAP7_75t_L g557 ( 
.A(n_407),
.B(n_344),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_430),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_383),
.B(n_221),
.Y(n_559)
);

OR2x2_ASAP7_75t_L g560 ( 
.A(n_407),
.B(n_297),
.Y(n_560)
);

OR2x6_ASAP7_75t_L g561 ( 
.A(n_405),
.B(n_240),
.Y(n_561)
);

INVx3_ASAP7_75t_L g562 ( 
.A(n_435),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_437),
.B(n_156),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_430),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_399),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_446),
.B(n_375),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_399),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_399),
.Y(n_568)
);

INVxp67_ASAP7_75t_SL g569 ( 
.A(n_395),
.Y(n_569)
);

BUFx4f_ASAP7_75t_L g570 ( 
.A(n_400),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_430),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_393),
.Y(n_572)
);

INVx4_ASAP7_75t_L g573 ( 
.A(n_386),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_386),
.B(n_156),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_446),
.B(n_250),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_400),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_432),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_432),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_426),
.B(n_163),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_399),
.Y(n_580)
);

INVx3_ASAP7_75t_L g581 ( 
.A(n_400),
.Y(n_581)
);

INVx3_ASAP7_75t_L g582 ( 
.A(n_400),
.Y(n_582)
);

NAND2xp33_ASAP7_75t_R g583 ( 
.A(n_390),
.B(n_314),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_405),
.B(n_324),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_R g585 ( 
.A(n_393),
.B(n_327),
.Y(n_585)
);

HB1xp67_ASAP7_75t_L g586 ( 
.A(n_412),
.Y(n_586)
);

AOI22xp33_ASAP7_75t_L g587 ( 
.A1(n_386),
.A2(n_276),
.B1(n_301),
.B2(n_293),
.Y(n_587)
);

INVxp67_ASAP7_75t_SL g588 ( 
.A(n_395),
.Y(n_588)
);

OAI21xp33_ASAP7_75t_SL g589 ( 
.A1(n_429),
.A2(n_242),
.B(n_296),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_403),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_403),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_432),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_434),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_426),
.B(n_163),
.Y(n_594)
);

OAI22xp5_ASAP7_75t_L g595 ( 
.A1(n_498),
.A2(n_415),
.B1(n_179),
.B2(n_177),
.Y(n_595)
);

AOI22xp5_ASAP7_75t_L g596 ( 
.A1(n_449),
.A2(n_405),
.B1(n_415),
.B2(n_391),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_569),
.B(n_391),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_449),
.B(n_391),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_588),
.B(n_391),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_511),
.B(n_439),
.Y(n_600)
);

AOI22xp33_ASAP7_75t_L g601 ( 
.A1(n_475),
.A2(n_388),
.B1(n_386),
.B2(n_439),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_470),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_475),
.B(n_171),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_511),
.B(n_439),
.Y(n_604)
);

NOR3xp33_ASAP7_75t_L g605 ( 
.A(n_465),
.B(n_161),
.C(n_160),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_489),
.B(n_498),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_499),
.B(n_386),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_SL g608 ( 
.A(n_566),
.B(n_406),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_456),
.B(n_455),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_499),
.B(n_386),
.Y(n_610)
);

O2A1O1Ixp33_ASAP7_75t_L g611 ( 
.A1(n_486),
.A2(n_445),
.B(n_438),
.C(n_439),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_470),
.Y(n_612)
);

BUFx3_ASAP7_75t_L g613 ( 
.A(n_519),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_502),
.B(n_388),
.Y(n_614)
);

BUFx12f_ASAP7_75t_SL g615 ( 
.A(n_549),
.Y(n_615)
);

INVx3_ASAP7_75t_L g616 ( 
.A(n_514),
.Y(n_616)
);

AOI22xp33_ASAP7_75t_L g617 ( 
.A1(n_475),
.A2(n_538),
.B1(n_529),
.B2(n_522),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_R g618 ( 
.A(n_583),
.B(n_332),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_538),
.B(n_439),
.Y(n_619)
);

AOI22xp33_ASAP7_75t_L g620 ( 
.A1(n_538),
.A2(n_388),
.B1(n_429),
.B2(n_445),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_502),
.B(n_388),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_479),
.B(n_388),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_471),
.Y(n_623)
);

INVx2_ASAP7_75t_SL g624 ( 
.A(n_532),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_462),
.B(n_388),
.Y(n_625)
);

AOI22xp5_ASAP7_75t_L g626 ( 
.A1(n_448),
.A2(n_171),
.B1(n_290),
.B2(n_173),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_561),
.B(n_458),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_514),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_462),
.B(n_429),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_462),
.B(n_478),
.Y(n_630)
);

INVx3_ASAP7_75t_L g631 ( 
.A(n_520),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_451),
.B(n_459),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_462),
.B(n_438),
.Y(n_633)
);

OAI22xp33_ASAP7_75t_L g634 ( 
.A1(n_561),
.A2(n_272),
.B1(n_164),
.B2(n_167),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_462),
.B(n_438),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_461),
.B(n_342),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_500),
.B(n_350),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_471),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_478),
.B(n_445),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_537),
.B(n_357),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_478),
.B(n_387),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_469),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_478),
.B(n_387),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_474),
.B(n_174),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_476),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_478),
.B(n_416),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_575),
.B(n_174),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_476),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_478),
.B(n_416),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_487),
.B(n_490),
.Y(n_650)
);

BUFx6f_ASAP7_75t_L g651 ( 
.A(n_452),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_481),
.Y(n_652)
);

INVxp67_ASAP7_75t_L g653 ( 
.A(n_557),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_491),
.B(n_416),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_528),
.B(n_507),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_528),
.B(n_416),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_507),
.B(n_434),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_469),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_507),
.B(n_176),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_472),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_484),
.B(n_160),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_L g662 ( 
.A(n_492),
.B(n_164),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_481),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_485),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_522),
.B(n_434),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_485),
.Y(n_666)
);

INVxp67_ASAP7_75t_SL g667 ( 
.A(n_452),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_501),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_505),
.B(n_512),
.Y(n_669)
);

AOI22xp5_ASAP7_75t_L g670 ( 
.A1(n_525),
.A2(n_181),
.B1(n_176),
.B2(n_290),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_529),
.B(n_181),
.Y(n_671)
);

AOI22xp5_ASAP7_75t_L g672 ( 
.A1(n_525),
.A2(n_224),
.B1(n_215),
.B2(n_225),
.Y(n_672)
);

INVx8_ASAP7_75t_L g673 ( 
.A(n_532),
.Y(n_673)
);

NOR3xp33_ASAP7_75t_L g674 ( 
.A(n_553),
.B(n_272),
.C(n_168),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_472),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_521),
.Y(n_676)
);

OAI221xp5_ASAP7_75t_L g677 ( 
.A1(n_550),
.A2(n_274),
.B1(n_168),
.B2(n_177),
.C(n_179),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_473),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_548),
.B(n_436),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_501),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_504),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_504),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_510),
.Y(n_683)
);

AOI22xp33_ASAP7_75t_L g684 ( 
.A1(n_542),
.A2(n_262),
.B1(n_443),
.B2(n_441),
.Y(n_684)
);

BUFx6f_ASAP7_75t_L g685 ( 
.A(n_452),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_559),
.B(n_436),
.Y(n_686)
);

INVxp33_ASAP7_75t_L g687 ( 
.A(n_557),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_555),
.B(n_167),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_473),
.Y(n_689)
);

AOI22xp33_ASAP7_75t_L g690 ( 
.A1(n_542),
.A2(n_262),
.B1(n_443),
.B2(n_441),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_555),
.B(n_269),
.Y(n_691)
);

OR2x2_ASAP7_75t_L g692 ( 
.A(n_560),
.B(n_269),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_510),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_519),
.B(n_436),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_561),
.B(n_443),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_555),
.B(n_274),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_536),
.B(n_441),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_477),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_515),
.Y(n_699)
);

AOI221xp5_ASAP7_75t_L g700 ( 
.A1(n_584),
.A2(n_275),
.B1(n_278),
.B2(n_292),
.C(n_288),
.Y(n_700)
);

AOI22xp5_ASAP7_75t_L g701 ( 
.A1(n_549),
.A2(n_235),
.B1(n_253),
.B2(n_260),
.Y(n_701)
);

HB1xp67_ASAP7_75t_L g702 ( 
.A(n_554),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_563),
.B(n_275),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_515),
.Y(n_704)
);

INVxp67_ASAP7_75t_L g705 ( 
.A(n_586),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_536),
.B(n_397),
.Y(n_706)
);

NAND2x1p5_ASAP7_75t_L g707 ( 
.A(n_542),
.B(n_266),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_573),
.B(n_278),
.Y(n_708)
);

AOI221xp5_ASAP7_75t_L g709 ( 
.A1(n_508),
.A2(n_279),
.B1(n_280),
.B2(n_292),
.C(n_288),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_573),
.B(n_279),
.Y(n_710)
);

NAND2xp33_ASAP7_75t_L g711 ( 
.A(n_452),
.B(n_187),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_483),
.B(n_573),
.Y(n_712)
);

OAI22xp5_ASAP7_75t_L g713 ( 
.A1(n_549),
.A2(n_280),
.B1(n_286),
.B2(n_285),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_520),
.B(n_397),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_477),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_520),
.B(n_397),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_518),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_480),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_560),
.B(n_281),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_480),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_482),
.Y(n_721)
);

INVxp33_ASAP7_75t_L g722 ( 
.A(n_585),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_579),
.B(n_281),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_482),
.Y(n_724)
);

INVx2_ASAP7_75t_SL g725 ( 
.A(n_532),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_534),
.B(n_398),
.Y(n_726)
);

BUFx3_ASAP7_75t_L g727 ( 
.A(n_532),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_534),
.B(n_398),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_594),
.B(n_283),
.Y(n_729)
);

INVxp67_ASAP7_75t_SL g730 ( 
.A(n_452),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_562),
.B(n_398),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_562),
.B(n_403),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_488),
.Y(n_733)
);

OAI22xp33_ASAP7_75t_L g734 ( 
.A1(n_561),
.A2(n_283),
.B1(n_285),
.B2(n_286),
.Y(n_734)
);

INVxp67_ASAP7_75t_L g735 ( 
.A(n_524),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_488),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_518),
.Y(n_737)
);

NAND3xp33_ASAP7_75t_L g738 ( 
.A(n_509),
.B(n_234),
.C(n_239),
.Y(n_738)
);

OAI22xp5_ASAP7_75t_L g739 ( 
.A1(n_549),
.A2(n_245),
.B1(n_251),
.B2(n_268),
.Y(n_739)
);

BUFx2_ASAP7_75t_L g740 ( 
.A(n_521),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_587),
.B(n_247),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_513),
.B(n_403),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_533),
.B(n_535),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_447),
.B(n_404),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_572),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_447),
.B(n_450),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_530),
.Y(n_747)
);

OR2x2_ASAP7_75t_L g748 ( 
.A(n_572),
.B(n_248),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_530),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_574),
.B(n_254),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_539),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_450),
.B(n_404),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_464),
.B(n_258),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_453),
.B(n_261),
.Y(n_754)
);

INVxp67_ASAP7_75t_L g755 ( 
.A(n_541),
.Y(n_755)
);

AND2x2_ASAP7_75t_L g756 ( 
.A(n_453),
.B(n_404),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_539),
.Y(n_757)
);

AOI22xp5_ASAP7_75t_L g758 ( 
.A1(n_543),
.A2(n_547),
.B1(n_468),
.B2(n_467),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_457),
.B(n_404),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_457),
.B(n_424),
.Y(n_760)
);

AND2x2_ASAP7_75t_L g761 ( 
.A(n_460),
.B(n_424),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_460),
.B(n_264),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_464),
.B(n_265),
.Y(n_763)
);

INVxp67_ASAP7_75t_L g764 ( 
.A(n_546),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_467),
.B(n_186),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_602),
.Y(n_766)
);

NAND2xp33_ASAP7_75t_L g767 ( 
.A(n_651),
.B(n_543),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_597),
.B(n_543),
.Y(n_768)
);

INVx3_ASAP7_75t_L g769 ( 
.A(n_673),
.Y(n_769)
);

AOI21xp5_ASAP7_75t_L g770 ( 
.A1(n_732),
.A2(n_463),
.B(n_570),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_599),
.B(n_543),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_653),
.B(n_463),
.Y(n_772)
);

AOI21x1_ASAP7_75t_L g773 ( 
.A1(n_629),
.A2(n_593),
.B(n_592),
.Y(n_773)
);

AOI22xp5_ASAP7_75t_L g774 ( 
.A1(n_598),
.A2(n_547),
.B1(n_543),
.B2(n_523),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_655),
.B(n_543),
.Y(n_775)
);

AOI21xp5_ASAP7_75t_L g776 ( 
.A1(n_667),
.A2(n_570),
.B(n_589),
.Y(n_776)
);

AOI21xp5_ASAP7_75t_L g777 ( 
.A1(n_730),
.A2(n_570),
.B(n_592),
.Y(n_777)
);

AOI21xp5_ASAP7_75t_L g778 ( 
.A1(n_714),
.A2(n_593),
.B(n_564),
.Y(n_778)
);

INVx4_ASAP7_75t_L g779 ( 
.A(n_673),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_606),
.B(n_547),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_755),
.B(n_547),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_764),
.B(n_547),
.Y(n_782)
);

OR2x2_ASAP7_75t_L g783 ( 
.A(n_692),
.B(n_454),
.Y(n_783)
);

OAI22xp5_ASAP7_75t_L g784 ( 
.A1(n_622),
.A2(n_564),
.B1(n_540),
.B2(n_571),
.Y(n_784)
);

AOI21xp5_ASAP7_75t_L g785 ( 
.A1(n_716),
.A2(n_577),
.B(n_540),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_687),
.B(n_526),
.Y(n_786)
);

BUFx6f_ASAP7_75t_L g787 ( 
.A(n_673),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_618),
.Y(n_788)
);

NOR3xp33_ASAP7_75t_L g789 ( 
.A(n_700),
.B(n_406),
.C(n_544),
.Y(n_789)
);

AOI21xp5_ASAP7_75t_L g790 ( 
.A1(n_712),
.A2(n_466),
.B(n_552),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_596),
.B(n_466),
.Y(n_791)
);

INVx3_ASAP7_75t_L g792 ( 
.A(n_673),
.Y(n_792)
);

NAND3xp33_ASAP7_75t_L g793 ( 
.A(n_705),
.B(n_545),
.C(n_551),
.Y(n_793)
);

AOI21xp5_ASAP7_75t_L g794 ( 
.A1(n_746),
.A2(n_526),
.B(n_552),
.Y(n_794)
);

AOI21xp5_ASAP7_75t_L g795 ( 
.A1(n_726),
.A2(n_556),
.B(n_571),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_600),
.B(n_547),
.Y(n_796)
);

AOI21xp5_ASAP7_75t_L g797 ( 
.A1(n_728),
.A2(n_556),
.B(n_577),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_642),
.Y(n_798)
);

AOI21xp5_ASAP7_75t_L g799 ( 
.A1(n_731),
.A2(n_578),
.B(n_576),
.Y(n_799)
);

AOI22xp5_ASAP7_75t_L g800 ( 
.A1(n_632),
.A2(n_609),
.B1(n_627),
.B2(n_669),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_624),
.B(n_578),
.Y(n_801)
);

AND2x4_ASAP7_75t_L g802 ( 
.A(n_727),
.B(n_624),
.Y(n_802)
);

AOI21xp5_ASAP7_75t_L g803 ( 
.A1(n_765),
.A2(n_576),
.B(n_581),
.Y(n_803)
);

AOI21xp5_ASAP7_75t_L g804 ( 
.A1(n_651),
.A2(n_576),
.B(n_581),
.Y(n_804)
);

AOI21xp5_ASAP7_75t_L g805 ( 
.A1(n_651),
.A2(n_581),
.B(n_582),
.Y(n_805)
);

A2O1A1Ixp33_ASAP7_75t_L g806 ( 
.A1(n_611),
.A2(n_558),
.B(n_493),
.C(n_496),
.Y(n_806)
);

BUFx2_ASAP7_75t_L g807 ( 
.A(n_702),
.Y(n_807)
);

AOI21xp5_ASAP7_75t_L g808 ( 
.A1(n_743),
.A2(n_494),
.B(n_495),
.Y(n_808)
);

NAND2x1p5_ASAP7_75t_L g809 ( 
.A(n_727),
.B(n_494),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_687),
.B(n_495),
.Y(n_810)
);

INVx3_ASAP7_75t_L g811 ( 
.A(n_631),
.Y(n_811)
);

O2A1O1Ixp5_ASAP7_75t_L g812 ( 
.A1(n_750),
.A2(n_763),
.B(n_753),
.C(n_644),
.Y(n_812)
);

O2A1O1Ixp33_ASAP7_75t_SL g813 ( 
.A1(n_612),
.A2(n_582),
.B(n_506),
.C(n_517),
.Y(n_813)
);

AND2x2_ASAP7_75t_L g814 ( 
.A(n_692),
.B(n_591),
.Y(n_814)
);

OAI21xp5_ASAP7_75t_L g815 ( 
.A1(n_758),
.A2(n_517),
.B(n_497),
.Y(n_815)
);

AOI21xp33_ASAP7_75t_L g816 ( 
.A1(n_703),
.A2(n_506),
.B(n_497),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_600),
.B(n_503),
.Y(n_817)
);

AOI21xp5_ASAP7_75t_L g818 ( 
.A1(n_612),
.A2(n_503),
.B(n_582),
.Y(n_818)
);

AOI21xp5_ASAP7_75t_L g819 ( 
.A1(n_623),
.A2(n_591),
.B(n_590),
.Y(n_819)
);

BUFx12f_ASAP7_75t_L g820 ( 
.A(n_676),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_604),
.B(n_565),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_637),
.B(n_590),
.Y(n_822)
);

NAND2x1p5_ASAP7_75t_L g823 ( 
.A(n_725),
.B(n_565),
.Y(n_823)
);

O2A1O1Ixp33_ASAP7_75t_L g824 ( 
.A1(n_634),
.A2(n_580),
.B(n_568),
.C(n_567),
.Y(n_824)
);

AOI21xp5_ASAP7_75t_L g825 ( 
.A1(n_623),
.A2(n_580),
.B(n_568),
.Y(n_825)
);

A2O1A1Ixp33_ASAP7_75t_L g826 ( 
.A1(n_645),
.A2(n_567),
.B(n_284),
.C(n_427),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_645),
.Y(n_827)
);

AOI22xp5_ASAP7_75t_L g828 ( 
.A1(n_627),
.A2(n_523),
.B1(n_527),
.B2(n_249),
.Y(n_828)
);

BUFx6f_ASAP7_75t_L g829 ( 
.A(n_613),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_725),
.B(n_531),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_658),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_604),
.B(n_523),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_648),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_619),
.B(n_523),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_648),
.A2(n_531),
.B(n_424),
.Y(n_835)
);

AOI21xp5_ASAP7_75t_L g836 ( 
.A1(n_652),
.A2(n_531),
.B(n_424),
.Y(n_836)
);

O2A1O1Ixp33_ASAP7_75t_L g837 ( 
.A1(n_734),
.A2(n_427),
.B(n_433),
.C(n_442),
.Y(n_837)
);

BUFx6f_ASAP7_75t_L g838 ( 
.A(n_613),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_619),
.B(n_523),
.Y(n_839)
);

OAI21xp5_ASAP7_75t_L g840 ( 
.A1(n_656),
.A2(n_531),
.B(n_527),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_640),
.B(n_735),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_652),
.A2(n_531),
.B(n_427),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_663),
.A2(n_427),
.B(n_433),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_658),
.Y(n_844)
);

BUFx6f_ASAP7_75t_L g845 ( 
.A(n_651),
.Y(n_845)
);

AOI21xp33_ASAP7_75t_L g846 ( 
.A1(n_723),
.A2(n_442),
.B(n_433),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_685),
.A2(n_252),
.B(n_197),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_617),
.B(n_199),
.Y(n_848)
);

AOI21xp5_ASAP7_75t_L g849 ( 
.A1(n_685),
.A2(n_256),
.B(n_200),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_754),
.B(n_523),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_762),
.B(n_527),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_685),
.A2(n_257),
.B(n_203),
.Y(n_852)
);

AOI21xp5_ASAP7_75t_L g853 ( 
.A1(n_685),
.A2(n_211),
.B(n_206),
.Y(n_853)
);

OAI21xp5_ASAP7_75t_L g854 ( 
.A1(n_711),
.A2(n_527),
.B(n_442),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_663),
.A2(n_433),
.B(n_442),
.Y(n_855)
);

NOR2xp67_ASAP7_75t_R g856 ( 
.A(n_740),
.B(n_527),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_680),
.A2(n_220),
.B(n_208),
.Y(n_857)
);

AOI21xp33_ASAP7_75t_L g858 ( 
.A1(n_729),
.A2(n_212),
.B(n_226),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_650),
.B(n_527),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_695),
.B(n_243),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_660),
.Y(n_861)
);

AOI21xp5_ASAP7_75t_L g862 ( 
.A1(n_680),
.A2(n_230),
.B(n_238),
.Y(n_862)
);

BUFx2_ASAP7_75t_L g863 ( 
.A(n_615),
.Y(n_863)
);

AND2x4_ASAP7_75t_SL g864 ( 
.A(n_695),
.B(n_396),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_636),
.B(n_8),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_601),
.B(n_228),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_L g867 ( 
.A(n_647),
.B(n_9),
.Y(n_867)
);

AND2x2_ASAP7_75t_L g868 ( 
.A(n_661),
.B(n_9),
.Y(n_868)
);

BUFx4f_ASAP7_75t_L g869 ( 
.A(n_740),
.Y(n_869)
);

A2O1A1Ixp33_ASAP7_75t_L g870 ( 
.A1(n_683),
.A2(n_699),
.B(n_757),
.C(n_751),
.Y(n_870)
);

A2O1A1Ixp33_ASAP7_75t_L g871 ( 
.A1(n_693),
.A2(n_413),
.B(n_400),
.C(n_402),
.Y(n_871)
);

BUFx2_ASAP7_75t_SL g872 ( 
.A(n_659),
.Y(n_872)
);

OAI22xp5_ASAP7_75t_L g873 ( 
.A1(n_693),
.A2(n_413),
.B1(n_400),
.B2(n_402),
.Y(n_873)
);

AND2x4_ASAP7_75t_L g874 ( 
.A(n_603),
.B(n_516),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_660),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_719),
.B(n_10),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_638),
.B(n_664),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_666),
.B(n_516),
.Y(n_878)
);

BUFx6f_ASAP7_75t_L g879 ( 
.A(n_628),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_704),
.A2(n_396),
.B(n_428),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_668),
.B(n_516),
.Y(n_881)
);

INVx5_ASAP7_75t_L g882 ( 
.A(n_616),
.Y(n_882)
);

INVx3_ASAP7_75t_L g883 ( 
.A(n_631),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_704),
.A2(n_396),
.B(n_428),
.Y(n_884)
);

BUFx2_ASAP7_75t_L g885 ( 
.A(n_615),
.Y(n_885)
);

AOI22xp33_ASAP7_75t_L g886 ( 
.A1(n_741),
.A2(n_516),
.B1(n_428),
.B2(n_419),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_717),
.A2(n_396),
.B(n_428),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_681),
.B(n_516),
.Y(n_888)
);

AOI21x1_ASAP7_75t_L g889 ( 
.A1(n_744),
.A2(n_516),
.B(n_396),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_682),
.B(n_11),
.Y(n_890)
);

NOR2xp33_ASAP7_75t_R g891 ( 
.A(n_745),
.B(n_91),
.Y(n_891)
);

NOR2xp33_ASAP7_75t_L g892 ( 
.A(n_662),
.B(n_11),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_675),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_717),
.A2(n_396),
.B(n_419),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_737),
.B(n_13),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_737),
.Y(n_896)
);

A2O1A1Ixp33_ASAP7_75t_L g897 ( 
.A1(n_747),
.A2(n_428),
.B(n_419),
.C(n_414),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_747),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_749),
.A2(n_396),
.B(n_419),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_749),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_748),
.B(n_13),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_751),
.B(n_15),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_757),
.B(n_15),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_SL g904 ( 
.A(n_670),
.B(n_428),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_631),
.B(n_16),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_742),
.B(n_20),
.Y(n_906)
);

OAI321xp33_ASAP7_75t_L g907 ( 
.A1(n_677),
.A2(n_428),
.A3(n_419),
.B1(n_414),
.B2(n_413),
.C(n_409),
.Y(n_907)
);

AND2x2_ASAP7_75t_L g908 ( 
.A(n_608),
.B(n_20),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_752),
.A2(n_419),
.B(n_414),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_742),
.B(n_22),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_679),
.B(n_22),
.Y(n_911)
);

AOI22xp5_ASAP7_75t_L g912 ( 
.A1(n_701),
.A2(n_672),
.B1(n_626),
.B2(n_713),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_686),
.B(n_616),
.Y(n_913)
);

HB1xp67_ASAP7_75t_L g914 ( 
.A(n_745),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_756),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_616),
.B(n_24),
.Y(n_916)
);

INVx3_ASAP7_75t_L g917 ( 
.A(n_628),
.Y(n_917)
);

A2O1A1Ixp33_ASAP7_75t_L g918 ( 
.A1(n_657),
.A2(n_419),
.B(n_414),
.C(n_413),
.Y(n_918)
);

AO21x1_ASAP7_75t_L g919 ( 
.A1(n_711),
.A2(n_187),
.B(n_414),
.Y(n_919)
);

CKINVDCx10_ASAP7_75t_R g920 ( 
.A(n_676),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_759),
.A2(n_419),
.B(n_414),
.Y(n_921)
);

HB1xp67_ASAP7_75t_L g922 ( 
.A(n_748),
.Y(n_922)
);

BUFx3_ASAP7_75t_L g923 ( 
.A(n_738),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_607),
.B(n_24),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_760),
.A2(n_419),
.B(n_414),
.Y(n_925)
);

AOI22xp5_ASAP7_75t_L g926 ( 
.A1(n_739),
.A2(n_414),
.B1(n_413),
.B2(n_409),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_610),
.B(n_25),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_595),
.B(n_29),
.Y(n_928)
);

HB1xp67_ASAP7_75t_L g929 ( 
.A(n_641),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_694),
.A2(n_414),
.B(n_413),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_614),
.B(n_30),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_621),
.B(n_30),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_722),
.B(n_31),
.Y(n_933)
);

OAI21xp5_ASAP7_75t_L g934 ( 
.A1(n_756),
.A2(n_413),
.B(n_409),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_761),
.Y(n_935)
);

BUFx6f_ASAP7_75t_L g936 ( 
.A(n_707),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_620),
.B(n_35),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_761),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_697),
.A2(n_413),
.B(n_409),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_706),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_654),
.B(n_42),
.Y(n_941)
);

OR2x6_ASAP7_75t_L g942 ( 
.A(n_707),
.B(n_413),
.Y(n_942)
);

OAI21xp5_ASAP7_75t_L g943 ( 
.A1(n_665),
.A2(n_413),
.B(n_409),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_722),
.B(n_43),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_772),
.B(n_709),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_784),
.A2(n_688),
.B(n_708),
.Y(n_946)
);

AO21x2_ASAP7_75t_L g947 ( 
.A1(n_773),
.A2(n_639),
.B(n_633),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_841),
.B(n_674),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_776),
.A2(n_696),
.B(n_691),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_822),
.B(n_605),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_800),
.B(n_643),
.Y(n_951)
);

A2O1A1Ixp33_ASAP7_75t_SL g952 ( 
.A1(n_892),
.A2(n_690),
.B(n_684),
.C(n_724),
.Y(n_952)
);

O2A1O1Ixp33_ASAP7_75t_L g953 ( 
.A1(n_901),
.A2(n_710),
.B(n_671),
.C(n_635),
.Y(n_953)
);

NOR2xp33_ASAP7_75t_R g954 ( 
.A(n_788),
.B(n_625),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_814),
.B(n_736),
.Y(n_955)
);

INVxp67_ASAP7_75t_L g956 ( 
.A(n_807),
.Y(n_956)
);

AOI22xp5_ASAP7_75t_L g957 ( 
.A1(n_789),
.A2(n_630),
.B1(n_646),
.B2(n_649),
.Y(n_957)
);

CKINVDCx20_ASAP7_75t_R g958 ( 
.A(n_869),
.Y(n_958)
);

BUFx6f_ASAP7_75t_L g959 ( 
.A(n_787),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_783),
.B(n_736),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_798),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_766),
.Y(n_962)
);

BUFx12f_ASAP7_75t_L g963 ( 
.A(n_820),
.Y(n_963)
);

A2O1A1Ixp33_ASAP7_75t_SL g964 ( 
.A1(n_933),
.A2(n_733),
.B(n_724),
.C(n_721),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_915),
.B(n_721),
.Y(n_965)
);

OAI22xp5_ASAP7_75t_L g966 ( 
.A1(n_912),
.A2(n_689),
.B1(n_718),
.B2(n_715),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_935),
.B(n_720),
.Y(n_967)
);

AOI21x1_ASAP7_75t_L g968 ( 
.A1(n_770),
.A2(n_720),
.B(n_718),
.Y(n_968)
);

AND2x6_ASAP7_75t_L g969 ( 
.A(n_787),
.B(n_715),
.Y(n_969)
);

O2A1O1Ixp5_ASAP7_75t_L g970 ( 
.A1(n_919),
.A2(n_812),
.B(n_776),
.C(n_850),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_922),
.B(n_698),
.Y(n_971)
);

NOR2xp67_ASAP7_75t_L g972 ( 
.A(n_914),
.B(n_689),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_938),
.B(n_678),
.Y(n_973)
);

INVx8_ASAP7_75t_L g974 ( 
.A(n_787),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_827),
.Y(n_975)
);

NOR2xp33_ASAP7_75t_L g976 ( 
.A(n_865),
.B(n_43),
.Y(n_976)
);

AOI22xp5_ASAP7_75t_L g977 ( 
.A1(n_868),
.A2(n_409),
.B1(n_402),
.B2(n_400),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_833),
.Y(n_978)
);

OAI221xp5_ASAP7_75t_L g979 ( 
.A1(n_876),
.A2(n_409),
.B1(n_402),
.B2(n_400),
.C(n_57),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_940),
.B(n_44),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_810),
.B(n_45),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_786),
.B(n_45),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_896),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_R g984 ( 
.A(n_920),
.B(n_105),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_770),
.A2(n_409),
.B(n_402),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_869),
.B(n_400),
.Y(n_986)
);

OAI22xp5_ASAP7_75t_L g987 ( 
.A1(n_877),
.A2(n_402),
.B1(n_400),
.B2(n_46),
.Y(n_987)
);

CKINVDCx8_ASAP7_75t_R g988 ( 
.A(n_872),
.Y(n_988)
);

O2A1O1Ixp33_ASAP7_75t_L g989 ( 
.A1(n_867),
.A2(n_58),
.B(n_187),
.C(n_402),
.Y(n_989)
);

OAI22xp5_ASAP7_75t_L g990 ( 
.A1(n_898),
.A2(n_402),
.B1(n_187),
.B2(n_70),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_790),
.A2(n_187),
.B(n_66),
.Y(n_991)
);

NOR3xp33_ASAP7_75t_L g992 ( 
.A(n_944),
.B(n_65),
.C(n_72),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_831),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_900),
.B(n_860),
.Y(n_994)
);

INVx3_ASAP7_75t_L g995 ( 
.A(n_779),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_870),
.A2(n_78),
.B(n_82),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_777),
.A2(n_84),
.B(n_94),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_895),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_802),
.B(n_97),
.Y(n_999)
);

O2A1O1Ixp33_ASAP7_75t_SL g1000 ( 
.A1(n_780),
.A2(n_98),
.B(n_101),
.C(n_104),
.Y(n_1000)
);

NOR2xp33_ASAP7_75t_R g1001 ( 
.A(n_863),
.B(n_107),
.Y(n_1001)
);

O2A1O1Ixp33_ASAP7_75t_L g1002 ( 
.A1(n_928),
.A2(n_116),
.B(n_117),
.C(n_123),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_777),
.A2(n_124),
.B(n_128),
.Y(n_1003)
);

OAI22xp5_ASAP7_75t_L g1004 ( 
.A1(n_796),
.A2(n_135),
.B1(n_141),
.B2(n_146),
.Y(n_1004)
);

OR2x2_ASAP7_75t_L g1005 ( 
.A(n_885),
.B(n_150),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_802),
.B(n_821),
.Y(n_1006)
);

OAI22xp5_ASAP7_75t_L g1007 ( 
.A1(n_768),
.A2(n_771),
.B1(n_817),
.B2(n_937),
.Y(n_1007)
);

HB1xp67_ASAP7_75t_L g1008 ( 
.A(n_829),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_829),
.B(n_838),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_844),
.Y(n_1010)
);

O2A1O1Ixp33_ASAP7_75t_L g1011 ( 
.A1(n_858),
.A2(n_911),
.B(n_941),
.C(n_806),
.Y(n_1011)
);

AOI22xp5_ASAP7_75t_L g1012 ( 
.A1(n_793),
.A2(n_782),
.B1(n_781),
.B2(n_908),
.Y(n_1012)
);

A2O1A1Ixp33_ASAP7_75t_L g1013 ( 
.A1(n_851),
.A2(n_907),
.B(n_775),
.C(n_906),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_891),
.Y(n_1014)
);

A2O1A1Ixp33_ASAP7_75t_L g1015 ( 
.A1(n_910),
.A2(n_902),
.B(n_903),
.C(n_824),
.Y(n_1015)
);

AOI22xp5_ASAP7_75t_L g1016 ( 
.A1(n_834),
.A2(n_839),
.B1(n_767),
.B2(n_791),
.Y(n_1016)
);

AND2x4_ASAP7_75t_L g1017 ( 
.A(n_779),
.B(n_769),
.Y(n_1017)
);

O2A1O1Ixp33_ASAP7_75t_L g1018 ( 
.A1(n_890),
.A2(n_924),
.B(n_932),
.C(n_931),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_838),
.B(n_913),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_SL g1020 ( 
.A(n_882),
.B(n_936),
.Y(n_1020)
);

O2A1O1Ixp33_ASAP7_75t_L g1021 ( 
.A1(n_927),
.A2(n_905),
.B(n_832),
.C(n_916),
.Y(n_1021)
);

OAI22xp5_ASAP7_75t_L g1022 ( 
.A1(n_811),
.A2(n_883),
.B1(n_866),
.B2(n_882),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_929),
.B(n_769),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_792),
.B(n_923),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_L g1025 ( 
.A(n_811),
.B(n_883),
.Y(n_1025)
);

AOI22xp5_ASAP7_75t_L g1026 ( 
.A1(n_801),
.A2(n_848),
.B1(n_774),
.B2(n_792),
.Y(n_1026)
);

AND2x2_ASAP7_75t_L g1027 ( 
.A(n_864),
.B(n_809),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_778),
.A2(n_785),
.B(n_813),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_SL g1029 ( 
.A(n_882),
.B(n_936),
.Y(n_1029)
);

BUFx3_ASAP7_75t_L g1030 ( 
.A(n_809),
.Y(n_1030)
);

CKINVDCx20_ASAP7_75t_R g1031 ( 
.A(n_936),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_861),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_917),
.B(n_882),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_SL g1034 ( 
.A(n_845),
.B(n_879),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_875),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_778),
.A2(n_785),
.B(n_818),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_893),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_818),
.A2(n_805),
.B(n_804),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_L g1039 ( 
.A(n_879),
.B(n_917),
.Y(n_1039)
);

NAND3xp33_ASAP7_75t_L g1040 ( 
.A(n_857),
.B(n_862),
.C(n_826),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_SL g1041 ( 
.A(n_845),
.B(n_828),
.Y(n_1041)
);

O2A1O1Ixp33_ASAP7_75t_L g1042 ( 
.A1(n_918),
.A2(n_871),
.B(n_897),
.C(n_859),
.Y(n_1042)
);

NOR3xp33_ASAP7_75t_SL g1043 ( 
.A(n_795),
.B(n_797),
.C(n_794),
.Y(n_1043)
);

AND2x4_ASAP7_75t_L g1044 ( 
.A(n_942),
.B(n_874),
.Y(n_1044)
);

O2A1O1Ixp33_ASAP7_75t_L g1045 ( 
.A1(n_837),
.A2(n_816),
.B(n_943),
.C(n_934),
.Y(n_1045)
);

HB1xp67_ASAP7_75t_L g1046 ( 
.A(n_823),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_823),
.B(n_808),
.Y(n_1047)
);

NOR2xp33_ASAP7_75t_L g1048 ( 
.A(n_830),
.B(n_846),
.Y(n_1048)
);

A2O1A1Ixp33_ASAP7_75t_L g1049 ( 
.A1(n_840),
.A2(n_819),
.B(n_825),
.C(n_835),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_808),
.A2(n_842),
.B(n_835),
.Y(n_1050)
);

OAI22xp5_ASAP7_75t_L g1051 ( 
.A1(n_942),
.A2(n_825),
.B1(n_819),
.B2(n_799),
.Y(n_1051)
);

NOR3xp33_ASAP7_75t_SL g1052 ( 
.A(n_847),
.B(n_849),
.C(n_853),
.Y(n_1052)
);

AO21x1_ASAP7_75t_L g1053 ( 
.A1(n_836),
.A2(n_842),
.B(n_930),
.Y(n_1053)
);

BUFx6f_ASAP7_75t_L g1054 ( 
.A(n_942),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_SL g1055 ( 
.A(n_852),
.B(n_815),
.Y(n_1055)
);

NOR3xp33_ASAP7_75t_SL g1056 ( 
.A(n_843),
.B(n_855),
.C(n_899),
.Y(n_1056)
);

NOR2xp33_ASAP7_75t_R g1057 ( 
.A(n_889),
.B(n_878),
.Y(n_1057)
);

NOR3xp33_ASAP7_75t_SL g1058 ( 
.A(n_843),
.B(n_855),
.C(n_899),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_856),
.B(n_939),
.Y(n_1059)
);

OAI22xp5_ASAP7_75t_L g1060 ( 
.A1(n_881),
.A2(n_888),
.B1(n_836),
.B2(n_939),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_873),
.Y(n_1061)
);

BUFx2_ASAP7_75t_L g1062 ( 
.A(n_854),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_930),
.B(n_925),
.Y(n_1063)
);

AOI22xp5_ASAP7_75t_L g1064 ( 
.A1(n_904),
.A2(n_926),
.B1(n_886),
.B2(n_884),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_803),
.A2(n_925),
.B(n_921),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_L g1066 ( 
.A(n_909),
.B(n_921),
.Y(n_1066)
);

BUFx6f_ASAP7_75t_L g1067 ( 
.A(n_880),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_909),
.A2(n_884),
.B(n_887),
.Y(n_1068)
);

INVxp67_ASAP7_75t_L g1069 ( 
.A(n_894),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_784),
.A2(n_776),
.B(n_730),
.Y(n_1070)
);

AND2x2_ASAP7_75t_L g1071 ( 
.A(n_841),
.B(n_653),
.Y(n_1071)
);

AOI22xp5_ASAP7_75t_L g1072 ( 
.A1(n_892),
.A2(n_640),
.B1(n_637),
.B2(n_566),
.Y(n_1072)
);

INVx3_ASAP7_75t_L g1073 ( 
.A(n_779),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_SL g1074 ( 
.A(n_788),
.B(n_676),
.Y(n_1074)
);

AND2x4_ASAP7_75t_L g1075 ( 
.A(n_779),
.B(n_787),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_784),
.A2(n_776),
.B(n_730),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_SL g1077 ( 
.A(n_841),
.B(n_449),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_L g1078 ( 
.A(n_841),
.B(n_312),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_772),
.B(n_449),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_784),
.A2(n_776),
.B(n_730),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_1071),
.B(n_1078),
.Y(n_1081)
);

OAI21x1_ASAP7_75t_SL g1082 ( 
.A1(n_1011),
.A2(n_994),
.B(n_946),
.Y(n_1082)
);

A2O1A1Ixp33_ASAP7_75t_L g1083 ( 
.A1(n_1072),
.A2(n_976),
.B(n_945),
.C(n_953),
.Y(n_1083)
);

BUFx3_ASAP7_75t_L g1084 ( 
.A(n_958),
.Y(n_1084)
);

AO31x2_ASAP7_75t_L g1085 ( 
.A1(n_1053),
.A2(n_1066),
.A3(n_1049),
.B(n_1050),
.Y(n_1085)
);

AOI22xp33_ASAP7_75t_L g1086 ( 
.A1(n_1077),
.A2(n_1079),
.B1(n_950),
.B2(n_998),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_962),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_971),
.B(n_948),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_956),
.B(n_1014),
.Y(n_1089)
);

AO31x2_ASAP7_75t_L g1090 ( 
.A1(n_1050),
.A2(n_1007),
.A3(n_1060),
.B(n_1036),
.Y(n_1090)
);

O2A1O1Ixp33_ASAP7_75t_SL g1091 ( 
.A1(n_1015),
.A2(n_980),
.B(n_986),
.C(n_1018),
.Y(n_1091)
);

AOI22xp33_ASAP7_75t_SL g1092 ( 
.A1(n_979),
.A2(n_982),
.B1(n_981),
.B2(n_1001),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_1080),
.A2(n_1076),
.B(n_1070),
.Y(n_1093)
);

AOI22xp5_ASAP7_75t_L g1094 ( 
.A1(n_1012),
.A2(n_951),
.B1(n_1006),
.B2(n_1044),
.Y(n_1094)
);

OAI21x1_ASAP7_75t_L g1095 ( 
.A1(n_968),
.A2(n_985),
.B(n_1036),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_1080),
.A2(n_1076),
.B(n_1070),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_SL g1097 ( 
.A(n_972),
.B(n_1024),
.Y(n_1097)
);

NOR2xp33_ASAP7_75t_L g1098 ( 
.A(n_1074),
.B(n_988),
.Y(n_1098)
);

CKINVDCx14_ASAP7_75t_R g1099 ( 
.A(n_984),
.Y(n_1099)
);

INVx3_ASAP7_75t_L g1100 ( 
.A(n_1017),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_975),
.B(n_978),
.Y(n_1101)
);

AOI221x1_ASAP7_75t_L g1102 ( 
.A1(n_996),
.A2(n_949),
.B1(n_946),
.B2(n_991),
.C(n_992),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_1028),
.A2(n_1021),
.B(n_1051),
.Y(n_1103)
);

NAND3xp33_ASAP7_75t_L g1104 ( 
.A(n_989),
.B(n_1002),
.C(n_949),
.Y(n_1104)
);

O2A1O1Ixp33_ASAP7_75t_L g1105 ( 
.A1(n_952),
.A2(n_987),
.B(n_964),
.C(n_1055),
.Y(n_1105)
);

CKINVDCx11_ASAP7_75t_R g1106 ( 
.A(n_963),
.Y(n_1106)
);

OAI21x1_ASAP7_75t_L g1107 ( 
.A1(n_985),
.A2(n_1038),
.B(n_1068),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_1028),
.A2(n_1063),
.B(n_1038),
.Y(n_1108)
);

AOI22xp5_ASAP7_75t_L g1109 ( 
.A1(n_1044),
.A2(n_1062),
.B1(n_1016),
.B2(n_1048),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_983),
.B(n_955),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_1008),
.B(n_1031),
.Y(n_1111)
);

AO31x2_ASAP7_75t_L g1112 ( 
.A1(n_1013),
.A2(n_1068),
.A3(n_1065),
.B(n_966),
.Y(n_1112)
);

O2A1O1Ixp33_ASAP7_75t_L g1113 ( 
.A1(n_990),
.A2(n_996),
.B(n_970),
.C(n_1019),
.Y(n_1113)
);

O2A1O1Ixp33_ASAP7_75t_L g1114 ( 
.A1(n_1059),
.A2(n_1022),
.B(n_1045),
.C(n_1042),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_1023),
.B(n_954),
.Y(n_1115)
);

AO21x2_ASAP7_75t_L g1116 ( 
.A1(n_1057),
.A2(n_1047),
.B(n_991),
.Y(n_1116)
);

BUFx10_ASAP7_75t_L g1117 ( 
.A(n_959),
.Y(n_1117)
);

OAI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_1069),
.A2(n_1040),
.B(n_1061),
.Y(n_1118)
);

BUFx6f_ASAP7_75t_L g1119 ( 
.A(n_974),
.Y(n_1119)
);

OAI21x1_ASAP7_75t_L g1120 ( 
.A1(n_997),
.A2(n_1003),
.B(n_1064),
.Y(n_1120)
);

HB1xp67_ASAP7_75t_L g1121 ( 
.A(n_1009),
.Y(n_1121)
);

INVx3_ASAP7_75t_L g1122 ( 
.A(n_1054),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_1035),
.Y(n_1123)
);

O2A1O1Ixp33_ASAP7_75t_L g1124 ( 
.A1(n_1025),
.A2(n_1000),
.B(n_1004),
.C(n_1005),
.Y(n_1124)
);

OAI22xp5_ASAP7_75t_L g1125 ( 
.A1(n_977),
.A2(n_1026),
.B1(n_957),
.B2(n_1054),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_1067),
.A2(n_1033),
.B(n_947),
.Y(n_1126)
);

AO22x2_ASAP7_75t_L g1127 ( 
.A1(n_1037),
.A2(n_993),
.B1(n_1010),
.B2(n_1032),
.Y(n_1127)
);

O2A1O1Ixp33_ASAP7_75t_L g1128 ( 
.A1(n_965),
.A2(n_967),
.B(n_973),
.C(n_1041),
.Y(n_1128)
);

AO31x2_ASAP7_75t_L g1129 ( 
.A1(n_960),
.A2(n_1039),
.A3(n_999),
.B(n_947),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1046),
.Y(n_1130)
);

INVx1_ASAP7_75t_SL g1131 ( 
.A(n_1027),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_974),
.Y(n_1132)
);

OAI21x1_ASAP7_75t_L g1133 ( 
.A1(n_1020),
.A2(n_1029),
.B(n_1034),
.Y(n_1133)
);

INVx3_ASAP7_75t_SL g1134 ( 
.A(n_974),
.Y(n_1134)
);

NAND2xp33_ASAP7_75t_SL g1135 ( 
.A(n_995),
.B(n_1073),
.Y(n_1135)
);

BUFx4_ASAP7_75t_SL g1136 ( 
.A(n_1030),
.Y(n_1136)
);

BUFx12f_ASAP7_75t_L g1137 ( 
.A(n_959),
.Y(n_1137)
);

O2A1O1Ixp33_ASAP7_75t_L g1138 ( 
.A1(n_1056),
.A2(n_1058),
.B(n_1043),
.C(n_1052),
.Y(n_1138)
);

NOR4xp25_ASAP7_75t_L g1139 ( 
.A(n_969),
.B(n_989),
.C(n_979),
.D(n_1011),
.Y(n_1139)
);

AOI22xp5_ASAP7_75t_L g1140 ( 
.A1(n_969),
.A2(n_1072),
.B1(n_892),
.B2(n_637),
.Y(n_1140)
);

AOI22xp33_ASAP7_75t_L g1141 ( 
.A1(n_969),
.A2(n_637),
.B1(n_640),
.B2(n_789),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_1080),
.A2(n_1076),
.B(n_1070),
.Y(n_1142)
);

A2O1A1Ixp33_ASAP7_75t_L g1143 ( 
.A1(n_1072),
.A2(n_892),
.B(n_976),
.C(n_945),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_1071),
.B(n_1078),
.Y(n_1144)
);

INVx2_ASAP7_75t_SL g1145 ( 
.A(n_958),
.Y(n_1145)
);

INVxp67_ASAP7_75t_L g1146 ( 
.A(n_1071),
.Y(n_1146)
);

A2O1A1Ixp33_ASAP7_75t_L g1147 ( 
.A1(n_1072),
.A2(n_892),
.B(n_976),
.C(n_945),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_1080),
.A2(n_1076),
.B(n_1070),
.Y(n_1148)
);

INVx1_ASAP7_75t_SL g1149 ( 
.A(n_1031),
.Y(n_1149)
);

AOI21x1_ASAP7_75t_L g1150 ( 
.A1(n_1028),
.A2(n_1050),
.B(n_1068),
.Y(n_1150)
);

OAI22xp33_ASAP7_75t_L g1151 ( 
.A1(n_1072),
.A2(n_945),
.B1(n_608),
.B2(n_912),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_962),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_1080),
.A2(n_1076),
.B(n_1070),
.Y(n_1153)
);

AO31x2_ASAP7_75t_L g1154 ( 
.A1(n_1053),
.A2(n_1066),
.A3(n_1049),
.B(n_1050),
.Y(n_1154)
);

AOI22xp5_ASAP7_75t_L g1155 ( 
.A1(n_1072),
.A2(n_892),
.B1(n_637),
.B2(n_640),
.Y(n_1155)
);

BUFx6f_ASAP7_75t_L g1156 ( 
.A(n_974),
.Y(n_1156)
);

OR2x2_ASAP7_75t_L g1157 ( 
.A(n_1071),
.B(n_653),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_1071),
.B(n_1078),
.Y(n_1158)
);

OA21x2_ASAP7_75t_L g1159 ( 
.A1(n_1050),
.A2(n_1036),
.B(n_1028),
.Y(n_1159)
);

BUFx4_ASAP7_75t_SL g1160 ( 
.A(n_958),
.Y(n_1160)
);

INVx2_ASAP7_75t_SL g1161 ( 
.A(n_958),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1071),
.B(n_1078),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1071),
.B(n_1078),
.Y(n_1163)
);

AO31x2_ASAP7_75t_L g1164 ( 
.A1(n_1053),
.A2(n_1066),
.A3(n_1049),
.B(n_1050),
.Y(n_1164)
);

HB1xp67_ASAP7_75t_L g1165 ( 
.A(n_956),
.Y(n_1165)
);

O2A1O1Ixp33_ASAP7_75t_L g1166 ( 
.A1(n_945),
.A2(n_892),
.B(n_948),
.C(n_1078),
.Y(n_1166)
);

AO31x2_ASAP7_75t_L g1167 ( 
.A1(n_1053),
.A2(n_1066),
.A3(n_1049),
.B(n_1050),
.Y(n_1167)
);

A2O1A1Ixp33_ASAP7_75t_L g1168 ( 
.A1(n_1072),
.A2(n_892),
.B(n_976),
.C(n_945),
.Y(n_1168)
);

INVx2_ASAP7_75t_SL g1169 ( 
.A(n_958),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_962),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1071),
.B(n_1078),
.Y(n_1171)
);

AOI221x1_ASAP7_75t_L g1172 ( 
.A1(n_976),
.A2(n_892),
.B1(n_996),
.B2(n_949),
.C(n_946),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_1080),
.A2(n_1076),
.B(n_1070),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_1080),
.A2(n_1076),
.B(n_1070),
.Y(n_1174)
);

AOI21x1_ASAP7_75t_SL g1175 ( 
.A1(n_1063),
.A2(n_941),
.B(n_902),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_961),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_1080),
.A2(n_1076),
.B(n_1070),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1071),
.B(n_1078),
.Y(n_1178)
);

AND2x4_ASAP7_75t_L g1179 ( 
.A(n_1075),
.B(n_779),
.Y(n_1179)
);

AOI22xp5_ASAP7_75t_L g1180 ( 
.A1(n_1072),
.A2(n_892),
.B1(n_637),
.B2(n_640),
.Y(n_1180)
);

BUFx3_ASAP7_75t_L g1181 ( 
.A(n_958),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_962),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1071),
.B(n_1078),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1071),
.B(n_1078),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1071),
.B(n_1078),
.Y(n_1185)
);

OA21x2_ASAP7_75t_L g1186 ( 
.A1(n_1050),
.A2(n_1036),
.B(n_1028),
.Y(n_1186)
);

OAI21x1_ASAP7_75t_L g1187 ( 
.A1(n_968),
.A2(n_985),
.B(n_1050),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1071),
.B(n_1078),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1071),
.B(n_1078),
.Y(n_1189)
);

CKINVDCx8_ASAP7_75t_R g1190 ( 
.A(n_1014),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_1080),
.A2(n_1076),
.B(n_1070),
.Y(n_1191)
);

AO21x1_ASAP7_75t_L g1192 ( 
.A1(n_1011),
.A2(n_892),
.B(n_989),
.Y(n_1192)
);

INVx3_ASAP7_75t_L g1193 ( 
.A(n_1017),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_962),
.Y(n_1194)
);

OAI21x1_ASAP7_75t_L g1195 ( 
.A1(n_968),
.A2(n_985),
.B(n_1050),
.Y(n_1195)
);

OAI21x1_ASAP7_75t_SL g1196 ( 
.A1(n_1011),
.A2(n_994),
.B(n_946),
.Y(n_1196)
);

CKINVDCx8_ASAP7_75t_R g1197 ( 
.A(n_1014),
.Y(n_1197)
);

OAI22xp5_ASAP7_75t_L g1198 ( 
.A1(n_1072),
.A2(n_945),
.B1(n_948),
.B2(n_912),
.Y(n_1198)
);

OR2x2_ASAP7_75t_L g1199 ( 
.A(n_1071),
.B(n_653),
.Y(n_1199)
);

AOI21x1_ASAP7_75t_L g1200 ( 
.A1(n_1028),
.A2(n_1050),
.B(n_1068),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1071),
.B(n_1078),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_SL g1202 ( 
.A(n_1072),
.B(n_1079),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1071),
.B(n_1078),
.Y(n_1203)
);

BUFx12f_ASAP7_75t_L g1204 ( 
.A(n_963),
.Y(n_1204)
);

BUFx12f_ASAP7_75t_L g1205 ( 
.A(n_963),
.Y(n_1205)
);

A2O1A1Ixp33_ASAP7_75t_L g1206 ( 
.A1(n_1072),
.A2(n_892),
.B(n_976),
.C(n_945),
.Y(n_1206)
);

OAI21x1_ASAP7_75t_L g1207 ( 
.A1(n_968),
.A2(n_985),
.B(n_1050),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_SL g1208 ( 
.A1(n_1007),
.A2(n_942),
.B(n_1015),
.Y(n_1208)
);

OAI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1072),
.A2(n_892),
.B(n_945),
.Y(n_1209)
);

INVx5_ASAP7_75t_L g1210 ( 
.A(n_969),
.Y(n_1210)
);

NOR2xp33_ASAP7_75t_L g1211 ( 
.A(n_1078),
.B(n_1072),
.Y(n_1211)
);

BUFx8_ASAP7_75t_L g1212 ( 
.A(n_963),
.Y(n_1212)
);

NOR4xp25_ASAP7_75t_L g1213 ( 
.A(n_989),
.B(n_979),
.C(n_1011),
.D(n_892),
.Y(n_1213)
);

O2A1O1Ixp33_ASAP7_75t_SL g1214 ( 
.A1(n_945),
.A2(n_870),
.B(n_1015),
.C(n_1079),
.Y(n_1214)
);

BUFx12f_ASAP7_75t_L g1215 ( 
.A(n_1106),
.Y(n_1215)
);

OAI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1211),
.A2(n_1147),
.B(n_1143),
.Y(n_1216)
);

HB1xp67_ASAP7_75t_L g1217 ( 
.A(n_1085),
.Y(n_1217)
);

AOI22xp33_ASAP7_75t_L g1218 ( 
.A1(n_1209),
.A2(n_1198),
.B1(n_1180),
.B2(n_1155),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1087),
.Y(n_1219)
);

AOI22xp33_ASAP7_75t_SL g1220 ( 
.A1(n_1125),
.A2(n_1088),
.B1(n_1151),
.B2(n_1144),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1152),
.Y(n_1221)
);

AOI22xp33_ASAP7_75t_L g1222 ( 
.A1(n_1155),
.A2(n_1180),
.B1(n_1141),
.B2(n_1140),
.Y(n_1222)
);

BUFx2_ASAP7_75t_L g1223 ( 
.A(n_1137),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1166),
.B(n_1168),
.Y(n_1224)
);

CKINVDCx11_ASAP7_75t_R g1225 ( 
.A(n_1204),
.Y(n_1225)
);

INVx8_ASAP7_75t_L g1226 ( 
.A(n_1205),
.Y(n_1226)
);

AOI22xp33_ASAP7_75t_L g1227 ( 
.A1(n_1140),
.A2(n_1092),
.B1(n_1202),
.B2(n_1192),
.Y(n_1227)
);

CKINVDCx11_ASAP7_75t_R g1228 ( 
.A(n_1190),
.Y(n_1228)
);

AOI22xp33_ASAP7_75t_L g1229 ( 
.A1(n_1081),
.A2(n_1184),
.B1(n_1158),
.B2(n_1162),
.Y(n_1229)
);

CKINVDCx11_ASAP7_75t_R g1230 ( 
.A(n_1197),
.Y(n_1230)
);

AOI22xp33_ASAP7_75t_SL g1231 ( 
.A1(n_1163),
.A2(n_1188),
.B1(n_1189),
.B2(n_1185),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1170),
.Y(n_1232)
);

AOI22xp5_ASAP7_75t_L g1233 ( 
.A1(n_1206),
.A2(n_1183),
.B1(n_1178),
.B2(n_1171),
.Y(n_1233)
);

OAI21xp33_ASAP7_75t_L g1234 ( 
.A1(n_1083),
.A2(n_1213),
.B(n_1201),
.Y(n_1234)
);

CKINVDCx8_ASAP7_75t_R g1235 ( 
.A(n_1132),
.Y(n_1235)
);

INVx1_ASAP7_75t_SL g1236 ( 
.A(n_1160),
.Y(n_1236)
);

INVx6_ASAP7_75t_L g1237 ( 
.A(n_1119),
.Y(n_1237)
);

BUFx4f_ASAP7_75t_SL g1238 ( 
.A(n_1212),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1182),
.Y(n_1239)
);

AOI22xp33_ASAP7_75t_L g1240 ( 
.A1(n_1203),
.A2(n_1176),
.B1(n_1086),
.B2(n_1131),
.Y(n_1240)
);

INVx6_ASAP7_75t_L g1241 ( 
.A(n_1119),
.Y(n_1241)
);

OAI22xp33_ASAP7_75t_L g1242 ( 
.A1(n_1146),
.A2(n_1109),
.B1(n_1199),
.B2(n_1157),
.Y(n_1242)
);

AOI22xp33_ASAP7_75t_SL g1243 ( 
.A1(n_1082),
.A2(n_1196),
.B1(n_1104),
.B2(n_1210),
.Y(n_1243)
);

OAI22xp5_ASAP7_75t_L g1244 ( 
.A1(n_1104),
.A2(n_1109),
.B1(n_1165),
.B2(n_1208),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1110),
.B(n_1131),
.Y(n_1245)
);

AOI22xp33_ASAP7_75t_L g1246 ( 
.A1(n_1094),
.A2(n_1127),
.B1(n_1123),
.B2(n_1130),
.Y(n_1246)
);

INVx6_ASAP7_75t_L g1247 ( 
.A(n_1119),
.Y(n_1247)
);

CKINVDCx20_ASAP7_75t_R g1248 ( 
.A(n_1212),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1194),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1121),
.Y(n_1250)
);

INVx5_ASAP7_75t_L g1251 ( 
.A(n_1210),
.Y(n_1251)
);

AOI22xp33_ASAP7_75t_L g1252 ( 
.A1(n_1094),
.A2(n_1127),
.B1(n_1084),
.B2(n_1181),
.Y(n_1252)
);

CKINVDCx11_ASAP7_75t_R g1253 ( 
.A(n_1149),
.Y(n_1253)
);

BUFx4f_ASAP7_75t_SL g1254 ( 
.A(n_1134),
.Y(n_1254)
);

OAI22xp5_ASAP7_75t_L g1255 ( 
.A1(n_1115),
.A2(n_1098),
.B1(n_1103),
.B2(n_1138),
.Y(n_1255)
);

INVx1_ASAP7_75t_SL g1256 ( 
.A(n_1149),
.Y(n_1256)
);

AND2x2_ASAP7_75t_L g1257 ( 
.A(n_1145),
.B(n_1161),
.Y(n_1257)
);

OAI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1089),
.A2(n_1124),
.B1(n_1193),
.B2(n_1100),
.Y(n_1258)
);

OAI22xp33_ASAP7_75t_L g1259 ( 
.A1(n_1172),
.A2(n_1210),
.B1(n_1102),
.B2(n_1193),
.Y(n_1259)
);

INVx3_ASAP7_75t_L g1260 ( 
.A(n_1179),
.Y(n_1260)
);

CKINVDCx20_ASAP7_75t_R g1261 ( 
.A(n_1099),
.Y(n_1261)
);

INVx2_ASAP7_75t_SL g1262 ( 
.A(n_1136),
.Y(n_1262)
);

INVx4_ASAP7_75t_L g1263 ( 
.A(n_1156),
.Y(n_1263)
);

AOI22xp33_ASAP7_75t_L g1264 ( 
.A1(n_1169),
.A2(n_1097),
.B1(n_1111),
.B2(n_1122),
.Y(n_1264)
);

AOI22xp33_ASAP7_75t_SL g1265 ( 
.A1(n_1213),
.A2(n_1139),
.B1(n_1120),
.B2(n_1118),
.Y(n_1265)
);

OAI22xp33_ASAP7_75t_L g1266 ( 
.A1(n_1100),
.A2(n_1122),
.B1(n_1191),
.B2(n_1177),
.Y(n_1266)
);

BUFx12f_ASAP7_75t_L g1267 ( 
.A(n_1117),
.Y(n_1267)
);

BUFx4f_ASAP7_75t_L g1268 ( 
.A(n_1156),
.Y(n_1268)
);

AOI22xp33_ASAP7_75t_L g1269 ( 
.A1(n_1116),
.A2(n_1139),
.B1(n_1126),
.B2(n_1174),
.Y(n_1269)
);

INVx2_ASAP7_75t_SL g1270 ( 
.A(n_1117),
.Y(n_1270)
);

OAI22xp33_ASAP7_75t_L g1271 ( 
.A1(n_1093),
.A2(n_1142),
.B1(n_1173),
.B2(n_1148),
.Y(n_1271)
);

INVxp67_ASAP7_75t_L g1272 ( 
.A(n_1133),
.Y(n_1272)
);

CKINVDCx5p33_ASAP7_75t_R g1273 ( 
.A(n_1135),
.Y(n_1273)
);

BUFx12f_ASAP7_75t_SL g1274 ( 
.A(n_1091),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1128),
.Y(n_1275)
);

AOI22xp33_ASAP7_75t_SL g1276 ( 
.A1(n_1214),
.A2(n_1153),
.B1(n_1096),
.B2(n_1186),
.Y(n_1276)
);

AOI22xp5_ASAP7_75t_L g1277 ( 
.A1(n_1159),
.A2(n_1186),
.B1(n_1108),
.B2(n_1095),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1129),
.Y(n_1278)
);

OAI21xp5_ASAP7_75t_SL g1279 ( 
.A1(n_1114),
.A2(n_1105),
.B(n_1113),
.Y(n_1279)
);

OAI22xp33_ASAP7_75t_L g1280 ( 
.A1(n_1159),
.A2(n_1200),
.B1(n_1150),
.B2(n_1175),
.Y(n_1280)
);

INVx3_ASAP7_75t_L g1281 ( 
.A(n_1085),
.Y(n_1281)
);

AND2x2_ASAP7_75t_L g1282 ( 
.A(n_1154),
.B(n_1167),
.Y(n_1282)
);

OAI22xp5_ASAP7_75t_L g1283 ( 
.A1(n_1090),
.A2(n_1164),
.B1(n_1167),
.B2(n_1112),
.Y(n_1283)
);

AOI22xp33_ASAP7_75t_L g1284 ( 
.A1(n_1107),
.A2(n_1187),
.B1(n_1195),
.B2(n_1207),
.Y(n_1284)
);

BUFx2_ASAP7_75t_L g1285 ( 
.A(n_1164),
.Y(n_1285)
);

OAI22xp5_ASAP7_75t_L g1286 ( 
.A1(n_1090),
.A2(n_1164),
.B1(n_1167),
.B2(n_1112),
.Y(n_1286)
);

OAI22xp33_ASAP7_75t_L g1287 ( 
.A1(n_1112),
.A2(n_1155),
.B1(n_1180),
.B2(n_1198),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1101),
.Y(n_1288)
);

AOI22xp33_ASAP7_75t_L g1289 ( 
.A1(n_1209),
.A2(n_1211),
.B1(n_1198),
.B2(n_1155),
.Y(n_1289)
);

AOI22xp5_ASAP7_75t_L g1290 ( 
.A1(n_1211),
.A2(n_1155),
.B1(n_1180),
.B2(n_1072),
.Y(n_1290)
);

OAI22xp5_ASAP7_75t_SL g1291 ( 
.A1(n_1211),
.A2(n_1072),
.B1(n_1180),
.B2(n_1155),
.Y(n_1291)
);

BUFx3_ASAP7_75t_L g1292 ( 
.A(n_1084),
.Y(n_1292)
);

CKINVDCx20_ASAP7_75t_R g1293 ( 
.A(n_1106),
.Y(n_1293)
);

AOI22xp33_ASAP7_75t_L g1294 ( 
.A1(n_1209),
.A2(n_1211),
.B1(n_1198),
.B2(n_1155),
.Y(n_1294)
);

BUFx3_ASAP7_75t_L g1295 ( 
.A(n_1084),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1101),
.Y(n_1296)
);

INVx5_ASAP7_75t_L g1297 ( 
.A(n_1210),
.Y(n_1297)
);

BUFx10_ASAP7_75t_L g1298 ( 
.A(n_1098),
.Y(n_1298)
);

AOI22xp33_ASAP7_75t_L g1299 ( 
.A1(n_1211),
.A2(n_640),
.B1(n_637),
.B2(n_1209),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1101),
.Y(n_1300)
);

OAI22xp5_ASAP7_75t_L g1301 ( 
.A1(n_1155),
.A2(n_1180),
.B1(n_1211),
.B2(n_1147),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1088),
.B(n_1198),
.Y(n_1302)
);

INVx4_ASAP7_75t_L g1303 ( 
.A(n_1134),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1101),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_SL g1305 ( 
.A(n_1211),
.B(n_1140),
.Y(n_1305)
);

AOI22xp33_ASAP7_75t_SL g1306 ( 
.A1(n_1211),
.A2(n_1209),
.B1(n_1198),
.B2(n_608),
.Y(n_1306)
);

BUFx3_ASAP7_75t_L g1307 ( 
.A(n_1084),
.Y(n_1307)
);

CKINVDCx6p67_ASAP7_75t_R g1308 ( 
.A(n_1106),
.Y(n_1308)
);

BUFx2_ASAP7_75t_L g1309 ( 
.A(n_1137),
.Y(n_1309)
);

INVx1_ASAP7_75t_SL g1310 ( 
.A(n_1160),
.Y(n_1310)
);

AOI22xp33_ASAP7_75t_L g1311 ( 
.A1(n_1211),
.A2(n_640),
.B1(n_637),
.B2(n_1209),
.Y(n_1311)
);

AOI22xp33_ASAP7_75t_L g1312 ( 
.A1(n_1209),
.A2(n_1211),
.B1(n_1198),
.B2(n_1155),
.Y(n_1312)
);

CKINVDCx5p33_ASAP7_75t_R g1313 ( 
.A(n_1106),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1081),
.B(n_1144),
.Y(n_1314)
);

BUFx2_ASAP7_75t_SL g1315 ( 
.A(n_1190),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_SL g1316 ( 
.A1(n_1211),
.A2(n_1209),
.B1(n_1198),
.B2(n_608),
.Y(n_1316)
);

AOI22xp33_ASAP7_75t_L g1317 ( 
.A1(n_1209),
.A2(n_1211),
.B1(n_1198),
.B2(n_1155),
.Y(n_1317)
);

AOI22xp33_ASAP7_75t_L g1318 ( 
.A1(n_1211),
.A2(n_640),
.B1(n_637),
.B2(n_1209),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1101),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1101),
.Y(n_1320)
);

AOI22xp33_ASAP7_75t_L g1321 ( 
.A1(n_1211),
.A2(n_640),
.B1(n_637),
.B2(n_1209),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1101),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1101),
.Y(n_1323)
);

OAI22xp5_ASAP7_75t_L g1324 ( 
.A1(n_1155),
.A2(n_1180),
.B1(n_1211),
.B2(n_1147),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1088),
.B(n_1198),
.Y(n_1325)
);

OAI21x1_ASAP7_75t_L g1326 ( 
.A1(n_1269),
.A2(n_1286),
.B(n_1283),
.Y(n_1326)
);

HB1xp67_ASAP7_75t_L g1327 ( 
.A(n_1250),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1217),
.Y(n_1328)
);

OAI21xp5_ASAP7_75t_L g1329 ( 
.A1(n_1301),
.A2(n_1324),
.B(n_1290),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1282),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1302),
.B(n_1325),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1289),
.B(n_1294),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1285),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1219),
.Y(n_1334)
);

OR2x2_ASAP7_75t_L g1335 ( 
.A(n_1305),
.B(n_1281),
.Y(n_1335)
);

AND2x4_ASAP7_75t_L g1336 ( 
.A(n_1251),
.B(n_1297),
.Y(n_1336)
);

OAI21x1_ASAP7_75t_L g1337 ( 
.A1(n_1269),
.A2(n_1284),
.B(n_1277),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1221),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1232),
.Y(n_1339)
);

AO21x1_ASAP7_75t_SL g1340 ( 
.A1(n_1218),
.A2(n_1289),
.B(n_1317),
.Y(n_1340)
);

CKINVDCx5p33_ASAP7_75t_R g1341 ( 
.A(n_1228),
.Y(n_1341)
);

INVx3_ASAP7_75t_L g1342 ( 
.A(n_1281),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1239),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1249),
.Y(n_1344)
);

AO21x2_ASAP7_75t_L g1345 ( 
.A1(n_1287),
.A2(n_1278),
.B(n_1280),
.Y(n_1345)
);

INVx1_ASAP7_75t_SL g1346 ( 
.A(n_1245),
.Y(n_1346)
);

AND2x4_ASAP7_75t_L g1347 ( 
.A(n_1251),
.B(n_1297),
.Y(n_1347)
);

OAI21x1_ASAP7_75t_L g1348 ( 
.A1(n_1244),
.A2(n_1279),
.B(n_1275),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1272),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1265),
.B(n_1216),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1272),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1266),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1265),
.B(n_1294),
.Y(n_1353)
);

NOR2xp33_ASAP7_75t_L g1354 ( 
.A(n_1291),
.B(n_1236),
.Y(n_1354)
);

OAI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1312),
.A2(n_1317),
.B(n_1218),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1266),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1280),
.Y(n_1357)
);

OA21x2_ASAP7_75t_L g1358 ( 
.A1(n_1224),
.A2(n_1234),
.B(n_1222),
.Y(n_1358)
);

BUFx2_ASAP7_75t_L g1359 ( 
.A(n_1274),
.Y(n_1359)
);

OAI22xp33_ASAP7_75t_L g1360 ( 
.A1(n_1233),
.A2(n_1287),
.B1(n_1242),
.B2(n_1255),
.Y(n_1360)
);

NOR2xp33_ASAP7_75t_L g1361 ( 
.A(n_1310),
.B(n_1253),
.Y(n_1361)
);

OAI21x1_ASAP7_75t_L g1362 ( 
.A1(n_1258),
.A2(n_1252),
.B(n_1227),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_SL g1363 ( 
.A(n_1312),
.B(n_1220),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1288),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1314),
.B(n_1296),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1300),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1304),
.B(n_1319),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1320),
.B(n_1322),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1323),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1271),
.Y(n_1370)
);

HB1xp67_ASAP7_75t_L g1371 ( 
.A(n_1256),
.Y(n_1371)
);

INVx3_ASAP7_75t_L g1372 ( 
.A(n_1273),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1271),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1276),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1276),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1259),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1259),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1243),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1242),
.B(n_1316),
.Y(n_1379)
);

INVxp33_ASAP7_75t_L g1380 ( 
.A(n_1230),
.Y(n_1380)
);

INVxp67_ASAP7_75t_SL g1381 ( 
.A(n_1246),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1243),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1220),
.Y(n_1383)
);

INVx2_ASAP7_75t_SL g1384 ( 
.A(n_1298),
.Y(n_1384)
);

BUFx2_ASAP7_75t_L g1385 ( 
.A(n_1267),
.Y(n_1385)
);

CKINVDCx20_ASAP7_75t_R g1386 ( 
.A(n_1293),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1240),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1306),
.B(n_1316),
.Y(n_1388)
);

OA21x2_ASAP7_75t_L g1389 ( 
.A1(n_1299),
.A2(n_1318),
.B(n_1311),
.Y(n_1389)
);

HB1xp67_ASAP7_75t_L g1390 ( 
.A(n_1260),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1229),
.B(n_1306),
.Y(n_1391)
);

INVx2_ASAP7_75t_L g1392 ( 
.A(n_1260),
.Y(n_1392)
);

AO31x2_ASAP7_75t_L g1393 ( 
.A1(n_1263),
.A2(n_1321),
.A3(n_1231),
.B(n_1309),
.Y(n_1393)
);

BUFx12f_ASAP7_75t_L g1394 ( 
.A(n_1225),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1229),
.B(n_1231),
.Y(n_1395)
);

BUFx2_ASAP7_75t_L g1396 ( 
.A(n_1270),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1327),
.B(n_1257),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1331),
.B(n_1264),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1334),
.Y(n_1399)
);

CKINVDCx8_ASAP7_75t_R g1400 ( 
.A(n_1341),
.Y(n_1400)
);

BUFx3_ASAP7_75t_L g1401 ( 
.A(n_1396),
.Y(n_1401)
);

AOI221xp5_ASAP7_75t_L g1402 ( 
.A1(n_1350),
.A2(n_1383),
.B1(n_1360),
.B2(n_1363),
.C(n_1388),
.Y(n_1402)
);

NOR2xp33_ASAP7_75t_R g1403 ( 
.A(n_1394),
.B(n_1238),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1365),
.B(n_1307),
.Y(n_1404)
);

AOI221xp5_ASAP7_75t_L g1405 ( 
.A1(n_1350),
.A2(n_1292),
.B1(n_1295),
.B2(n_1313),
.C(n_1262),
.Y(n_1405)
);

O2A1O1Ixp33_ASAP7_75t_L g1406 ( 
.A1(n_1329),
.A2(n_1223),
.B(n_1261),
.C(n_1248),
.Y(n_1406)
);

OAI21xp5_ASAP7_75t_L g1407 ( 
.A1(n_1348),
.A2(n_1268),
.B(n_1303),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1371),
.B(n_1315),
.Y(n_1408)
);

INVxp67_ASAP7_75t_L g1409 ( 
.A(n_1349),
.Y(n_1409)
);

OA21x2_ASAP7_75t_L g1410 ( 
.A1(n_1337),
.A2(n_1241),
.B(n_1247),
.Y(n_1410)
);

AND2x2_ASAP7_75t_SL g1411 ( 
.A(n_1353),
.B(n_1308),
.Y(n_1411)
);

AND2x6_ASAP7_75t_L g1412 ( 
.A(n_1336),
.B(n_1347),
.Y(n_1412)
);

OAI21xp5_ASAP7_75t_L g1413 ( 
.A1(n_1348),
.A2(n_1254),
.B(n_1235),
.Y(n_1413)
);

INVxp67_ASAP7_75t_L g1414 ( 
.A(n_1349),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1331),
.B(n_1237),
.Y(n_1415)
);

INVx1_ASAP7_75t_SL g1416 ( 
.A(n_1359),
.Y(n_1416)
);

AOI22xp5_ASAP7_75t_L g1417 ( 
.A1(n_1383),
.A2(n_1215),
.B1(n_1241),
.B2(n_1247),
.Y(n_1417)
);

OAI22xp5_ASAP7_75t_L g1418 ( 
.A1(n_1332),
.A2(n_1226),
.B1(n_1238),
.B2(n_1355),
.Y(n_1418)
);

NOR2xp33_ASAP7_75t_L g1419 ( 
.A(n_1389),
.B(n_1332),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1354),
.B(n_1359),
.Y(n_1420)
);

O2A1O1Ixp33_ASAP7_75t_L g1421 ( 
.A1(n_1355),
.A2(n_1388),
.B(n_1379),
.C(n_1389),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1346),
.B(n_1358),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1390),
.B(n_1392),
.Y(n_1423)
);

INVxp67_ASAP7_75t_L g1424 ( 
.A(n_1351),
.Y(n_1424)
);

AO32x2_ASAP7_75t_L g1425 ( 
.A1(n_1384),
.A2(n_1330),
.A3(n_1393),
.B1(n_1381),
.B2(n_1335),
.Y(n_1425)
);

OAI22xp5_ASAP7_75t_L g1426 ( 
.A1(n_1379),
.A2(n_1358),
.B1(n_1391),
.B2(n_1378),
.Y(n_1426)
);

OAI221xp5_ASAP7_75t_L g1427 ( 
.A1(n_1358),
.A2(n_1391),
.B1(n_1377),
.B2(n_1376),
.C(n_1395),
.Y(n_1427)
);

AOI22xp33_ASAP7_75t_L g1428 ( 
.A1(n_1395),
.A2(n_1340),
.B1(n_1387),
.B2(n_1362),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1367),
.B(n_1368),
.Y(n_1429)
);

AOI221xp5_ASAP7_75t_L g1430 ( 
.A1(n_1376),
.A2(n_1377),
.B1(n_1374),
.B2(n_1375),
.C(n_1369),
.Y(n_1430)
);

A2O1A1Ixp33_ASAP7_75t_L g1431 ( 
.A1(n_1362),
.A2(n_1378),
.B(n_1382),
.C(n_1375),
.Y(n_1431)
);

AO32x1_ASAP7_75t_L g1432 ( 
.A1(n_1382),
.A2(n_1374),
.A3(n_1357),
.B1(n_1333),
.B2(n_1328),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1367),
.B(n_1368),
.Y(n_1433)
);

CKINVDCx20_ASAP7_75t_R g1434 ( 
.A(n_1386),
.Y(n_1434)
);

A2O1A1Ixp33_ASAP7_75t_L g1435 ( 
.A1(n_1326),
.A2(n_1356),
.B(n_1352),
.C(n_1340),
.Y(n_1435)
);

OAI21xp33_ASAP7_75t_L g1436 ( 
.A1(n_1370),
.A2(n_1373),
.B(n_1352),
.Y(n_1436)
);

CKINVDCx14_ASAP7_75t_R g1437 ( 
.A(n_1394),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1372),
.B(n_1338),
.Y(n_1438)
);

CKINVDCx5p33_ASAP7_75t_R g1439 ( 
.A(n_1394),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1399),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1438),
.B(n_1345),
.Y(n_1441)
);

AOI22xp33_ASAP7_75t_L g1442 ( 
.A1(n_1402),
.A2(n_1387),
.B1(n_1345),
.B2(n_1364),
.Y(n_1442)
);

BUFx3_ASAP7_75t_L g1443 ( 
.A(n_1412),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1425),
.B(n_1345),
.Y(n_1444)
);

OR2x2_ASAP7_75t_L g1445 ( 
.A(n_1429),
.B(n_1393),
.Y(n_1445)
);

AND2x4_ASAP7_75t_L g1446 ( 
.A(n_1412),
.B(n_1342),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1425),
.B(n_1337),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1425),
.B(n_1337),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1425),
.B(n_1326),
.Y(n_1449)
);

OR2x2_ASAP7_75t_L g1450 ( 
.A(n_1433),
.B(n_1393),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1423),
.B(n_1326),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1419),
.B(n_1366),
.Y(n_1452)
);

OAI21xp5_ASAP7_75t_SL g1453 ( 
.A1(n_1421),
.A2(n_1380),
.B(n_1372),
.Y(n_1453)
);

OAI22xp5_ASAP7_75t_SL g1454 ( 
.A1(n_1437),
.A2(n_1372),
.B1(n_1361),
.B2(n_1385),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1409),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1409),
.Y(n_1456)
);

AND2x2_ASAP7_75t_SL g1457 ( 
.A(n_1419),
.B(n_1347),
.Y(n_1457)
);

OR2x2_ASAP7_75t_L g1458 ( 
.A(n_1422),
.B(n_1393),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1414),
.B(n_1424),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1410),
.B(n_1344),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1414),
.Y(n_1461)
);

AOI22xp33_ASAP7_75t_L g1462 ( 
.A1(n_1428),
.A2(n_1426),
.B1(n_1427),
.B2(n_1411),
.Y(n_1462)
);

NAND2x1_ASAP7_75t_L g1463 ( 
.A(n_1446),
.B(n_1412),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1441),
.B(n_1451),
.Y(n_1464)
);

OR2x2_ASAP7_75t_L g1465 ( 
.A(n_1445),
.B(n_1393),
.Y(n_1465)
);

AOI21xp5_ASAP7_75t_L g1466 ( 
.A1(n_1453),
.A2(n_1432),
.B(n_1435),
.Y(n_1466)
);

OR2x2_ASAP7_75t_L g1467 ( 
.A(n_1445),
.B(n_1401),
.Y(n_1467)
);

OAI22xp5_ASAP7_75t_L g1468 ( 
.A1(n_1462),
.A2(n_1428),
.B1(n_1435),
.B2(n_1431),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1440),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1440),
.Y(n_1470)
);

HB1xp67_ASAP7_75t_L g1471 ( 
.A(n_1455),
.Y(n_1471)
);

AOI22xp33_ASAP7_75t_L g1472 ( 
.A1(n_1442),
.A2(n_1411),
.B1(n_1430),
.B2(n_1398),
.Y(n_1472)
);

OAI21xp5_ASAP7_75t_L g1473 ( 
.A1(n_1453),
.A2(n_1431),
.B(n_1418),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1460),
.Y(n_1474)
);

AND2x4_ASAP7_75t_L g1475 ( 
.A(n_1443),
.B(n_1412),
.Y(n_1475)
);

INVx3_ASAP7_75t_L g1476 ( 
.A(n_1443),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1452),
.B(n_1339),
.Y(n_1477)
);

HB1xp67_ASAP7_75t_L g1478 ( 
.A(n_1455),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1440),
.Y(n_1479)
);

INVx3_ASAP7_75t_L g1480 ( 
.A(n_1443),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1452),
.B(n_1339),
.Y(n_1481)
);

OAI221xp5_ASAP7_75t_L g1482 ( 
.A1(n_1462),
.A2(n_1436),
.B1(n_1405),
.B2(n_1413),
.C(n_1417),
.Y(n_1482)
);

INVxp67_ASAP7_75t_L g1483 ( 
.A(n_1455),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1451),
.B(n_1397),
.Y(n_1484)
);

AOI22xp33_ASAP7_75t_SL g1485 ( 
.A1(n_1444),
.A2(n_1437),
.B1(n_1420),
.B2(n_1404),
.Y(n_1485)
);

AO21x2_ASAP7_75t_L g1486 ( 
.A1(n_1444),
.A2(n_1447),
.B(n_1448),
.Y(n_1486)
);

NAND3xp33_ASAP7_75t_L g1487 ( 
.A(n_1444),
.B(n_1415),
.C(n_1406),
.Y(n_1487)
);

HB1xp67_ASAP7_75t_L g1488 ( 
.A(n_1456),
.Y(n_1488)
);

NAND3xp33_ASAP7_75t_L g1489 ( 
.A(n_1449),
.B(n_1442),
.C(n_1448),
.Y(n_1489)
);

OR2x2_ASAP7_75t_L g1490 ( 
.A(n_1445),
.B(n_1343),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1456),
.B(n_1344),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1464),
.B(n_1449),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1469),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1469),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1470),
.Y(n_1495)
);

BUFx3_ASAP7_75t_L g1496 ( 
.A(n_1463),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1490),
.B(n_1461),
.Y(n_1497)
);

OR2x2_ASAP7_75t_L g1498 ( 
.A(n_1490),
.B(n_1450),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1464),
.B(n_1457),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1470),
.Y(n_1500)
);

INVx2_ASAP7_75t_SL g1501 ( 
.A(n_1463),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1483),
.B(n_1461),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1479),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1483),
.B(n_1461),
.Y(n_1504)
);

INVx1_ASAP7_75t_SL g1505 ( 
.A(n_1467),
.Y(n_1505)
);

BUFx2_ASAP7_75t_L g1506 ( 
.A(n_1476),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1477),
.B(n_1459),
.Y(n_1507)
);

NOR2xp33_ASAP7_75t_L g1508 ( 
.A(n_1487),
.B(n_1416),
.Y(n_1508)
);

INVx2_ASAP7_75t_SL g1509 ( 
.A(n_1475),
.Y(n_1509)
);

HB1xp67_ASAP7_75t_L g1510 ( 
.A(n_1471),
.Y(n_1510)
);

OR2x2_ASAP7_75t_L g1511 ( 
.A(n_1486),
.B(n_1477),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1479),
.Y(n_1512)
);

INVxp67_ASAP7_75t_L g1513 ( 
.A(n_1487),
.Y(n_1513)
);

BUFx3_ASAP7_75t_L g1514 ( 
.A(n_1475),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1481),
.B(n_1459),
.Y(n_1515)
);

INVx2_ASAP7_75t_SL g1516 ( 
.A(n_1475),
.Y(n_1516)
);

INVx3_ASAP7_75t_L g1517 ( 
.A(n_1475),
.Y(n_1517)
);

INVx3_ASAP7_75t_L g1518 ( 
.A(n_1474),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1493),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1513),
.B(n_1484),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1518),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1493),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1493),
.Y(n_1523)
);

OAI22xp5_ASAP7_75t_L g1524 ( 
.A1(n_1513),
.A2(n_1473),
.B1(n_1466),
.B2(n_1468),
.Y(n_1524)
);

NOR2xp33_ASAP7_75t_L g1525 ( 
.A(n_1508),
.B(n_1439),
.Y(n_1525)
);

OR2x2_ASAP7_75t_L g1526 ( 
.A(n_1507),
.B(n_1481),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1499),
.B(n_1476),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1494),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1499),
.B(n_1476),
.Y(n_1529)
);

INVx3_ASAP7_75t_L g1530 ( 
.A(n_1496),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1494),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1508),
.B(n_1484),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1494),
.Y(n_1533)
);

AOI31xp33_ASAP7_75t_L g1534 ( 
.A1(n_1501),
.A2(n_1473),
.A3(n_1439),
.B(n_1466),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1495),
.Y(n_1535)
);

INVx2_ASAP7_75t_SL g1536 ( 
.A(n_1514),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1495),
.Y(n_1537)
);

OR2x2_ASAP7_75t_L g1538 ( 
.A(n_1507),
.B(n_1471),
.Y(n_1538)
);

OR2x2_ASAP7_75t_L g1539 ( 
.A(n_1515),
.B(n_1478),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1495),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1500),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1500),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1499),
.B(n_1476),
.Y(n_1543)
);

AND2x4_ASAP7_75t_L g1544 ( 
.A(n_1514),
.B(n_1476),
.Y(n_1544)
);

HB1xp67_ASAP7_75t_L g1545 ( 
.A(n_1505),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1514),
.B(n_1480),
.Y(n_1546)
);

OR2x2_ASAP7_75t_L g1547 ( 
.A(n_1515),
.B(n_1478),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1505),
.B(n_1484),
.Y(n_1548)
);

OR2x2_ASAP7_75t_L g1549 ( 
.A(n_1498),
.B(n_1488),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1503),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1503),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1512),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1512),
.Y(n_1553)
);

OR2x2_ASAP7_75t_L g1554 ( 
.A(n_1498),
.B(n_1488),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1514),
.B(n_1480),
.Y(n_1555)
);

INVx2_ASAP7_75t_L g1556 ( 
.A(n_1518),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1518),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1518),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1519),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1521),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1527),
.B(n_1529),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1519),
.Y(n_1562)
);

HB1xp67_ASAP7_75t_L g1563 ( 
.A(n_1545),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1527),
.B(n_1517),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1528),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1529),
.B(n_1517),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1524),
.B(n_1510),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1521),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1543),
.B(n_1517),
.Y(n_1569)
);

NOR2x1p5_ASAP7_75t_SL g1570 ( 
.A(n_1556),
.B(n_1511),
.Y(n_1570)
);

NOR3xp33_ASAP7_75t_SL g1571 ( 
.A(n_1525),
.B(n_1454),
.C(n_1482),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1528),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1520),
.B(n_1510),
.Y(n_1573)
);

INVx2_ASAP7_75t_SL g1574 ( 
.A(n_1544),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1526),
.B(n_1502),
.Y(n_1575)
);

INVx3_ASAP7_75t_L g1576 ( 
.A(n_1544),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1531),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1526),
.B(n_1502),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1543),
.B(n_1517),
.Y(n_1579)
);

INVx1_ASAP7_75t_SL g1580 ( 
.A(n_1530),
.Y(n_1580)
);

INVx3_ASAP7_75t_L g1581 ( 
.A(n_1544),
.Y(n_1581)
);

INVxp67_ASAP7_75t_L g1582 ( 
.A(n_1536),
.Y(n_1582)
);

AOI21xp5_ASAP7_75t_L g1583 ( 
.A1(n_1534),
.A2(n_1468),
.B(n_1489),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1531),
.Y(n_1584)
);

O2A1O1Ixp5_ASAP7_75t_R g1585 ( 
.A1(n_1532),
.A2(n_1504),
.B(n_1497),
.C(n_1491),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1533),
.Y(n_1586)
);

OR2x2_ASAP7_75t_L g1587 ( 
.A(n_1538),
.B(n_1539),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1546),
.B(n_1517),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1546),
.B(n_1517),
.Y(n_1589)
);

HB1xp67_ASAP7_75t_L g1590 ( 
.A(n_1533),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1535),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1555),
.B(n_1509),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1556),
.Y(n_1593)
);

OAI221xp5_ASAP7_75t_SL g1594 ( 
.A1(n_1567),
.A2(n_1482),
.B1(n_1472),
.B2(n_1511),
.C(n_1554),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1563),
.B(n_1536),
.Y(n_1595)
);

OAI221xp5_ASAP7_75t_L g1596 ( 
.A1(n_1583),
.A2(n_1571),
.B1(n_1567),
.B2(n_1489),
.C(n_1585),
.Y(n_1596)
);

AND2x4_ASAP7_75t_SL g1597 ( 
.A(n_1571),
.B(n_1434),
.Y(n_1597)
);

AOI22xp5_ASAP7_75t_L g1598 ( 
.A1(n_1583),
.A2(n_1472),
.B1(n_1447),
.B2(n_1448),
.Y(n_1598)
);

AOI21xp5_ASAP7_75t_L g1599 ( 
.A1(n_1585),
.A2(n_1563),
.B(n_1575),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1582),
.B(n_1538),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1564),
.Y(n_1601)
);

OAI22xp5_ASAP7_75t_L g1602 ( 
.A1(n_1561),
.A2(n_1509),
.B1(n_1516),
.B2(n_1485),
.Y(n_1602)
);

OAI22xp5_ASAP7_75t_L g1603 ( 
.A1(n_1561),
.A2(n_1509),
.B1(n_1516),
.B2(n_1485),
.Y(n_1603)
);

INVxp67_ASAP7_75t_L g1604 ( 
.A(n_1580),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1590),
.Y(n_1605)
);

AO22x1_ASAP7_75t_L g1606 ( 
.A1(n_1576),
.A2(n_1530),
.B1(n_1555),
.B2(n_1496),
.Y(n_1606)
);

AOI21xp5_ASAP7_75t_L g1607 ( 
.A1(n_1575),
.A2(n_1504),
.B(n_1530),
.Y(n_1607)
);

OAI31xp33_ASAP7_75t_L g1608 ( 
.A1(n_1587),
.A2(n_1511),
.A3(n_1465),
.B(n_1447),
.Y(n_1608)
);

OAI322xp33_ASAP7_75t_SL g1609 ( 
.A1(n_1578),
.A2(n_1548),
.A3(n_1540),
.B1(n_1537),
.B2(n_1553),
.C1(n_1552),
.C2(n_1551),
.Y(n_1609)
);

OAI21xp33_ASAP7_75t_L g1610 ( 
.A1(n_1570),
.A2(n_1547),
.B(n_1539),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1582),
.B(n_1547),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1590),
.Y(n_1612)
);

NOR2xp33_ASAP7_75t_L g1613 ( 
.A(n_1587),
.B(n_1434),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1587),
.B(n_1492),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1559),
.Y(n_1615)
);

OAI221xp5_ASAP7_75t_L g1616 ( 
.A1(n_1578),
.A2(n_1465),
.B1(n_1458),
.B2(n_1509),
.C(n_1516),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1561),
.B(n_1492),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1559),
.Y(n_1618)
);

OR2x2_ASAP7_75t_L g1619 ( 
.A(n_1614),
.B(n_1573),
.Y(n_1619)
);

NOR2xp33_ASAP7_75t_L g1620 ( 
.A(n_1613),
.B(n_1574),
.Y(n_1620)
);

OAI21xp5_ASAP7_75t_SL g1621 ( 
.A1(n_1596),
.A2(n_1592),
.B(n_1566),
.Y(n_1621)
);

AOI22xp5_ASAP7_75t_L g1622 ( 
.A1(n_1598),
.A2(n_1486),
.B1(n_1465),
.B2(n_1574),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1613),
.B(n_1592),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1615),
.Y(n_1624)
);

AOI22xp33_ASAP7_75t_L g1625 ( 
.A1(n_1608),
.A2(n_1597),
.B1(n_1610),
.B2(n_1603),
.Y(n_1625)
);

OAI22xp5_ASAP7_75t_L g1626 ( 
.A1(n_1594),
.A2(n_1573),
.B1(n_1454),
.B2(n_1580),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1618),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1604),
.B(n_1574),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1601),
.B(n_1592),
.Y(n_1629)
);

INVx1_ASAP7_75t_SL g1630 ( 
.A(n_1595),
.Y(n_1630)
);

OAI32xp33_ASAP7_75t_L g1631 ( 
.A1(n_1602),
.A2(n_1576),
.A3(n_1581),
.B1(n_1554),
.B2(n_1549),
.Y(n_1631)
);

OAI32xp33_ASAP7_75t_L g1632 ( 
.A1(n_1594),
.A2(n_1576),
.A3(n_1581),
.B1(n_1549),
.B2(n_1566),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1604),
.B(n_1570),
.Y(n_1633)
);

OR2x2_ASAP7_75t_L g1634 ( 
.A(n_1600),
.B(n_1562),
.Y(n_1634)
);

OAI22xp5_ASAP7_75t_L g1635 ( 
.A1(n_1599),
.A2(n_1454),
.B1(n_1576),
.B2(n_1581),
.Y(n_1635)
);

A2O1A1Ixp33_ASAP7_75t_L g1636 ( 
.A1(n_1616),
.A2(n_1570),
.B(n_1496),
.C(n_1458),
.Y(n_1636)
);

OAI221xp5_ASAP7_75t_L g1637 ( 
.A1(n_1607),
.A2(n_1576),
.B1(n_1581),
.B2(n_1562),
.C(n_1565),
.Y(n_1637)
);

CKINVDCx14_ASAP7_75t_R g1638 ( 
.A(n_1620),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1626),
.B(n_1605),
.Y(n_1639)
);

OAI21xp5_ASAP7_75t_SL g1640 ( 
.A1(n_1626),
.A2(n_1611),
.B(n_1589),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1629),
.B(n_1612),
.Y(n_1641)
);

A2O1A1Ixp33_ASAP7_75t_L g1642 ( 
.A1(n_1632),
.A2(n_1609),
.B(n_1496),
.C(n_1617),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1623),
.B(n_1588),
.Y(n_1643)
);

AOI221xp5_ASAP7_75t_L g1644 ( 
.A1(n_1635),
.A2(n_1586),
.B1(n_1572),
.B2(n_1591),
.C(n_1584),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1634),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1628),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1624),
.Y(n_1647)
);

NAND3xp33_ASAP7_75t_L g1648 ( 
.A(n_1635),
.B(n_1606),
.C(n_1572),
.Y(n_1648)
);

NOR2xp33_ASAP7_75t_L g1649 ( 
.A(n_1638),
.B(n_1630),
.Y(n_1649)
);

INVx1_ASAP7_75t_SL g1650 ( 
.A(n_1643),
.Y(n_1650)
);

OAI22xp5_ASAP7_75t_L g1651 ( 
.A1(n_1640),
.A2(n_1625),
.B1(n_1621),
.B2(n_1622),
.Y(n_1651)
);

NAND4xp25_ASAP7_75t_L g1652 ( 
.A(n_1644),
.B(n_1633),
.C(n_1631),
.D(n_1637),
.Y(n_1652)
);

NOR2xp33_ASAP7_75t_L g1653 ( 
.A(n_1645),
.B(n_1619),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1641),
.Y(n_1654)
);

NOR2xp33_ASAP7_75t_L g1655 ( 
.A(n_1646),
.B(n_1581),
.Y(n_1655)
);

AOI21xp5_ASAP7_75t_L g1656 ( 
.A1(n_1639),
.A2(n_1636),
.B(n_1627),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1647),
.Y(n_1657)
);

INVx1_ASAP7_75t_SL g1658 ( 
.A(n_1639),
.Y(n_1658)
);

AOI22xp5_ASAP7_75t_L g1659 ( 
.A1(n_1658),
.A2(n_1648),
.B1(n_1642),
.B2(n_1565),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1650),
.B(n_1564),
.Y(n_1660)
);

NAND2xp33_ASAP7_75t_L g1661 ( 
.A(n_1654),
.B(n_1403),
.Y(n_1661)
);

A2O1A1Ixp33_ASAP7_75t_L g1662 ( 
.A1(n_1656),
.A2(n_1577),
.B(n_1591),
.C(n_1584),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1649),
.B(n_1564),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1663),
.Y(n_1664)
);

AOI22xp5_ASAP7_75t_L g1665 ( 
.A1(n_1661),
.A2(n_1651),
.B1(n_1653),
.B2(n_1652),
.Y(n_1665)
);

OAI22xp5_ASAP7_75t_L g1666 ( 
.A1(n_1659),
.A2(n_1655),
.B1(n_1657),
.B2(n_1577),
.Y(n_1666)
);

OAI211xp5_ASAP7_75t_SL g1667 ( 
.A1(n_1662),
.A2(n_1593),
.B(n_1560),
.C(n_1568),
.Y(n_1667)
);

OAI221xp5_ASAP7_75t_L g1668 ( 
.A1(n_1660),
.A2(n_1586),
.B1(n_1568),
.B2(n_1593),
.C(n_1560),
.Y(n_1668)
);

OAI22xp33_ASAP7_75t_L g1669 ( 
.A1(n_1659),
.A2(n_1568),
.B1(n_1560),
.B2(n_1593),
.Y(n_1669)
);

NAND4xp75_ASAP7_75t_L g1670 ( 
.A(n_1665),
.B(n_1664),
.C(n_1669),
.D(n_1666),
.Y(n_1670)
);

INVxp67_ASAP7_75t_L g1671 ( 
.A(n_1668),
.Y(n_1671)
);

HB1xp67_ASAP7_75t_L g1672 ( 
.A(n_1667),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1664),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1664),
.Y(n_1674)
);

NOR3xp33_ASAP7_75t_L g1675 ( 
.A(n_1670),
.B(n_1385),
.C(n_1403),
.Y(n_1675)
);

OAI322xp33_ASAP7_75t_L g1676 ( 
.A1(n_1671),
.A2(n_1551),
.A3(n_1537),
.B1(n_1540),
.B2(n_1550),
.C1(n_1535),
.C2(n_1552),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1673),
.B(n_1588),
.Y(n_1677)
);

OA22x2_ASAP7_75t_L g1678 ( 
.A1(n_1677),
.A2(n_1674),
.B1(n_1672),
.B2(n_1670),
.Y(n_1678)
);

AND4x2_ASAP7_75t_L g1679 ( 
.A(n_1678),
.B(n_1676),
.C(n_1675),
.D(n_1400),
.Y(n_1679)
);

XNOR2xp5_ASAP7_75t_L g1680 ( 
.A(n_1679),
.B(n_1408),
.Y(n_1680)
);

XNOR2xp5_ASAP7_75t_L g1681 ( 
.A(n_1679),
.B(n_1566),
.Y(n_1681)
);

OAI321xp33_ASAP7_75t_L g1682 ( 
.A1(n_1681),
.A2(n_1589),
.A3(n_1588),
.B1(n_1579),
.B2(n_1569),
.C(n_1550),
.Y(n_1682)
);

AOI22x1_ASAP7_75t_L g1683 ( 
.A1(n_1680),
.A2(n_1589),
.B1(n_1579),
.B2(n_1569),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1682),
.Y(n_1684)
);

AOI21xp5_ASAP7_75t_L g1685 ( 
.A1(n_1683),
.A2(n_1579),
.B(n_1569),
.Y(n_1685)
);

OAI21x1_ASAP7_75t_L g1686 ( 
.A1(n_1685),
.A2(n_1558),
.B(n_1557),
.Y(n_1686)
);

NOR2xp33_ASAP7_75t_L g1687 ( 
.A(n_1686),
.B(n_1684),
.Y(n_1687)
);

OAI31xp33_ASAP7_75t_L g1688 ( 
.A1(n_1687),
.A2(n_1553),
.A3(n_1523),
.B(n_1522),
.Y(n_1688)
);

OAI221xp5_ASAP7_75t_R g1689 ( 
.A1(n_1688),
.A2(n_1506),
.B1(n_1557),
.B2(n_1558),
.C(n_1501),
.Y(n_1689)
);

AOI211xp5_ASAP7_75t_L g1690 ( 
.A1(n_1689),
.A2(n_1407),
.B(n_1542),
.C(n_1541),
.Y(n_1690)
);


endmodule