module fake_jpeg_26493_n_325 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_325);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_325;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx5p33_ASAP7_75t_R g22 ( 
.A(n_16),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_8),
.B(n_7),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_3),
.B(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx4f_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx2_ASAP7_75t_SL g52 ( 
.A(n_35),
.Y(n_52)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_27),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_37),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_27),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_22),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_20),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_44),
.Y(n_51)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_22),
.B(n_9),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_31),
.C(n_34),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_45),
.B(n_32),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_40),
.A2(n_31),
.B1(n_20),
.B2(n_34),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_48),
.A2(n_67),
.B1(n_40),
.B2(n_17),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_19),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_49),
.B(n_35),
.Y(n_78)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_53),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_39),
.Y(n_53)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_59),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_40),
.A2(n_34),
.B1(n_33),
.B2(n_17),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_60),
.A2(n_33),
.B1(n_21),
.B2(n_18),
.Y(n_85)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_37),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_64),
.Y(n_76)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_40),
.A2(n_33),
.B1(n_17),
.B2(n_18),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_55),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_71),
.B(n_75),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_72),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_73),
.B(n_78),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_55),
.Y(n_75)
);

AO22x1_ASAP7_75t_SL g77 ( 
.A1(n_52),
.A2(n_35),
.B1(n_39),
.B2(n_36),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_77),
.A2(n_52),
.B1(n_61),
.B2(n_46),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g79 ( 
.A(n_67),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_79),
.B(n_80),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_50),
.B(n_42),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_51),
.B(n_38),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_83),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_51),
.B(n_38),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_51),
.B(n_35),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_84),
.B(n_87),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_85),
.A2(n_21),
.B1(n_22),
.B2(n_29),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_58),
.A2(n_39),
.B(n_25),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_86),
.A2(n_53),
.B(n_23),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_64),
.B(n_35),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_45),
.A2(n_36),
.B1(n_35),
.B2(n_32),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_89),
.A2(n_94),
.B1(n_52),
.B2(n_46),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_47),
.B(n_26),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_90),
.B(n_91),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_47),
.B(n_26),
.Y(n_91)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_92),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_48),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_93),
.B(n_57),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_71),
.B(n_24),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_96),
.B(n_105),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_56),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_97),
.B(n_104),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_98),
.A2(n_112),
.B1(n_114),
.B2(n_115),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_100),
.B(n_107),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_103),
.B(n_110),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_76),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

INVx1_ASAP7_75t_SL g106 ( 
.A(n_84),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_106),
.B(n_111),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_75),
.B(n_56),
.Y(n_110)
);

INVxp33_ASAP7_75t_L g111 ( 
.A(n_68),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_79),
.A2(n_61),
.B1(n_65),
.B2(n_63),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_78),
.B(n_57),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_113),
.B(n_117),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_93),
.A2(n_66),
.B1(n_54),
.B2(n_28),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_94),
.A2(n_54),
.B1(n_28),
.B2(n_23),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_32),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_118),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_73),
.A2(n_32),
.B1(n_30),
.B2(n_29),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_119),
.B(n_77),
.Y(n_146)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_88),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_120),
.B(n_121),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_88),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_95),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_123),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_116),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_124),
.B(n_127),
.Y(n_168)
);

INVxp33_ASAP7_75t_L g127 ( 
.A(n_95),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_110),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_129),
.B(n_130),
.Y(n_158)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_113),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_112),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_131),
.B(n_138),
.Y(n_173)
);

NAND2x1_ASAP7_75t_SL g135 ( 
.A(n_98),
.B(n_77),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_135),
.A2(n_68),
.B(n_86),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_121),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_137),
.Y(n_159)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_100),
.Y(n_138)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_116),
.Y(n_140)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_140),
.Y(n_169)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_100),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_141),
.B(n_142),
.Y(n_174)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_114),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_108),
.B(n_76),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_143),
.B(n_145),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_120),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_144),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_99),
.B(n_83),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_146),
.A2(n_131),
.B1(n_150),
.B2(n_128),
.Y(n_175)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_122),
.Y(n_147)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_147),
.Y(n_179)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_122),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_148),
.A2(n_69),
.B1(n_92),
.B2(n_81),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_101),
.B(n_74),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_149),
.B(n_151),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_99),
.B(n_74),
.Y(n_151)
);

BUFx5_ASAP7_75t_L g152 ( 
.A(n_124),
.Y(n_152)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_152),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_139),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_153),
.B(n_165),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_125),
.A2(n_122),
.B1(n_105),
.B2(n_119),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_154),
.A2(n_156),
.B1(n_170),
.B2(n_175),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_134),
.B(n_97),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_155),
.B(n_178),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_128),
.A2(n_108),
.B1(n_106),
.B2(n_118),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_142),
.A2(n_101),
.B1(n_103),
.B2(n_107),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_160),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_140),
.Y(n_162)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_162),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_147),
.B(n_109),
.C(n_117),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_163),
.B(n_133),
.C(n_136),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_138),
.A2(n_109),
.B(n_115),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_164),
.A2(n_172),
.B(n_143),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_139),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_137),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_166),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_144),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_167),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_135),
.A2(n_102),
.B1(n_89),
.B2(n_69),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_176),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_148),
.B(n_102),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_177),
.B(n_183),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_126),
.B(n_80),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_123),
.A2(n_92),
.B1(n_69),
.B2(n_81),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_180),
.A2(n_70),
.B1(n_77),
.B2(n_30),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_144),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_182),
.B(n_70),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_126),
.B(n_91),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_168),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_189),
.B(n_191),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_190),
.B(n_209),
.C(n_211),
.Y(n_219)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_173),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_192),
.B(n_178),
.Y(n_217)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_173),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_194),
.B(n_199),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_172),
.A2(n_141),
.B(n_136),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_195),
.A2(n_197),
.B(n_156),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_174),
.A2(n_129),
.B(n_133),
.Y(n_197)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_174),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_170),
.A2(n_130),
.B1(n_135),
.B2(n_146),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_200),
.A2(n_205),
.B1(n_206),
.B2(n_160),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_171),
.B(n_132),
.Y(n_201)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_201),
.Y(n_216)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_203),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_181),
.B(n_151),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_204),
.B(n_10),
.Y(n_235)
);

OAI22xp33_ASAP7_75t_L g205 ( 
.A1(n_171),
.A2(n_150),
.B1(n_81),
.B2(n_132),
.Y(n_205)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_158),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_208),
.B(n_210),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_155),
.B(n_145),
.C(n_90),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_180),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_163),
.B(n_30),
.C(n_29),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_187),
.B(n_177),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_212),
.B(n_217),
.Y(n_243)
);

O2A1O1Ixp33_ASAP7_75t_L g242 ( 
.A1(n_213),
.A2(n_236),
.B(n_222),
.C(n_216),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_214),
.A2(n_223),
.B1(n_229),
.B2(n_188),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_185),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_215),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_193),
.B(n_152),
.Y(n_218)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_218),
.Y(n_239)
);

MAJx2_ASAP7_75t_L g220 ( 
.A(n_190),
.B(n_183),
.C(n_157),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_220),
.B(n_232),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_187),
.B(n_164),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_221),
.B(n_230),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_196),
.A2(n_165),
.B1(n_179),
.B2(n_159),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_202),
.A2(n_179),
.B1(n_154),
.B2(n_161),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_224),
.B(n_225),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_202),
.A2(n_169),
.B1(n_30),
.B2(n_29),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_192),
.B(n_169),
.C(n_24),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_227),
.B(n_233),
.C(n_237),
.Y(n_238)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_201),
.Y(n_228)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_228),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_196),
.A2(n_24),
.B1(n_1),
.B2(n_0),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_207),
.B(n_9),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_200),
.B(n_9),
.Y(n_231)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_231),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_207),
.B(n_10),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_195),
.B(n_10),
.C(n_15),
.Y(n_233)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_235),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_198),
.B(n_8),
.Y(n_237)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_242),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_219),
.B(n_211),
.C(n_194),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_244),
.B(n_245),
.C(n_251),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_219),
.B(n_199),
.C(n_198),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g246 ( 
.A(n_234),
.Y(n_246)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_246),
.Y(n_265)
);

AO21x1_ASAP7_75t_L g250 ( 
.A1(n_223),
.A2(n_197),
.B(n_205),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_250),
.B(n_0),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_221),
.B(n_212),
.C(n_220),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_227),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_252),
.B(n_254),
.Y(n_273)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_229),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_256),
.A2(n_11),
.B1(n_15),
.B2(n_3),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_233),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_257),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_217),
.B(n_209),
.C(n_184),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_258),
.B(n_237),
.Y(n_260)
);

OA21x2_ASAP7_75t_SL g259 ( 
.A1(n_240),
.A2(n_230),
.B(n_232),
.Y(n_259)
);

NOR2xp67_ASAP7_75t_L g285 ( 
.A(n_259),
.B(n_253),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_260),
.A2(n_238),
.B(n_244),
.Y(n_283)
);

NAND4xp25_ASAP7_75t_SL g261 ( 
.A(n_255),
.B(n_186),
.C(n_226),
.D(n_184),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_261),
.B(n_275),
.Y(n_282)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_242),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_262),
.B(n_263),
.Y(n_287)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_250),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_251),
.B(n_206),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_266),
.B(n_267),
.Y(n_276)
);

OAI21xp33_ASAP7_75t_L g267 ( 
.A1(n_241),
.A2(n_239),
.B(n_247),
.Y(n_267)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_268),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_253),
.B(n_12),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_270),
.B(n_271),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_258),
.B(n_12),
.Y(n_271)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_272),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_238),
.Y(n_275)
);

NAND3xp33_ASAP7_75t_L g278 ( 
.A(n_271),
.B(n_249),
.C(n_270),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_278),
.B(n_283),
.Y(n_291)
);

INVxp33_ASAP7_75t_L g281 ( 
.A(n_267),
.Y(n_281)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_281),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_266),
.B(n_243),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_284),
.B(n_6),
.Y(n_299)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_285),
.Y(n_294)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_273),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_286),
.B(n_269),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_274),
.B(n_245),
.C(n_243),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_288),
.B(n_289),
.C(n_264),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_274),
.B(n_248),
.C(n_12),
.Y(n_289)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_290),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_287),
.A2(n_263),
.B1(n_262),
.B2(n_272),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_292),
.A2(n_284),
.B1(n_288),
.B2(n_0),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_281),
.B(n_265),
.Y(n_293)
);

OR2x2_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_295),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_289),
.B(n_261),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_296),
.B(n_297),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_282),
.B(n_279),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_299),
.B(n_279),
.Y(n_305)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_276),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_300),
.B(n_301),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_277),
.B(n_13),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_291),
.A2(n_280),
.B(n_276),
.Y(n_302)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_302),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_305),
.B(n_309),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_307),
.B(n_310),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_298),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_294),
.A2(n_4),
.B(n_5),
.Y(n_310)
);

A2O1A1Ixp33_ASAP7_75t_L g312 ( 
.A1(n_303),
.A2(n_295),
.B(n_298),
.C(n_292),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_312),
.B(n_16),
.C(n_1),
.Y(n_320)
);

NOR3xp33_ASAP7_75t_SL g314 ( 
.A(n_308),
.B(n_299),
.C(n_4),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_314),
.B(n_315),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_304),
.B(n_13),
.Y(n_315)
);

NOR2x1_ASAP7_75t_L g316 ( 
.A(n_306),
.B(n_14),
.Y(n_316)
);

NOR4xp25_ASAP7_75t_L g318 ( 
.A(n_316),
.B(n_309),
.C(n_14),
.D(n_15),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_318),
.A2(n_320),
.B(n_311),
.Y(n_321)
);

AOI31xp33_ASAP7_75t_L g322 ( 
.A1(n_321),
.A2(n_317),
.A3(n_319),
.B(n_313),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_322),
.B(n_317),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_323),
.B(n_1),
.Y(n_324)
);

BUFx24_ASAP7_75t_SL g325 ( 
.A(n_324),
.Y(n_325)
);


endmodule