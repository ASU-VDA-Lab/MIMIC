module fake_jpeg_10749_n_476 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_476);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_476;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx6_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_6),
.B(n_0),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_4),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_5),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g113 ( 
.A(n_46),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_12),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_47),
.B(n_73),
.Y(n_102)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

CKINVDCx6p67_ASAP7_75t_R g135 ( 
.A(n_48),
.Y(n_135)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_49),
.Y(n_105)
);

INVx4_ASAP7_75t_SL g50 ( 
.A(n_38),
.Y(n_50)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_50),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_51),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_52),
.Y(n_134)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_53),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_12),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_54),
.B(n_92),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_55),
.Y(n_117)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g125 ( 
.A(n_56),
.Y(n_125)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_57),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_58),
.Y(n_136)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_59),
.Y(n_152)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_60),
.Y(n_119)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_61),
.Y(n_123)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_62),
.Y(n_104)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_63),
.Y(n_124)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_17),
.Y(n_64)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_64),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_29),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_65),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_66),
.Y(n_148)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_14),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g139 ( 
.A(n_67),
.Y(n_139)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_17),
.Y(n_68)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_68),
.Y(n_138)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_24),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g142 ( 
.A(n_69),
.Y(n_142)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_70),
.Y(n_144)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_71),
.Y(n_110)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_24),
.Y(n_72)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_72),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_16),
.B(n_12),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_74),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_37),
.B(n_11),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_75),
.B(n_89),
.Y(n_107)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_28),
.Y(n_76)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_76),
.Y(n_151)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_34),
.Y(n_77)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_77),
.Y(n_116)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_38),
.Y(n_78)
);

BUFx10_ASAP7_75t_L g103 ( 
.A(n_78),
.Y(n_103)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_24),
.Y(n_79)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_79),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_23),
.Y(n_80)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_80),
.Y(n_157)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_28),
.Y(n_81)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_81),
.Y(n_155)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_20),
.Y(n_82)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_82),
.Y(n_141)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_24),
.Y(n_83)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_83),
.Y(n_111)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_28),
.Y(n_84)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_84),
.Y(n_146)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_34),
.Y(n_85)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_85),
.Y(n_133)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_23),
.Y(n_86)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_86),
.Y(n_158)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_13),
.Y(n_87)
);

BUFx10_ASAP7_75t_L g122 ( 
.A(n_87),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_23),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_88),
.B(n_90),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_38),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_32),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_20),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_93),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_16),
.B(n_11),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_21),
.B(n_11),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_14),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_94),
.B(n_98),
.Y(n_114)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_14),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_95),
.B(n_96),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_32),
.Y(n_96)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_38),
.Y(n_97)
);

CKINVDCx14_ASAP7_75t_SL g112 ( 
.A(n_97),
.Y(n_112)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_13),
.Y(n_98)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_38),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_99),
.Y(n_140)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_13),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_100),
.B(n_101),
.Y(n_115)
);

INVx11_ASAP7_75t_L g101 ( 
.A(n_43),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_75),
.A2(n_15),
.B1(n_32),
.B2(n_36),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_120),
.A2(n_130),
.B1(n_137),
.B2(n_143),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_87),
.B(n_30),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_121),
.B(n_129),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_49),
.A2(n_15),
.B1(n_36),
.B2(n_32),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_126),
.A2(n_43),
.B1(n_86),
.B2(n_90),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_87),
.B(n_21),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_56),
.A2(n_27),
.B1(n_15),
.B2(n_43),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_57),
.B(n_25),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_131),
.B(n_106),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_77),
.A2(n_27),
.B1(n_43),
.B2(n_36),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_53),
.A2(n_36),
.B1(n_27),
.B2(n_45),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_50),
.B(n_33),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g190 ( 
.A(n_149),
.B(n_150),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_67),
.B(n_45),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_160),
.A2(n_174),
.B1(n_182),
.B2(n_157),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_161),
.B(n_165),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_110),
.A2(n_85),
.B1(n_46),
.B2(n_55),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_162),
.Y(n_223)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_106),
.Y(n_163)
);

BUFx2_ASAP7_75t_L g206 ( 
.A(n_163),
.Y(n_206)
);

OA22x2_ASAP7_75t_L g164 ( 
.A1(n_140),
.A2(n_137),
.B1(n_130),
.B2(n_104),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_164),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_102),
.B(n_35),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_109),
.B(n_35),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_166),
.B(n_172),
.Y(n_235)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_158),
.Y(n_167)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_167),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_107),
.B(n_114),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_168),
.B(n_142),
.C(n_135),
.Y(n_214)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_145),
.Y(n_169)
);

BUFx2_ASAP7_75t_L g233 ( 
.A(n_169),
.Y(n_233)
);

AO22x1_ASAP7_75t_SL g170 ( 
.A1(n_119),
.A2(n_101),
.B1(n_99),
.B2(n_97),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_170),
.B(n_194),
.Y(n_216)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_155),
.Y(n_171)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_171),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_128),
.B(n_31),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_122),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g210 ( 
.A(n_173),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_153),
.A2(n_96),
.B1(n_51),
.B2(n_88),
.Y(n_174)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_141),
.Y(n_176)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_176),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_113),
.Y(n_177)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_177),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_122),
.Y(n_178)
);

INVx13_ASAP7_75t_L g219 ( 
.A(n_178),
.Y(n_219)
);

INVx8_ASAP7_75t_L g179 ( 
.A(n_116),
.Y(n_179)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_179),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_154),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_180),
.Y(n_208)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_145),
.Y(n_181)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_181),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_123),
.A2(n_52),
.B1(n_80),
.B2(n_66),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_108),
.Y(n_183)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_183),
.Y(n_209)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_124),
.Y(n_184)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_184),
.Y(n_217)
);

INVxp67_ASAP7_75t_SL g185 ( 
.A(n_122),
.Y(n_185)
);

INVx11_ASAP7_75t_L g232 ( 
.A(n_185),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_127),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_186),
.A2(n_187),
.B1(n_200),
.B2(n_202),
.Y(n_218)
);

OA22x2_ASAP7_75t_L g187 ( 
.A1(n_110),
.A2(n_95),
.B1(n_144),
.B2(n_138),
.Y(n_187)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_156),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_189),
.B(n_191),
.Y(n_205)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_146),
.Y(n_191)
);

HAxp5_ASAP7_75t_SL g192 ( 
.A(n_135),
.B(n_43),
.CON(n_192),
.SN(n_192)
);

OR2x4_ASAP7_75t_L g227 ( 
.A(n_192),
.B(n_201),
.Y(n_227)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_142),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_193),
.B(n_196),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_118),
.B(n_31),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_115),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_195),
.Y(n_231)
);

BUFx2_ASAP7_75t_L g196 ( 
.A(n_133),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_139),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_197),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_132),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_198),
.B(n_199),
.Y(n_234)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_156),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_127),
.Y(n_200)
);

AO22x1_ASAP7_75t_L g201 ( 
.A1(n_135),
.A2(n_78),
.B1(n_48),
.B2(n_43),
.Y(n_201)
);

INVx2_ASAP7_75t_SL g202 ( 
.A(n_151),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_139),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_203),
.A2(n_159),
.B1(n_117),
.B2(n_136),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_111),
.B(n_30),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_204),
.B(n_33),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_214),
.B(n_225),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_168),
.B(n_152),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_220),
.B(n_229),
.C(n_187),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_224),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_228),
.A2(n_157),
.B1(n_202),
.B2(n_134),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_168),
.B(n_151),
.Y(n_229)
);

OAI21xp33_ASAP7_75t_SL g230 ( 
.A1(n_195),
.A2(n_125),
.B(n_103),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_230),
.A2(n_201),
.B(n_192),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_175),
.B(n_26),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_238),
.B(n_26),
.Y(n_259)
);

A2O1A1Ixp33_ASAP7_75t_L g239 ( 
.A1(n_216),
.A2(n_190),
.B(n_164),
.C(n_188),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_239),
.B(n_266),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_220),
.B(n_190),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_240),
.B(n_252),
.C(n_258),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_234),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_241),
.B(n_245),
.Y(n_288)
);

XOR2x2_ASAP7_75t_L g242 ( 
.A(n_229),
.B(n_174),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_242),
.B(n_211),
.Y(n_272)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_207),
.Y(n_243)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_243),
.Y(n_277)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_207),
.Y(n_244)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_244),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_234),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_208),
.B(n_193),
.Y(n_247)
);

CKINVDCx14_ASAP7_75t_R g276 ( 
.A(n_247),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_248),
.A2(n_232),
.B1(n_221),
.B2(n_159),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_208),
.B(n_163),
.Y(n_249)
);

CKINVDCx14_ASAP7_75t_R g278 ( 
.A(n_249),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_SL g269 ( 
.A(n_250),
.B(n_225),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_231),
.B(n_167),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_251),
.B(n_257),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_214),
.B(n_164),
.C(n_187),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_222),
.Y(n_253)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_253),
.Y(n_285)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_209),
.Y(n_255)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_255),
.Y(n_289)
);

AOI32xp33_ASAP7_75t_L g256 ( 
.A1(n_226),
.A2(n_164),
.A3(n_187),
.B1(n_202),
.B2(n_103),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_256),
.A2(n_264),
.B(n_254),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_231),
.B(n_169),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_226),
.B(n_170),
.C(n_196),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_259),
.B(n_235),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_216),
.A2(n_228),
.B1(n_227),
.B2(n_223),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_260),
.A2(n_263),
.B1(n_236),
.B2(n_116),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_218),
.A2(n_160),
.B1(n_182),
.B2(n_170),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_261),
.A2(n_262),
.B1(n_210),
.B2(n_179),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_227),
.A2(n_105),
.B1(n_147),
.B2(n_134),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_223),
.A2(n_178),
.B(n_173),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_209),
.Y(n_265)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_265),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_212),
.B(n_189),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_268),
.A2(n_256),
.B1(n_263),
.B2(n_258),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_SL g311 ( 
.A(n_269),
.B(n_272),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_266),
.B(n_238),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_270),
.B(n_275),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_271),
.A2(n_280),
.B(n_272),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_240),
.B(n_234),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_273),
.B(n_287),
.C(n_293),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_249),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_250),
.A2(n_211),
.B(n_212),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_281),
.A2(n_286),
.B1(n_205),
.B2(n_233),
.Y(n_313)
);

NAND3xp33_ASAP7_75t_L g306 ( 
.A(n_283),
.B(n_259),
.C(n_247),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_284),
.A2(n_264),
.B(n_232),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_260),
.A2(n_235),
.B1(n_221),
.B2(n_148),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_240),
.B(n_211),
.Y(n_287)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_243),
.Y(n_291)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_291),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_252),
.A2(n_205),
.B1(n_222),
.B2(n_236),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_292),
.A2(n_260),
.B1(n_263),
.B2(n_258),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_246),
.B(n_205),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_281),
.A2(n_286),
.B1(n_261),
.B2(n_252),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_295),
.A2(n_309),
.B1(n_313),
.B2(n_320),
.Y(n_333)
);

CKINVDCx16_ASAP7_75t_R g296 ( 
.A(n_267),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_296),
.B(n_285),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_297),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_298),
.A2(n_299),
.B1(n_304),
.B2(n_305),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_267),
.A2(n_239),
.B1(n_250),
.B2(n_241),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_300),
.A2(n_310),
.B(n_314),
.Y(n_347)
);

INVxp33_ASAP7_75t_L g302 ( 
.A(n_274),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_302),
.B(n_316),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_275),
.B(n_242),
.Y(n_303)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_303),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_268),
.A2(n_239),
.B1(n_245),
.B2(n_242),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_292),
.A2(n_246),
.B1(n_257),
.B2(n_251),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_306),
.B(n_206),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_282),
.A2(n_262),
.B1(n_265),
.B2(n_255),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_307),
.A2(n_312),
.B1(n_317),
.B2(n_213),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_278),
.A2(n_282),
.B1(n_276),
.B2(n_280),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_271),
.A2(n_288),
.B(n_274),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_288),
.A2(n_244),
.B1(n_248),
.B2(n_253),
.Y(n_312)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_277),
.Y(n_315)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_315),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_270),
.B(n_217),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_269),
.A2(n_293),
.B1(n_291),
.B2(n_290),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_287),
.B(n_217),
.C(n_213),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_318),
.B(n_181),
.C(n_147),
.Y(n_342)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_277),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_319),
.B(n_289),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_279),
.A2(n_233),
.B1(n_186),
.B2(n_200),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_308),
.B(n_273),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_322),
.B(n_331),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_310),
.A2(n_290),
.B(n_289),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_324),
.Y(n_364)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_326),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_316),
.B(n_279),
.Y(n_327)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_327),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_294),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_329),
.B(n_346),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_330),
.A2(n_337),
.B1(n_313),
.B2(n_315),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_308),
.B(n_197),
.Y(n_331)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_332),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_308),
.B(n_237),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_334),
.B(n_336),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_295),
.A2(n_285),
.B1(n_215),
.B2(n_206),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_335),
.A2(n_299),
.B1(n_307),
.B2(n_298),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_311),
.B(n_103),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_314),
.A2(n_125),
.B(n_177),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_338),
.B(n_345),
.Y(n_348)
);

AO21x1_ASAP7_75t_L g339 ( 
.A1(n_304),
.A2(n_237),
.B(n_203),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_339),
.A2(n_133),
.B1(n_117),
.B2(n_58),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_SL g340 ( 
.A(n_311),
.B(n_219),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_SL g370 ( 
.A(n_340),
.B(n_136),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_342),
.B(n_343),
.C(n_344),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_311),
.B(n_219),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_309),
.B(n_317),
.C(n_318),
.Y(n_344)
);

AND2x2_ASAP7_75t_L g345 ( 
.A(n_312),
.B(n_215),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_305),
.B(n_111),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_349),
.A2(n_339),
.B1(n_323),
.B2(n_325),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_322),
.B(n_318),
.C(n_300),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_353),
.B(n_358),
.C(n_363),
.Y(n_376)
);

FAx1_ASAP7_75t_SL g354 ( 
.A(n_347),
.B(n_303),
.CI(n_296),
.CON(n_354),
.SN(n_354)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_354),
.B(n_369),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_SL g355 ( 
.A1(n_341),
.A2(n_300),
.B(n_306),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_355),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_334),
.B(n_331),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_356),
.B(n_368),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_344),
.B(n_294),
.C(n_319),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_360),
.A2(n_361),
.B1(n_367),
.B2(n_372),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_321),
.A2(n_313),
.B1(n_301),
.B2(n_297),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_336),
.B(n_347),
.C(n_342),
.Y(n_363)
);

INVx2_ASAP7_75t_SL g365 ( 
.A(n_328),
.Y(n_365)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_365),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_321),
.A2(n_301),
.B1(n_320),
.B2(n_148),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_324),
.B(n_337),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_343),
.B(n_105),
.C(n_112),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_370),
.B(n_368),
.Y(n_389)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_326),
.Y(n_371)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_371),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_356),
.B(n_333),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_377),
.B(n_379),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_351),
.B(n_333),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_SL g380 ( 
.A1(n_364),
.A2(n_341),
.B(n_358),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_380),
.B(n_385),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_382),
.A2(n_370),
.B1(n_357),
.B2(n_113),
.Y(n_400)
);

A2O1A1Ixp33_ASAP7_75t_SL g383 ( 
.A1(n_354),
.A2(n_345),
.B(n_335),
.C(n_338),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_SL g408 ( 
.A1(n_383),
.A2(n_41),
.B(n_42),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_349),
.A2(n_325),
.B1(n_327),
.B2(n_345),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_365),
.Y(n_386)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_386),
.Y(n_398)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_350),
.Y(n_387)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_387),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_351),
.B(n_340),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_388),
.B(n_389),
.Y(n_412)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_352),
.Y(n_390)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_390),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_367),
.A2(n_364),
.B1(n_348),
.B2(n_362),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g395 ( 
.A1(n_391),
.A2(n_354),
.B1(n_363),
.B2(n_369),
.Y(n_395)
);

BUFx4f_ASAP7_75t_SL g392 ( 
.A(n_348),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_392),
.B(n_0),
.Y(n_407)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_366),
.Y(n_393)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_393),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_348),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_394),
.B(n_113),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_395),
.A2(n_413),
.B1(n_383),
.B2(n_375),
.Y(n_420)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_373),
.A2(n_353),
.B(n_359),
.Y(n_396)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_396),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_376),
.B(n_357),
.C(n_359),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_399),
.B(n_402),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_400),
.A2(n_378),
.B1(n_384),
.B2(n_391),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_381),
.B(n_11),
.Y(n_401)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_401),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_376),
.B(n_112),
.C(n_39),
.Y(n_402)
);

AOI21xp33_ASAP7_75t_L g405 ( 
.A1(n_373),
.A2(n_41),
.B(n_25),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_SL g430 ( 
.A1(n_405),
.A2(n_404),
.B(n_398),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_406),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_407),
.B(n_411),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_408),
.B(n_22),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_379),
.B(n_42),
.C(n_39),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_374),
.A2(n_22),
.B1(n_14),
.B2(n_3),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_SL g415 ( 
.A(n_412),
.B(n_389),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_415),
.B(n_416),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_397),
.A2(n_383),
.B1(n_392),
.B2(n_377),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_417),
.B(n_418),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_400),
.A2(n_383),
.B1(n_392),
.B2(n_375),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_420),
.B(n_428),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_423),
.B(n_425),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_411),
.B(n_388),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_410),
.B(n_1),
.C(n_2),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_426),
.B(n_427),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_410),
.B(n_412),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_408),
.A2(n_10),
.B1(n_2),
.B2(n_3),
.Y(n_428)
);

CKINVDCx16_ASAP7_75t_R g429 ( 
.A(n_401),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_429),
.B(n_430),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_427),
.B(n_399),
.C(n_396),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_432),
.B(n_433),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_419),
.B(n_404),
.Y(n_433)
);

AOI21xp5_ASAP7_75t_L g434 ( 
.A1(n_422),
.A2(n_402),
.B(n_403),
.Y(n_434)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_434),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_421),
.B(n_409),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_435),
.B(n_440),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_414),
.B(n_416),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_420),
.B(n_403),
.C(n_413),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_441),
.B(n_444),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_425),
.B(n_1),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_443),
.B(n_428),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_L g444 ( 
.A1(n_418),
.A2(n_3),
.B(n_4),
.Y(n_444)
);

NOR2x1_ASAP7_75t_L g445 ( 
.A(n_436),
.B(n_437),
.Y(n_445)
);

NOR3xp33_ASAP7_75t_L g462 ( 
.A(n_445),
.B(n_6),
.C(n_7),
.Y(n_462)
);

OAI21x1_ASAP7_75t_L g460 ( 
.A1(n_446),
.A2(n_6),
.B(n_7),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_432),
.B(n_415),
.C(n_426),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_449),
.B(n_450),
.Y(n_456)
);

INVx6_ASAP7_75t_L g450 ( 
.A(n_431),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_SL g451 ( 
.A(n_438),
.B(n_424),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_451),
.B(n_443),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_L g453 ( 
.A1(n_441),
.A2(n_423),
.B1(n_4),
.B2(n_5),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_453),
.B(n_455),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_439),
.B(n_3),
.Y(n_455)
);

AOI21xp5_ASAP7_75t_L g457 ( 
.A1(n_452),
.A2(n_442),
.B(n_437),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_SL g464 ( 
.A1(n_457),
.A2(n_459),
.B(n_447),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_458),
.B(n_461),
.Y(n_468)
);

AOI21x1_ASAP7_75t_SL g459 ( 
.A1(n_454),
.A2(n_5),
.B(n_6),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_460),
.B(n_462),
.Y(n_465)
);

NOR2x1_ASAP7_75t_L g461 ( 
.A(n_448),
.B(n_8),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_464),
.B(n_466),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_456),
.B(n_449),
.C(n_450),
.Y(n_466)
);

INVxp67_ASAP7_75t_L g467 ( 
.A(n_463),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_467),
.B(n_446),
.Y(n_471)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_468),
.A2(n_445),
.B(n_455),
.Y(n_470)
);

OAI21xp5_ASAP7_75t_SL g472 ( 
.A1(n_470),
.A2(n_465),
.B(n_8),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_471),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_L g474 ( 
.A1(n_472),
.A2(n_469),
.B(n_8),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_SL g475 ( 
.A(n_474),
.B(n_473),
.Y(n_475)
);

BUFx24_ASAP7_75t_SL g476 ( 
.A(n_475),
.Y(n_476)
);


endmodule