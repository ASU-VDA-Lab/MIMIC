module fake_jpeg_16301_n_213 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_213);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_213;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx6_ASAP7_75t_SL g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_0),
.B(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx6_ASAP7_75t_SL g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_31),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_35),
.B(n_20),
.Y(n_57)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_26),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_32),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

CKINVDCx6p67_ASAP7_75t_R g47 ( 
.A(n_39),
.Y(n_47)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_26),
.B(n_27),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_30),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_27),
.B(n_2),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_42),
.B(n_32),
.Y(n_60)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_41),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_46),
.B(n_54),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_48),
.B(n_50),
.Y(n_80)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_37),
.Y(n_49)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_34),
.Y(n_54)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_57),
.B(n_59),
.Y(n_85)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_60),
.B(n_19),
.Y(n_73)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_36),
.B(n_20),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_62),
.B(n_39),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_45),
.A2(n_35),
.B1(n_30),
.B2(n_23),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_64),
.A2(n_69),
.B1(n_74),
.B2(n_51),
.Y(n_89)
);

O2A1O1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_45),
.A2(n_23),
.B(n_40),
.C(n_44),
.Y(n_65)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_65),
.Y(n_92)
);

OR2x2_ASAP7_75t_SL g66 ( 
.A(n_48),
.B(n_42),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_66),
.B(n_83),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_63),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_67),
.B(n_71),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_51),
.A2(n_44),
.B1(n_39),
.B2(n_34),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_48),
.A2(n_38),
.B(n_31),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_72),
.B(n_25),
.C(n_16),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_73),
.B(n_76),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_56),
.A2(n_33),
.B1(n_21),
.B2(n_36),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_50),
.B(n_17),
.Y(n_76)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_79),
.Y(n_104)
);

O2A1O1Ixp33_ASAP7_75t_SL g81 ( 
.A1(n_47),
.A2(n_44),
.B(n_39),
.C(n_34),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_81),
.A2(n_52),
.B1(n_58),
.B2(n_47),
.Y(n_91)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_49),
.B(n_17),
.Y(n_86)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_83),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_93),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_89),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_90),
.B(n_106),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_91),
.A2(n_96),
.B1(n_99),
.B2(n_84),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_63),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_80),
.B(n_19),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_95),
.B(n_97),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_77),
.A2(n_52),
.B1(n_59),
.B2(n_47),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_85),
.B(n_82),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_72),
.A2(n_25),
.B1(n_33),
.B2(n_21),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_100),
.A2(n_65),
.B(n_81),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_79),
.B(n_53),
.Y(n_101)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_101),
.Y(n_119)
);

BUFx5_ASAP7_75t_L g106 ( 
.A(n_75),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_70),
.B(n_53),
.Y(n_107)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_107),
.Y(n_125)
);

INVx2_ASAP7_75t_SL g108 ( 
.A(n_81),
.Y(n_108)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_108),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_70),
.B(n_78),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_109),
.A2(n_68),
.B(n_47),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_110),
.B(n_116),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_104),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_111),
.B(n_114),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_113),
.A2(n_109),
.B(n_101),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_104),
.Y(n_114)
);

AND2x6_ASAP7_75t_L g116 ( 
.A(n_102),
.B(n_88),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_106),
.Y(n_117)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_117),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_105),
.B(n_84),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_118),
.B(n_120),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_98),
.Y(n_120)
);

INVx13_ASAP7_75t_L g121 ( 
.A(n_90),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_129),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_98),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_122),
.B(n_126),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_124),
.A2(n_111),
.B(n_114),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_94),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_108),
.A2(n_68),
.B1(n_66),
.B2(n_4),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_127),
.A2(n_102),
.B1(n_92),
.B2(n_130),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_87),
.B(n_24),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_133),
.B(n_110),
.Y(n_151)
);

AND2x2_ASAP7_75t_SL g135 ( 
.A(n_125),
.B(n_93),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_135),
.A2(n_145),
.B(n_147),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_128),
.A2(n_108),
.B1(n_92),
.B2(n_102),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_136),
.A2(n_143),
.B1(n_121),
.B2(n_3),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_137),
.B(n_148),
.Y(n_158)
);

NAND2x1p5_ASAP7_75t_L g140 ( 
.A(n_128),
.B(n_112),
.Y(n_140)
);

OR2x2_ASAP7_75t_L g165 ( 
.A(n_140),
.B(n_2),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_112),
.B(n_109),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_141),
.B(n_150),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_125),
.A2(n_91),
.B1(n_100),
.B2(n_107),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_117),
.B(n_96),
.Y(n_144)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_144),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_115),
.B(n_103),
.Y(n_146)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_146),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_113),
.A2(n_53),
.B(n_37),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_124),
.A2(n_37),
.B(n_29),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_116),
.B(n_119),
.C(n_127),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_149),
.B(n_119),
.C(n_122),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_123),
.B(n_28),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_SL g173 ( 
.A(n_151),
.B(n_152),
.C(n_156),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_149),
.B(n_120),
.C(n_67),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_154),
.B(n_155),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_137),
.B(n_135),
.C(n_132),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_135),
.B(n_16),
.C(n_24),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_157),
.B(n_164),
.Y(n_176)
);

NOR3xp33_ASAP7_75t_L g159 ( 
.A(n_138),
.B(n_9),
.C(n_15),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_159),
.B(n_165),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_142),
.B(n_2),
.Y(n_162)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_162),
.Y(n_174)
);

MAJx2_ASAP7_75t_L g164 ( 
.A(n_140),
.B(n_28),
.C(n_29),
.Y(n_164)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_131),
.Y(n_166)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_166),
.Y(n_178)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_163),
.Y(n_167)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_167),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_160),
.B(n_139),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_170),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_153),
.B(n_131),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_171),
.B(n_177),
.C(n_157),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_155),
.A2(n_140),
.B1(n_136),
.B2(n_133),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g183 ( 
.A(n_172),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_161),
.B(n_134),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_175),
.B(n_179),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_154),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_152),
.A2(n_143),
.B1(n_141),
.B2(n_147),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_181),
.B(n_182),
.C(n_186),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_168),
.B(n_158),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_168),
.B(n_158),
.C(n_145),
.Y(n_186)
);

MAJx2_ASAP7_75t_L g187 ( 
.A(n_179),
.B(n_164),
.C(n_148),
.Y(n_187)
);

NOR2xp67_ASAP7_75t_SL g189 ( 
.A(n_187),
.B(n_173),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_172),
.B(n_165),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_188),
.B(n_176),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_189),
.A2(n_196),
.B(n_176),
.Y(n_202)
);

A2O1A1Ixp33_ASAP7_75t_L g190 ( 
.A1(n_183),
.A2(n_167),
.B(n_169),
.C(n_173),
.Y(n_190)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_190),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_180),
.B(n_174),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_191),
.B(n_194),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_183),
.A2(n_185),
.B1(n_187),
.B2(n_188),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_193),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_184),
.B(n_178),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_195),
.B(n_192),
.Y(n_197)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_188),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_197),
.B(n_202),
.C(n_199),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_192),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_201),
.B(n_7),
.Y(n_204)
);

OR2x2_ASAP7_75t_L g203 ( 
.A(n_198),
.B(n_190),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_203),
.B(n_204),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_205),
.B(n_15),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_200),
.A2(n_7),
.B1(n_13),
.B2(n_10),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_206),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_208),
.B(n_209),
.C(n_203),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_210),
.B(n_211),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_208),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_212),
.B(n_207),
.Y(n_213)
);


endmodule