module fake_ariane_2843_n_4997 (n_295, n_356, n_556, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_516, n_332, n_294, n_197, n_463, n_176, n_34, n_404, n_172, n_347, n_423, n_183, n_469, n_479, n_373, n_299, n_541, n_499, n_12, n_564, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_421, n_96, n_549, n_522, n_319, n_49, n_20, n_416, n_283, n_50, n_187, n_525, n_367, n_345, n_374, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_443, n_57, n_424, n_528, n_387, n_406, n_117, n_139, n_524, n_85, n_130, n_349, n_391, n_466, n_346, n_214, n_348, n_552, n_2, n_462, n_32, n_410, n_379, n_445, n_515, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_441, n_568, n_385, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_23, n_399, n_554, n_520, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_473, n_186, n_202, n_145, n_193, n_500, n_59, n_336, n_315, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_339, n_487, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_446, n_553, n_143, n_566, n_152, n_405, n_557, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_559, n_401, n_485, n_267, n_495, n_504, n_483, n_335, n_435, n_350, n_291, n_344, n_381, n_426, n_433, n_481, n_398, n_62, n_210, n_200, n_529, n_502, n_166, n_253, n_561, n_218, n_79, n_3, n_271, n_465, n_486, n_507, n_247, n_569, n_567, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_547, n_420, n_562, n_518, n_439, n_222, n_478, n_510, n_256, n_326, n_227, n_48, n_188, n_323, n_550, n_330, n_400, n_11, n_129, n_126, n_282, n_328, n_368, n_277, n_248, n_301, n_467, n_432, n_545, n_536, n_293, n_228, n_325, n_276, n_93, n_427, n_108, n_497, n_303, n_442, n_168, n_81, n_1, n_206, n_352, n_538, n_511, n_238, n_365, n_429, n_455, n_136, n_334, n_192, n_488, n_300, n_533, n_505, n_14, n_163, n_88, n_141, n_390, n_498, n_104, n_501, n_438, n_314, n_16, n_440, n_273, n_305, n_539, n_312, n_233, n_56, n_60, n_388, n_333, n_449, n_413, n_392, n_376, n_512, n_459, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_237, n_175, n_453, n_74, n_491, n_19, n_40, n_181, n_570, n_53, n_260, n_362, n_543, n_310, n_236, n_565, n_281, n_24, n_7, n_461, n_209, n_262, n_490, n_17, n_225, n_235, n_464, n_575, n_546, n_297, n_503, n_290, n_527, n_46, n_84, n_371, n_199, n_107, n_217, n_452, n_178, n_42, n_551, n_308, n_417, n_201, n_70, n_572, n_343, n_10, n_414, n_571, n_287, n_302, n_380, n_6, n_94, n_284, n_4, n_448, n_249, n_534, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_278, n_255, n_560, n_450, n_257, n_148, n_451, n_475, n_135, n_409, n_171, n_519, n_384, n_468, n_61, n_526, n_102, n_182, n_482, n_316, n_196, n_125, n_43, n_407, n_13, n_27, n_254, n_476, n_460, n_219, n_55, n_535, n_231, n_366, n_555, n_234, n_492, n_574, n_280, n_215, n_252, n_161, n_454, n_298, n_532, n_68, n_415, n_78, n_63, n_99, n_540, n_216, n_544, n_5, n_514, n_418, n_537, n_223, n_403, n_25, n_83, n_389, n_513, n_288, n_179, n_395, n_195, n_213, n_110, n_304, n_67, n_509, n_306, n_313, n_92, n_430, n_493, n_203, n_378, n_436, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_337, n_437, n_111, n_21, n_274, n_472, n_296, n_265, n_208, n_456, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_521, n_51, n_496, n_76, n_342, n_26, n_246, n_517, n_530, n_0, n_428, n_159, n_358, n_105, n_30, n_494, n_131, n_263, n_434, n_360, n_563, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_542, n_548, n_523, n_268, n_266, n_470, n_457, n_164, n_157, n_184, n_177, n_477, n_364, n_258, n_425, n_431, n_508, n_118, n_121, n_411, n_484, n_353, n_22, n_241, n_29, n_357, n_412, n_447, n_191, n_382, n_489, n_80, n_480, n_211, n_97, n_408, n_322, n_251, n_506, n_558, n_116, n_397, n_471, n_351, n_39, n_393, n_474, n_359, n_155, n_573, n_127, n_531, n_4997);

input n_295;
input n_356;
input n_556;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_516;
input n_332;
input n_294;
input n_197;
input n_463;
input n_176;
input n_34;
input n_404;
input n_172;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_373;
input n_299;
input n_541;
input n_499;
input n_12;
input n_564;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_549;
input n_522;
input n_319;
input n_49;
input n_20;
input n_416;
input n_283;
input n_50;
input n_187;
input n_525;
input n_367;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_443;
input n_57;
input n_424;
input n_528;
input n_387;
input n_406;
input n_117;
input n_139;
input n_524;
input n_85;
input n_130;
input n_349;
input n_391;
input n_466;
input n_346;
input n_214;
input n_348;
input n_552;
input n_2;
input n_462;
input n_32;
input n_410;
input n_379;
input n_445;
input n_515;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_568;
input n_385;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_23;
input n_399;
input n_554;
input n_520;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_202;
input n_145;
input n_193;
input n_500;
input n_59;
input n_336;
input n_315;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_487;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_446;
input n_553;
input n_143;
input n_566;
input n_152;
input n_405;
input n_557;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_559;
input n_401;
input n_485;
input n_267;
input n_495;
input n_504;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_344;
input n_381;
input n_426;
input n_433;
input n_481;
input n_398;
input n_62;
input n_210;
input n_200;
input n_529;
input n_502;
input n_166;
input n_253;
input n_561;
input n_218;
input n_79;
input n_3;
input n_271;
input n_465;
input n_486;
input n_507;
input n_247;
input n_569;
input n_567;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_547;
input n_420;
input n_562;
input n_518;
input n_439;
input n_222;
input n_478;
input n_510;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_550;
input n_330;
input n_400;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_545;
input n_536;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_427;
input n_108;
input n_497;
input n_303;
input n_442;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_538;
input n_511;
input n_238;
input n_365;
input n_429;
input n_455;
input n_136;
input n_334;
input n_192;
input n_488;
input n_300;
input n_533;
input n_505;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_498;
input n_104;
input n_501;
input n_438;
input n_314;
input n_16;
input n_440;
input n_273;
input n_305;
input n_539;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_449;
input n_413;
input n_392;
input n_376;
input n_512;
input n_459;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_237;
input n_175;
input n_453;
input n_74;
input n_491;
input n_19;
input n_40;
input n_181;
input n_570;
input n_53;
input n_260;
input n_362;
input n_543;
input n_310;
input n_236;
input n_565;
input n_281;
input n_24;
input n_7;
input n_461;
input n_209;
input n_262;
input n_490;
input n_17;
input n_225;
input n_235;
input n_464;
input n_575;
input n_546;
input n_297;
input n_503;
input n_290;
input n_527;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_217;
input n_452;
input n_178;
input n_42;
input n_551;
input n_308;
input n_417;
input n_201;
input n_70;
input n_572;
input n_343;
input n_10;
input n_414;
input n_571;
input n_287;
input n_302;
input n_380;
input n_6;
input n_94;
input n_284;
input n_4;
input n_448;
input n_249;
input n_534;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_278;
input n_255;
input n_560;
input n_450;
input n_257;
input n_148;
input n_451;
input n_475;
input n_135;
input n_409;
input n_171;
input n_519;
input n_384;
input n_468;
input n_61;
input n_526;
input n_102;
input n_182;
input n_482;
input n_316;
input n_196;
input n_125;
input n_43;
input n_407;
input n_13;
input n_27;
input n_254;
input n_476;
input n_460;
input n_219;
input n_55;
input n_535;
input n_231;
input n_366;
input n_555;
input n_234;
input n_492;
input n_574;
input n_280;
input n_215;
input n_252;
input n_161;
input n_454;
input n_298;
input n_532;
input n_68;
input n_415;
input n_78;
input n_63;
input n_99;
input n_540;
input n_216;
input n_544;
input n_5;
input n_514;
input n_418;
input n_537;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_513;
input n_288;
input n_179;
input n_395;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_509;
input n_306;
input n_313;
input n_92;
input n_430;
input n_493;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_472;
input n_296;
input n_265;
input n_208;
input n_456;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_521;
input n_51;
input n_496;
input n_76;
input n_342;
input n_26;
input n_246;
input n_517;
input n_530;
input n_0;
input n_428;
input n_159;
input n_358;
input n_105;
input n_30;
input n_494;
input n_131;
input n_263;
input n_434;
input n_360;
input n_563;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_542;
input n_548;
input n_523;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_425;
input n_431;
input n_508;
input n_118;
input n_121;
input n_411;
input n_484;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_412;
input n_447;
input n_191;
input n_382;
input n_489;
input n_80;
input n_480;
input n_211;
input n_97;
input n_408;
input n_322;
input n_251;
input n_506;
input n_558;
input n_116;
input n_397;
input n_471;
input n_351;
input n_39;
input n_393;
input n_474;
input n_359;
input n_155;
input n_573;
input n_127;
input n_531;

output n_4997;

wire n_2752;
wire n_3527;
wire n_4474;
wire n_4030;
wire n_4770;
wire n_3152;
wire n_4586;
wire n_3056;
wire n_3500;
wire n_2679;
wire n_2182;
wire n_2680;
wire n_3264;
wire n_1250;
wire n_2993;
wire n_4283;
wire n_2879;
wire n_4403;
wire n_4962;
wire n_1430;
wire n_2002;
wire n_1238;
wire n_2729;
wire n_4302;
wire n_4547;
wire n_3765;
wire n_864;
wire n_1096;
wire n_1379;
wire n_2376;
wire n_2790;
wire n_2207;
wire n_3954;
wire n_4982;
wire n_2042;
wire n_1131;
wire n_2646;
wire n_737;
wire n_2653;
wire n_4610;
wire n_3115;
wire n_4028;
wire n_2482;
wire n_1682;
wire n_958;
wire n_2554;
wire n_4321;
wire n_1985;
wire n_2621;
wire n_4853;
wire n_1909;
wire n_4260;
wire n_903;
wire n_3348;
wire n_3261;
wire n_1761;
wire n_1690;
wire n_2807;
wire n_1018;
wire n_4512;
wire n_4132;
wire n_1364;
wire n_2390;
wire n_4500;
wire n_625;
wire n_2322;
wire n_1107;
wire n_2663;
wire n_4824;
wire n_3545;
wire n_1428;
wire n_1284;
wire n_4741;
wire n_1241;
wire n_4143;
wire n_4273;
wire n_901;
wire n_4136;
wire n_3144;
wire n_2359;
wire n_1519;
wire n_4567;
wire n_786;
wire n_3552;
wire n_2950;
wire n_3639;
wire n_3254;
wire n_2227;
wire n_2301;
wire n_3121;
wire n_2847;
wire n_3015;
wire n_3870;
wire n_3749;
wire n_1676;
wire n_1085;
wire n_3482;
wire n_823;
wire n_1900;
wire n_620;
wire n_4268;
wire n_587;
wire n_863;
wire n_3960;
wire n_2433;
wire n_899;
wire n_3975;
wire n_2004;
wire n_4018;
wire n_1495;
wire n_3325;
wire n_661;
wire n_4227;
wire n_1917;
wire n_2456;
wire n_1924;
wire n_1811;
wire n_3612;
wire n_4505;
wire n_1840;
wire n_4476;
wire n_579;
wire n_844;
wire n_1267;
wire n_2956;
wire n_1213;
wire n_2382;
wire n_780;
wire n_1918;
wire n_4119;
wire n_4443;
wire n_4000;
wire n_2686;
wire n_1949;
wire n_1140;
wire n_3458;
wire n_3511;
wire n_2077;
wire n_1121;
wire n_3012;
wire n_1947;
wire n_4529;
wire n_3850;
wire n_1216;
wire n_4908;
wire n_3754;
wire n_4432;
wire n_2263;
wire n_3518;
wire n_2800;
wire n_2116;
wire n_4530;
wire n_1432;
wire n_2245;
wire n_3359;
wire n_3841;
wire n_851;
wire n_3900;
wire n_3413;
wire n_3539;
wire n_2134;
wire n_3862;
wire n_930;
wire n_4912;
wire n_4226;
wire n_4311;
wire n_3284;
wire n_1386;
wire n_3506;
wire n_4827;
wire n_1842;
wire n_4993;
wire n_3678;
wire n_2791;
wire n_1661;
wire n_3212;
wire n_4871;
wire n_3529;
wire n_4405;
wire n_992;
wire n_966;
wire n_3549;
wire n_3914;
wire n_1692;
wire n_2611;
wire n_3029;
wire n_4745;
wire n_2398;
wire n_4233;
wire n_4791;
wire n_1178;
wire n_2015;
wire n_2877;
wire n_4951;
wire n_4959;
wire n_3000;
wire n_2930;
wire n_2745;
wire n_2087;
wire n_619;
wire n_2161;
wire n_746;
wire n_1357;
wire n_1787;
wire n_1389;
wire n_3172;
wire n_2659;
wire n_4033;
wire n_3747;
wire n_4905;
wire n_4508;
wire n_4045;
wire n_4894;
wire n_3651;
wire n_1812;
wire n_3614;
wire n_959;
wire n_2257;
wire n_1101;
wire n_1343;
wire n_3116;
wire n_4141;
wire n_3784;
wire n_3372;
wire n_3891;
wire n_4422;
wire n_1623;
wire n_3559;
wire n_2435;
wire n_1932;
wire n_1780;
wire n_2825;
wire n_1087;
wire n_632;
wire n_2388;
wire n_2273;
wire n_1911;
wire n_3496;
wire n_4364;
wire n_3493;
wire n_3700;
wire n_4307;
wire n_2795;
wire n_1841;
wire n_1680;
wire n_2954;
wire n_4438;
wire n_974;
wire n_3814;
wire n_4367;
wire n_2467;
wire n_4195;
wire n_4866;
wire n_1447;
wire n_1220;
wire n_2019;
wire n_698;
wire n_3010;
wire n_2160;
wire n_1992;
wire n_1209;
wire n_4254;
wire n_646;
wire n_3438;
wire n_2625;
wire n_1578;
wire n_3147;
wire n_3661;
wire n_3320;
wire n_4179;
wire n_2144;
wire n_1029;
wire n_2649;
wire n_1247;
wire n_1568;
wire n_2919;
wire n_3108;
wire n_2632;
wire n_4314;
wire n_2980;
wire n_1728;
wire n_4315;
wire n_3239;
wire n_2631;
wire n_3311;
wire n_3516;
wire n_4442;
wire n_4857;
wire n_1651;
wire n_3087;
wire n_4637;
wire n_2697;
wire n_1263;
wire n_1817;
wire n_3704;
wire n_670;
wire n_2677;
wire n_4296;
wire n_2483;
wire n_1032;
wire n_1592;
wire n_4714;
wire n_3074;
wire n_2655;
wire n_3589;
wire n_1743;
wire n_720;
wire n_1943;
wire n_4588;
wire n_1163;
wire n_3054;
wire n_4970;
wire n_4153;
wire n_1868;
wire n_3601;
wire n_2373;
wire n_3881;
wire n_2099;
wire n_3759;
wire n_3323;
wire n_4643;
wire n_2617;
wire n_808;
wire n_2476;
wire n_2814;
wire n_4133;
wire n_2636;
wire n_1439;
wire n_3466;
wire n_2074;
wire n_1665;
wire n_2122;
wire n_4543;
wire n_4337;
wire n_4788;
wire n_1414;
wire n_2067;
wire n_4555;
wire n_1901;
wire n_4486;
wire n_3465;
wire n_2117;
wire n_1053;
wire n_1906;
wire n_2194;
wire n_4780;
wire n_4640;
wire n_1828;
wire n_1304;
wire n_3335;
wire n_3007;
wire n_2267;
wire n_604;
wire n_1349;
wire n_1061;
wire n_2102;
wire n_4157;
wire n_3477;
wire n_3370;
wire n_874;
wire n_3949;
wire n_2286;
wire n_4247;
wire n_707;
wire n_3036;
wire n_2783;
wire n_4583;
wire n_1015;
wire n_1162;
wire n_4292;
wire n_2118;
wire n_688;
wire n_636;
wire n_1490;
wire n_3764;
wire n_1553;
wire n_4773;
wire n_1760;
wire n_1086;
wire n_3025;
wire n_3051;
wire n_986;
wire n_1104;
wire n_2802;
wire n_887;
wire n_2125;
wire n_1156;
wire n_4974;
wire n_2861;
wire n_4344;
wire n_3130;
wire n_1188;
wire n_1498;
wire n_4856;
wire n_2618;
wire n_4216;
wire n_957;
wire n_1242;
wire n_2707;
wire n_2849;
wire n_1489;
wire n_2756;
wire n_3781;
wire n_2217;
wire n_4864;
wire n_2226;
wire n_4313;
wire n_4460;
wire n_4670;
wire n_1119;
wire n_3713;
wire n_1863;
wire n_4798;
wire n_1500;
wire n_616;
wire n_4946;
wire n_4848;
wire n_4297;
wire n_4941;
wire n_4229;
wire n_3337;
wire n_1189;
wire n_3750;
wire n_3424;
wire n_3356;
wire n_1523;
wire n_2190;
wire n_3931;
wire n_2516;
wire n_4991;
wire n_3070;
wire n_1005;
wire n_3275;
wire n_3245;
wire n_2894;
wire n_2452;
wire n_4182;
wire n_2827;
wire n_3214;
wire n_3085;
wire n_3373;
wire n_4252;
wire n_3710;
wire n_1844;
wire n_1957;
wire n_1953;
wire n_1219;
wire n_710;
wire n_3944;
wire n_4729;
wire n_1793;
wire n_4446;
wire n_4662;
wire n_4800;
wire n_1373;
wire n_1540;
wire n_4440;
wire n_1797;
wire n_4425;
wire n_832;
wire n_744;
wire n_2821;
wire n_3696;
wire n_1331;
wire n_4781;
wire n_1529;
wire n_3531;
wire n_655;
wire n_4237;
wire n_4828;
wire n_3333;
wire n_4652;
wire n_4114;
wire n_1007;
wire n_1580;
wire n_3135;
wire n_4925;
wire n_2448;
wire n_2211;
wire n_951;
wire n_2424;
wire n_4697;
wire n_4765;
wire n_722;
wire n_3277;
wire n_4863;
wire n_1766;
wire n_1338;
wire n_2978;
wire n_4859;
wire n_4568;
wire n_3617;
wire n_704;
wire n_2958;
wire n_1044;
wire n_1714;
wire n_4429;
wire n_3340;
wire n_1243;
wire n_3486;
wire n_608;
wire n_2457;
wire n_2992;
wire n_3197;
wire n_3256;
wire n_1878;
wire n_3646;
wire n_2520;
wire n_811;
wire n_791;
wire n_3864;
wire n_4694;
wire n_1025;
wire n_4664;
wire n_3450;
wire n_687;
wire n_4633;
wire n_2026;
wire n_4050;
wire n_3173;
wire n_642;
wire n_1406;
wire n_4306;
wire n_2684;
wire n_2726;
wire n_4006;
wire n_3266;
wire n_3102;
wire n_1499;
wire n_4288;
wire n_3452;
wire n_4098;
wire n_2691;
wire n_4511;
wire n_3422;
wire n_4675;
wire n_695;
wire n_2991;
wire n_1596;
wire n_4289;
wire n_4972;
wire n_2723;
wire n_1476;
wire n_2016;
wire n_3925;
wire n_4689;
wire n_678;
wire n_651;
wire n_2850;
wire n_1874;
wire n_3780;
wire n_1657;
wire n_3753;
wire n_1488;
wire n_4846;
wire n_1330;
wire n_906;
wire n_2295;
wire n_4076;
wire n_3142;
wire n_3129;
wire n_3495;
wire n_3843;
wire n_4805;
wire n_2606;
wire n_2386;
wire n_4822;
wire n_1829;
wire n_4635;
wire n_1450;
wire n_3740;
wire n_2417;
wire n_1815;
wire n_1493;
wire n_2911;
wire n_3313;
wire n_2354;
wire n_4281;
wire n_3945;
wire n_3726;
wire n_4419;
wire n_1256;
wire n_3560;
wire n_3345;
wire n_3421;
wire n_1448;
wire n_1009;
wire n_3548;
wire n_4906;
wire n_4630;
wire n_4829;
wire n_2612;
wire n_3236;
wire n_1995;
wire n_1397;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_4966;
wire n_2250;
wire n_1117;
wire n_3321;
wire n_1303;
wire n_4188;
wire n_2001;
wire n_2506;
wire n_2413;
wire n_4825;
wire n_1593;
wire n_2610;
wire n_3715;
wire n_2626;
wire n_2892;
wire n_2605;
wire n_2804;
wire n_4882;
wire n_3206;
wire n_1035;
wire n_3475;
wire n_4878;
wire n_2070;
wire n_3842;
wire n_1367;
wire n_4202;
wire n_2044;
wire n_3886;
wire n_825;
wire n_732;
wire n_2619;
wire n_1192;
wire n_3098;
wire n_4503;
wire n_1291;
wire n_3987;
wire n_4249;
wire n_3160;
wire n_1160;
wire n_2968;
wire n_1882;
wire n_1976;
wire n_2711;
wire n_3223;
wire n_3386;
wire n_3921;
wire n_2177;
wire n_2766;
wire n_4196;
wire n_1197;
wire n_2613;
wire n_1517;
wire n_2647;
wire n_3920;
wire n_3444;
wire n_3851;
wire n_1671;
wire n_1048;
wire n_2343;
wire n_775;
wire n_667;
wire n_3380;
wire n_2826;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_2411;
wire n_4631;
wire n_1504;
wire n_2110;
wire n_3822;
wire n_889;
wire n_4355;
wire n_3818;
wire n_3587;
wire n_2608;
wire n_1948;
wire n_4155;
wire n_810;
wire n_4278;
wire n_4710;
wire n_1959;
wire n_3497;
wire n_4542;
wire n_3243;
wire n_4326;
wire n_2121;
wire n_3865;
wire n_4685;
wire n_3927;
wire n_2068;
wire n_3595;
wire n_1194;
wire n_4060;
wire n_1647;
wire n_1454;
wire n_2459;
wire n_941;
wire n_3396;
wire n_4093;
wire n_4123;
wire n_4294;
wire n_1521;
wire n_1940;
wire n_3683;
wire n_4452;
wire n_3887;
wire n_3195;
wire n_4722;
wire n_3048;
wire n_3339;
wire n_4164;
wire n_4126;
wire n_2963;
wire n_2561;
wire n_1056;
wire n_674;
wire n_3168;
wire n_4079;
wire n_1749;
wire n_1653;
wire n_4088;
wire n_2669;
wire n_3911;
wire n_3802;
wire n_4366;
wire n_1584;
wire n_848;
wire n_4922;
wire n_629;
wire n_4733;
wire n_1814;
wire n_2441;
wire n_4041;
wire n_2688;
wire n_4208;
wire n_4623;
wire n_4935;
wire n_4509;
wire n_2073;
wire n_4004;
wire n_750;
wire n_834;
wire n_3630;
wire n_1612;
wire n_800;
wire n_1910;
wire n_2189;
wire n_4194;
wire n_2672;
wire n_2018;
wire n_2602;
wire n_724;
wire n_2931;
wire n_3433;
wire n_3597;
wire n_1956;
wire n_1589;
wire n_4111;
wire n_3786;
wire n_875;
wire n_2828;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_4204;
wire n_3553;
wire n_3645;
wire n_793;
wire n_4996;
wire n_1485;
wire n_2883;
wire n_4411;
wire n_4317;
wire n_3550;
wire n_4785;
wire n_2870;
wire n_1494;
wire n_1893;
wire n_1805;
wire n_4068;
wire n_2270;
wire n_4163;
wire n_3294;
wire n_2443;
wire n_3610;
wire n_1554;
wire n_3279;
wire n_972;
wire n_4262;
wire n_2923;
wire n_2843;
wire n_3714;
wire n_4832;
wire n_3676;
wire n_2010;
wire n_1679;
wire n_3109;
wire n_1952;
wire n_2394;
wire n_3125;
wire n_2356;
wire n_4672;
wire n_2564;
wire n_3558;
wire n_3034;
wire n_3502;
wire n_783;
wire n_4053;
wire n_1127;
wire n_1008;
wire n_3963;
wire n_581;
wire n_3091;
wire n_1024;
wire n_4496;
wire n_2518;
wire n_936;
wire n_4596;
wire n_3105;
wire n_1525;
wire n_4628;
wire n_1775;
wire n_908;
wire n_1036;
wire n_4083;
wire n_1270;
wire n_1272;
wire n_2794;
wire n_2901;
wire n_3940;
wire n_3225;
wire n_3621;
wire n_3473;
wire n_3680;
wire n_3565;
wire n_2453;
wire n_3331;
wire n_1788;
wire n_2138;
wire n_3040;
wire n_4230;
wire n_3360;
wire n_1930;
wire n_1809;
wire n_3585;
wire n_1843;
wire n_2000;
wire n_4037;
wire n_3804;
wire n_4659;
wire n_3211;
wire n_917;
wire n_2096;
wire n_2440;
wire n_2556;
wire n_2215;
wire n_3847;
wire n_4073;
wire n_1261;
wire n_3633;
wire n_857;
wire n_1235;
wire n_2584;
wire n_4001;
wire n_1462;
wire n_1064;
wire n_633;
wire n_1446;
wire n_1701;
wire n_3111;
wire n_731;
wire n_1813;
wire n_2997;
wire n_1573;
wire n_3258;
wire n_758;
wire n_3691;
wire n_2252;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_784;
wire n_4339;
wire n_4690;
wire n_2987;
wire n_1473;
wire n_1076;
wire n_1348;
wire n_2651;
wire n_753;
wire n_2733;
wire n_2445;
wire n_2103;
wire n_4024;
wire n_4169;
wire n_3316;
wire n_4023;
wire n_4253;
wire n_2522;
wire n_3632;
wire n_1344;
wire n_4064;
wire n_3351;
wire n_1141;
wire n_3457;
wire n_2324;
wire n_840;
wire n_3454;
wire n_2139;
wire n_2521;
wire n_2740;
wire n_1991;
wire n_614;
wire n_4066;
wire n_4681;
wire n_3303;
wire n_4414;
wire n_2541;
wire n_3232;
wire n_1113;
wire n_3768;
wire n_4295;
wire n_1615;
wire n_4100;
wire n_1265;
wire n_2372;
wire n_2105;
wire n_3445;
wire n_1806;
wire n_4087;
wire n_1409;
wire n_1684;
wire n_1588;
wire n_1148;
wire n_1673;
wire n_4473;
wire n_4619;
wire n_2290;
wire n_4398;
wire n_2856;
wire n_3235;
wire n_3265;
wire n_3018;
wire n_1875;
wire n_2429;
wire n_4449;
wire n_3285;
wire n_4607;
wire n_1039;
wire n_1150;
wire n_4266;
wire n_1628;
wire n_2971;
wire n_4407;
wire n_4695;
wire n_1136;
wire n_1190;
wire n_3628;
wire n_4777;
wire n_3941;
wire n_1915;
wire n_658;
wire n_2846;
wire n_3371;
wire n_4918;
wire n_3872;
wire n_4415;
wire n_1964;
wire n_3659;
wire n_3928;
wire n_1777;
wire n_3366;
wire n_3441;
wire n_3020;
wire n_4146;
wire n_4947;
wire n_708;
wire n_2545;
wire n_2513;
wire n_4408;
wire n_2115;
wire n_2017;
wire n_1810;
wire n_1347;
wire n_4976;
wire n_860;
wire n_3555;
wire n_3534;
wire n_4548;
wire n_2670;
wire n_3556;
wire n_896;
wire n_4574;
wire n_2644;
wire n_4557;
wire n_3071;
wire n_1698;
wire n_1337;
wire n_774;
wire n_2148;
wire n_1168;
wire n_4663;
wire n_3296;
wire n_3762;
wire n_3794;
wire n_4624;
wire n_656;
wire n_4963;
wire n_4205;
wire n_3293;
wire n_4902;
wire n_1683;
wire n_4686;
wire n_2384;
wire n_1705;
wire n_768;
wire n_3707;
wire n_1091;
wire n_3895;
wire n_3149;
wire n_3934;
wire n_4338;
wire n_2058;
wire n_3231;
wire n_1846;
wire n_4161;
wire n_1581;
wire n_3058;
wire n_757;
wire n_2047;
wire n_946;
wire n_1655;
wire n_3398;
wire n_3709;
wire n_1146;
wire n_998;
wire n_3592;
wire n_2536;
wire n_1604;
wire n_3399;
wire n_4772;
wire n_1368;
wire n_963;
wire n_4120;
wire n_925;
wire n_2880;
wire n_1313;
wire n_3722;
wire n_1001;
wire n_4716;
wire n_4654;
wire n_1115;
wire n_1339;
wire n_1051;
wire n_3771;
wire n_719;
wire n_3158;
wire n_3221;
wire n_2316;
wire n_1010;
wire n_2830;
wire n_4622;
wire n_4757;
wire n_803;
wire n_1871;
wire n_4016;
wire n_3334;
wire n_2940;
wire n_3427;
wire n_3162;
wire n_4591;
wire n_3083;
wire n_4570;
wire n_2491;
wire n_1931;
wire n_2259;
wire n_849;
wire n_4655;
wire n_1820;
wire n_1233;
wire n_4493;
wire n_1808;
wire n_1635;
wire n_1704;
wire n_4896;
wire n_4851;
wire n_2479;
wire n_886;
wire n_1308;
wire n_1451;
wire n_1487;
wire n_675;
wire n_3432;
wire n_2163;
wire n_1938;
wire n_2484;
wire n_1469;
wire n_4901;
wire n_3480;
wire n_1355;
wire n_4213;
wire n_4127;
wire n_2500;
wire n_2334;
wire n_1169;
wire n_789;
wire n_3181;
wire n_1916;
wire n_610;
wire n_4602;
wire n_1713;
wire n_1436;
wire n_2818;
wire n_4900;
wire n_3578;
wire n_1109;
wire n_2537;
wire n_3745;
wire n_3487;
wire n_3668;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1566;
wire n_2837;
wire n_717;
wire n_952;
wire n_2446;
wire n_4116;
wire n_2671;
wire n_2702;
wire n_4363;
wire n_3561;
wire n_1839;
wire n_1138;
wire n_4103;
wire n_2529;
wire n_2374;
wire n_1225;
wire n_3154;
wire n_1366;
wire n_3938;
wire n_2278;
wire n_1424;
wire n_4736;
wire n_2976;
wire n_4842;
wire n_4416;
wire n_4439;
wire n_870;
wire n_4985;
wire n_3382;
wire n_3930;
wire n_3808;
wire n_2248;
wire n_813;
wire n_4660;
wire n_3081;
wire n_995;
wire n_2579;
wire n_1961;
wire n_1535;
wire n_2960;
wire n_3270;
wire n_871;
wire n_2844;
wire n_1979;
wire n_829;
wire n_4814;
wire n_2221;
wire n_1283;
wire n_2317;
wire n_2838;
wire n_1736;
wire n_2200;
wire n_2781;
wire n_2442;
wire n_3657;
wire n_2634;
wire n_2746;
wire n_645;
wire n_721;
wire n_1084;
wire n_1276;
wire n_2878;
wire n_3830;
wire n_3252;
wire n_1528;
wire n_3315;
wire n_3523;
wire n_3999;
wire n_3420;
wire n_3859;
wire n_868;
wire n_3474;
wire n_2458;
wire n_3150;
wire n_1542;
wire n_4831;
wire n_4782;
wire n_1539;
wire n_2859;
wire n_3412;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1636;
wire n_4597;
wire n_4546;
wire n_4031;
wire n_1254;
wire n_4147;
wire n_1703;
wire n_3073;
wire n_3571;
wire n_4576;
wire n_3297;
wire n_3003;
wire n_4340;
wire n_3136;
wire n_2867;
wire n_1560;
wire n_2899;
wire n_4284;
wire n_3274;
wire n_3877;
wire n_3817;
wire n_2722;
wire n_3728;
wire n_612;
wire n_4680;
wire n_1012;
wire n_2061;
wire n_2685;
wire n_2512;
wire n_1790;
wire n_2788;
wire n_1443;
wire n_2595;
wire n_1465;
wire n_3084;
wire n_705;
wire n_4593;
wire n_4562;
wire n_3860;
wire n_2909;
wire n_3554;
wire n_2717;
wire n_1391;
wire n_2981;
wire n_1006;
wire n_4995;
wire n_1159;
wire n_4498;
wire n_772;
wire n_1245;
wire n_2743;
wire n_1669;
wire n_2969;
wire n_3429;
wire n_1675;
wire n_2466;
wire n_676;
wire n_3758;
wire n_2568;
wire n_2271;
wire n_2326;
wire n_3485;
wire n_1594;
wire n_4109;
wire n_1935;
wire n_3777;
wire n_1872;
wire n_1585;
wire n_3767;
wire n_3692;
wire n_1351;
wire n_3234;
wire n_2216;
wire n_2426;
wire n_652;
wire n_4850;
wire n_1260;
wire n_3716;
wire n_2926;
wire n_4937;
wire n_798;
wire n_3391;
wire n_912;
wire n_4786;
wire n_4354;
wire n_4235;
wire n_3159;
wire n_2855;
wire n_794;
wire n_2848;
wire n_3306;
wire n_2185;
wire n_4345;
wire n_1292;
wire n_1026;
wire n_3460;
wire n_1610;
wire n_2202;
wire n_2952;
wire n_3530;
wire n_2693;
wire n_3240;
wire n_931;
wire n_3362;
wire n_4992;
wire n_4130;
wire n_967;
wire n_4175;
wire n_1079;
wire n_3393;
wire n_2836;
wire n_2864;
wire n_4456;
wire n_1717;
wire n_2172;
wire n_2601;
wire n_2365;
wire n_1880;
wire n_1399;
wire n_1855;
wire n_2333;
wire n_3629;
wire n_4948;
wire n_1903;
wire n_2147;
wire n_4020;
wire n_2224;
wire n_1226;
wire n_1970;
wire n_3724;
wire n_3287;
wire n_2167;
wire n_3046;
wire n_2293;
wire n_2921;
wire n_1240;
wire n_4984;
wire n_4055;
wire n_4410;
wire n_3980;
wire n_3257;
wire n_3730;
wire n_3979;
wire n_2695;
wire n_2598;
wire n_3727;
wire n_976;
wire n_4003;
wire n_1832;
wire n_767;
wire n_2302;
wire n_3014;
wire n_2294;
wire n_2274;
wire n_3342;
wire n_2895;
wire n_3796;
wire n_3884;
wire n_4492;
wire n_3625;
wire n_3375;
wire n_2768;
wire n_3760;
wire n_4975;
wire n_3515;
wire n_2363;
wire n_2728;
wire n_2025;
wire n_3744;
wire n_4022;
wire n_1020;
wire n_2495;
wire n_1058;
wire n_4336;
wire n_2223;
wire n_1279;
wire n_2511;
wire n_3981;
wire n_2681;
wire n_1689;
wire n_2535;
wire n_1255;
wire n_3031;
wire n_2335;
wire n_3215;
wire n_1401;
wire n_3138;
wire n_776;
wire n_2860;
wire n_2041;
wire n_1933;
wire n_4494;
wire n_4201;
wire n_4719;
wire n_3577;
wire n_4074;
wire n_3994;
wire n_4636;
wire n_4983;
wire n_3185;
wire n_1217;
wire n_2662;
wire n_4386;
wire n_3917;
wire n_1231;
wire n_4275;
wire n_3774;
wire n_926;
wire n_2296;
wire n_2178;
wire n_4243;
wire n_2765;
wire n_4225;
wire n_4658;
wire n_4186;
wire n_1501;
wire n_2241;
wire n_4699;
wire n_4096;
wire n_2531;
wire n_1570;
wire n_3377;
wire n_1518;
wire n_4907;
wire n_3961;
wire n_855;
wire n_2059;
wire n_4713;
wire n_1287;
wire n_1611;
wire n_3374;
wire n_4870;
wire n_4818;
wire n_4916;
wire n_4323;
wire n_1899;
wire n_3508;
wire n_4129;
wire n_1105;
wire n_3599;
wire n_4480;
wire n_3734;
wire n_3401;
wire n_983;
wire n_699;
wire n_3542;
wire n_3263;
wire n_2523;
wire n_1945;
wire n_2418;
wire n_1377;
wire n_1614;
wire n_3819;
wire n_3222;
wire n_1740;
wire n_4616;
wire n_1092;
wire n_3205;
wire n_4374;
wire n_2225;
wire n_1963;
wire n_3868;
wire n_729;
wire n_2218;
wire n_1122;
wire n_1408;
wire n_2593;
wire n_1693;
wire n_2741;
wire n_2184;
wire n_2714;
wire n_2754;
wire n_4580;
wire n_1218;
wire n_3611;
wire n_4826;
wire n_3959;
wire n_3338;
wire n_2962;
wire n_4514;
wire n_1543;
wire n_877;
wire n_3995;
wire n_3908;
wire n_1055;
wire n_1395;
wire n_3892;
wire n_1346;
wire n_1089;
wire n_1502;
wire n_3501;
wire n_1478;
wire n_2555;
wire n_3216;
wire n_3568;
wire n_2708;
wire n_735;
wire n_4844;
wire n_1294;
wire n_4049;
wire n_2661;
wire n_845;
wire n_1649;
wire n_2470;
wire n_1297;
wire n_3551;
wire n_1708;
wire n_4677;
wire n_4525;
wire n_3364;
wire n_2643;
wire n_755;
wire n_3766;
wire n_3985;
wire n_4369;
wire n_3826;
wire n_2266;
wire n_4324;
wire n_842;
wire n_1898;
wire n_1741;
wire n_1907;
wire n_742;
wire n_1719;
wire n_2742;
wire n_769;
wire n_3671;
wire n_2366;
wire n_1753;
wire n_1372;
wire n_1895;
wire n_4104;
wire n_982;
wire n_3791;
wire n_915;
wire n_2008;
wire n_4989;
wire n_3064;
wire n_3199;
wire n_2127;
wire n_3151;
wire n_3016;
wire n_2460;
wire n_1319;
wire n_3367;
wire n_3669;
wire n_3956;
wire n_4898;
wire n_4081;
wire n_2292;
wire n_2480;
wire n_606;
wire n_4528;
wire n_2772;
wire n_1700;
wire n_659;
wire n_1332;
wire n_1747;
wire n_3990;
wire n_1171;
wire n_4069;
wire n_3582;
wire n_4280;
wire n_1867;
wire n_3993;
wire n_2576;
wire n_3459;
wire n_4811;
wire n_2696;
wire n_4779;
wire n_2140;
wire n_2157;
wire n_1966;
wire n_1400;
wire n_3735;
wire n_1527;
wire n_1513;
wire n_3656;
wire n_4524;
wire n_2831;
wire n_3069;
wire n_4657;
wire n_4891;
wire n_2629;
wire n_3369;
wire n_1257;
wire n_1954;
wire n_3964;
wire n_3302;
wire n_2486;
wire n_1897;
wire n_2137;
wire n_3685;
wire n_4977;
wire n_2492;
wire n_2939;
wire n_3425;
wire n_4876;
wire n_1449;
wire n_2900;
wire n_797;
wire n_2912;
wire n_595;
wire n_1405;
wire n_3813;
wire n_2622;
wire n_3447;
wire n_1757;
wire n_2264;
wire n_1950;
wire n_805;
wire n_2032;
wire n_2090;
wire n_3124;
wire n_3811;
wire n_4200;
wire n_2249;
wire n_3411;
wire n_3463;
wire n_2785;
wire n_730;
wire n_4938;
wire n_1281;
wire n_2574;
wire n_2364;
wire n_1856;
wire n_1524;
wire n_2928;
wire n_1118;
wire n_4604;
wire n_2905;
wire n_2884;
wire n_3408;
wire n_1293;
wire n_961;
wire n_726;
wire n_878;
wire n_4118;
wire n_3857;
wire n_3110;
wire n_4239;
wire n_3157;
wire n_1180;
wire n_1697;
wire n_2730;
wire n_806;
wire n_1350;
wire n_4704;
wire n_2720;
wire n_649;
wire n_1561;
wire n_2405;
wire n_2700;
wire n_1616;
wire n_2416;
wire n_2064;
wire n_3640;
wire n_1557;
wire n_4744;
wire n_4706;
wire n_3879;
wire n_2022;
wire n_4343;
wire n_1505;
wire n_2408;
wire n_4764;
wire n_4990;
wire n_2986;
wire n_949;
wire n_2454;
wire n_3591;
wire n_2760;
wire n_4919;
wire n_1208;
wire n_3317;
wire n_4835;
wire n_1151;
wire n_4420;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_4251;
wire n_4559;
wire n_4742;
wire n_3566;
wire n_1133;
wire n_883;
wire n_4372;
wire n_4097;
wire n_4162;
wire n_779;
wire n_4790;
wire n_594;
wire n_4173;
wire n_3573;
wire n_2943;
wire n_3319;
wire n_2247;
wire n_2230;
wire n_1269;
wire n_4727;
wire n_1547;
wire n_1438;
wire n_3654;
wire n_1047;
wire n_3783;
wire n_4008;
wire n_2158;
wire n_3643;
wire n_2285;
wire n_3184;
wire n_1288;
wire n_2173;
wire n_3982;
wire n_3647;
wire n_1143;
wire n_3973;
wire n_4799;
wire n_4534;
wire n_4960;
wire n_1153;
wire n_1103;
wire n_3738;
wire n_894;
wire n_1380;
wire n_2020;
wire n_2310;
wire n_3600;
wire n_1023;
wire n_914;
wire n_689;
wire n_4327;
wire n_3190;
wire n_3027;
wire n_4011;
wire n_3695;
wire n_3800;
wire n_3462;
wire n_3906;
wire n_3011;
wire n_3395;
wire n_2820;
wire n_3733;
wire n_1165;
wire n_3967;
wire n_588;
wire n_638;
wire n_4370;
wire n_4816;
wire n_4091;
wire n_1417;
wire n_3096;
wire n_4166;
wire n_2777;
wire n_2234;
wire n_1341;
wire n_3233;
wire n_2431;
wire n_3322;
wire n_1603;
wire n_4478;
wire n_2935;
wire n_4246;
wire n_715;
wire n_1066;
wire n_2863;
wire n_2331;
wire n_4632;
wire n_685;
wire n_4061;
wire n_2920;
wire n_1712;
wire n_3344;
wire n_4754;
wire n_1534;
wire n_1290;
wire n_4375;
wire n_617;
wire n_2396;
wire n_3368;
wire n_1559;
wire n_3117;
wire n_4684;
wire n_743;
wire n_1546;
wire n_3384;
wire n_2592;
wire n_3490;
wire n_962;
wire n_4241;
wire n_1622;
wire n_2751;
wire n_3113;
wire n_4183;
wire n_1968;
wire n_918;
wire n_639;
wire n_673;
wire n_2842;
wire n_2196;
wire n_3603;
wire n_2371;
wire n_1978;
wire n_3720;
wire n_2560;
wire n_4256;
wire n_1164;
wire n_1193;
wire n_1345;
wire n_3037;
wire n_1336;
wire n_1033;
wire n_4333;
wire n_1166;
wire n_2007;
wire n_3363;
wire n_1158;
wire n_1803;
wire n_872;
wire n_3522;
wire n_4455;
wire n_3241;
wire n_3899;
wire n_3481;
wire n_2236;
wire n_692;
wire n_4457;
wire n_2150;
wire n_1816;
wire n_2803;
wire n_2887;
wire n_2648;
wire n_4735;
wire n_3305;
wire n_3810;
wire n_4062;
wire n_2093;
wire n_3354;
wire n_2204;
wire n_1481;
wire n_2040;
wire n_2151;
wire n_2455;
wire n_827;
wire n_3437;
wire n_2231;
wire n_4212;
wire n_622;
wire n_4584;
wire n_3574;
wire n_2530;
wire n_2289;
wire n_2299;
wire n_751;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_4477;
wire n_4110;
wire n_1221;
wire n_4217;
wire n_1262;
wire n_792;
wire n_1942;
wire n_2951;
wire n_3807;
wire n_4048;
wire n_1579;
wire n_4949;
wire n_2181;
wire n_2014;
wire n_2974;
wire n_923;
wire n_1124;
wire n_1326;
wire n_3969;
wire n_2282;
wire n_4605;
wire n_981;
wire n_3873;
wire n_4649;
wire n_1204;
wire n_994;
wire n_2428;
wire n_1360;
wire n_2858;
wire n_3076;
wire n_3410;
wire n_856;
wire n_4592;
wire n_1564;
wire n_2872;
wire n_3701;
wire n_3706;
wire n_4820;
wire n_1858;
wire n_1678;
wire n_2589;
wire n_4086;
wire n_1482;
wire n_1361;
wire n_4656;
wire n_1520;
wire n_4862;
wire n_1411;
wire n_1359;
wire n_3536;
wire n_1721;
wire n_3782;
wire n_1317;
wire n_3594;
wire n_2385;
wire n_1980;
wire n_4177;
wire n_2501;
wire n_1385;
wire n_1998;
wire n_2675;
wire n_2604;
wire n_3521;
wire n_3855;
wire n_2985;
wire n_2630;
wire n_2028;
wire n_919;
wire n_3114;
wire n_2092;
wire n_3622;
wire n_2817;
wire n_2773;
wire n_2402;
wire n_1458;
wire n_679;
wire n_3047;
wire n_3163;
wire n_1550;
wire n_1358;
wire n_1200;
wire n_826;
wire n_2808;
wire n_2344;
wire n_3520;
wire n_2392;
wire n_3272;
wire n_3122;
wire n_607;
wire n_3687;
wire n_2787;
wire n_3799;
wire n_3133;
wire n_2805;
wire n_1268;
wire n_2676;
wire n_2770;
wire n_4550;
wire n_4347;
wire n_702;
wire n_4933;
wire n_968;
wire n_4144;
wire n_2375;
wire n_3278;
wire n_4167;
wire n_3608;
wire n_4895;
wire n_1282;
wire n_4726;
wire n_1755;
wire n_2212;
wire n_4434;
wire n_2569;
wire n_4019;
wire n_4199;
wire n_816;
wire n_1322;
wire n_3829;
wire n_4510;
wire n_2469;
wire n_1125;
wire n_2358;
wire n_1710;
wire n_3546;
wire n_2355;
wire n_1390;
wire n_3068;
wire n_1629;
wire n_1094;
wire n_1510;
wire n_3002;
wire n_1099;
wire n_4899;
wire n_3146;
wire n_3038;
wire n_759;
wire n_4156;
wire n_1727;
wire n_3693;
wire n_3132;
wire n_831;
wire n_3681;
wire n_3970;
wire n_778;
wire n_2351;
wire n_1619;
wire n_3188;
wire n_4448;
wire n_3218;
wire n_1152;
wire n_2447;
wire n_2101;
wire n_4193;
wire n_1236;
wire n_4579;
wire n_4776;
wire n_671;
wire n_2704;
wire n_1334;
wire n_3729;
wire n_4471;
wire n_4392;
wire n_3103;
wire n_2048;
wire n_3028;
wire n_4691;
wire n_3148;
wire n_3775;
wire n_684;
wire n_3966;
wire n_4397;
wire n_3616;
wire n_4753;
wire n_4803;
wire n_1289;
wire n_1831;
wire n_3874;
wire n_2191;
wire n_4165;
wire n_2056;
wire n_2852;
wire n_2515;
wire n_1600;
wire n_1144;
wire n_838;
wire n_1941;
wire n_3637;
wire n_1017;
wire n_734;
wire n_4893;
wire n_2240;
wire n_4258;
wire n_709;
wire n_2917;
wire n_3194;
wire n_2085;
wire n_2432;
wire n_1686;
wire n_4232;
wire n_2097;
wire n_662;
wire n_3461;
wire n_1410;
wire n_939;
wire n_2297;
wire n_4203;
wire n_1325;
wire n_1223;
wire n_2957;
wire n_1983;
wire n_4767;
wire n_4569;
wire n_948;
wire n_3820;
wire n_3072;
wire n_2961;
wire n_4468;
wire n_1923;
wire n_3848;
wire n_3631;
wire n_4885;
wire n_1479;
wire n_4698;
wire n_1031;
wire n_3674;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_3763;
wire n_933;
wire n_3499;
wire n_1821;
wire n_3910;
wire n_3947;
wire n_2585;
wire n_3361;
wire n_2995;
wire n_4533;
wire n_4287;
wire n_3228;
wire n_2164;
wire n_1732;
wire n_2678;
wire n_1186;
wire n_2052;
wire n_4761;
wire n_4627;
wire n_4556;
wire n_2205;
wire n_2183;
wire n_1724;
wire n_3088;
wire n_1707;
wire n_2080;
wire n_3590;
wire n_1126;
wire n_2761;
wire n_2357;
wire n_4520;
wire n_895;
wire n_1639;
wire n_2421;
wire n_1302;
wire n_3295;
wire n_626;
wire n_3849;
wire n_4263;
wire n_4444;
wire n_1818;
wire n_4265;
wire n_3557;
wire n_1598;
wire n_2269;
wire n_1583;
wire n_4612;
wire n_1264;
wire n_4149;
wire n_1827;
wire n_4958;
wire n_1752;
wire n_2361;
wire n_4538;
wire n_3030;
wire n_3505;
wire n_3075;
wire n_1102;
wire n_2239;
wire n_1296;
wire n_4730;
wire n_4421;
wire n_2464;
wire n_3697;
wire n_882;
wire n_2304;
wire n_2514;
wire n_1299;
wire n_3430;
wire n_2063;
wire n_3489;
wire n_2079;
wire n_2152;
wire n_4967;
wire n_2517;
wire n_4696;
wire n_3484;
wire n_4971;
wire n_2095;
wire n_2738;
wire n_2590;
wire n_4661;
wire n_2797;
wire n_3041;
wire n_1421;
wire n_2208;
wire n_2423;
wire n_4376;
wire n_3832;
wire n_3525;
wire n_3712;
wire n_1069;
wire n_4305;
wire n_2037;
wire n_2953;
wire n_2823;
wire n_3684;
wire n_913;
wire n_1681;
wire n_4834;
wire n_1507;
wire n_589;
wire n_2866;
wire n_3153;
wire n_1174;
wire n_2346;
wire n_4692;
wire n_1353;
wire n_3268;
wire n_2559;
wire n_1383;
wire n_603;
wire n_4259;
wire n_2030;
wire n_850;
wire n_4299;
wire n_2407;
wire n_690;
wire n_2243;
wire n_2694;
wire n_3742;
wire n_4965;
wire n_1837;
wire n_4178;
wire n_2006;
wire n_4953;
wire n_4813;
wire n_3352;
wire n_2367;
wire n_2731;
wire n_3703;
wire n_1246;
wire n_2123;
wire n_2238;
wire n_4802;
wire n_4793;
wire n_1196;
wire n_3435;
wire n_2380;
wire n_1187;
wire n_4897;
wire n_1298;
wire n_1745;
wire n_4674;
wire n_4796;
wire n_1088;
wire n_766;
wire n_2750;
wire n_2547;
wire n_945;
wire n_4575;
wire n_3665;
wire n_3063;
wire n_3281;
wire n_3535;
wire n_2288;
wire n_3858;
wire n_4653;
wire n_4589;
wire n_3220;
wire n_4581;
wire n_665;
wire n_4625;
wire n_2107;
wire n_4845;
wire n_4148;
wire n_3679;
wire n_738;
wire n_672;
wire n_4968;
wire n_2342;
wire n_4590;
wire n_3856;
wire n_4038;
wire n_2735;
wire n_953;
wire n_4214;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_2709;
wire n_3419;
wire n_989;
wire n_2233;
wire n_795;
wire n_4892;
wire n_1936;
wire n_3890;
wire n_821;
wire n_770;
wire n_1514;
wire n_2782;
wire n_3929;
wire n_971;
wire n_4353;
wire n_2201;
wire n_4950;
wire n_1650;
wire n_4176;
wire n_4124;
wire n_4431;
wire n_1404;
wire n_3347;
wire n_4797;
wire n_4823;
wire n_4488;
wire n_2779;
wire n_3627;
wire n_3596;
wire n_3756;
wire n_4077;
wire n_3209;
wire n_4608;
wire n_3948;
wire n_4839;
wire n_1074;
wire n_1765;
wire n_1977;
wire n_2650;
wire n_4454;
wire n_4184;
wire n_2332;
wire n_2391;
wire n_611;
wire n_1295;
wire n_2060;
wire n_3883;
wire n_1013;
wire n_4032;
wire n_2571;
wire n_4929;
wire n_2874;
wire n_4117;
wire n_3049;
wire n_3634;
wire n_2341;
wire n_1654;
wire n_3066;
wire n_2045;
wire n_3913;
wire n_2575;
wire n_3739;
wire n_1230;
wire n_1597;
wire n_2942;
wire n_1771;
wire n_4541;
wire n_3271;
wire n_3164;
wire n_3861;
wire n_2043;
wire n_4171;
wire n_4815;
wire n_4665;
wire n_4884;
wire n_3580;
wire n_1437;
wire n_4276;
wire n_1378;
wire n_1461;
wire n_1876;
wire n_1830;
wire n_1112;
wire n_700;
wire n_4174;
wire n_2145;
wire n_4801;
wire n_680;
wire n_4582;
wire n_4774;
wire n_4108;
wire n_3119;
wire n_4740;
wire n_1108;
wire n_1274;
wire n_4394;
wire n_4920;
wire n_3909;
wire n_4220;
wire n_2703;
wire n_577;
wire n_916;
wire n_2810;
wire n_1884;
wire n_1555;
wire n_762;
wire n_1253;
wire n_4378;
wire n_1468;
wire n_2683;
wire n_4180;
wire n_4459;
wire n_3624;
wire n_1182;
wire n_4594;
wire n_2748;
wire n_4642;
wire n_1376;
wire n_2925;
wire n_1435;
wire n_1750;
wire n_1506;
wire n_3544;
wire n_2072;
wire n_3852;
wire n_1491;
wire n_2628;
wire n_3219;
wire n_1083;
wire n_4914;
wire n_3510;
wire n_4587;
wire n_1139;
wire n_3688;
wire n_1312;
wire n_3871;
wire n_892;
wire n_3757;
wire n_1567;
wire n_2219;
wire n_2100;
wire n_3666;
wire n_990;
wire n_867;
wire n_3479;
wire n_944;
wire n_749;
wire n_2888;
wire n_3998;
wire n_4150;
wire n_1920;
wire n_4285;
wire n_2668;
wire n_2701;
wire n_2400;
wire n_650;
wire n_3741;
wire n_2567;
wire n_2557;
wire n_1908;
wire n_1155;
wire n_2755;
wire n_1071;
wire n_712;
wire n_909;
wire n_1392;
wire n_2066;
wire n_2762;
wire n_964;
wire n_2220;
wire n_4433;
wire n_2829;
wire n_1914;
wire n_2253;
wire n_2130;
wire n_4861;
wire n_2021;
wire n_1563;
wire n_3673;
wire n_3052;
wire n_2507;
wire n_1633;
wire n_4621;
wire n_3187;
wire n_4451;
wire n_2328;
wire n_2434;
wire n_1234;
wire n_3936;
wire n_2261;
wire n_3082;
wire n_2473;
wire n_4784;
wire n_2438;
wire n_3210;
wire n_3867;
wire n_3397;
wire n_1646;
wire n_2262;
wire n_4613;
wire n_2565;
wire n_1237;
wire n_1095;
wire n_3078;
wire n_3971;
wire n_4979;
wire n_3869;
wire n_1531;
wire n_2113;
wire n_1387;
wire n_3711;
wire n_3171;
wire n_4751;
wire n_4242;
wire n_1951;
wire n_2490;
wire n_2558;
wire n_1496;
wire n_2812;
wire n_3300;
wire n_3104;
wire n_4122;
wire n_2132;
wire n_4522;
wire n_4952;
wire n_4426;
wire n_4362;
wire n_3267;
wire n_3946;
wire n_2112;
wire n_2640;
wire n_4634;
wire n_4932;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2983;
wire n_4089;
wire n_3513;
wire n_1173;
wire n_3498;
wire n_2350;
wire n_1068;
wire n_1198;
wire n_4506;
wire n_4728;
wire n_1886;
wire n_4346;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2481;
wire n_3863;
wire n_2327;
wire n_3882;
wire n_3916;
wire n_1365;
wire n_3968;
wire n_3675;
wire n_2437;
wire n_2841;
wire n_3332;
wire n_2055;
wire n_2998;
wire n_1423;
wire n_4359;
wire n_1609;
wire n_2822;
wire n_2308;
wire n_1939;
wire n_2242;
wire n_4447;
wire n_2937;
wire n_4293;
wire n_4039;
wire n_1798;
wire n_3057;
wire n_1608;
wire n_677;
wire n_3983;
wire n_703;
wire n_3318;
wire n_3385;
wire n_3773;
wire n_3494;
wire n_1278;
wire n_3788;
wire n_3939;
wire n_590;
wire n_727;
wire n_3569;
wire n_3837;
wire n_4942;
wire n_3835;
wire n_2496;
wire n_3260;
wire n_3349;
wire n_4348;
wire n_1602;
wire n_3139;
wire n_3801;
wire n_2338;
wire n_1080;
wire n_3636;
wire n_3653;
wire n_3823;
wire n_3403;
wire n_2057;
wire n_1205;
wire n_2716;
wire n_2944;
wire n_2780;
wire n_3439;
wire n_1120;
wire n_1202;
wire n_4084;
wire n_627;
wire n_1371;
wire n_4240;
wire n_2033;
wire n_4121;
wire n_3602;
wire n_2774;
wire n_2799;
wire n_4393;
wire n_3984;
wire n_1586;
wire n_1431;
wire n_4389;
wire n_1763;
wire n_4461;
wire n_2763;
wire n_3156;
wire n_1859;
wire n_2660;
wire n_3426;
wire n_4615;
wire n_3044;
wire n_3492;
wire n_3737;
wire n_2379;
wire n_3579;
wire n_1667;
wire n_888;
wire n_3896;
wire n_2300;
wire n_4067;
wire n_1677;
wire n_4551;
wire n_4521;
wire n_2284;
wire n_3005;
wire n_2283;
wire n_582;
wire n_2526;
wire n_1097;
wire n_1711;
wire n_4387;
wire n_2508;
wire n_3186;
wire n_2594;
wire n_1239;
wire n_3417;
wire n_890;
wire n_3626;
wire n_4598;
wire n_4464;
wire n_4789;
wire n_3180;
wire n_3423;
wire n_1081;
wire n_2119;
wire n_2493;
wire n_4565;
wire n_3392;
wire n_1800;
wire n_2904;
wire n_3353;
wire n_2946;
wire n_3512;
wire n_1860;
wire n_1734;
wire n_4552;
wire n_2840;
wire n_4482;
wire n_837;
wire n_812;
wire n_4172;
wire n_4040;
wire n_3024;
wire n_4328;
wire n_1854;
wire n_666;
wire n_1206;
wire n_1729;
wire n_1508;
wire n_2893;
wire n_4940;
wire n_785;
wire n_3161;
wire n_2389;
wire n_1309;
wire n_999;
wire n_2280;
wire n_1394;
wire n_3365;
wire n_4113;
wire n_873;
wire n_3977;
wire n_2468;
wire n_2171;
wire n_4112;
wire n_2035;
wire n_4928;
wire n_2614;
wire n_2494;
wire n_1538;
wire n_4865;
wire n_2128;
wire n_4071;
wire n_4436;
wire n_3586;
wire n_4160;
wire n_1668;
wire n_4137;
wire n_1078;
wire n_4545;
wire n_4758;
wire n_1161;
wire n_4840;
wire n_3097;
wire n_4395;
wire n_4873;
wire n_3507;
wire n_618;
wire n_1191;
wire n_4535;
wire n_4385;
wire n_1215;
wire n_3748;
wire n_4731;
wire n_2337;
wire n_1786;
wire n_3732;
wire n_1804;
wire n_4671;
wire n_2272;
wire n_4766;
wire n_592;
wire n_4558;
wire n_1318;
wire n_1632;
wire n_1769;
wire n_1929;
wire n_4319;
wire n_2929;
wire n_4358;
wire n_1526;
wire n_4874;
wire n_2656;
wire n_4904;
wire n_1997;
wire n_1137;
wire n_1258;
wire n_640;
wire n_1733;
wire n_4651;
wire n_943;
wire n_3167;
wire n_4748;
wire n_1807;
wire n_1123;
wire n_2857;
wire n_1784;
wire n_4618;
wire n_3787;
wire n_4025;
wire n_1321;
wire n_3050;
wire n_3919;
wire n_752;
wire n_985;
wire n_2412;
wire n_3298;
wire n_3107;
wire n_1352;
wire n_643;
wire n_2383;
wire n_2764;
wire n_1441;
wire n_1822;
wire n_682;
wire n_2633;
wire n_3708;
wire n_2907;
wire n_1429;
wire n_2353;
wire n_2528;
wire n_1778;
wire n_686;
wire n_1154;
wire n_584;
wire n_4910;
wire n_1759;
wire n_2325;
wire n_4724;
wire n_1130;
wire n_3718;
wire n_756;
wire n_3390;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_4666;
wire n_4082;
wire n_2320;
wire n_3140;
wire n_979;
wire n_3976;
wire n_2813;
wire n_897;
wire n_2546;
wire n_3381;
wire n_3736;
wire n_4466;
wire n_891;
wire n_885;
wire n_1659;
wire n_3955;
wire n_1864;
wire n_3086;
wire n_1887;
wire n_3165;
wire n_3336;
wire n_3635;
wire n_3541;
wire n_2502;
wire n_714;
wire n_3605;
wire n_2170;
wire n_4721;
wire n_725;
wire n_1577;
wire n_3840;
wire n_2198;
wire n_3067;
wire n_3809;
wire n_4921;
wire n_1852;
wire n_801;
wire n_4377;
wire n_818;
wire n_2410;
wire n_2314;
wire n_3468;
wire n_1877;
wire n_4301;
wire n_2133;
wire n_2497;
wire n_879;
wire n_4561;
wire n_1541;
wire n_597;
wire n_3291;
wire n_1472;
wire n_1050;
wire n_2578;
wire n_1201;
wire n_1185;
wire n_2475;
wire n_4715;
wire n_2715;
wire n_2665;
wire n_4879;
wire n_3755;
wire n_1090;
wire n_4536;
wire n_4304;
wire n_4927;
wire n_4078;
wire n_1624;
wire n_1801;
wire n_2854;
wire n_4418;
wire n_3341;
wire n_4125;
wire n_1116;
wire n_3043;
wire n_2747;
wire n_1511;
wire n_3226;
wire n_3378;
wire n_1641;
wire n_3731;
wire n_4527;
wire n_4291;
wire n_2845;
wire n_4151;
wire n_4412;
wire n_2036;
wire n_843;
wire n_3358;
wire n_2003;
wire n_2533;
wire n_1307;
wire n_4682;
wire n_1128;
wire n_2419;
wire n_2330;
wire n_4810;
wire n_3189;
wire n_2309;
wire n_4957;
wire n_4855;
wire n_1955;
wire n_3289;
wire n_1440;
wire n_1370;
wire n_1549;
wire n_2658;
wire n_3620;
wire n_4601;
wire n_1065;
wire n_4518;
wire n_2767;
wire n_3376;
wire n_1362;
wire n_3123;
wire n_2692;
wire n_683;
wire n_1300;
wire n_1960;
wire n_4102;
wire n_4308;
wire n_2862;
wire n_4325;
wire n_1420;
wire n_2645;
wire n_2553;
wire n_4711;
wire n_2749;
wire n_660;
wire n_4413;
wire n_1210;
wire n_3307;
wire n_1885;
wire n_3251;
wire n_3288;
wire n_2833;
wire n_1038;
wire n_3723;
wire n_4135;
wire n_3880;
wire n_3904;
wire n_3008;
wire n_4821;
wire n_3242;
wire n_3405;
wire n_2313;
wire n_613;
wire n_1022;
wire n_3532;
wire n_2609;
wire n_1767;
wire n_4138;
wire n_1040;
wire n_3131;
wire n_1973;
wire n_1444;
wire n_820;
wire n_2882;
wire n_2303;
wire n_4384;
wire n_4639;
wire n_1664;
wire n_4577;
wire n_2154;
wire n_1986;
wire n_2624;
wire n_2054;
wire n_1857;
wire n_3926;
wire n_4481;
wire n_984;
wire n_1552;
wire n_2938;
wire n_2498;
wire n_3992;
wire n_621;
wire n_1772;
wire n_1311;
wire n_3106;
wire n_2881;
wire n_3092;
wire n_4270;
wire n_697;
wire n_4620;
wire n_4924;
wire n_4044;
wire n_2305;
wire n_880;
wire n_3304;
wire n_4388;
wire n_3247;
wire n_739;
wire n_1028;
wire n_4271;
wire n_2180;
wire n_4406;
wire n_2809;
wire n_975;
wire n_1645;
wire n_932;
wire n_2276;
wire n_3301;
wire n_2910;
wire n_2503;
wire n_3785;
wire n_2465;
wire n_2972;
wire n_4401;
wire n_2586;
wire n_2989;
wire n_3178;
wire n_2251;
wire n_3100;
wire n_3721;
wire n_3389;
wire n_2126;
wire n_2425;
wire n_4973;
wire n_4792;
wire n_1601;
wire n_3537;
wire n_4402;
wire n_2487;
wire n_1834;
wire n_1011;
wire n_2534;
wire n_2941;
wire n_4286;
wire n_3638;
wire n_3576;
wire n_4858;
wire n_1445;
wire n_4435;
wire n_3248;
wire n_2387;
wire n_4318;
wire n_830;
wire n_987;
wire n_2510;
wire n_3570;
wire n_3227;
wire n_4673;
wire n_2793;
wire n_2639;
wire n_4738;
wire n_2603;
wire n_1167;
wire n_4554;
wire n_4526;
wire n_4105;
wire n_969;
wire n_3663;
wire n_1663;
wire n_2086;
wire n_1926;
wire n_1630;
wire n_663;
wire n_1720;
wire n_2409;
wire n_2966;
wire n_3431;
wire n_3355;
wire n_1738;
wire n_3897;
wire n_1735;
wire n_4005;
wire n_4181;
wire n_2543;
wire n_2321;
wire n_1077;
wire n_2597;
wire n_956;
wire n_765;
wire n_4092;
wire n_4875;
wire n_4255;
wire n_2758;
wire n_1271;
wire n_2186;
wire n_4647;
wire n_3575;
wire n_2471;
wire n_3042;
wire n_1067;
wire n_1323;
wire n_1937;
wire n_4142;
wire n_900;
wire n_3004;
wire n_1551;
wire n_4849;
wire n_2039;
wire n_1285;
wire n_733;
wire n_761;
wire n_3838;
wire n_4059;
wire n_2734;
wire n_4499;
wire n_4504;
wire n_3598;
wire n_4917;
wire n_2420;
wire n_648;
wire n_3273;
wire n_2918;
wire n_835;
wire n_1865;
wire n_2641;
wire n_2463;
wire n_2580;
wire n_1792;
wire n_2062;
wire n_4489;
wire n_822;
wire n_1459;
wire n_2153;
wire n_839;
wire n_1754;
wire n_4833;
wire n_3394;
wire n_2235;
wire n_1575;
wire n_4564;
wire n_1848;
wire n_1172;
wire n_3776;
wire n_2775;
wire n_3903;
wire n_3581;
wire n_3778;
wire n_4322;
wire n_2260;
wire n_1660;
wire n_1315;
wire n_4080;
wire n_2206;
wire n_997;
wire n_635;
wire n_1643;
wire n_4185;
wire n_1320;
wire n_3001;
wire n_4981;
wire n_2347;
wire n_4676;
wire n_2657;
wire n_2990;
wire n_2538;
wire n_2034;
wire n_3932;
wire n_1934;
wire n_2577;
wire n_2362;
wire n_4507;
wire n_4756;
wire n_1576;
wire n_2422;
wire n_654;
wire n_2933;
wire n_3387;
wire n_3952;
wire n_4365;
wire n_3584;
wire n_4349;
wire n_3446;
wire n_1059;
wire n_2736;
wire n_3825;
wire n_4198;
wire n_977;
wire n_2339;
wire n_2532;
wire n_4373;
wire n_1866;
wire n_2664;
wire n_4154;
wire n_4390;
wire n_1782;
wire n_4107;
wire n_1558;
wire n_2519;
wire n_4380;
wire n_4361;
wire n_4609;
wire n_2360;
wire n_4453;
wire n_723;
wire n_1393;
wire n_4571;
wire n_3137;
wire n_2544;
wire n_809;
wire n_3032;
wire n_4886;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1982;
wire n_641;
wire n_910;
wire n_4964;
wire n_4700;
wire n_4002;
wire n_1114;
wire n_1742;
wire n_4679;
wire n_3815;
wire n_1768;
wire n_2193;
wire n_2369;
wire n_1199;
wire n_1273;
wire n_2982;
wire n_4483;
wire n_3061;
wire n_2587;
wire n_3504;
wire n_4693;
wire n_1043;
wire n_4956;
wire n_2869;
wire n_4487;
wire n_2674;
wire n_1737;
wire n_1613;
wire n_3026;
wire n_2979;
wire n_4329;
wire n_4010;
wire n_4501;
wire n_4808;
wire n_3902;
wire n_3244;
wire n_1779;
wire n_2562;
wire n_3112;
wire n_954;
wire n_2051;
wire n_3196;
wire n_2673;
wire n_4678;
wire n_664;
wire n_1591;
wire n_2548;
wire n_3488;
wire n_2381;
wire n_2744;
wire n_1967;
wire n_2179;
wire n_1280;
wire n_3779;
wire n_599;
wire n_1063;
wire n_991;
wire n_2275;
wire n_4606;
wire n_3834;
wire n_4303;
wire n_2029;
wire n_1912;
wire n_3923;
wire n_938;
wire n_1891;
wire n_583;
wire n_1000;
wire n_4868;
wire n_4072;
wire n_2792;
wire n_4465;
wire n_2596;
wire n_3986;
wire n_3725;
wire n_4026;
wire n_4245;
wire n_2524;
wire n_3894;
wire n_1702;
wire n_4852;
wire n_3202;
wire n_4290;
wire n_4945;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1082;
wire n_1725;
wire n_2318;
wire n_866;
wire n_2819;
wire n_1722;
wire n_2229;
wire n_1644;
wire n_3547;
wire n_4014;
wire n_2551;
wire n_2255;
wire n_1252;
wire n_3045;
wire n_773;
wire n_4599;
wire n_2706;
wire n_4222;
wire n_718;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_2573;
wire n_2336;
wire n_1662;
wire n_3249;
wire n_3483;
wire n_4046;
wire n_4701;
wire n_1925;
wire n_782;
wire n_2915;
wire n_4869;
wire n_3213;
wire n_4047;
wire n_1244;
wire n_1796;
wire n_2719;
wire n_2876;
wire n_4063;
wire n_2778;
wire n_1574;
wire n_3033;
wire n_893;
wire n_1582;
wire n_1981;
wire n_2824;
wire n_4417;
wire n_796;
wire n_1374;
wire n_2089;
wire n_4688;
wire n_4939;
wire n_1486;
wire n_3619;
wire n_4013;
wire n_3434;
wire n_4342;
wire n_691;
wire n_4903;
wire n_2131;
wire n_3853;
wire n_4382;
wire n_2509;
wire n_4085;
wire n_2135;
wire n_4475;
wire n_1463;
wire n_4626;
wire n_924;
wire n_781;
wire n_2013;
wire n_4638;
wire n_2786;
wire n_4058;
wire n_4090;
wire n_4819;
wire n_2436;
wire n_3517;
wire n_1706;
wire n_2461;
wire n_3719;
wire n_634;
wire n_1214;
wire n_3526;
wire n_3888;
wire n_3198;
wire n_1853;
wire n_764;
wire n_1503;
wire n_1181;
wire n_1999;
wire n_4841;
wire n_4683;
wire n_2873;
wire n_2084;
wire n_3330;
wire n_3514;
wire n_3383;
wire n_1835;
wire n_3965;
wire n_1457;
wire n_3905;
wire n_3797;
wire n_1836;
wire n_3416;
wire n_4600;
wire n_1453;
wire n_3943;
wire n_3145;
wire n_2908;
wire n_4106;
wire n_2156;
wire n_1184;
wire n_754;
wire n_2323;
wire n_1073;
wire n_4549;
wire n_1277;
wire n_1746;
wire n_1062;
wire n_4702;
wire n_4954;
wire n_740;
wire n_1974;
wire n_4491;
wire n_2906;
wire n_3283;
wire n_4331;
wire n_4159;
wire n_3451;
wire n_4734;
wire n_2832;
wire n_1688;
wire n_2370;
wire n_1944;
wire n_2914;
wire n_1988;
wire n_1718;
wire n_4515;
wire n_2149;
wire n_2277;
wire n_2539;
wire n_2078;
wire n_1145;
wire n_4809;
wire n_787;
wire n_4012;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_4760;
wire n_1207;
wire n_3606;
wire n_2232;
wire n_1847;
wire n_4320;
wire n_1314;
wire n_1512;
wire n_884;
wire n_4980;
wire n_3324;
wire n_2192;
wire n_2988;
wire n_4560;
wire n_3230;
wire n_3793;
wire n_859;
wire n_4768;
wire n_1889;
wire n_693;
wire n_929;
wire n_3207;
wire n_3641;
wire n_3828;
wire n_1850;
wire n_3183;
wire n_3607;
wire n_1637;
wire n_2427;
wire n_3613;
wire n_2885;
wire n_2098;
wire n_2616;
wire n_1751;
wire n_2769;
wire n_1548;
wire n_4987;
wire n_3013;
wire n_4572;
wire n_1396;
wire n_2739;
wire n_3962;
wire n_4988;
wire n_2902;
wire n_4360;
wire n_1544;
wire n_4540;
wire n_2094;
wire n_3854;
wire n_1354;
wire n_2349;
wire n_3652;
wire n_3449;
wire n_1021;
wire n_3089;
wire n_4854;
wire n_1595;
wire n_1142;
wire n_2727;
wire n_942;
wire n_1416;
wire n_1599;
wire n_4747;
wire n_3472;
wire n_2527;
wire n_3126;
wire n_2759;
wire n_4881;
wire n_2038;
wire n_3958;
wire n_4495;
wire n_4737;
wire n_1838;
wire n_4357;
wire n_2806;
wire n_4502;
wire n_3191;
wire n_1716;
wire n_3562;
wire n_2281;
wire n_3588;
wire n_1590;
wire n_3280;
wire n_4115;
wire n_1819;
wire n_3095;
wire n_947;
wire n_3698;
wire n_4513;
wire n_1179;
wire n_696;
wire n_1442;
wire n_4775;
wire n_2620;
wire n_1833;
wire n_1691;
wire n_2499;
wire n_2549;
wire n_804;
wire n_1656;
wire n_1382;
wire n_3093;
wire n_2970;
wire n_3885;
wire n_955;
wire n_4264;
wire n_2166;
wire n_3192;
wire n_4709;
wire n_1562;
wire n_3250;
wire n_4223;
wire n_3538;
wire n_3915;
wire n_3839;
wire n_1972;
wire n_4718;
wire n_3717;
wire n_3407;
wire n_3875;
wire n_4029;
wire n_4206;
wire n_2415;
wire n_4099;
wire n_3120;
wire n_2922;
wire n_3193;
wire n_2871;
wire n_4794;
wire n_4843;
wire n_669;
wire n_3937;
wire n_4763;
wire n_1418;
wire n_4170;
wire n_2462;
wire n_2155;
wire n_615;
wire n_2439;
wire n_4838;
wire n_4795;
wire n_3604;
wire n_824;
wire n_4272;
wire n_3176;
wire n_3792;
wire n_4267;
wire n_2083;
wire n_815;
wire n_2753;
wire n_1340;
wire n_3021;
wire n_4352;
wire n_2712;
wire n_1433;
wire n_3805;
wire n_3912;
wire n_3950;
wire n_2898;
wire n_1825;
wire n_3567;
wire n_2682;
wire n_1627;
wire n_2903;
wire n_3812;
wire n_3127;
wire n_1731;
wire n_799;
wire n_1147;
wire n_2378;
wire n_965;
wire n_934;
wire n_2213;
wire n_4056;
wire n_4806;
wire n_1674;
wire n_4015;
wire n_2924;
wire n_4445;
wire n_4462;
wire n_4219;
wire n_4484;
wire n_4723;
wire n_2142;
wire n_4517;
wire n_2896;
wire n_1913;
wire n_2069;
wire n_4043;
wire n_1042;
wire n_3170;
wire n_2311;
wire n_1455;
wire n_2287;
wire n_836;
wire n_3415;
wire n_3464;
wire n_3414;
wire n_4234;
wire n_760;
wire n_1483;
wire n_1363;
wire n_1111;
wire n_970;
wire n_3467;
wire n_713;
wire n_3179;
wire n_598;
wire n_4836;
wire n_3889;
wire n_3262;
wire n_927;
wire n_3699;
wire n_2120;
wire n_706;
wire n_1419;
wire n_3816;
wire n_3528;
wire n_4207;
wire n_2404;
wire n_2168;
wire n_2757;
wire n_4725;
wire n_2312;
wire n_1826;
wire n_4880;
wire n_2834;
wire n_4051;
wire n_3660;
wire n_4563;
wire n_2996;
wire n_637;
wire n_1259;
wire n_2801;
wire n_1177;
wire n_4334;
wire n_4978;
wire n_3246;
wire n_3299;
wire n_980;
wire n_1618;
wire n_1869;
wire n_3623;
wire n_905;
wire n_2718;
wire n_4707;
wire n_2687;
wire n_4923;
wire n_4911;
wire n_3876;
wire n_3615;
wire n_1802;
wire n_2811;
wire n_3019;
wire n_3200;
wire n_3642;
wire n_2146;
wire n_4274;
wire n_3276;
wire n_3682;
wire n_4007;
wire n_1456;
wire n_1879;
wire n_2129;
wire n_814;
wire n_578;
wire n_3572;
wire n_2975;
wire n_2399;
wire n_1134;
wire n_3471;
wire n_4075;
wire n_1484;
wire n_647;
wire n_2027;
wire n_2932;
wire n_600;
wire n_3118;
wire n_4441;
wire n_3039;
wire n_3922;
wire n_2195;
wire n_1467;
wire n_4458;
wire n_2159;
wire n_4889;
wire n_3831;
wire n_1744;
wire n_4523;
wire n_3618;
wire n_3705;
wire n_3022;
wire n_1709;
wire n_681;
wire n_3286;
wire n_2023;
wire n_3974;
wire n_3443;
wire n_2599;
wire n_3988;
wire n_2075;
wire n_1726;
wire n_2031;
wire n_3761;
wire n_3996;
wire n_4771;
wire n_2853;
wire n_3350;
wire n_1098;
wire n_3009;
wire n_777;
wire n_920;
wire n_3951;
wire n_3035;
wire n_4261;
wire n_1132;
wire n_1823;
wire n_4236;
wire n_3942;
wire n_3023;
wire n_2254;
wire n_3290;
wire n_1402;
wire n_3957;
wire n_3418;
wire n_1607;
wire n_861;
wire n_1666;
wire n_4648;
wire n_2214;
wire n_2256;
wire n_3326;
wire n_2732;
wire n_1883;
wire n_4094;
wire n_2776;
wire n_3224;
wire n_1969;
wire n_2949;
wire n_4269;
wire n_1927;
wire n_1222;
wire n_3803;
wire n_1919;
wire n_2994;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_4913;
wire n_2449;
wire n_4428;
wire n_745;
wire n_1572;
wire n_4463;
wire n_3648;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_4396;
wire n_1990;
wire n_3491;
wire n_2690;
wire n_3090;
wire n_2474;
wire n_2623;
wire n_1075;
wire n_1890;
wire n_4034;
wire n_4228;
wire n_1227;
wire n_3166;
wire n_3649;
wire n_3065;
wire n_657;
wire n_3924;
wire n_3997;
wire n_3564;
wire n_862;
wire n_2637;
wire n_3795;
wire n_4931;
wire n_2306;
wire n_2071;
wire n_3953;
wire n_4400;
wire n_2414;
wire n_2082;
wire n_2959;
wire n_1532;
wire n_1030;
wire n_3208;
wire n_1342;
wire n_2737;
wire n_3282;
wire n_852;
wire n_2916;
wire n_1060;
wire n_4424;
wire n_4351;
wire n_4192;
wire n_1748;
wire n_1301;
wire n_3400;
wire n_1466;
wire n_2581;
wire n_1783;
wire n_4646;
wire n_4221;
wire n_1037;
wire n_3650;
wire n_1329;
wire n_1993;
wire n_1545;
wire n_4035;
wire n_1480;
wire n_3670;
wire n_2540;
wire n_4190;
wire n_1605;
wire n_3060;
wire n_2984;
wire n_4009;
wire n_2489;
wire n_4145;
wire n_624;
wire n_876;
wire n_736;
wire n_2265;
wire n_3524;
wire n_2627;
wire n_1327;
wire n_1475;
wire n_2106;
wire n_4717;
wire n_4739;
wire n_3174;
wire n_3314;
wire n_602;
wire n_854;
wire n_2091;
wire n_4312;
wire n_3789;
wire n_1658;
wire n_1072;
wire n_1305;
wire n_4750;
wire n_2348;
wire n_1873;
wire n_2725;
wire n_2667;
wire n_3746;
wire n_4537;
wire n_1046;
wire n_3694;
wire n_771;
wire n_3893;
wire n_4847;
wire n_2307;
wire n_3702;
wire n_1984;
wire n_3453;
wire n_1556;
wire n_2815;
wire n_4427;
wire n_1824;
wire n_1492;
wire n_4065;
wire n_4705;
wire n_819;
wire n_1971;
wire n_2945;
wire n_586;
wire n_1324;
wire n_3543;
wire n_1776;
wire n_3448;
wire n_4279;
wire n_605;
wire n_2936;
wire n_3609;
wire n_4330;
wire n_4152;
wire n_2698;
wire n_4783;
wire n_3017;
wire n_2329;
wire n_2570;
wire n_1642;
wire n_2789;
wire n_2525;
wire n_2890;
wire n_4539;
wire n_3455;
wire n_807;
wire n_3907;
wire n_4603;
wire n_4332;
wire n_1987;
wire n_4052;
wire n_3357;
wire n_3388;
wire n_2368;
wire n_802;
wire n_4595;
wire n_960;
wire n_2352;
wire n_790;
wire n_4404;
wire n_2377;
wire n_2652;
wire n_4054;
wire n_1286;
wire n_4617;
wire n_1685;
wire n_2477;
wire n_4611;
wire n_2279;
wire n_3169;
wire n_2222;
wire n_1052;
wire n_4732;
wire n_2203;
wire n_2076;
wire n_1426;
wire n_4969;
wire n_4641;
wire n_4399;
wire n_4140;
wire n_2607;
wire n_3343;
wire n_4712;
wire n_3309;
wire n_2796;
wire n_858;
wire n_4817;
wire n_2136;
wire n_3134;
wire n_4909;
wire n_4755;
wire n_2771;
wire n_2403;
wire n_2947;
wire n_928;
wire n_3769;
wire n_1565;
wire n_4437;
wire n_3055;
wire n_4070;
wire n_748;
wire n_1045;
wire n_1881;
wire n_2635;
wire n_2999;
wire n_988;
wire n_4139;
wire n_4769;
wire n_1958;
wire n_4867;
wire n_3667;
wire n_2713;
wire n_1422;
wire n_1965;
wire n_644;
wire n_4450;
wire n_2934;
wire n_576;
wire n_2210;
wire n_4368;
wire n_3141;
wire n_2053;
wire n_3476;
wire n_1049;
wire n_4430;
wire n_3238;
wire n_2450;
wire n_1356;
wire n_1773;
wire n_3175;
wire n_4544;
wire n_2666;
wire n_728;
wire n_4191;
wire n_4409;
wire n_2401;
wire n_3255;
wire n_2588;
wire n_935;
wire n_2886;
wire n_4961;
wire n_3827;
wire n_2478;
wire n_911;
wire n_623;
wire n_3509;
wire n_1403;
wire n_3006;
wire n_4531;
wire n_3770;
wire n_3456;
wire n_4532;
wire n_601;
wire n_628;
wire n_3790;
wire n_907;
wire n_847;
wire n_747;
wire n_1135;
wire n_2566;
wire n_3101;
wire n_3662;
wire n_4257;
wire n_4282;
wire n_4341;
wire n_1694;
wire n_593;
wire n_1695;
wire n_4027;
wire n_4309;
wire n_4650;
wire n_609;
wire n_3077;
wire n_4944;
wire n_3478;
wire n_3062;
wire n_1774;
wire n_4994;
wire n_3533;
wire n_1994;
wire n_3978;
wire n_3836;
wire n_3409;
wire n_4381;
wire n_3583;
wire n_4316;
wire n_4860;
wire n_4469;
wire n_3540;
wire n_4930;
wire n_1157;
wire n_3563;
wire n_1739;
wire n_2642;
wire n_3310;
wire n_4423;
wire n_3689;
wire n_1789;
wire n_763;
wire n_2174;
wire n_3442;
wire n_3972;
wire n_2315;
wire n_4209;
wire n_4703;
wire n_1687;
wire n_4934;
wire n_2638;
wire n_2046;
wire n_1756;
wire n_4350;
wire n_1606;
wire n_1587;
wire n_2340;
wire n_4804;
wire n_2444;
wire n_4888;
wire n_1014;
wire n_1427;
wire n_2977;
wire n_3991;
wire n_4936;
wire n_2199;
wire n_4669;
wire n_1100;
wire n_585;
wire n_1617;
wire n_2600;
wire n_3436;
wire n_1962;
wire n_3806;
wire n_4759;
wire n_2114;
wire n_3329;
wire n_2927;
wire n_3833;
wire n_1175;
wire n_4887;
wire n_3751;
wire n_3402;
wire n_1621;
wire n_4585;
wire n_1785;
wire n_3406;
wire n_580;
wire n_3664;
wire n_4218;
wire n_4687;
wire n_1381;
wire n_3686;
wire n_1183;
wire n_4720;
wire n_2889;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_3470;
wire n_1407;
wire n_2865;
wire n_973;
wire n_4762;
wire n_3844;
wire n_3259;
wire n_2572;
wire n_4490;
wire n_1248;
wire n_1176;
wire n_3677;
wire n_1054;
wire n_3292;
wire n_3989;
wire n_4644;
wire n_4752;
wire n_4746;
wire n_1057;
wire n_4131;
wire n_4215;
wire n_978;
wire n_2488;
wire n_1509;
wire n_828;
wire n_4158;
wire n_3079;
wire n_3269;
wire n_4231;
wire n_2591;
wire n_653;
wire n_4926;
wire n_2050;
wire n_2197;
wire n_4872;
wire n_4778;
wire n_2550;
wire n_1536;
wire n_3177;
wire n_4667;
wire n_1471;
wire n_3440;
wire n_3658;
wire n_3404;
wire n_2291;
wire n_3346;
wire n_2816;
wire n_1620;
wire n_2542;
wire n_2165;
wire n_4837;
wire n_4210;
wire n_788;
wire n_2169;
wire n_591;
wire n_2175;
wire n_1625;
wire n_4578;
wire n_3644;
wire n_2176;
wire n_1412;
wire n_3059;
wire n_1922;
wire n_940;
wire n_1537;
wire n_4877;
wire n_2065;
wire n_4470;
wire n_4187;
wire n_1904;
wire n_2395;
wire n_2868;
wire n_1530;
wire n_4057;
wire n_631;
wire n_1170;
wire n_2724;
wire n_2258;
wire n_898;
wire n_3328;
wire n_2012;
wire n_3182;
wire n_2967;
wire n_1093;
wire n_4021;
wire n_3379;
wire n_4379;
wire n_2268;
wire n_3469;
wire n_1452;
wire n_2835;
wire n_668;
wire n_2111;
wire n_3743;
wire n_2948;
wire n_3099;
wire n_2897;
wire n_4812;
wire n_4497;
wire n_2583;
wire n_3155;
wire n_4300;
wire n_2024;
wire n_1770;
wire n_701;
wire n_1003;
wire n_4472;
wire n_2699;
wire n_3901;
wire n_1640;
wire n_2973;
wire n_2710;
wire n_2505;
wire n_4519;
wire n_2397;
wire n_3878;
wire n_4197;
wire n_2721;
wire n_1892;
wire n_2615;
wire n_4787;
wire n_1212;
wire n_4310;
wire n_4566;
wire n_3933;
wire n_4371;
wire n_1902;
wire n_2784;
wire n_3898;
wire n_694;
wire n_4749;
wire n_1845;
wire n_921;
wire n_2104;
wire n_2552;
wire n_1470;
wire n_1533;
wire n_3253;
wire n_2088;
wire n_1275;
wire n_4238;
wire n_904;
wire n_2005;
wire n_1696;
wire n_2108;
wire n_3824;
wire n_2246;
wire n_3846;
wire n_1497;
wire n_4189;
wire n_2472;
wire n_2705;
wire n_4479;
wire n_3845;
wire n_3203;
wire n_4986;
wire n_1316;
wire n_4668;
wire n_950;
wire n_711;
wire n_630;
wire n_4168;
wire n_1369;
wire n_4298;
wire n_4743;
wire n_1781;
wire n_4250;
wire n_3143;
wire n_3690;
wire n_3229;
wire n_2188;
wire n_2430;
wire n_2504;
wire n_4211;
wire n_3094;
wire n_741;
wire n_2964;
wire n_865;
wire n_3312;
wire n_1041;
wire n_2451;
wire n_2913;
wire n_993;
wire n_1862;
wire n_3752;
wire n_3672;
wire n_922;
wire n_1004;
wire n_2839;
wire n_3237;
wire n_4128;
wire n_4036;
wire n_3655;
wire n_2955;
wire n_1764;
wire n_4807;
wire n_902;
wire n_1723;
wire n_3918;
wire n_4101;
wire n_4915;
wire n_3866;
wire n_1946;
wire n_4383;
wire n_4830;
wire n_4391;
wire n_596;
wire n_4095;
wire n_1310;
wire n_4485;
wire n_3593;
wire n_1229;
wire n_2582;
wire n_3327;
wire n_4356;
wire n_1896;
wire n_1516;
wire n_4890;
wire n_2485;
wire n_2563;
wire n_4224;
wire n_1670;
wire n_1799;
wire n_4573;
wire n_1328;
wire n_4943;
wire n_2875;
wire n_3519;
wire n_2209;
wire n_4042;
wire n_4244;
wire n_1928;
wire n_4708;
wire n_4883;
wire n_4553;
wire n_1634;
wire n_1203;
wire n_1699;
wire n_2081;
wire n_937;
wire n_1474;
wire n_1631;
wire n_1794;
wire n_1375;
wire n_3053;
wire n_3772;
wire n_2891;
wire n_4335;
wire n_3128;
wire n_4277;
wire n_4614;
wire n_4629;
wire n_1002;
wire n_4516;
wire n_1129;
wire n_1464;
wire n_2798;
wire n_3217;
wire n_1249;
wire n_3821;
wire n_3201;
wire n_3503;
wire n_1870;
wire n_4467;
wire n_2654;
wire n_3935;
wire n_1861;
wire n_1228;
wire n_2319;
wire n_2965;
wire n_4955;
wire n_1251;
wire n_1989;
wire n_2689;
wire n_1762;
wire n_3798;
wire n_3080;
wire n_4248;
wire n_1672;
wire n_2228;
wire n_4645;
wire n_3308;
wire n_841;
wire n_3204;
wire n_4134;
wire n_3428;
wire n_2851;
wire n_4017;
wire n_2345;
wire n_1730;

INVx3_ASAP7_75t_L g576 ( 
.A(n_40),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_381),
.Y(n_577)
);

BUFx6f_ASAP7_75t_L g578 ( 
.A(n_521),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_44),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_187),
.Y(n_580)
);

BUFx3_ASAP7_75t_L g581 ( 
.A(n_217),
.Y(n_581)
);

CKINVDCx20_ASAP7_75t_R g582 ( 
.A(n_7),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_59),
.Y(n_583)
);

CKINVDCx20_ASAP7_75t_R g584 ( 
.A(n_202),
.Y(n_584)
);

BUFx10_ASAP7_75t_L g585 ( 
.A(n_506),
.Y(n_585)
);

INVx1_ASAP7_75t_SL g586 ( 
.A(n_527),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_118),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_249),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_363),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_48),
.Y(n_590)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_108),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_257),
.Y(n_592)
);

CKINVDCx20_ASAP7_75t_R g593 ( 
.A(n_376),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_86),
.Y(n_594)
);

CKINVDCx20_ASAP7_75t_R g595 ( 
.A(n_463),
.Y(n_595)
);

BUFx5_ASAP7_75t_L g596 ( 
.A(n_56),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_358),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_575),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_399),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_571),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_322),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_53),
.Y(n_602)
);

CKINVDCx20_ASAP7_75t_R g603 ( 
.A(n_38),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_475),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_293),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_333),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_139),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_327),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_75),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_547),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_205),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_334),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_255),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_562),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_410),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_206),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_211),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_398),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_253),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_551),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_265),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_566),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_248),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_148),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_520),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_280),
.Y(n_626)
);

INVxp67_ASAP7_75t_L g627 ( 
.A(n_125),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_359),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_82),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_532),
.Y(n_630)
);

CKINVDCx20_ASAP7_75t_R g631 ( 
.A(n_331),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_429),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_322),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_573),
.Y(n_634)
);

CKINVDCx20_ASAP7_75t_R g635 ( 
.A(n_310),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_344),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_394),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_305),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_427),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_8),
.Y(n_640)
);

CKINVDCx20_ASAP7_75t_R g641 ( 
.A(n_557),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_533),
.Y(n_642)
);

CKINVDCx16_ASAP7_75t_R g643 ( 
.A(n_312),
.Y(n_643)
);

INVx1_ASAP7_75t_SL g644 ( 
.A(n_574),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_290),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_77),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_221),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_231),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_508),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_176),
.Y(n_650)
);

BUFx10_ASAP7_75t_L g651 ( 
.A(n_204),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_522),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_50),
.Y(n_653)
);

CKINVDCx20_ASAP7_75t_R g654 ( 
.A(n_287),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_229),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_89),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_433),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_497),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_505),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_145),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_205),
.Y(n_661)
);

CKINVDCx20_ASAP7_75t_R g662 ( 
.A(n_199),
.Y(n_662)
);

CKINVDCx20_ASAP7_75t_R g663 ( 
.A(n_428),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_111),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_217),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_507),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_510),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_124),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_65),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_420),
.Y(n_670)
);

CKINVDCx20_ASAP7_75t_R g671 ( 
.A(n_158),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_387),
.Y(n_672)
);

INVx3_ASAP7_75t_L g673 ( 
.A(n_518),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_480),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_157),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_530),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_487),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_561),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_572),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_95),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_316),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_324),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_418),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_346),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_336),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_385),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_102),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_473),
.Y(n_688)
);

INVx1_ASAP7_75t_SL g689 ( 
.A(n_187),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_119),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_130),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_244),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_514),
.Y(n_693)
);

INVx1_ASAP7_75t_SL g694 ( 
.A(n_94),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_460),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_374),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_257),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_19),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_47),
.Y(n_699)
);

INVx1_ASAP7_75t_SL g700 ( 
.A(n_537),
.Y(n_700)
);

INVxp33_ASAP7_75t_R g701 ( 
.A(n_523),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_280),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_16),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_78),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_472),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_305),
.Y(n_706)
);

CKINVDCx16_ASAP7_75t_R g707 ( 
.A(n_165),
.Y(n_707)
);

INVx1_ASAP7_75t_SL g708 ( 
.A(n_216),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_502),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_147),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_315),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_84),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_259),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_459),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_403),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_139),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_91),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_395),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_52),
.Y(n_719)
);

INVx2_ASAP7_75t_SL g720 ( 
.A(n_206),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_199),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_509),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_434),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_220),
.Y(n_724)
);

CKINVDCx20_ASAP7_75t_R g725 ( 
.A(n_445),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_264),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_563),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_138),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_143),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_152),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_119),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_170),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_474),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_467),
.Y(n_734)
);

CKINVDCx12_ASAP7_75t_R g735 ( 
.A(n_504),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_365),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_12),
.Y(n_737)
);

CKINVDCx20_ASAP7_75t_R g738 ( 
.A(n_155),
.Y(n_738)
);

INVx1_ASAP7_75t_SL g739 ( 
.A(n_8),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_44),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_339),
.Y(n_741)
);

CKINVDCx16_ASAP7_75t_R g742 ( 
.A(n_221),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_456),
.Y(n_743)
);

CKINVDCx16_ASAP7_75t_R g744 ( 
.A(n_278),
.Y(n_744)
);

HB1xp67_ASAP7_75t_L g745 ( 
.A(n_155),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_416),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_179),
.Y(n_747)
);

INVx1_ASAP7_75t_SL g748 ( 
.A(n_421),
.Y(n_748)
);

CKINVDCx16_ASAP7_75t_R g749 ( 
.A(n_481),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_347),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_181),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_109),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_274),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_477),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_336),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_32),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_355),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_345),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_313),
.Y(n_759)
);

CKINVDCx16_ASAP7_75t_R g760 ( 
.A(n_540),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_417),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_337),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_107),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_525),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_24),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_343),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_307),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_35),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_454),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_17),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_301),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_470),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_435),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_478),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_483),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_362),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_564),
.Y(n_777)
);

INVxp67_ASAP7_75t_L g778 ( 
.A(n_270),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_378),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_260),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_26),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_531),
.Y(n_782)
);

BUFx3_ASAP7_75t_L g783 ( 
.A(n_344),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_267),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_382),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_248),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_545),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_392),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_431),
.Y(n_789)
);

BUFx10_ASAP7_75t_L g790 ( 
.A(n_330),
.Y(n_790)
);

BUFx6f_ASAP7_75t_L g791 ( 
.A(n_436),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_13),
.Y(n_792)
);

CKINVDCx20_ASAP7_75t_R g793 ( 
.A(n_182),
.Y(n_793)
);

CKINVDCx20_ASAP7_75t_R g794 ( 
.A(n_161),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_488),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_102),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_235),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_83),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_450),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_565),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_499),
.Y(n_801)
);

CKINVDCx20_ASAP7_75t_R g802 ( 
.A(n_494),
.Y(n_802)
);

INVx1_ASAP7_75t_SL g803 ( 
.A(n_283),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_311),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_4),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_173),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_47),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_282),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_73),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_401),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_489),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_457),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_300),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_142),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_295),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_289),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_560),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_64),
.Y(n_818)
);

CKINVDCx20_ASAP7_75t_R g819 ( 
.A(n_110),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_441),
.Y(n_820)
);

CKINVDCx16_ASAP7_75t_R g821 ( 
.A(n_24),
.Y(n_821)
);

BUFx6f_ASAP7_75t_L g822 ( 
.A(n_0),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_405),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_141),
.Y(n_824)
);

BUFx3_ASAP7_75t_L g825 ( 
.A(n_301),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_235),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_388),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_328),
.Y(n_828)
);

BUFx6f_ASAP7_75t_L g829 ( 
.A(n_116),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_106),
.Y(n_830)
);

BUFx3_ASAP7_75t_L g831 ( 
.A(n_135),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_259),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_193),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_449),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_285),
.Y(n_835)
);

BUFx3_ASAP7_75t_L g836 ( 
.A(n_101),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_425),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_89),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_201),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_19),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_2),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_486),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_141),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_372),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_340),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_146),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_16),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_105),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_127),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_383),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_517),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_134),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_498),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_361),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_183),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_462),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_274),
.Y(n_857)
);

INVxp67_ASAP7_75t_L g858 ( 
.A(n_27),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_348),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_229),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_115),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_461),
.Y(n_862)
);

BUFx5_ASAP7_75t_L g863 ( 
.A(n_1),
.Y(n_863)
);

INVx2_ASAP7_75t_SL g864 ( 
.A(n_237),
.Y(n_864)
);

INVx2_ASAP7_75t_SL g865 ( 
.A(n_21),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_261),
.Y(n_866)
);

BUFx5_ASAP7_75t_L g867 ( 
.A(n_233),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_111),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_287),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_207),
.Y(n_870)
);

CKINVDCx20_ASAP7_75t_R g871 ( 
.A(n_559),
.Y(n_871)
);

CKINVDCx20_ASAP7_75t_R g872 ( 
.A(n_30),
.Y(n_872)
);

BUFx6f_ASAP7_75t_L g873 ( 
.A(n_75),
.Y(n_873)
);

BUFx10_ASAP7_75t_L g874 ( 
.A(n_0),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_237),
.Y(n_875)
);

CKINVDCx20_ASAP7_75t_R g876 ( 
.A(n_538),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_80),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_476),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_179),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_151),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_175),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_264),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_511),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_379),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_328),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_275),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_72),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_269),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_4),
.Y(n_889)
);

CKINVDCx16_ASAP7_75t_R g890 ( 
.A(n_354),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_430),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_496),
.Y(n_892)
);

CKINVDCx16_ASAP7_75t_R g893 ( 
.A(n_424),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_315),
.Y(n_894)
);

BUFx3_ASAP7_75t_L g895 ( 
.A(n_440),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_299),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_15),
.Y(n_897)
);

BUFx10_ASAP7_75t_L g898 ( 
.A(n_178),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_281),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_26),
.Y(n_900)
);

CKINVDCx20_ASAP7_75t_R g901 ( 
.A(n_302),
.Y(n_901)
);

CKINVDCx20_ASAP7_75t_R g902 ( 
.A(n_128),
.Y(n_902)
);

BUFx10_ASAP7_75t_L g903 ( 
.A(n_377),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_569),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_567),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_99),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_101),
.Y(n_907)
);

BUFx3_ASAP7_75t_L g908 ( 
.A(n_240),
.Y(n_908)
);

BUFx10_ASAP7_75t_L g909 ( 
.A(n_212),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_149),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_162),
.Y(n_911)
);

CKINVDCx20_ASAP7_75t_R g912 ( 
.A(n_72),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_14),
.Y(n_913)
);

INVx1_ASAP7_75t_SL g914 ( 
.A(n_138),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_154),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_98),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_183),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_234),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_412),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_113),
.Y(n_920)
);

BUFx5_ASAP7_75t_L g921 ( 
.A(n_369),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_400),
.Y(n_922)
);

BUFx6f_ASAP7_75t_L g923 ( 
.A(n_318),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_338),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_549),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_3),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_352),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_33),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_297),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_171),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_413),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_316),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_339),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_150),
.Y(n_934)
);

CKINVDCx20_ASAP7_75t_R g935 ( 
.A(n_335),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_512),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_539),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_367),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_314),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_351),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_70),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_161),
.Y(n_942)
);

BUFx2_ASAP7_75t_L g943 ( 
.A(n_53),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_332),
.Y(n_944)
);

BUFx10_ASAP7_75t_L g945 ( 
.A(n_251),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_10),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_201),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_337),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_92),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_34),
.Y(n_950)
);

BUFx5_ASAP7_75t_L g951 ( 
.A(n_260),
.Y(n_951)
);

INVx1_ASAP7_75t_SL g952 ( 
.A(n_61),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_360),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_196),
.Y(n_954)
);

HB1xp67_ASAP7_75t_L g955 ( 
.A(n_9),
.Y(n_955)
);

HB1xp67_ASAP7_75t_L g956 ( 
.A(n_108),
.Y(n_956)
);

CKINVDCx20_ASAP7_75t_R g957 ( 
.A(n_304),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_546),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_110),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_225),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_94),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_31),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_558),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_11),
.Y(n_964)
);

BUFx5_ASAP7_75t_L g965 ( 
.A(n_366),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_271),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_529),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_127),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_33),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_182),
.Y(n_970)
);

BUFx3_ASAP7_75t_L g971 ( 
.A(n_224),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_544),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_312),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_342),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_31),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_130),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_373),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_552),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_28),
.Y(n_979)
);

BUFx6f_ASAP7_75t_L g980 ( 
.A(n_296),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_335),
.Y(n_981)
);

INVx1_ASAP7_75t_SL g982 ( 
.A(n_384),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_570),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_28),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_326),
.Y(n_985)
);

CKINVDCx20_ASAP7_75t_R g986 ( 
.A(n_169),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_389),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_135),
.Y(n_988)
);

CKINVDCx20_ASAP7_75t_R g989 ( 
.A(n_438),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_256),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_164),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_137),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_41),
.Y(n_993)
);

CKINVDCx16_ASAP7_75t_R g994 ( 
.A(n_302),
.Y(n_994)
);

INVx1_ASAP7_75t_SL g995 ( 
.A(n_295),
.Y(n_995)
);

CKINVDCx20_ASAP7_75t_R g996 ( 
.A(n_464),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_185),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_303),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_226),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_32),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_568),
.Y(n_1001)
);

BUFx10_ASAP7_75t_L g1002 ( 
.A(n_169),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_1),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_324),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_554),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_501),
.Y(n_1006)
);

INVx2_ASAP7_75t_SL g1007 ( 
.A(n_5),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_5),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_371),
.Y(n_1009)
);

INVx1_ASAP7_75t_SL g1010 ( 
.A(n_582),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_749),
.Y(n_1011)
);

INVxp33_ASAP7_75t_SL g1012 ( 
.A(n_745),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_596),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_576),
.Y(n_1014)
);

INVxp67_ASAP7_75t_SL g1015 ( 
.A(n_576),
.Y(n_1015)
);

BUFx6f_ASAP7_75t_L g1016 ( 
.A(n_578),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_760),
.Y(n_1017)
);

CKINVDCx20_ASAP7_75t_R g1018 ( 
.A(n_584),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_576),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_581),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_581),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_783),
.Y(n_1022)
);

INVxp67_ASAP7_75t_L g1023 ( 
.A(n_943),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_890),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_783),
.Y(n_1025)
);

AND2x4_ASAP7_75t_L g1026 ( 
.A(n_825),
.B(n_2),
.Y(n_1026)
);

CKINVDCx20_ASAP7_75t_R g1027 ( 
.A(n_603),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_825),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_831),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_831),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_836),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_836),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_893),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_908),
.Y(n_1034)
);

CKINVDCx16_ASAP7_75t_R g1035 ( 
.A(n_643),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_908),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_971),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_971),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_596),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_596),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_596),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_596),
.Y(n_1042)
);

INVxp67_ASAP7_75t_L g1043 ( 
.A(n_955),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_596),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_596),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_863),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_863),
.Y(n_1047)
);

INVxp67_ASAP7_75t_SL g1048 ( 
.A(n_591),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_863),
.Y(n_1049)
);

CKINVDCx20_ASAP7_75t_R g1050 ( 
.A(n_631),
.Y(n_1050)
);

BUFx6f_ASAP7_75t_L g1051 ( 
.A(n_578),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_863),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_863),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_863),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_863),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_863),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_867),
.Y(n_1057)
);

CKINVDCx16_ASAP7_75t_R g1058 ( 
.A(n_707),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_585),
.Y(n_1059)
);

BUFx3_ASAP7_75t_L g1060 ( 
.A(n_895),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_867),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_867),
.Y(n_1062)
);

NOR2xp67_ASAP7_75t_L g1063 ( 
.A(n_720),
.B(n_3),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_867),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_867),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_867),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_951),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_951),
.Y(n_1068)
);

CKINVDCx16_ASAP7_75t_R g1069 ( 
.A(n_742),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_585),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_951),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_951),
.Y(n_1072)
);

CKINVDCx20_ASAP7_75t_R g1073 ( 
.A(n_635),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_951),
.Y(n_1074)
);

INVxp67_ASAP7_75t_SL g1075 ( 
.A(n_591),
.Y(n_1075)
);

INVxp67_ASAP7_75t_SL g1076 ( 
.A(n_591),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_951),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_951),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_951),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_579),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_591),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_580),
.Y(n_1082)
);

CKINVDCx20_ASAP7_75t_R g1083 ( 
.A(n_654),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_583),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_606),
.Y(n_1085)
);

BUFx6f_ASAP7_75t_L g1086 ( 
.A(n_578),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_608),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_609),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_585),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_613),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_617),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_903),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_619),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_591),
.Y(n_1094)
);

CKINVDCx20_ASAP7_75t_R g1095 ( 
.A(n_662),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_621),
.Y(n_1096)
);

CKINVDCx16_ASAP7_75t_R g1097 ( 
.A(n_744),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_903),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_624),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_633),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_638),
.Y(n_1101)
);

BUFx2_ASAP7_75t_L g1102 ( 
.A(n_956),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_645),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_665),
.Y(n_1104)
);

INVxp33_ASAP7_75t_SL g1105 ( 
.A(n_587),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_675),
.Y(n_1106)
);

INVxp33_ASAP7_75t_L g1107 ( 
.A(n_590),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_903),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_577),
.Y(n_1109)
);

INVxp67_ASAP7_75t_SL g1110 ( 
.A(n_822),
.Y(n_1110)
);

CKINVDCx20_ASAP7_75t_R g1111 ( 
.A(n_671),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_822),
.Y(n_1112)
);

BUFx6f_ASAP7_75t_L g1113 ( 
.A(n_578),
.Y(n_1113)
);

INVxp33_ASAP7_75t_SL g1114 ( 
.A(n_587),
.Y(n_1114)
);

BUFx6f_ASAP7_75t_L g1115 ( 
.A(n_578),
.Y(n_1115)
);

INVxp67_ASAP7_75t_SL g1116 ( 
.A(n_822),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_822),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_691),
.Y(n_1118)
);

INVx1_ASAP7_75t_SL g1119 ( 
.A(n_738),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_697),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_698),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_822),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_728),
.Y(n_1123)
);

CKINVDCx20_ASAP7_75t_R g1124 ( 
.A(n_793),
.Y(n_1124)
);

INVxp67_ASAP7_75t_L g1125 ( 
.A(n_720),
.Y(n_1125)
);

CKINVDCx16_ASAP7_75t_R g1126 ( 
.A(n_821),
.Y(n_1126)
);

BUFx6f_ASAP7_75t_L g1127 ( 
.A(n_791),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_577),
.Y(n_1128)
);

INVxp33_ASAP7_75t_L g1129 ( 
.A(n_590),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_732),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_741),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_751),
.Y(n_1132)
);

CKINVDCx16_ASAP7_75t_R g1133 ( 
.A(n_994),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_755),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_759),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_829),
.Y(n_1136)
);

CKINVDCx20_ASAP7_75t_R g1137 ( 
.A(n_794),
.Y(n_1137)
);

BUFx2_ASAP7_75t_L g1138 ( 
.A(n_588),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_762),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_768),
.Y(n_1140)
);

INVx2_ASAP7_75t_L g1141 ( 
.A(n_829),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_589),
.Y(n_1142)
);

BUFx3_ASAP7_75t_L g1143 ( 
.A(n_895),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_780),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_589),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_786),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_798),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_804),
.Y(n_1148)
);

BUFx6f_ASAP7_75t_L g1149 ( 
.A(n_791),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_599),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_806),
.Y(n_1151)
);

CKINVDCx14_ASAP7_75t_R g1152 ( 
.A(n_593),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_807),
.Y(n_1153)
);

CKINVDCx20_ASAP7_75t_R g1154 ( 
.A(n_819),
.Y(n_1154)
);

CKINVDCx20_ASAP7_75t_R g1155 ( 
.A(n_872),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_814),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_815),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_828),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_841),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_599),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_845),
.Y(n_1161)
);

INVx1_ASAP7_75t_SL g1162 ( 
.A(n_901),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_846),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_604),
.Y(n_1164)
);

CKINVDCx16_ASAP7_75t_R g1165 ( 
.A(n_651),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_849),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_829),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_852),
.Y(n_1168)
);

INVxp67_ASAP7_75t_SL g1169 ( 
.A(n_829),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_855),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_877),
.Y(n_1171)
);

INVxp67_ASAP7_75t_SL g1172 ( 
.A(n_829),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_887),
.Y(n_1173)
);

INVx2_ASAP7_75t_SL g1174 ( 
.A(n_651),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_897),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_907),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_604),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_911),
.Y(n_1178)
);

BUFx2_ASAP7_75t_L g1179 ( 
.A(n_588),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_915),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_926),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_928),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_610),
.Y(n_1183)
);

INVxp67_ASAP7_75t_SL g1184 ( 
.A(n_873),
.Y(n_1184)
);

INVxp67_ASAP7_75t_SL g1185 ( 
.A(n_873),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_929),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_932),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_610),
.Y(n_1188)
);

CKINVDCx20_ASAP7_75t_R g1189 ( 
.A(n_902),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_934),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_950),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_962),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_974),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_873),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_985),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_873),
.Y(n_1196)
);

INVxp67_ASAP7_75t_L g1197 ( 
.A(n_864),
.Y(n_1197)
);

INVxp67_ASAP7_75t_SL g1198 ( 
.A(n_873),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_993),
.Y(n_1199)
);

CKINVDCx16_ASAP7_75t_R g1200 ( 
.A(n_651),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_997),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_660),
.Y(n_1202)
);

BUFx2_ASAP7_75t_L g1203 ( 
.A(n_592),
.Y(n_1203)
);

CKINVDCx20_ASAP7_75t_R g1204 ( 
.A(n_912),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_614),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_614),
.Y(n_1206)
);

BUFx10_ASAP7_75t_L g1207 ( 
.A(n_923),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_660),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_668),
.Y(n_1209)
);

CKINVDCx16_ASAP7_75t_R g1210 ( 
.A(n_790),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_668),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_684),
.Y(n_1212)
);

NOR2xp67_ASAP7_75t_L g1213 ( 
.A(n_864),
.B(n_6),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_923),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_684),
.Y(n_1215)
);

BUFx3_ASAP7_75t_L g1216 ( 
.A(n_597),
.Y(n_1216)
);

CKINVDCx16_ASAP7_75t_R g1217 ( 
.A(n_790),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_618),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_685),
.Y(n_1219)
);

CKINVDCx16_ASAP7_75t_R g1220 ( 
.A(n_790),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_685),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_721),
.Y(n_1222)
);

CKINVDCx20_ASAP7_75t_R g1223 ( 
.A(n_935),
.Y(n_1223)
);

INVxp67_ASAP7_75t_SL g1224 ( 
.A(n_923),
.Y(n_1224)
);

INVx2_ASAP7_75t_L g1225 ( 
.A(n_923),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_721),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_726),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_726),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_731),
.Y(n_1229)
);

BUFx3_ASAP7_75t_L g1230 ( 
.A(n_598),
.Y(n_1230)
);

INVx1_ASAP7_75t_SL g1231 ( 
.A(n_957),
.Y(n_1231)
);

INVx2_ASAP7_75t_L g1232 ( 
.A(n_923),
.Y(n_1232)
);

INVxp33_ASAP7_75t_SL g1233 ( 
.A(n_592),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_731),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_618),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_770),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_770),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_816),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_980),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_620),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_816),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_980),
.Y(n_1242)
);

INVxp33_ASAP7_75t_L g1243 ( 
.A(n_818),
.Y(n_1243)
);

INVxp67_ASAP7_75t_SL g1244 ( 
.A(n_980),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_818),
.Y(n_1245)
);

CKINVDCx20_ASAP7_75t_R g1246 ( 
.A(n_986),
.Y(n_1246)
);

CKINVDCx20_ASAP7_75t_R g1247 ( 
.A(n_874),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_839),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_839),
.Y(n_1249)
);

HB1xp67_ASAP7_75t_L g1250 ( 
.A(n_594),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_843),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_980),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_843),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_848),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_980),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_848),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_941),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_941),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_865),
.Y(n_1259)
);

INVx2_ASAP7_75t_SL g1260 ( 
.A(n_874),
.Y(n_1260)
);

BUFx2_ASAP7_75t_L g1261 ( 
.A(n_594),
.Y(n_1261)
);

CKINVDCx14_ASAP7_75t_R g1262 ( 
.A(n_595),
.Y(n_1262)
);

INVxp67_ASAP7_75t_SL g1263 ( 
.A(n_865),
.Y(n_1263)
);

INVxp33_ASAP7_75t_SL g1264 ( 
.A(n_601),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1007),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1007),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_620),
.Y(n_1267)
);

INVxp33_ASAP7_75t_L g1268 ( 
.A(n_600),
.Y(n_1268)
);

INVx2_ASAP7_75t_L g1269 ( 
.A(n_615),
.Y(n_1269)
);

INVx1_ASAP7_75t_SL g1270 ( 
.A(n_689),
.Y(n_1270)
);

INVx1_ASAP7_75t_SL g1271 ( 
.A(n_694),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_622),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_874),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_898),
.Y(n_1274)
);

CKINVDCx5p33_ASAP7_75t_R g1275 ( 
.A(n_622),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_898),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_625),
.Y(n_1277)
);

CKINVDCx14_ASAP7_75t_R g1278 ( 
.A(n_641),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_898),
.Y(n_1279)
);

CKINVDCx20_ASAP7_75t_R g1280 ( 
.A(n_909),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_625),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_909),
.Y(n_1282)
);

INVxp33_ASAP7_75t_L g1283 ( 
.A(n_600),
.Y(n_1283)
);

INVxp67_ASAP7_75t_L g1284 ( 
.A(n_909),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_945),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_628),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_945),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_945),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1002),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_639),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1002),
.Y(n_1291)
);

INVxp67_ASAP7_75t_SL g1292 ( 
.A(n_627),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1002),
.Y(n_1293)
);

INVxp33_ASAP7_75t_L g1294 ( 
.A(n_667),
.Y(n_1294)
);

NOR2xp33_ASAP7_75t_L g1295 ( 
.A(n_673),
.B(n_6),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_649),
.Y(n_1296)
);

CKINVDCx20_ASAP7_75t_R g1297 ( 
.A(n_663),
.Y(n_1297)
);

BUFx3_ASAP7_75t_L g1298 ( 
.A(n_666),
.Y(n_1298)
);

INVxp33_ASAP7_75t_L g1299 ( 
.A(n_667),
.Y(n_1299)
);

NOR2xp33_ASAP7_75t_L g1300 ( 
.A(n_673),
.B(n_7),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_677),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_688),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_693),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_695),
.Y(n_1304)
);

INVxp67_ASAP7_75t_L g1305 ( 
.A(n_601),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_714),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_733),
.Y(n_1307)
);

CKINVDCx5p33_ASAP7_75t_R g1308 ( 
.A(n_628),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_736),
.Y(n_1309)
);

HB1xp67_ASAP7_75t_L g1310 ( 
.A(n_602),
.Y(n_1310)
);

BUFx6f_ASAP7_75t_L g1311 ( 
.A(n_791),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_746),
.Y(n_1312)
);

INVx2_ASAP7_75t_L g1313 ( 
.A(n_757),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_769),
.Y(n_1314)
);

CKINVDCx20_ASAP7_75t_R g1315 ( 
.A(n_725),
.Y(n_1315)
);

INVx1_ASAP7_75t_SL g1316 ( 
.A(n_708),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_776),
.Y(n_1317)
);

INVxp33_ASAP7_75t_SL g1318 ( 
.A(n_602),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_779),
.Y(n_1319)
);

INVxp67_ASAP7_75t_L g1320 ( 
.A(n_605),
.Y(n_1320)
);

CKINVDCx5p33_ASAP7_75t_R g1321 ( 
.A(n_630),
.Y(n_1321)
);

CKINVDCx5p33_ASAP7_75t_R g1322 ( 
.A(n_630),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_789),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_801),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_632),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_820),
.Y(n_1326)
);

BUFx3_ASAP7_75t_L g1327 ( 
.A(n_827),
.Y(n_1327)
);

BUFx6f_ASAP7_75t_L g1328 ( 
.A(n_791),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_632),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_834),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_844),
.Y(n_1331)
);

INVxp33_ASAP7_75t_SL g1332 ( 
.A(n_605),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_850),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_851),
.Y(n_1334)
);

BUFx2_ASAP7_75t_L g1335 ( 
.A(n_607),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_856),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_883),
.Y(n_1337)
);

CKINVDCx20_ASAP7_75t_R g1338 ( 
.A(n_802),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_891),
.Y(n_1339)
);

INVxp67_ASAP7_75t_L g1340 ( 
.A(n_607),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_936),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_937),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_953),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_963),
.Y(n_1344)
);

INVxp33_ASAP7_75t_L g1345 ( 
.A(n_686),
.Y(n_1345)
);

CKINVDCx5p33_ASAP7_75t_R g1346 ( 
.A(n_634),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_978),
.Y(n_1347)
);

BUFx10_ASAP7_75t_L g1348 ( 
.A(n_634),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1006),
.Y(n_1349)
);

CKINVDCx16_ASAP7_75t_R g1350 ( 
.A(n_871),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1009),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_686),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_735),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_778),
.Y(n_1354)
);

INVxp67_ASAP7_75t_SL g1355 ( 
.A(n_858),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_727),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_611),
.Y(n_1357)
);

INVxp33_ASAP7_75t_L g1358 ( 
.A(n_727),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_837),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_611),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_612),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_837),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_612),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_616),
.Y(n_1364)
);

INVx2_ASAP7_75t_SL g1365 ( 
.A(n_616),
.Y(n_1365)
);

INVx2_ASAP7_75t_SL g1366 ( 
.A(n_623),
.Y(n_1366)
);

CKINVDCx5p33_ASAP7_75t_R g1367 ( 
.A(n_637),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_623),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_626),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_626),
.Y(n_1370)
);

CKINVDCx16_ASAP7_75t_R g1371 ( 
.A(n_876),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_919),
.Y(n_1372)
);

INVxp33_ASAP7_75t_L g1373 ( 
.A(n_919),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_629),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_629),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_636),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_636),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_640),
.Y(n_1378)
);

INVxp67_ASAP7_75t_SL g1379 ( 
.A(n_673),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_640),
.Y(n_1380)
);

INVxp67_ASAP7_75t_L g1381 ( 
.A(n_646),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_646),
.Y(n_1382)
);

CKINVDCx5p33_ASAP7_75t_R g1383 ( 
.A(n_637),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_647),
.Y(n_1384)
);

OR2x2_ASAP7_75t_L g1385 ( 
.A(n_739),
.B(n_9),
.Y(n_1385)
);

CKINVDCx20_ASAP7_75t_R g1386 ( 
.A(n_989),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_647),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_648),
.Y(n_1388)
);

CKINVDCx16_ASAP7_75t_R g1389 ( 
.A(n_996),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_648),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_650),
.Y(n_1391)
);

CKINVDCx14_ASAP7_75t_R g1392 ( 
.A(n_642),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_650),
.Y(n_1393)
);

INVxp67_ASAP7_75t_SL g1394 ( 
.A(n_977),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_977),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1379),
.B(n_586),
.Y(n_1396)
);

NOR2xp33_ASAP7_75t_L g1397 ( 
.A(n_1392),
.B(n_644),
.Y(n_1397)
);

AND2x4_ASAP7_75t_L g1398 ( 
.A(n_1060),
.B(n_700),
.Y(n_1398)
);

INVx2_ASAP7_75t_SL g1399 ( 
.A(n_1348),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1081),
.Y(n_1400)
);

INVx5_ASAP7_75t_L g1401 ( 
.A(n_1016),
.Y(n_1401)
);

BUFx8_ASAP7_75t_SL g1402 ( 
.A(n_1018),
.Y(n_1402)
);

NOR2xp33_ASAP7_75t_SL g1403 ( 
.A(n_1270),
.B(n_701),
.Y(n_1403)
);

BUFx3_ASAP7_75t_L g1404 ( 
.A(n_1207),
.Y(n_1404)
);

INVx3_ASAP7_75t_L g1405 ( 
.A(n_1207),
.Y(n_1405)
);

INVx5_ASAP7_75t_L g1406 ( 
.A(n_1016),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1107),
.B(n_653),
.Y(n_1407)
);

INVx5_ASAP7_75t_L g1408 ( 
.A(n_1016),
.Y(n_1408)
);

BUFx12f_ASAP7_75t_L g1409 ( 
.A(n_1348),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1107),
.B(n_1129),
.Y(n_1410)
);

BUFx6f_ASAP7_75t_L g1411 ( 
.A(n_1051),
.Y(n_1411)
);

BUFx6f_ASAP7_75t_L g1412 ( 
.A(n_1051),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1081),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1094),
.Y(n_1414)
);

AND2x4_ASAP7_75t_L g1415 ( 
.A(n_1060),
.B(n_748),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1048),
.Y(n_1416)
);

BUFx12f_ASAP7_75t_L g1417 ( 
.A(n_1348),
.Y(n_1417)
);

BUFx6f_ASAP7_75t_L g1418 ( 
.A(n_1051),
.Y(n_1418)
);

AND2x4_ASAP7_75t_L g1419 ( 
.A(n_1143),
.B(n_982),
.Y(n_1419)
);

INVx2_ASAP7_75t_L g1420 ( 
.A(n_1094),
.Y(n_1420)
);

AND2x4_ASAP7_75t_L g1421 ( 
.A(n_1143),
.B(n_803),
.Y(n_1421)
);

HB1xp67_ASAP7_75t_L g1422 ( 
.A(n_1271),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1015),
.B(n_670),
.Y(n_1423)
);

NOR2xp33_ASAP7_75t_L g1424 ( 
.A(n_1392),
.B(n_642),
.Y(n_1424)
);

BUFx6f_ASAP7_75t_L g1425 ( 
.A(n_1051),
.Y(n_1425)
);

AND2x4_ASAP7_75t_L g1426 ( 
.A(n_1026),
.B(n_914),
.Y(n_1426)
);

CKINVDCx5p33_ASAP7_75t_R g1427 ( 
.A(n_1152),
.Y(n_1427)
);

BUFx3_ASAP7_75t_L g1428 ( 
.A(n_1207),
.Y(n_1428)
);

INVxp67_ASAP7_75t_L g1429 ( 
.A(n_1316),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1268),
.B(n_672),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1112),
.Y(n_1431)
);

BUFx6f_ASAP7_75t_L g1432 ( 
.A(n_1113),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1112),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1075),
.Y(n_1434)
);

INVx5_ASAP7_75t_L g1435 ( 
.A(n_1016),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1268),
.B(n_674),
.Y(n_1436)
);

HB1xp67_ASAP7_75t_L g1437 ( 
.A(n_1035),
.Y(n_1437)
);

BUFx12f_ASAP7_75t_L g1438 ( 
.A(n_1011),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1129),
.B(n_1243),
.Y(n_1439)
);

HB1xp67_ASAP7_75t_L g1440 ( 
.A(n_1058),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1283),
.B(n_1294),
.Y(n_1441)
);

NOR2xp33_ASAP7_75t_L g1442 ( 
.A(n_1353),
.B(n_652),
.Y(n_1442)
);

AND2x4_ASAP7_75t_L g1443 ( 
.A(n_1026),
.B(n_1263),
.Y(n_1443)
);

INVx3_ASAP7_75t_L g1444 ( 
.A(n_1352),
.Y(n_1444)
);

BUFx12f_ASAP7_75t_L g1445 ( 
.A(n_1011),
.Y(n_1445)
);

NOR2x1_ASAP7_75t_L g1446 ( 
.A(n_1216),
.B(n_791),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1283),
.B(n_1294),
.Y(n_1447)
);

INVx3_ASAP7_75t_L g1448 ( 
.A(n_1352),
.Y(n_1448)
);

BUFx3_ASAP7_75t_L g1449 ( 
.A(n_1039),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1076),
.Y(n_1450)
);

BUFx12f_ASAP7_75t_L g1451 ( 
.A(n_1017),
.Y(n_1451)
);

BUFx8_ASAP7_75t_L g1452 ( 
.A(n_1138),
.Y(n_1452)
);

BUFx12f_ASAP7_75t_L g1453 ( 
.A(n_1017),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1299),
.B(n_676),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1299),
.B(n_678),
.Y(n_1455)
);

AND2x4_ASAP7_75t_L g1456 ( 
.A(n_1026),
.B(n_952),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1243),
.B(n_653),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1110),
.Y(n_1458)
);

INVx6_ASAP7_75t_L g1459 ( 
.A(n_1216),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1345),
.B(n_679),
.Y(n_1460)
);

INVxp67_ASAP7_75t_L g1461 ( 
.A(n_1179),
.Y(n_1461)
);

NOR2xp33_ASAP7_75t_SL g1462 ( 
.A(n_1024),
.B(n_995),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1117),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_SL g1464 ( 
.A(n_1059),
.B(n_652),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1345),
.B(n_655),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1358),
.B(n_683),
.Y(n_1466)
);

AND2x4_ASAP7_75t_L g1467 ( 
.A(n_1230),
.B(n_1298),
.Y(n_1467)
);

INVx5_ASAP7_75t_L g1468 ( 
.A(n_1086),
.Y(n_1468)
);

BUFx8_ASAP7_75t_SL g1469 ( 
.A(n_1018),
.Y(n_1469)
);

NOR2xp33_ASAP7_75t_L g1470 ( 
.A(n_1109),
.B(n_657),
.Y(n_1470)
);

NOR2xp33_ASAP7_75t_L g1471 ( 
.A(n_1109),
.B(n_657),
.Y(n_1471)
);

BUFx6f_ASAP7_75t_L g1472 ( 
.A(n_1113),
.Y(n_1472)
);

BUFx12f_ASAP7_75t_L g1473 ( 
.A(n_1024),
.Y(n_1473)
);

INVx3_ASAP7_75t_L g1474 ( 
.A(n_1356),
.Y(n_1474)
);

BUFx12f_ASAP7_75t_L g1475 ( 
.A(n_1033),
.Y(n_1475)
);

BUFx3_ASAP7_75t_L g1476 ( 
.A(n_1040),
.Y(n_1476)
);

BUFx6f_ASAP7_75t_L g1477 ( 
.A(n_1113),
.Y(n_1477)
);

HB1xp67_ASAP7_75t_L g1478 ( 
.A(n_1069),
.Y(n_1478)
);

HB1xp67_ASAP7_75t_L g1479 ( 
.A(n_1097),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1116),
.Y(n_1480)
);

BUFx8_ASAP7_75t_L g1481 ( 
.A(n_1203),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1358),
.B(n_696),
.Y(n_1482)
);

HB1xp67_ASAP7_75t_L g1483 ( 
.A(n_1126),
.Y(n_1483)
);

INVx5_ASAP7_75t_L g1484 ( 
.A(n_1086),
.Y(n_1484)
);

BUFx6f_ASAP7_75t_L g1485 ( 
.A(n_1113),
.Y(n_1485)
);

BUFx12f_ASAP7_75t_L g1486 ( 
.A(n_1033),
.Y(n_1486)
);

BUFx6f_ASAP7_75t_L g1487 ( 
.A(n_1115),
.Y(n_1487)
);

AND2x4_ASAP7_75t_L g1488 ( 
.A(n_1230),
.B(n_658),
.Y(n_1488)
);

CKINVDCx6p67_ASAP7_75t_R g1489 ( 
.A(n_1133),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1373),
.B(n_655),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1117),
.Y(n_1491)
);

INVx5_ASAP7_75t_L g1492 ( 
.A(n_1086),
.Y(n_1492)
);

NOR2xp33_ASAP7_75t_L g1493 ( 
.A(n_1128),
.B(n_658),
.Y(n_1493)
);

INVx5_ASAP7_75t_L g1494 ( 
.A(n_1086),
.Y(n_1494)
);

NOR2xp33_ASAP7_75t_L g1495 ( 
.A(n_1128),
.B(n_659),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1373),
.B(n_1394),
.Y(n_1496)
);

BUFx12f_ASAP7_75t_L g1497 ( 
.A(n_1059),
.Y(n_1497)
);

AND2x4_ASAP7_75t_L g1498 ( 
.A(n_1298),
.B(n_659),
.Y(n_1498)
);

BUFx6f_ASAP7_75t_L g1499 ( 
.A(n_1115),
.Y(n_1499)
);

INVx5_ASAP7_75t_L g1500 ( 
.A(n_1127),
.Y(n_1500)
);

AND2x4_ASAP7_75t_L g1501 ( 
.A(n_1327),
.B(n_754),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1169),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_1122),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1172),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1020),
.B(n_656),
.Y(n_1505)
);

INVx3_ASAP7_75t_L g1506 ( 
.A(n_1356),
.Y(n_1506)
);

BUFx6f_ASAP7_75t_L g1507 ( 
.A(n_1115),
.Y(n_1507)
);

INVxp33_ASAP7_75t_SL g1508 ( 
.A(n_1142),
.Y(n_1508)
);

AND2x4_ASAP7_75t_L g1509 ( 
.A(n_1327),
.B(n_1273),
.Y(n_1509)
);

HB1xp67_ASAP7_75t_L g1510 ( 
.A(n_1010),
.Y(n_1510)
);

INVx2_ASAP7_75t_SL g1511 ( 
.A(n_1142),
.Y(n_1511)
);

BUFx3_ASAP7_75t_L g1512 ( 
.A(n_1041),
.Y(n_1512)
);

BUFx6f_ASAP7_75t_L g1513 ( 
.A(n_1115),
.Y(n_1513)
);

BUFx6f_ASAP7_75t_L g1514 ( 
.A(n_1127),
.Y(n_1514)
);

INVx3_ASAP7_75t_L g1515 ( 
.A(n_1359),
.Y(n_1515)
);

BUFx8_ASAP7_75t_L g1516 ( 
.A(n_1261),
.Y(n_1516)
);

BUFx3_ASAP7_75t_L g1517 ( 
.A(n_1042),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1357),
.B(n_705),
.Y(n_1518)
);

INVx5_ASAP7_75t_L g1519 ( 
.A(n_1127),
.Y(n_1519)
);

BUFx6f_ASAP7_75t_L g1520 ( 
.A(n_1127),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1122),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1292),
.B(n_656),
.Y(n_1522)
);

NOR2xp33_ASAP7_75t_L g1523 ( 
.A(n_1145),
.B(n_754),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_SL g1524 ( 
.A(n_1070),
.B(n_884),
.Y(n_1524)
);

BUFx6f_ASAP7_75t_L g1525 ( 
.A(n_1127),
.Y(n_1525)
);

INVx1_ASAP7_75t_SL g1526 ( 
.A(n_1119),
.Y(n_1526)
);

NOR2xp33_ASAP7_75t_L g1527 ( 
.A(n_1145),
.B(n_884),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1360),
.B(n_709),
.Y(n_1528)
);

NOR2xp33_ASAP7_75t_L g1529 ( 
.A(n_1150),
.B(n_892),
.Y(n_1529)
);

HB1xp67_ASAP7_75t_L g1530 ( 
.A(n_1162),
.Y(n_1530)
);

BUFx8_ASAP7_75t_SL g1531 ( 
.A(n_1027),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1361),
.B(n_1363),
.Y(n_1532)
);

BUFx2_ASAP7_75t_L g1533 ( 
.A(n_1150),
.Y(n_1533)
);

HB1xp67_ASAP7_75t_L g1534 ( 
.A(n_1231),
.Y(n_1534)
);

INVx3_ASAP7_75t_L g1535 ( 
.A(n_1359),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1364),
.B(n_715),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1368),
.B(n_718),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1369),
.B(n_722),
.Y(n_1538)
);

INVxp33_ASAP7_75t_SL g1539 ( 
.A(n_1160),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1184),
.Y(n_1540)
);

NOR2xp33_ASAP7_75t_L g1541 ( 
.A(n_1160),
.B(n_892),
.Y(n_1541)
);

BUFx6f_ASAP7_75t_L g1542 ( 
.A(n_1149),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1136),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1185),
.Y(n_1544)
);

AND2x4_ASAP7_75t_SL g1545 ( 
.A(n_1247),
.B(n_1280),
.Y(n_1545)
);

NOR2xp33_ASAP7_75t_L g1546 ( 
.A(n_1164),
.B(n_904),
.Y(n_1546)
);

INVxp67_ASAP7_75t_L g1547 ( 
.A(n_1335),
.Y(n_1547)
);

BUFx3_ASAP7_75t_L g1548 ( 
.A(n_1044),
.Y(n_1548)
);

HB1xp67_ASAP7_75t_L g1549 ( 
.A(n_1305),
.Y(n_1549)
);

BUFx6f_ASAP7_75t_L g1550 ( 
.A(n_1149),
.Y(n_1550)
);

BUFx6f_ASAP7_75t_L g1551 ( 
.A(n_1149),
.Y(n_1551)
);

CKINVDCx5p33_ASAP7_75t_R g1552 ( 
.A(n_1152),
.Y(n_1552)
);

AND2x6_ASAP7_75t_L g1553 ( 
.A(n_1295),
.B(n_921),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1198),
.Y(n_1554)
);

BUFx12f_ASAP7_75t_L g1555 ( 
.A(n_1070),
.Y(n_1555)
);

AND2x4_ASAP7_75t_L g1556 ( 
.A(n_1274),
.B(n_904),
.Y(n_1556)
);

NOR2xp33_ASAP7_75t_L g1557 ( 
.A(n_1164),
.B(n_905),
.Y(n_1557)
);

INVx5_ASAP7_75t_L g1558 ( 
.A(n_1149),
.Y(n_1558)
);

INVx5_ASAP7_75t_L g1559 ( 
.A(n_1149),
.Y(n_1559)
);

INVx3_ASAP7_75t_L g1560 ( 
.A(n_1362),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1021),
.B(n_880),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1370),
.B(n_723),
.Y(n_1562)
);

BUFx3_ASAP7_75t_L g1563 ( 
.A(n_1045),
.Y(n_1563)
);

BUFx12f_ASAP7_75t_L g1564 ( 
.A(n_1089),
.Y(n_1564)
);

INVx2_ASAP7_75t_SL g1565 ( 
.A(n_1177),
.Y(n_1565)
);

BUFx6f_ASAP7_75t_L g1566 ( 
.A(n_1311),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1224),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1136),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1244),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_SL g1570 ( 
.A(n_1089),
.B(n_905),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1374),
.B(n_734),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1022),
.B(n_880),
.Y(n_1572)
);

BUFx6f_ASAP7_75t_L g1573 ( 
.A(n_1311),
.Y(n_1573)
);

BUFx6f_ASAP7_75t_L g1574 ( 
.A(n_1311),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1014),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1025),
.B(n_1028),
.Y(n_1576)
);

NOR2xp33_ASAP7_75t_SL g1577 ( 
.A(n_1165),
.B(n_922),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1141),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1029),
.B(n_881),
.Y(n_1579)
);

BUFx8_ASAP7_75t_SL g1580 ( 
.A(n_1027),
.Y(n_1580)
);

BUFx6f_ASAP7_75t_L g1581 ( 
.A(n_1311),
.Y(n_1581)
);

BUFx2_ASAP7_75t_L g1582 ( 
.A(n_1177),
.Y(n_1582)
);

HB1xp67_ASAP7_75t_L g1583 ( 
.A(n_1320),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1030),
.B(n_881),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1031),
.B(n_1032),
.Y(n_1585)
);

BUFx6f_ASAP7_75t_L g1586 ( 
.A(n_1311),
.Y(n_1586)
);

NOR2xp33_ASAP7_75t_L g1587 ( 
.A(n_1183),
.B(n_922),
.Y(n_1587)
);

BUFx12f_ASAP7_75t_L g1588 ( 
.A(n_1092),
.Y(n_1588)
);

BUFx6f_ASAP7_75t_L g1589 ( 
.A(n_1328),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1375),
.B(n_743),
.Y(n_1590)
);

BUFx8_ASAP7_75t_SL g1591 ( 
.A(n_1050),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1034),
.B(n_882),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1036),
.B(n_882),
.Y(n_1593)
);

BUFx8_ASAP7_75t_SL g1594 ( 
.A(n_1050),
.Y(n_1594)
);

BUFx12f_ASAP7_75t_L g1595 ( 
.A(n_1092),
.Y(n_1595)
);

INVx5_ASAP7_75t_L g1596 ( 
.A(n_1328),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1037),
.B(n_885),
.Y(n_1597)
);

NOR2xp33_ASAP7_75t_L g1598 ( 
.A(n_1183),
.B(n_925),
.Y(n_1598)
);

CKINVDCx5p33_ASAP7_75t_R g1599 ( 
.A(n_1262),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1141),
.Y(n_1600)
);

BUFx6f_ASAP7_75t_L g1601 ( 
.A(n_1328),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1376),
.B(n_761),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1019),
.Y(n_1603)
);

INVx3_ASAP7_75t_L g1604 ( 
.A(n_1362),
.Y(n_1604)
);

BUFx3_ASAP7_75t_L g1605 ( 
.A(n_1046),
.Y(n_1605)
);

INVx5_ASAP7_75t_L g1606 ( 
.A(n_1328),
.Y(n_1606)
);

INVx5_ASAP7_75t_L g1607 ( 
.A(n_1328),
.Y(n_1607)
);

BUFx3_ASAP7_75t_L g1608 ( 
.A(n_1047),
.Y(n_1608)
);

BUFx12f_ASAP7_75t_L g1609 ( 
.A(n_1098),
.Y(n_1609)
);

BUFx12f_ASAP7_75t_L g1610 ( 
.A(n_1098),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1080),
.Y(n_1611)
);

INVx5_ASAP7_75t_L g1612 ( 
.A(n_1013),
.Y(n_1612)
);

BUFx8_ASAP7_75t_L g1613 ( 
.A(n_1102),
.Y(n_1613)
);

BUFx8_ASAP7_75t_SL g1614 ( 
.A(n_1073),
.Y(n_1614)
);

NOR2x1_ASAP7_75t_L g1615 ( 
.A(n_1296),
.B(n_764),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1377),
.B(n_772),
.Y(n_1616)
);

BUFx6f_ASAP7_75t_L g1617 ( 
.A(n_1167),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_SL g1618 ( 
.A(n_1108),
.B(n_1188),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1167),
.Y(n_1619)
);

BUFx12f_ASAP7_75t_L g1620 ( 
.A(n_1108),
.Y(n_1620)
);

INVx3_ASAP7_75t_L g1621 ( 
.A(n_1372),
.Y(n_1621)
);

INVx3_ASAP7_75t_L g1622 ( 
.A(n_1372),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1378),
.B(n_773),
.Y(n_1623)
);

BUFx2_ASAP7_75t_L g1624 ( 
.A(n_1188),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1082),
.Y(n_1625)
);

AND2x4_ASAP7_75t_L g1626 ( 
.A(n_1276),
.B(n_925),
.Y(n_1626)
);

BUFx2_ASAP7_75t_L g1627 ( 
.A(n_1205),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1380),
.B(n_774),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1084),
.Y(n_1629)
);

BUFx6f_ASAP7_75t_L g1630 ( 
.A(n_1194),
.Y(n_1630)
);

HB1xp67_ASAP7_75t_L g1631 ( 
.A(n_1340),
.Y(n_1631)
);

INVxp67_ASAP7_75t_L g1632 ( 
.A(n_1250),
.Y(n_1632)
);

CKINVDCx11_ASAP7_75t_R g1633 ( 
.A(n_1073),
.Y(n_1633)
);

BUFx6f_ASAP7_75t_L g1634 ( 
.A(n_1194),
.Y(n_1634)
);

NOR2xp33_ASAP7_75t_L g1635 ( 
.A(n_1205),
.B(n_927),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1085),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1382),
.B(n_775),
.Y(n_1637)
);

CKINVDCx16_ASAP7_75t_R g1638 ( 
.A(n_1200),
.Y(n_1638)
);

BUFx3_ASAP7_75t_L g1639 ( 
.A(n_1049),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1038),
.B(n_885),
.Y(n_1640)
);

BUFx12f_ASAP7_75t_L g1641 ( 
.A(n_1206),
.Y(n_1641)
);

BUFx6f_ASAP7_75t_L g1642 ( 
.A(n_1196),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1087),
.Y(n_1643)
);

NOR2xp33_ASAP7_75t_L g1644 ( 
.A(n_1206),
.B(n_927),
.Y(n_1644)
);

BUFx6f_ASAP7_75t_L g1645 ( 
.A(n_1196),
.Y(n_1645)
);

BUFx6f_ASAP7_75t_L g1646 ( 
.A(n_1214),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1125),
.B(n_886),
.Y(n_1647)
);

INVx2_ASAP7_75t_L g1648 ( 
.A(n_1214),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_SL g1649 ( 
.A(n_1218),
.B(n_931),
.Y(n_1649)
);

HB1xp67_ASAP7_75t_L g1650 ( 
.A(n_1381),
.Y(n_1650)
);

BUFx8_ASAP7_75t_SL g1651 ( 
.A(n_1083),
.Y(n_1651)
);

AND2x4_ASAP7_75t_L g1652 ( 
.A(n_1279),
.B(n_931),
.Y(n_1652)
);

INVx2_ASAP7_75t_SL g1653 ( 
.A(n_1218),
.Y(n_1653)
);

AND2x4_ASAP7_75t_L g1654 ( 
.A(n_1282),
.B(n_938),
.Y(n_1654)
);

INVx3_ASAP7_75t_L g1655 ( 
.A(n_1395),
.Y(n_1655)
);

BUFx12f_ASAP7_75t_L g1656 ( 
.A(n_1235),
.Y(n_1656)
);

AND2x4_ASAP7_75t_L g1657 ( 
.A(n_1285),
.B(n_938),
.Y(n_1657)
);

BUFx8_ASAP7_75t_SL g1658 ( 
.A(n_1083),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1197),
.B(n_886),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1088),
.Y(n_1660)
);

NOR2xp33_ASAP7_75t_L g1661 ( 
.A(n_1235),
.B(n_1001),
.Y(n_1661)
);

BUFx12f_ASAP7_75t_L g1662 ( 
.A(n_1240),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1384),
.B(n_777),
.Y(n_1663)
);

BUFx3_ASAP7_75t_L g1664 ( 
.A(n_1052),
.Y(n_1664)
);

BUFx2_ASAP7_75t_L g1665 ( 
.A(n_1240),
.Y(n_1665)
);

NOR2xp33_ASAP7_75t_L g1666 ( 
.A(n_1267),
.B(n_1001),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1090),
.Y(n_1667)
);

BUFx6f_ASAP7_75t_L g1668 ( 
.A(n_1225),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1091),
.Y(n_1669)
);

BUFx12f_ASAP7_75t_L g1670 ( 
.A(n_1267),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1093),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1301),
.B(n_888),
.Y(n_1672)
);

BUFx6f_ASAP7_75t_L g1673 ( 
.A(n_1225),
.Y(n_1673)
);

NOR2xp33_ASAP7_75t_L g1674 ( 
.A(n_1272),
.B(n_1005),
.Y(n_1674)
);

BUFx3_ASAP7_75t_L g1675 ( 
.A(n_1053),
.Y(n_1675)
);

INVx2_ASAP7_75t_L g1676 ( 
.A(n_1232),
.Y(n_1676)
);

BUFx6f_ASAP7_75t_L g1677 ( 
.A(n_1232),
.Y(n_1677)
);

BUFx6f_ASAP7_75t_L g1678 ( 
.A(n_1239),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_1239),
.Y(n_1679)
);

INVx2_ASAP7_75t_L g1680 ( 
.A(n_1242),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1387),
.B(n_782),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_SL g1682 ( 
.A(n_1272),
.B(n_1005),
.Y(n_1682)
);

NOR2xp33_ASAP7_75t_L g1683 ( 
.A(n_1275),
.B(n_785),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1388),
.B(n_787),
.Y(n_1684)
);

INVx4_ASAP7_75t_L g1685 ( 
.A(n_1395),
.Y(n_1685)
);

INVxp33_ASAP7_75t_SL g1686 ( 
.A(n_1275),
.Y(n_1686)
);

BUFx2_ASAP7_75t_L g1687 ( 
.A(n_1277),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1390),
.B(n_788),
.Y(n_1688)
);

BUFx6f_ASAP7_75t_L g1689 ( 
.A(n_1242),
.Y(n_1689)
);

INVxp67_ASAP7_75t_L g1690 ( 
.A(n_1310),
.Y(n_1690)
);

BUFx2_ASAP7_75t_L g1691 ( 
.A(n_1277),
.Y(n_1691)
);

BUFx3_ASAP7_75t_L g1692 ( 
.A(n_1054),
.Y(n_1692)
);

BUFx12f_ASAP7_75t_L g1693 ( 
.A(n_1281),
.Y(n_1693)
);

AND2x4_ASAP7_75t_L g1694 ( 
.A(n_1287),
.B(n_661),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_SL g1695 ( 
.A(n_1281),
.B(n_795),
.Y(n_1695)
);

INVx2_ASAP7_75t_L g1696 ( 
.A(n_1252),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1391),
.B(n_799),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1393),
.B(n_800),
.Y(n_1698)
);

AND2x4_ASAP7_75t_L g1699 ( 
.A(n_1288),
.B(n_664),
.Y(n_1699)
);

CKINVDCx5p33_ASAP7_75t_R g1700 ( 
.A(n_1262),
.Y(n_1700)
);

BUFx2_ASAP7_75t_L g1701 ( 
.A(n_1286),
.Y(n_1701)
);

BUFx6f_ASAP7_75t_L g1702 ( 
.A(n_1252),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1302),
.B(n_1303),
.Y(n_1703)
);

BUFx3_ASAP7_75t_L g1704 ( 
.A(n_1055),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1304),
.B(n_810),
.Y(n_1705)
);

BUFx3_ASAP7_75t_L g1706 ( 
.A(n_1056),
.Y(n_1706)
);

AND2x4_ASAP7_75t_L g1707 ( 
.A(n_1289),
.B(n_669),
.Y(n_1707)
);

BUFx12f_ASAP7_75t_L g1708 ( 
.A(n_1286),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1306),
.B(n_811),
.Y(n_1709)
);

NOR2xp33_ASAP7_75t_L g1710 ( 
.A(n_1308),
.B(n_812),
.Y(n_1710)
);

BUFx2_ASAP7_75t_L g1711 ( 
.A(n_1308),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1096),
.Y(n_1712)
);

AND2x4_ASAP7_75t_L g1713 ( 
.A(n_1291),
.B(n_680),
.Y(n_1713)
);

HB1xp67_ASAP7_75t_L g1714 ( 
.A(n_1023),
.Y(n_1714)
);

BUFx6f_ASAP7_75t_L g1715 ( 
.A(n_1255),
.Y(n_1715)
);

BUFx12f_ASAP7_75t_L g1716 ( 
.A(n_1321),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1307),
.B(n_888),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1099),
.Y(n_1718)
);

INVx4_ASAP7_75t_L g1719 ( 
.A(n_1074),
.Y(n_1719)
);

AND2x4_ASAP7_75t_L g1720 ( 
.A(n_1293),
.B(n_1309),
.Y(n_1720)
);

NOR2xp33_ASAP7_75t_L g1721 ( 
.A(n_1321),
.B(n_817),
.Y(n_1721)
);

NOR2xp33_ASAP7_75t_L g1722 ( 
.A(n_1322),
.B(n_823),
.Y(n_1722)
);

BUFx3_ASAP7_75t_L g1723 ( 
.A(n_1057),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1100),
.Y(n_1724)
);

INVx3_ASAP7_75t_L g1725 ( 
.A(n_1269),
.Y(n_1725)
);

INVx4_ASAP7_75t_L g1726 ( 
.A(n_1074),
.Y(n_1726)
);

BUFx6f_ASAP7_75t_L g1727 ( 
.A(n_1255),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1101),
.Y(n_1728)
);

BUFx6f_ASAP7_75t_L g1729 ( 
.A(n_1617),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1575),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1603),
.Y(n_1731)
);

NOR2xp33_ASAP7_75t_L g1732 ( 
.A(n_1518),
.B(n_1322),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1719),
.Y(n_1733)
);

INVx3_ASAP7_75t_L g1734 ( 
.A(n_1719),
.Y(n_1734)
);

BUFx2_ASAP7_75t_L g1735 ( 
.A(n_1429),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1611),
.Y(n_1736)
);

INVx6_ASAP7_75t_L g1737 ( 
.A(n_1459),
.Y(n_1737)
);

INVx2_ASAP7_75t_L g1738 ( 
.A(n_1719),
.Y(n_1738)
);

INVx2_ASAP7_75t_L g1739 ( 
.A(n_1726),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1625),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1629),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_SL g1742 ( 
.A(n_1443),
.B(n_1399),
.Y(n_1742)
);

AND2x6_ASAP7_75t_L g1743 ( 
.A(n_1443),
.B(n_1300),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1410),
.B(n_1269),
.Y(n_1744)
);

BUFx2_ASAP7_75t_L g1745 ( 
.A(n_1422),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1636),
.Y(n_1746)
);

INVx2_ASAP7_75t_L g1747 ( 
.A(n_1726),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1726),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1410),
.B(n_1290),
.Y(n_1749)
);

INVxp67_ASAP7_75t_L g1750 ( 
.A(n_1510),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1643),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_1400),
.Y(n_1752)
);

BUFx3_ASAP7_75t_L g1753 ( 
.A(n_1404),
.Y(n_1753)
);

INVx2_ASAP7_75t_L g1754 ( 
.A(n_1400),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1441),
.B(n_1325),
.Y(n_1755)
);

INVx2_ASAP7_75t_L g1756 ( 
.A(n_1413),
.Y(n_1756)
);

BUFx6f_ASAP7_75t_L g1757 ( 
.A(n_1617),
.Y(n_1757)
);

INVx3_ASAP7_75t_L g1758 ( 
.A(n_1449),
.Y(n_1758)
);

INVx3_ASAP7_75t_L g1759 ( 
.A(n_1449),
.Y(n_1759)
);

OA21x2_ASAP7_75t_L g1760 ( 
.A1(n_1705),
.A2(n_1062),
.B(n_1061),
.Y(n_1760)
);

INVx2_ASAP7_75t_L g1761 ( 
.A(n_1413),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1660),
.Y(n_1762)
);

BUFx6f_ASAP7_75t_L g1763 ( 
.A(n_1617),
.Y(n_1763)
);

INVx2_ASAP7_75t_L g1764 ( 
.A(n_1414),
.Y(n_1764)
);

INVx2_ASAP7_75t_L g1765 ( 
.A(n_1414),
.Y(n_1765)
);

BUFx6f_ASAP7_75t_L g1766 ( 
.A(n_1617),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1667),
.Y(n_1767)
);

BUFx6f_ASAP7_75t_L g1768 ( 
.A(n_1630),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1669),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1420),
.Y(n_1770)
);

BUFx8_ASAP7_75t_L g1771 ( 
.A(n_1438),
.Y(n_1771)
);

INVx2_ASAP7_75t_L g1772 ( 
.A(n_1420),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1431),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1671),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1712),
.Y(n_1775)
);

INVx3_ASAP7_75t_L g1776 ( 
.A(n_1476),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1718),
.Y(n_1777)
);

AND2x4_ASAP7_75t_L g1778 ( 
.A(n_1443),
.B(n_1174),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1724),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1728),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1447),
.B(n_1325),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_SL g1782 ( 
.A(n_1399),
.B(n_1367),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1576),
.Y(n_1783)
);

BUFx6f_ASAP7_75t_L g1784 ( 
.A(n_1630),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1576),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1397),
.B(n_1439),
.Y(n_1786)
);

INVxp67_ASAP7_75t_L g1787 ( 
.A(n_1530),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1585),
.Y(n_1788)
);

BUFx6f_ASAP7_75t_L g1789 ( 
.A(n_1630),
.Y(n_1789)
);

INVx2_ASAP7_75t_L g1790 ( 
.A(n_1431),
.Y(n_1790)
);

INVx2_ASAP7_75t_L g1791 ( 
.A(n_1433),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_1433),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1585),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1465),
.B(n_1490),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1416),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1496),
.B(n_1329),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1434),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1450),
.Y(n_1798)
);

INVx2_ASAP7_75t_L g1799 ( 
.A(n_1463),
.Y(n_1799)
);

BUFx6f_ASAP7_75t_L g1800 ( 
.A(n_1630),
.Y(n_1800)
);

BUFx2_ASAP7_75t_L g1801 ( 
.A(n_1534),
.Y(n_1801)
);

INVx2_ASAP7_75t_L g1802 ( 
.A(n_1463),
.Y(n_1802)
);

BUFx6f_ASAP7_75t_L g1803 ( 
.A(n_1634),
.Y(n_1803)
);

NOR2xp33_ASAP7_75t_SL g1804 ( 
.A(n_1497),
.B(n_1210),
.Y(n_1804)
);

INVxp33_ASAP7_75t_L g1805 ( 
.A(n_1714),
.Y(n_1805)
);

AND2x4_ASAP7_75t_L g1806 ( 
.A(n_1467),
.B(n_1174),
.Y(n_1806)
);

INVx3_ASAP7_75t_L g1807 ( 
.A(n_1476),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_1405),
.B(n_1329),
.Y(n_1808)
);

INVx2_ASAP7_75t_L g1809 ( 
.A(n_1491),
.Y(n_1809)
);

BUFx6f_ASAP7_75t_L g1810 ( 
.A(n_1634),
.Y(n_1810)
);

CKINVDCx16_ASAP7_75t_R g1811 ( 
.A(n_1638),
.Y(n_1811)
);

OA21x2_ASAP7_75t_L g1812 ( 
.A1(n_1709),
.A2(n_1065),
.B(n_1064),
.Y(n_1812)
);

AND2x4_ASAP7_75t_L g1813 ( 
.A(n_1467),
.B(n_1260),
.Y(n_1813)
);

AND2x4_ASAP7_75t_L g1814 ( 
.A(n_1467),
.B(n_1260),
.Y(n_1814)
);

CKINVDCx20_ASAP7_75t_R g1815 ( 
.A(n_1402),
.Y(n_1815)
);

AND2x4_ASAP7_75t_L g1816 ( 
.A(n_1426),
.B(n_1365),
.Y(n_1816)
);

BUFx8_ASAP7_75t_L g1817 ( 
.A(n_1438),
.Y(n_1817)
);

BUFx6f_ASAP7_75t_L g1818 ( 
.A(n_1634),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1458),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1480),
.Y(n_1820)
);

BUFx8_ASAP7_75t_L g1821 ( 
.A(n_1445),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1405),
.B(n_1346),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1502),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1405),
.B(n_1346),
.Y(n_1824)
);

BUFx6f_ASAP7_75t_L g1825 ( 
.A(n_1634),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1491),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1504),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1540),
.Y(n_1828)
);

AND2x4_ASAP7_75t_L g1829 ( 
.A(n_1426),
.B(n_1365),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1544),
.Y(n_1830)
);

BUFx6f_ASAP7_75t_L g1831 ( 
.A(n_1642),
.Y(n_1831)
);

BUFx6f_ASAP7_75t_L g1832 ( 
.A(n_1642),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1554),
.Y(n_1833)
);

INVx6_ASAP7_75t_L g1834 ( 
.A(n_1459),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1567),
.Y(n_1835)
);

INVx2_ASAP7_75t_L g1836 ( 
.A(n_1503),
.Y(n_1836)
);

INVx2_ASAP7_75t_L g1837 ( 
.A(n_1503),
.Y(n_1837)
);

HB1xp67_ASAP7_75t_L g1838 ( 
.A(n_1526),
.Y(n_1838)
);

INVx3_ASAP7_75t_L g1839 ( 
.A(n_1512),
.Y(n_1839)
);

BUFx2_ASAP7_75t_L g1840 ( 
.A(n_1437),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1569),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1703),
.Y(n_1842)
);

INVx1_ASAP7_75t_SL g1843 ( 
.A(n_1440),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_SL g1844 ( 
.A(n_1470),
.B(n_1367),
.Y(n_1844)
);

BUFx2_ASAP7_75t_L g1845 ( 
.A(n_1478),
.Y(n_1845)
);

INVx3_ASAP7_75t_L g1846 ( 
.A(n_1512),
.Y(n_1846)
);

AND3x2_ASAP7_75t_L g1847 ( 
.A(n_1577),
.B(n_1403),
.C(n_1462),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1703),
.Y(n_1848)
);

INVx1_ASAP7_75t_SL g1849 ( 
.A(n_1479),
.Y(n_1849)
);

OAI22xp5_ASAP7_75t_SL g1850 ( 
.A1(n_1508),
.A2(n_1095),
.B1(n_1124),
.B2(n_1111),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1725),
.Y(n_1851)
);

INVx3_ASAP7_75t_L g1852 ( 
.A(n_1517),
.Y(n_1852)
);

INVx2_ASAP7_75t_L g1853 ( 
.A(n_1521),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1396),
.B(n_1383),
.Y(n_1854)
);

CKINVDCx5p33_ASAP7_75t_R g1855 ( 
.A(n_1497),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1725),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1725),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1465),
.B(n_1290),
.Y(n_1858)
);

AND2x4_ASAP7_75t_L g1859 ( 
.A(n_1426),
.B(n_1366),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1685),
.Y(n_1860)
);

BUFx6f_ASAP7_75t_L g1861 ( 
.A(n_1642),
.Y(n_1861)
);

BUFx6f_ASAP7_75t_L g1862 ( 
.A(n_1642),
.Y(n_1862)
);

INVx2_ASAP7_75t_L g1863 ( 
.A(n_1521),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1685),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1685),
.Y(n_1865)
);

BUFx6f_ASAP7_75t_L g1866 ( 
.A(n_1645),
.Y(n_1866)
);

BUFx6f_ASAP7_75t_L g1867 ( 
.A(n_1645),
.Y(n_1867)
);

BUFx8_ASAP7_75t_L g1868 ( 
.A(n_1445),
.Y(n_1868)
);

AND2x2_ASAP7_75t_L g1869 ( 
.A(n_1490),
.B(n_1313),
.Y(n_1869)
);

CKINVDCx5p33_ASAP7_75t_R g1870 ( 
.A(n_1555),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1424),
.B(n_1383),
.Y(n_1871)
);

BUFx6f_ASAP7_75t_L g1872 ( 
.A(n_1645),
.Y(n_1872)
);

BUFx6f_ASAP7_75t_L g1873 ( 
.A(n_1645),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1398),
.B(n_1415),
.Y(n_1874)
);

BUFx2_ASAP7_75t_L g1875 ( 
.A(n_1483),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1517),
.Y(n_1876)
);

AND2x2_ASAP7_75t_L g1877 ( 
.A(n_1407),
.B(n_1457),
.Y(n_1877)
);

AND2x4_ASAP7_75t_L g1878 ( 
.A(n_1456),
.B(n_1366),
.Y(n_1878)
);

INVxp33_ASAP7_75t_SL g1879 ( 
.A(n_1427),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1548),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1548),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1563),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1563),
.Y(n_1883)
);

INVx2_ASAP7_75t_L g1884 ( 
.A(n_1543),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1398),
.B(n_1312),
.Y(n_1885)
);

BUFx6f_ASAP7_75t_L g1886 ( 
.A(n_1646),
.Y(n_1886)
);

BUFx6f_ASAP7_75t_L g1887 ( 
.A(n_1646),
.Y(n_1887)
);

AND2x4_ASAP7_75t_L g1888 ( 
.A(n_1456),
.B(n_1063),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1407),
.B(n_1313),
.Y(n_1889)
);

BUFx2_ASAP7_75t_L g1890 ( 
.A(n_1427),
.Y(n_1890)
);

AND2x4_ASAP7_75t_L g1891 ( 
.A(n_1456),
.B(n_1213),
.Y(n_1891)
);

INVx2_ASAP7_75t_L g1892 ( 
.A(n_1543),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1398),
.B(n_1314),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1605),
.Y(n_1894)
);

INVx3_ASAP7_75t_L g1895 ( 
.A(n_1605),
.Y(n_1895)
);

INVx2_ASAP7_75t_L g1896 ( 
.A(n_1568),
.Y(n_1896)
);

INVx2_ASAP7_75t_L g1897 ( 
.A(n_1568),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1608),
.Y(n_1898)
);

INVx3_ASAP7_75t_L g1899 ( 
.A(n_1608),
.Y(n_1899)
);

AND2x2_ASAP7_75t_L g1900 ( 
.A(n_1457),
.B(n_1323),
.Y(n_1900)
);

AND2x2_ASAP7_75t_L g1901 ( 
.A(n_1672),
.B(n_1323),
.Y(n_1901)
);

INVx2_ASAP7_75t_L g1902 ( 
.A(n_1578),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1639),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1639),
.Y(n_1904)
);

CKINVDCx16_ASAP7_75t_R g1905 ( 
.A(n_1409),
.Y(n_1905)
);

INVx2_ASAP7_75t_L g1906 ( 
.A(n_1578),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_L g1907 ( 
.A(n_1415),
.B(n_1317),
.Y(n_1907)
);

AND2x4_ASAP7_75t_L g1908 ( 
.A(n_1415),
.B(n_1103),
.Y(n_1908)
);

BUFx6f_ASAP7_75t_L g1909 ( 
.A(n_1646),
.Y(n_1909)
);

AND2x2_ASAP7_75t_L g1910 ( 
.A(n_1672),
.B(n_1319),
.Y(n_1910)
);

INVx2_ASAP7_75t_L g1911 ( 
.A(n_1600),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1664),
.Y(n_1912)
);

INVx2_ASAP7_75t_L g1913 ( 
.A(n_1600),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1664),
.Y(n_1914)
);

INVx2_ASAP7_75t_L g1915 ( 
.A(n_1619),
.Y(n_1915)
);

INVx2_ASAP7_75t_L g1916 ( 
.A(n_1619),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_SL g1917 ( 
.A(n_1471),
.B(n_1105),
.Y(n_1917)
);

BUFx6f_ASAP7_75t_L g1918 ( 
.A(n_1646),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1675),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1675),
.Y(n_1920)
);

AND2x4_ASAP7_75t_L g1921 ( 
.A(n_1419),
.B(n_1104),
.Y(n_1921)
);

INVx3_ASAP7_75t_L g1922 ( 
.A(n_1692),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1692),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1704),
.Y(n_1924)
);

INVx2_ASAP7_75t_L g1925 ( 
.A(n_1648),
.Y(n_1925)
);

NOR2xp33_ASAP7_75t_L g1926 ( 
.A(n_1528),
.B(n_1105),
.Y(n_1926)
);

HB1xp67_ASAP7_75t_L g1927 ( 
.A(n_1461),
.Y(n_1927)
);

INVx2_ASAP7_75t_L g1928 ( 
.A(n_1648),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_L g1929 ( 
.A(n_1419),
.B(n_1324),
.Y(n_1929)
);

AND2x2_ASAP7_75t_L g1930 ( 
.A(n_1717),
.B(n_1326),
.Y(n_1930)
);

INVx2_ASAP7_75t_L g1931 ( 
.A(n_1676),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1704),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_L g1933 ( 
.A(n_1419),
.B(n_1430),
.Y(n_1933)
);

INVx2_ASAP7_75t_L g1934 ( 
.A(n_1676),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1706),
.Y(n_1935)
);

INVx2_ASAP7_75t_L g1936 ( 
.A(n_1679),
.Y(n_1936)
);

BUFx8_ASAP7_75t_L g1937 ( 
.A(n_1451),
.Y(n_1937)
);

INVx2_ASAP7_75t_L g1938 ( 
.A(n_1679),
.Y(n_1938)
);

INVx3_ASAP7_75t_L g1939 ( 
.A(n_1706),
.Y(n_1939)
);

INVx2_ASAP7_75t_L g1940 ( 
.A(n_1680),
.Y(n_1940)
);

NOR2xp33_ASAP7_75t_L g1941 ( 
.A(n_1536),
.B(n_1114),
.Y(n_1941)
);

INVxp67_ASAP7_75t_L g1942 ( 
.A(n_1493),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_L g1943 ( 
.A(n_1436),
.B(n_1330),
.Y(n_1943)
);

INVx2_ASAP7_75t_L g1944 ( 
.A(n_1680),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_L g1945 ( 
.A(n_1454),
.B(n_1331),
.Y(n_1945)
);

INVx2_ASAP7_75t_L g1946 ( 
.A(n_1696),
.Y(n_1946)
);

BUFx3_ASAP7_75t_L g1947 ( 
.A(n_1404),
.Y(n_1947)
);

BUFx6f_ASAP7_75t_L g1948 ( 
.A(n_1668),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1723),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1723),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_L g1951 ( 
.A(n_1455),
.B(n_1333),
.Y(n_1951)
);

AND2x4_ASAP7_75t_L g1952 ( 
.A(n_1720),
.B(n_1509),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1444),
.Y(n_1953)
);

OAI22xp5_ASAP7_75t_SL g1954 ( 
.A1(n_1508),
.A2(n_1095),
.B1(n_1124),
.B2(n_1111),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1460),
.B(n_1334),
.Y(n_1955)
);

INVx3_ASAP7_75t_L g1956 ( 
.A(n_1668),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1444),
.Y(n_1957)
);

INVx3_ASAP7_75t_L g1958 ( 
.A(n_1668),
.Y(n_1958)
);

AND2x6_ASAP7_75t_L g1959 ( 
.A(n_1717),
.B(n_1556),
.Y(n_1959)
);

INVx4_ASAP7_75t_L g1960 ( 
.A(n_1612),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1444),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1448),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1448),
.Y(n_1963)
);

AND2x4_ASAP7_75t_L g1964 ( 
.A(n_1720),
.B(n_1106),
.Y(n_1964)
);

CKINVDCx16_ASAP7_75t_R g1965 ( 
.A(n_1409),
.Y(n_1965)
);

AND2x2_ASAP7_75t_L g1966 ( 
.A(n_1488),
.B(n_1336),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1448),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1474),
.Y(n_1968)
);

NOR2xp33_ASAP7_75t_L g1969 ( 
.A(n_1537),
.B(n_1114),
.Y(n_1969)
);

INVxp67_ASAP7_75t_L g1970 ( 
.A(n_1495),
.Y(n_1970)
);

CKINVDCx16_ASAP7_75t_R g1971 ( 
.A(n_1417),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1474),
.Y(n_1972)
);

AND2x2_ASAP7_75t_L g1973 ( 
.A(n_1488),
.B(n_1337),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_L g1974 ( 
.A(n_1466),
.B(n_1339),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1474),
.Y(n_1975)
);

INVx2_ASAP7_75t_L g1976 ( 
.A(n_1696),
.Y(n_1976)
);

INVx3_ASAP7_75t_L g1977 ( 
.A(n_1668),
.Y(n_1977)
);

INVx2_ASAP7_75t_L g1978 ( 
.A(n_1673),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1506),
.Y(n_1979)
);

HB1xp67_ASAP7_75t_L g1980 ( 
.A(n_1547),
.Y(n_1980)
);

BUFx6f_ASAP7_75t_L g1981 ( 
.A(n_1673),
.Y(n_1981)
);

AND2x2_ASAP7_75t_L g1982 ( 
.A(n_1488),
.B(n_1341),
.Y(n_1982)
);

INVx2_ASAP7_75t_L g1983 ( 
.A(n_1673),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1506),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1506),
.Y(n_1985)
);

NAND2xp5_ASAP7_75t_L g1986 ( 
.A(n_1482),
.B(n_1342),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_L g1987 ( 
.A(n_1683),
.B(n_1343),
.Y(n_1987)
);

BUFx8_ASAP7_75t_L g1988 ( 
.A(n_1451),
.Y(n_1988)
);

NOR2xp33_ASAP7_75t_L g1989 ( 
.A(n_1538),
.B(n_1233),
.Y(n_1989)
);

CKINVDCx8_ASAP7_75t_R g1990 ( 
.A(n_1552),
.Y(n_1990)
);

INVx2_ASAP7_75t_L g1991 ( 
.A(n_1673),
.Y(n_1991)
);

BUFx6f_ASAP7_75t_L g1992 ( 
.A(n_1677),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1515),
.Y(n_1993)
);

INVx2_ASAP7_75t_L g1994 ( 
.A(n_1677),
.Y(n_1994)
);

INVx2_ASAP7_75t_L g1995 ( 
.A(n_1677),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1515),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1515),
.Y(n_1997)
);

AND2x2_ASAP7_75t_L g1998 ( 
.A(n_1498),
.B(n_1344),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1535),
.Y(n_1999)
);

INVx3_ASAP7_75t_L g2000 ( 
.A(n_1677),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1535),
.Y(n_2001)
);

AND2x6_ASAP7_75t_L g2002 ( 
.A(n_1556),
.B(n_1347),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1535),
.Y(n_2003)
);

HB1xp67_ASAP7_75t_L g2004 ( 
.A(n_1498),
.Y(n_2004)
);

BUFx6f_ASAP7_75t_L g2005 ( 
.A(n_1678),
.Y(n_2005)
);

OAI22xp5_ASAP7_75t_SL g2006 ( 
.A1(n_1539),
.A2(n_1137),
.B1(n_1155),
.B2(n_1154),
.Y(n_2006)
);

AND2x2_ASAP7_75t_L g2007 ( 
.A(n_1498),
.B(n_1349),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1560),
.Y(n_2008)
);

BUFx6f_ASAP7_75t_L g2009 ( 
.A(n_1678),
.Y(n_2009)
);

INVx2_ASAP7_75t_L g2010 ( 
.A(n_1678),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1560),
.Y(n_2011)
);

AND2x2_ASAP7_75t_L g2012 ( 
.A(n_1501),
.B(n_1351),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1560),
.Y(n_2013)
);

BUFx6f_ASAP7_75t_L g2014 ( 
.A(n_1678),
.Y(n_2014)
);

INVx2_ASAP7_75t_L g2015 ( 
.A(n_1689),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_L g2016 ( 
.A(n_1710),
.B(n_1721),
.Y(n_2016)
);

INVx3_ASAP7_75t_L g2017 ( 
.A(n_1689),
.Y(n_2017)
);

BUFx6f_ASAP7_75t_L g2018 ( 
.A(n_1689),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1604),
.Y(n_2019)
);

OA21x2_ASAP7_75t_L g2020 ( 
.A1(n_1562),
.A2(n_1067),
.B(n_1066),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1604),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1604),
.Y(n_2022)
);

INVxp67_ASAP7_75t_L g2023 ( 
.A(n_1523),
.Y(n_2023)
);

HB1xp67_ASAP7_75t_L g2024 ( 
.A(n_1501),
.Y(n_2024)
);

AND2x4_ASAP7_75t_L g2025 ( 
.A(n_1720),
.B(n_1118),
.Y(n_2025)
);

BUFx6f_ASAP7_75t_L g2026 ( 
.A(n_1689),
.Y(n_2026)
);

AND2x2_ASAP7_75t_L g2027 ( 
.A(n_1501),
.B(n_1355),
.Y(n_2027)
);

BUFx6f_ASAP7_75t_L g2028 ( 
.A(n_1702),
.Y(n_2028)
);

OA21x2_ASAP7_75t_L g2029 ( 
.A1(n_1571),
.A2(n_1071),
.B(n_1068),
.Y(n_2029)
);

CKINVDCx6p67_ASAP7_75t_R g2030 ( 
.A(n_1489),
.Y(n_2030)
);

INVx3_ASAP7_75t_L g2031 ( 
.A(n_1702),
.Y(n_2031)
);

CKINVDCx20_ASAP7_75t_R g2032 ( 
.A(n_1402),
.Y(n_2032)
);

AND2x4_ASAP7_75t_L g2033 ( 
.A(n_1509),
.B(n_1120),
.Y(n_2033)
);

OA21x2_ASAP7_75t_L g2034 ( 
.A1(n_1590),
.A2(n_1078),
.B(n_1072),
.Y(n_2034)
);

AND2x4_ASAP7_75t_L g2035 ( 
.A(n_1509),
.B(n_1121),
.Y(n_2035)
);

CKINVDCx11_ASAP7_75t_R g2036 ( 
.A(n_1641),
.Y(n_2036)
);

AND2x4_ASAP7_75t_L g2037 ( 
.A(n_1421),
.B(n_1123),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1621),
.Y(n_2038)
);

AND2x6_ASAP7_75t_L g2039 ( 
.A(n_1556),
.B(n_1077),
.Y(n_2039)
);

INVx3_ASAP7_75t_L g2040 ( 
.A(n_1702),
.Y(n_2040)
);

AND2x4_ASAP7_75t_L g2041 ( 
.A(n_1421),
.B(n_1130),
.Y(n_2041)
);

BUFx2_ASAP7_75t_L g2042 ( 
.A(n_1533),
.Y(n_2042)
);

XOR2xp5_ASAP7_75t_L g2043 ( 
.A(n_1552),
.B(n_1297),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_L g2044 ( 
.A(n_1722),
.B(n_1079),
.Y(n_2044)
);

AND2x4_ASAP7_75t_L g2045 ( 
.A(n_1421),
.B(n_1131),
.Y(n_2045)
);

NAND2xp5_ASAP7_75t_L g2046 ( 
.A(n_1423),
.B(n_1284),
.Y(n_2046)
);

BUFx2_ASAP7_75t_L g2047 ( 
.A(n_1582),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1621),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1621),
.Y(n_2049)
);

BUFx6f_ASAP7_75t_L g2050 ( 
.A(n_1702),
.Y(n_2050)
);

INVx2_ASAP7_75t_L g2051 ( 
.A(n_1715),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_1622),
.Y(n_2052)
);

AND2x6_ASAP7_75t_L g2053 ( 
.A(n_1626),
.B(n_1077),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_1622),
.Y(n_2054)
);

NAND2x1p5_ASAP7_75t_L g2055 ( 
.A(n_1511),
.B(n_1385),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_1622),
.Y(n_2056)
);

HB1xp67_ASAP7_75t_L g2057 ( 
.A(n_1632),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_1655),
.Y(n_2058)
);

HB1xp67_ASAP7_75t_L g2059 ( 
.A(n_1690),
.Y(n_2059)
);

INVx2_ASAP7_75t_L g2060 ( 
.A(n_1715),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_1655),
.Y(n_2061)
);

BUFx6f_ASAP7_75t_L g2062 ( 
.A(n_1715),
.Y(n_2062)
);

INVx1_ASAP7_75t_SL g2063 ( 
.A(n_1624),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_1655),
.Y(n_2064)
);

INVx6_ASAP7_75t_L g2065 ( 
.A(n_1459),
.Y(n_2065)
);

BUFx6f_ASAP7_75t_L g2066 ( 
.A(n_1715),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_1446),
.Y(n_2067)
);

NOR2x1_ASAP7_75t_L g2068 ( 
.A(n_1527),
.B(n_1354),
.Y(n_2068)
);

INVx2_ASAP7_75t_L g2069 ( 
.A(n_1727),
.Y(n_2069)
);

INVx3_ASAP7_75t_L g2070 ( 
.A(n_1727),
.Y(n_2070)
);

BUFx6f_ASAP7_75t_L g2071 ( 
.A(n_1727),
.Y(n_2071)
);

INVx3_ASAP7_75t_L g2072 ( 
.A(n_1727),
.Y(n_2072)
);

INVx1_ASAP7_75t_SL g2073 ( 
.A(n_1627),
.Y(n_2073)
);

BUFx6f_ASAP7_75t_L g2074 ( 
.A(n_1411),
.Y(n_2074)
);

NAND2xp5_ASAP7_75t_L g2075 ( 
.A(n_1532),
.B(n_1318),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_1505),
.Y(n_2076)
);

INVx3_ASAP7_75t_L g2077 ( 
.A(n_1411),
.Y(n_2077)
);

BUFx8_ASAP7_75t_L g2078 ( 
.A(n_1453),
.Y(n_2078)
);

HB1xp67_ASAP7_75t_L g2079 ( 
.A(n_1665),
.Y(n_2079)
);

INVx2_ASAP7_75t_L g2080 ( 
.A(n_1514),
.Y(n_2080)
);

INVx2_ASAP7_75t_L g2081 ( 
.A(n_1514),
.Y(n_2081)
);

BUFx6f_ASAP7_75t_L g2082 ( 
.A(n_1411),
.Y(n_2082)
);

AND3x2_ASAP7_75t_L g2083 ( 
.A(n_1687),
.B(n_1043),
.C(n_1278),
.Y(n_2083)
);

BUFx2_ASAP7_75t_L g2084 ( 
.A(n_1691),
.Y(n_2084)
);

AND2x2_ASAP7_75t_L g2085 ( 
.A(n_1505),
.B(n_1561),
.Y(n_2085)
);

NAND2xp5_ASAP7_75t_L g2086 ( 
.A(n_1529),
.B(n_1318),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_1561),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_1572),
.Y(n_2088)
);

BUFx6f_ASAP7_75t_L g2089 ( 
.A(n_1411),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_1572),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_1579),
.Y(n_2091)
);

INVx2_ASAP7_75t_L g2092 ( 
.A(n_1514),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_1579),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_1584),
.Y(n_2094)
);

BUFx6f_ASAP7_75t_L g2095 ( 
.A(n_1412),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_1795),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_1797),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_SL g2098 ( 
.A(n_1942),
.B(n_1511),
.Y(n_2098)
);

INVx2_ASAP7_75t_L g2099 ( 
.A(n_1752),
.Y(n_2099)
);

AND2x2_ASAP7_75t_L g2100 ( 
.A(n_1794),
.B(n_1584),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_1798),
.Y(n_2101)
);

AOI21x1_ASAP7_75t_L g2102 ( 
.A1(n_2044),
.A2(n_1616),
.B(n_1602),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_1819),
.Y(n_2103)
);

INVx5_ASAP7_75t_L g2104 ( 
.A(n_1960),
.Y(n_2104)
);

INVx3_ASAP7_75t_L g2105 ( 
.A(n_1758),
.Y(n_2105)
);

NOR2xp33_ASAP7_75t_L g2106 ( 
.A(n_1970),
.B(n_1539),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_1820),
.Y(n_2107)
);

NAND3xp33_ASAP7_75t_L g2108 ( 
.A(n_2075),
.B(n_1546),
.C(n_1541),
.Y(n_2108)
);

BUFx6f_ASAP7_75t_SL g2109 ( 
.A(n_1959),
.Y(n_2109)
);

BUFx6f_ASAP7_75t_SL g2110 ( 
.A(n_1959),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_1823),
.Y(n_2111)
);

AND2x2_ASAP7_75t_L g2112 ( 
.A(n_1794),
.B(n_1592),
.Y(n_2112)
);

AOI21x1_ASAP7_75t_L g2113 ( 
.A1(n_1752),
.A2(n_1628),
.B(n_1623),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_1827),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_1828),
.Y(n_2115)
);

INVx2_ASAP7_75t_L g2116 ( 
.A(n_1754),
.Y(n_2116)
);

INVx2_ASAP7_75t_L g2117 ( 
.A(n_1754),
.Y(n_2117)
);

NAND2xp33_ASAP7_75t_L g2118 ( 
.A(n_1743),
.B(n_1553),
.Y(n_2118)
);

NAND2xp5_ASAP7_75t_SL g2119 ( 
.A(n_2023),
.B(n_1565),
.Y(n_2119)
);

NAND2xp5_ASAP7_75t_SL g2120 ( 
.A(n_1778),
.B(n_1565),
.Y(n_2120)
);

INVx2_ASAP7_75t_L g2121 ( 
.A(n_1756),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_SL g2122 ( 
.A(n_1778),
.B(n_1653),
.Y(n_2122)
);

NAND2xp5_ASAP7_75t_L g2123 ( 
.A(n_2016),
.B(n_1557),
.Y(n_2123)
);

INVx2_ASAP7_75t_L g2124 ( 
.A(n_1756),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_1830),
.Y(n_2125)
);

AOI21x1_ASAP7_75t_L g2126 ( 
.A1(n_1761),
.A2(n_1697),
.B(n_1688),
.Y(n_2126)
);

AOI22xp5_ASAP7_75t_L g2127 ( 
.A1(n_1743),
.A2(n_1653),
.B1(n_1686),
.B2(n_1618),
.Y(n_2127)
);

INVx2_ASAP7_75t_L g2128 ( 
.A(n_1761),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_1833),
.Y(n_2129)
);

INVx2_ASAP7_75t_L g2130 ( 
.A(n_1764),
.Y(n_2130)
);

INVx2_ASAP7_75t_L g2131 ( 
.A(n_1764),
.Y(n_2131)
);

INVx2_ASAP7_75t_L g2132 ( 
.A(n_1765),
.Y(n_2132)
);

INVx3_ASAP7_75t_L g2133 ( 
.A(n_1758),
.Y(n_2133)
);

BUFx10_ASAP7_75t_L g2134 ( 
.A(n_1855),
.Y(n_2134)
);

NAND2xp5_ASAP7_75t_SL g2135 ( 
.A(n_1778),
.B(n_1686),
.Y(n_2135)
);

INVx2_ASAP7_75t_L g2136 ( 
.A(n_1765),
.Y(n_2136)
);

INVx2_ASAP7_75t_L g2137 ( 
.A(n_1770),
.Y(n_2137)
);

BUFx6f_ASAP7_75t_L g2138 ( 
.A(n_1729),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_1835),
.Y(n_2139)
);

INVx2_ASAP7_75t_SL g2140 ( 
.A(n_1735),
.Y(n_2140)
);

BUFx6f_ASAP7_75t_L g2141 ( 
.A(n_1729),
.Y(n_2141)
);

BUFx2_ASAP7_75t_L g2142 ( 
.A(n_1745),
.Y(n_2142)
);

NAND2xp5_ASAP7_75t_L g2143 ( 
.A(n_1987),
.B(n_1587),
.Y(n_2143)
);

NOR2xp33_ASAP7_75t_L g2144 ( 
.A(n_2086),
.B(n_1701),
.Y(n_2144)
);

INVx1_ASAP7_75t_L g2145 ( 
.A(n_1841),
.Y(n_2145)
);

CKINVDCx20_ASAP7_75t_R g2146 ( 
.A(n_1850),
.Y(n_2146)
);

INVx2_ASAP7_75t_L g2147 ( 
.A(n_1770),
.Y(n_2147)
);

INVx2_ASAP7_75t_L g2148 ( 
.A(n_1772),
.Y(n_2148)
);

INVx2_ASAP7_75t_L g2149 ( 
.A(n_1772),
.Y(n_2149)
);

INVx3_ASAP7_75t_L g2150 ( 
.A(n_1758),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_1860),
.Y(n_2151)
);

INVx2_ASAP7_75t_L g2152 ( 
.A(n_1773),
.Y(n_2152)
);

INVx8_ASAP7_75t_L g2153 ( 
.A(n_2002),
.Y(n_2153)
);

INVx2_ASAP7_75t_L g2154 ( 
.A(n_1773),
.Y(n_2154)
);

NAND2xp5_ASAP7_75t_SL g2155 ( 
.A(n_1926),
.B(n_1711),
.Y(n_2155)
);

NAND2xp5_ASAP7_75t_L g2156 ( 
.A(n_1732),
.B(n_1598),
.Y(n_2156)
);

INVx3_ASAP7_75t_L g2157 ( 
.A(n_1759),
.Y(n_2157)
);

INVx2_ASAP7_75t_L g2158 ( 
.A(n_1790),
.Y(n_2158)
);

INVx2_ASAP7_75t_L g2159 ( 
.A(n_1790),
.Y(n_2159)
);

NOR2xp33_ASAP7_75t_L g2160 ( 
.A(n_1786),
.B(n_1735),
.Y(n_2160)
);

INVxp33_ASAP7_75t_L g2161 ( 
.A(n_1838),
.Y(n_2161)
);

NAND2xp5_ASAP7_75t_L g2162 ( 
.A(n_1732),
.B(n_1926),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_1864),
.Y(n_2163)
);

BUFx10_ASAP7_75t_L g2164 ( 
.A(n_1855),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_1865),
.Y(n_2165)
);

AOI22xp5_ASAP7_75t_L g2166 ( 
.A1(n_1743),
.A2(n_1618),
.B1(n_1661),
.B2(n_1644),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_1736),
.Y(n_2167)
);

NAND2xp33_ASAP7_75t_SL g2168 ( 
.A(n_1871),
.B(n_1464),
.Y(n_2168)
);

NAND2xp5_ASAP7_75t_L g2169 ( 
.A(n_1941),
.B(n_1635),
.Y(n_2169)
);

BUFx6f_ASAP7_75t_L g2170 ( 
.A(n_1729),
.Y(n_2170)
);

INVx2_ASAP7_75t_L g2171 ( 
.A(n_1791),
.Y(n_2171)
);

NOR2xp33_ASAP7_75t_L g2172 ( 
.A(n_1941),
.B(n_1278),
.Y(n_2172)
);

INVx2_ASAP7_75t_L g2173 ( 
.A(n_1791),
.Y(n_2173)
);

INVx1_ASAP7_75t_L g2174 ( 
.A(n_1740),
.Y(n_2174)
);

BUFx10_ASAP7_75t_L g2175 ( 
.A(n_1870),
.Y(n_2175)
);

INVx2_ASAP7_75t_L g2176 ( 
.A(n_1792),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_1741),
.Y(n_2177)
);

INVx3_ASAP7_75t_L g2178 ( 
.A(n_1759),
.Y(n_2178)
);

INVx2_ASAP7_75t_L g2179 ( 
.A(n_1792),
.Y(n_2179)
);

BUFx6f_ASAP7_75t_L g2180 ( 
.A(n_1729),
.Y(n_2180)
);

INVx2_ASAP7_75t_SL g2181 ( 
.A(n_1816),
.Y(n_2181)
);

NAND2xp5_ASAP7_75t_SL g2182 ( 
.A(n_1969),
.B(n_1666),
.Y(n_2182)
);

AND2x2_ASAP7_75t_L g2183 ( 
.A(n_1877),
.B(n_1593),
.Y(n_2183)
);

NOR2xp33_ASAP7_75t_L g2184 ( 
.A(n_1969),
.B(n_1989),
.Y(n_2184)
);

INVx8_ASAP7_75t_L g2185 ( 
.A(n_2002),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_1746),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_1751),
.Y(n_2187)
);

INVx2_ASAP7_75t_L g2188 ( 
.A(n_1799),
.Y(n_2188)
);

NAND2xp5_ASAP7_75t_SL g2189 ( 
.A(n_1989),
.B(n_1674),
.Y(n_2189)
);

INVx2_ASAP7_75t_L g2190 ( 
.A(n_1799),
.Y(n_2190)
);

INVx2_ASAP7_75t_SL g2191 ( 
.A(n_1816),
.Y(n_2191)
);

NOR2x1p5_ASAP7_75t_L g2192 ( 
.A(n_1870),
.B(n_1555),
.Y(n_2192)
);

INVx3_ASAP7_75t_L g2193 ( 
.A(n_1759),
.Y(n_2193)
);

INVx2_ASAP7_75t_L g2194 ( 
.A(n_1802),
.Y(n_2194)
);

INVx3_ASAP7_75t_L g2195 ( 
.A(n_1776),
.Y(n_2195)
);

BUFx3_ASAP7_75t_L g2196 ( 
.A(n_1737),
.Y(n_2196)
);

NAND3xp33_ASAP7_75t_L g2197 ( 
.A(n_1755),
.B(n_1781),
.C(n_1796),
.Y(n_2197)
);

CKINVDCx5p33_ASAP7_75t_R g2198 ( 
.A(n_2036),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_1762),
.Y(n_2199)
);

NAND3xp33_ASAP7_75t_L g2200 ( 
.A(n_1854),
.B(n_1682),
.C(n_1649),
.Y(n_2200)
);

INVx2_ASAP7_75t_L g2201 ( 
.A(n_1802),
.Y(n_2201)
);

INVxp67_ASAP7_75t_SL g2202 ( 
.A(n_1776),
.Y(n_2202)
);

INVx1_ASAP7_75t_L g2203 ( 
.A(n_1767),
.Y(n_2203)
);

CKINVDCx5p33_ASAP7_75t_R g2204 ( 
.A(n_2036),
.Y(n_2204)
);

INVx8_ASAP7_75t_L g2205 ( 
.A(n_2002),
.Y(n_2205)
);

INVx2_ASAP7_75t_L g2206 ( 
.A(n_1809),
.Y(n_2206)
);

BUFx3_ASAP7_75t_L g2207 ( 
.A(n_1737),
.Y(n_2207)
);

BUFx10_ASAP7_75t_L g2208 ( 
.A(n_2083),
.Y(n_2208)
);

NAND3xp33_ASAP7_75t_L g2209 ( 
.A(n_2046),
.B(n_1682),
.C(n_1649),
.Y(n_2209)
);

NOR2xp33_ASAP7_75t_L g2210 ( 
.A(n_1844),
.B(n_1464),
.Y(n_2210)
);

NAND2xp5_ASAP7_75t_SL g2211 ( 
.A(n_1816),
.B(n_1829),
.Y(n_2211)
);

BUFx6f_ASAP7_75t_SL g2212 ( 
.A(n_1959),
.Y(n_2212)
);

NAND2xp33_ASAP7_75t_SL g2213 ( 
.A(n_1877),
.B(n_1524),
.Y(n_2213)
);

NAND2xp5_ASAP7_75t_SL g2214 ( 
.A(n_1829),
.B(n_1626),
.Y(n_2214)
);

NAND2xp5_ASAP7_75t_SL g2215 ( 
.A(n_1829),
.B(n_1626),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_1769),
.Y(n_2216)
);

NOR2xp33_ASAP7_75t_L g2217 ( 
.A(n_1844),
.B(n_1524),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_1774),
.Y(n_2218)
);

BUFx3_ASAP7_75t_L g2219 ( 
.A(n_1737),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_1775),
.Y(n_2220)
);

INVx2_ASAP7_75t_L g2221 ( 
.A(n_1809),
.Y(n_2221)
);

NAND2xp5_ASAP7_75t_L g2222 ( 
.A(n_1933),
.B(n_1592),
.Y(n_2222)
);

INVx2_ASAP7_75t_L g2223 ( 
.A(n_1826),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_1777),
.Y(n_2224)
);

INVx2_ASAP7_75t_L g2225 ( 
.A(n_1826),
.Y(n_2225)
);

AOI21x1_ASAP7_75t_L g2226 ( 
.A1(n_1836),
.A2(n_1853),
.B(n_1837),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_1779),
.Y(n_2227)
);

INVx2_ASAP7_75t_L g2228 ( 
.A(n_1836),
.Y(n_2228)
);

INVx2_ASAP7_75t_L g2229 ( 
.A(n_1837),
.Y(n_2229)
);

INVx1_ASAP7_75t_SL g2230 ( 
.A(n_1801),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_1780),
.Y(n_2231)
);

INVx5_ASAP7_75t_L g2232 ( 
.A(n_1960),
.Y(n_2232)
);

NAND2xp33_ASAP7_75t_SL g2233 ( 
.A(n_1917),
.B(n_1570),
.Y(n_2233)
);

NAND2xp5_ASAP7_75t_SL g2234 ( 
.A(n_1859),
.B(n_1878),
.Y(n_2234)
);

NAND2xp5_ASAP7_75t_L g2235 ( 
.A(n_1858),
.B(n_1869),
.Y(n_2235)
);

INVx3_ASAP7_75t_L g2236 ( 
.A(n_1776),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_1730),
.Y(n_2237)
);

INVx2_ASAP7_75t_L g2238 ( 
.A(n_1853),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_1731),
.Y(n_2239)
);

INVx2_ASAP7_75t_L g2240 ( 
.A(n_1863),
.Y(n_2240)
);

AO21x2_ASAP7_75t_L g2241 ( 
.A1(n_1742),
.A2(n_1695),
.B(n_1663),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_1851),
.Y(n_2242)
);

BUFx3_ASAP7_75t_L g2243 ( 
.A(n_1834),
.Y(n_2243)
);

INVx2_ASAP7_75t_SL g2244 ( 
.A(n_1859),
.Y(n_2244)
);

NAND2xp33_ASAP7_75t_SL g2245 ( 
.A(n_1917),
.B(n_1570),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_1856),
.Y(n_2246)
);

BUFx6f_ASAP7_75t_L g2247 ( 
.A(n_1757),
.Y(n_2247)
);

INVx2_ASAP7_75t_L g2248 ( 
.A(n_1863),
.Y(n_2248)
);

CKINVDCx5p33_ASAP7_75t_R g2249 ( 
.A(n_2030),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_1857),
.Y(n_2250)
);

INVx2_ASAP7_75t_L g2251 ( 
.A(n_1884),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_1953),
.Y(n_2252)
);

NOR2xp33_ASAP7_75t_L g2253 ( 
.A(n_1750),
.B(n_1549),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_1957),
.Y(n_2254)
);

INVx3_ASAP7_75t_L g2255 ( 
.A(n_1807),
.Y(n_2255)
);

NOR2xp33_ASAP7_75t_L g2256 ( 
.A(n_1787),
.B(n_1583),
.Y(n_2256)
);

INVxp33_ASAP7_75t_L g2257 ( 
.A(n_1801),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_1961),
.Y(n_2258)
);

INVx2_ASAP7_75t_L g2259 ( 
.A(n_1884),
.Y(n_2259)
);

INVxp33_ASAP7_75t_L g2260 ( 
.A(n_1745),
.Y(n_2260)
);

INVx2_ASAP7_75t_L g2261 ( 
.A(n_1892),
.Y(n_2261)
);

INVx2_ASAP7_75t_L g2262 ( 
.A(n_1892),
.Y(n_2262)
);

INVx1_ASAP7_75t_L g2263 ( 
.A(n_1962),
.Y(n_2263)
);

INVx2_ASAP7_75t_L g2264 ( 
.A(n_1896),
.Y(n_2264)
);

AND2x2_ASAP7_75t_L g2265 ( 
.A(n_2085),
.B(n_1593),
.Y(n_2265)
);

AND3x1_ASAP7_75t_L g2266 ( 
.A(n_2079),
.B(n_1522),
.C(n_1647),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_1963),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_1967),
.Y(n_2268)
);

NAND3xp33_ASAP7_75t_L g2269 ( 
.A(n_1742),
.B(n_1650),
.C(n_1631),
.Y(n_2269)
);

NAND2xp33_ASAP7_75t_SL g2270 ( 
.A(n_1782),
.B(n_1808),
.Y(n_2270)
);

INVx2_ASAP7_75t_L g2271 ( 
.A(n_1896),
.Y(n_2271)
);

INVx3_ASAP7_75t_L g2272 ( 
.A(n_1807),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_1968),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_1972),
.Y(n_2274)
);

INVx1_ASAP7_75t_L g2275 ( 
.A(n_1975),
.Y(n_2275)
);

INVx1_ASAP7_75t_L g2276 ( 
.A(n_1979),
.Y(n_2276)
);

INVxp33_ASAP7_75t_SL g2277 ( 
.A(n_2063),
.Y(n_2277)
);

INVx1_ASAP7_75t_L g2278 ( 
.A(n_1984),
.Y(n_2278)
);

INVx2_ASAP7_75t_L g2279 ( 
.A(n_1897),
.Y(n_2279)
);

AO22x1_ASAP7_75t_L g2280 ( 
.A1(n_1743),
.A2(n_1553),
.B1(n_1654),
.B2(n_1652),
.Y(n_2280)
);

INVx5_ASAP7_75t_L g2281 ( 
.A(n_1960),
.Y(n_2281)
);

NAND2xp5_ASAP7_75t_SL g2282 ( 
.A(n_1859),
.B(n_1652),
.Y(n_2282)
);

INVx2_ASAP7_75t_L g2283 ( 
.A(n_1897),
.Y(n_2283)
);

INVx2_ASAP7_75t_L g2284 ( 
.A(n_1902),
.Y(n_2284)
);

INVx2_ASAP7_75t_L g2285 ( 
.A(n_1902),
.Y(n_2285)
);

INVx2_ASAP7_75t_L g2286 ( 
.A(n_1906),
.Y(n_2286)
);

AND2x2_ASAP7_75t_L g2287 ( 
.A(n_2085),
.B(n_1597),
.Y(n_2287)
);

NAND2xp5_ASAP7_75t_SL g2288 ( 
.A(n_1878),
.B(n_1652),
.Y(n_2288)
);

AND2x4_ASAP7_75t_L g2289 ( 
.A(n_1952),
.B(n_1597),
.Y(n_2289)
);

CKINVDCx11_ASAP7_75t_R g2290 ( 
.A(n_1815),
.Y(n_2290)
);

NAND2xp5_ASAP7_75t_SL g2291 ( 
.A(n_1878),
.B(n_1657),
.Y(n_2291)
);

INVx2_ASAP7_75t_L g2292 ( 
.A(n_1906),
.Y(n_2292)
);

INVx2_ASAP7_75t_L g2293 ( 
.A(n_1911),
.Y(n_2293)
);

AO21x2_ASAP7_75t_L g2294 ( 
.A1(n_1874),
.A2(n_1983),
.B(n_1978),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_1985),
.Y(n_2295)
);

NAND2xp5_ASAP7_75t_SL g2296 ( 
.A(n_1952),
.B(n_1657),
.Y(n_2296)
);

INVx2_ASAP7_75t_L g2297 ( 
.A(n_1911),
.Y(n_2297)
);

BUFx6f_ASAP7_75t_L g2298 ( 
.A(n_1757),
.Y(n_2298)
);

INVx4_ASAP7_75t_L g2299 ( 
.A(n_1734),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_1993),
.Y(n_2300)
);

BUFx6f_ASAP7_75t_L g2301 ( 
.A(n_1757),
.Y(n_2301)
);

NAND2xp5_ASAP7_75t_L g2302 ( 
.A(n_1858),
.B(n_1640),
.Y(n_2302)
);

AND2x2_ASAP7_75t_L g2303 ( 
.A(n_1869),
.B(n_1640),
.Y(n_2303)
);

INVx3_ASAP7_75t_L g2304 ( 
.A(n_1807),
.Y(n_2304)
);

INVx2_ASAP7_75t_L g2305 ( 
.A(n_1913),
.Y(n_2305)
);

INVx2_ASAP7_75t_L g2306 ( 
.A(n_1913),
.Y(n_2306)
);

INVx5_ASAP7_75t_L g2307 ( 
.A(n_1734),
.Y(n_2307)
);

INVx1_ASAP7_75t_L g2308 ( 
.A(n_1996),
.Y(n_2308)
);

OR2x2_ASAP7_75t_L g2309 ( 
.A(n_2073),
.B(n_1350),
.Y(n_2309)
);

INVx2_ASAP7_75t_L g2310 ( 
.A(n_1915),
.Y(n_2310)
);

AND2x2_ASAP7_75t_L g2311 ( 
.A(n_1889),
.B(n_1900),
.Y(n_2311)
);

NOR2xp33_ASAP7_75t_SL g2312 ( 
.A(n_1879),
.B(n_1610),
.Y(n_2312)
);

NAND2xp5_ASAP7_75t_SL g2313 ( 
.A(n_1952),
.B(n_1654),
.Y(n_2313)
);

AND2x2_ASAP7_75t_L g2314 ( 
.A(n_1889),
.B(n_1647),
.Y(n_2314)
);

NAND2xp33_ASAP7_75t_L g2315 ( 
.A(n_1743),
.B(n_2002),
.Y(n_2315)
);

OR2x2_ASAP7_75t_L g2316 ( 
.A(n_1843),
.B(n_1371),
.Y(n_2316)
);

NAND2x1p5_ASAP7_75t_L g2317 ( 
.A(n_1839),
.B(n_1612),
.Y(n_2317)
);

NAND2xp5_ASAP7_75t_L g2318 ( 
.A(n_1900),
.B(n_1654),
.Y(n_2318)
);

AOI22xp33_ASAP7_75t_L g2319 ( 
.A1(n_1959),
.A2(n_1743),
.B1(n_1891),
.B2(n_1888),
.Y(n_2319)
);

BUFx2_ASAP7_75t_L g2320 ( 
.A(n_1840),
.Y(n_2320)
);

NAND2xp5_ASAP7_75t_SL g2321 ( 
.A(n_1753),
.B(n_1657),
.Y(n_2321)
);

NAND3xp33_ASAP7_75t_L g2322 ( 
.A(n_2068),
.B(n_1695),
.C(n_1442),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_1997),
.Y(n_2323)
);

NAND2xp5_ASAP7_75t_L g2324 ( 
.A(n_1943),
.B(n_1945),
.Y(n_2324)
);

NAND2xp5_ASAP7_75t_L g2325 ( 
.A(n_1951),
.B(n_1694),
.Y(n_2325)
);

CKINVDCx20_ASAP7_75t_R g2326 ( 
.A(n_1954),
.Y(n_2326)
);

BUFx6f_ASAP7_75t_L g2327 ( 
.A(n_1757),
.Y(n_2327)
);

NAND2xp5_ASAP7_75t_SL g2328 ( 
.A(n_1753),
.B(n_1417),
.Y(n_2328)
);

INVx2_ASAP7_75t_L g2329 ( 
.A(n_1915),
.Y(n_2329)
);

NAND2xp5_ASAP7_75t_SL g2330 ( 
.A(n_1947),
.B(n_1694),
.Y(n_2330)
);

INVx1_ASAP7_75t_L g2331 ( 
.A(n_1999),
.Y(n_2331)
);

INVx2_ASAP7_75t_L g2332 ( 
.A(n_1916),
.Y(n_2332)
);

INVx2_ASAP7_75t_L g2333 ( 
.A(n_1916),
.Y(n_2333)
);

INVx1_ASAP7_75t_L g2334 ( 
.A(n_2001),
.Y(n_2334)
);

NAND2xp5_ASAP7_75t_SL g2335 ( 
.A(n_1947),
.B(n_1694),
.Y(n_2335)
);

INVx2_ASAP7_75t_SL g2336 ( 
.A(n_1908),
.Y(n_2336)
);

NAND2xp5_ASAP7_75t_SL g2337 ( 
.A(n_1822),
.B(n_1699),
.Y(n_2337)
);

INVx2_ASAP7_75t_L g2338 ( 
.A(n_1925),
.Y(n_2338)
);

BUFx2_ASAP7_75t_L g2339 ( 
.A(n_1840),
.Y(n_2339)
);

NAND2xp33_ASAP7_75t_L g2340 ( 
.A(n_2002),
.B(n_1553),
.Y(n_2340)
);

INVx1_ASAP7_75t_L g2341 ( 
.A(n_2003),
.Y(n_2341)
);

CKINVDCx5p33_ASAP7_75t_R g2342 ( 
.A(n_2030),
.Y(n_2342)
);

NAND2xp5_ASAP7_75t_SL g2343 ( 
.A(n_1824),
.B(n_1699),
.Y(n_2343)
);

INVx1_ASAP7_75t_L g2344 ( 
.A(n_2008),
.Y(n_2344)
);

NAND2xp33_ASAP7_75t_L g2345 ( 
.A(n_2002),
.B(n_1553),
.Y(n_2345)
);

NAND2xp5_ASAP7_75t_SL g2346 ( 
.A(n_2055),
.B(n_1699),
.Y(n_2346)
);

INVx2_ASAP7_75t_SL g2347 ( 
.A(n_1908),
.Y(n_2347)
);

INVx2_ASAP7_75t_L g2348 ( 
.A(n_1925),
.Y(n_2348)
);

INVx2_ASAP7_75t_L g2349 ( 
.A(n_1928),
.Y(n_2349)
);

NAND2xp5_ASAP7_75t_L g2350 ( 
.A(n_1955),
.B(n_1707),
.Y(n_2350)
);

INVxp33_ASAP7_75t_L g2351 ( 
.A(n_2043),
.Y(n_2351)
);

AOI22xp33_ASAP7_75t_L g2352 ( 
.A1(n_1959),
.A2(n_1012),
.B1(n_1553),
.B2(n_1707),
.Y(n_2352)
);

INVx4_ASAP7_75t_L g2353 ( 
.A(n_1734),
.Y(n_2353)
);

NAND2xp5_ASAP7_75t_SL g2354 ( 
.A(n_2055),
.B(n_1806),
.Y(n_2354)
);

INVx2_ASAP7_75t_L g2355 ( 
.A(n_1928),
.Y(n_2355)
);

BUFx3_ASAP7_75t_L g2356 ( 
.A(n_1834),
.Y(n_2356)
);

NAND2xp5_ASAP7_75t_SL g2357 ( 
.A(n_1806),
.B(n_1707),
.Y(n_2357)
);

INVx11_ASAP7_75t_L g2358 ( 
.A(n_1771),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_2011),
.Y(n_2359)
);

NAND2xp5_ASAP7_75t_L g2360 ( 
.A(n_1974),
.B(n_1713),
.Y(n_2360)
);

AND2x4_ASAP7_75t_L g2361 ( 
.A(n_1908),
.B(n_1713),
.Y(n_2361)
);

AOI22xp33_ASAP7_75t_L g2362 ( 
.A1(n_1959),
.A2(n_1012),
.B1(n_1553),
.B2(n_1713),
.Y(n_2362)
);

NAND2xp5_ASAP7_75t_SL g2363 ( 
.A(n_1806),
.B(n_1428),
.Y(n_2363)
);

AND2x4_ASAP7_75t_L g2364 ( 
.A(n_1921),
.B(n_1615),
.Y(n_2364)
);

INVxp67_ASAP7_75t_L g2365 ( 
.A(n_2042),
.Y(n_2365)
);

INVx2_ASAP7_75t_L g2366 ( 
.A(n_1931),
.Y(n_2366)
);

NAND2xp33_ASAP7_75t_SL g2367 ( 
.A(n_1782),
.B(n_1599),
.Y(n_2367)
);

INVx1_ASAP7_75t_L g2368 ( 
.A(n_2013),
.Y(n_2368)
);

BUFx6f_ASAP7_75t_L g2369 ( 
.A(n_1763),
.Y(n_2369)
);

INVx2_ASAP7_75t_L g2370 ( 
.A(n_1931),
.Y(n_2370)
);

INVx2_ASAP7_75t_SL g2371 ( 
.A(n_1921),
.Y(n_2371)
);

INVx2_ASAP7_75t_L g2372 ( 
.A(n_1934),
.Y(n_2372)
);

INVx2_ASAP7_75t_L g2373 ( 
.A(n_1934),
.Y(n_2373)
);

OR2x2_ASAP7_75t_L g2374 ( 
.A(n_1849),
.B(n_1389),
.Y(n_2374)
);

INVx8_ASAP7_75t_L g2375 ( 
.A(n_2039),
.Y(n_2375)
);

INVx2_ASAP7_75t_L g2376 ( 
.A(n_1936),
.Y(n_2376)
);

AND2x2_ASAP7_75t_L g2377 ( 
.A(n_1744),
.B(n_1749),
.Y(n_2377)
);

NAND2xp33_ASAP7_75t_SL g2378 ( 
.A(n_2004),
.B(n_1599),
.Y(n_2378)
);

INVx1_ASAP7_75t_L g2379 ( 
.A(n_2019),
.Y(n_2379)
);

INVx5_ASAP7_75t_L g2380 ( 
.A(n_2074),
.Y(n_2380)
);

NAND2xp5_ASAP7_75t_SL g2381 ( 
.A(n_1813),
.B(n_1428),
.Y(n_2381)
);

AND3x1_ASAP7_75t_L g2382 ( 
.A(n_2027),
.B(n_1659),
.C(n_1265),
.Y(n_2382)
);

INVx2_ASAP7_75t_L g2383 ( 
.A(n_1936),
.Y(n_2383)
);

INVx2_ASAP7_75t_L g2384 ( 
.A(n_1938),
.Y(n_2384)
);

XNOR2xp5_ASAP7_75t_L g2385 ( 
.A(n_2006),
.B(n_1137),
.Y(n_2385)
);

INVx2_ASAP7_75t_L g2386 ( 
.A(n_1938),
.Y(n_2386)
);

NOR2xp33_ASAP7_75t_L g2387 ( 
.A(n_1805),
.B(n_1233),
.Y(n_2387)
);

INVx3_ASAP7_75t_L g2388 ( 
.A(n_1839),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_2021),
.Y(n_2389)
);

BUFx6f_ASAP7_75t_L g2390 ( 
.A(n_1763),
.Y(n_2390)
);

NOR2xp33_ASAP7_75t_L g2391 ( 
.A(n_1805),
.B(n_1264),
.Y(n_2391)
);

INVx2_ASAP7_75t_L g2392 ( 
.A(n_1940),
.Y(n_2392)
);

INVx8_ASAP7_75t_L g2393 ( 
.A(n_2039),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_2022),
.Y(n_2394)
);

INVx1_ASAP7_75t_L g2395 ( 
.A(n_2038),
.Y(n_2395)
);

NOR2xp33_ASAP7_75t_L g2396 ( 
.A(n_2057),
.B(n_1264),
.Y(n_2396)
);

NAND2xp5_ASAP7_75t_L g2397 ( 
.A(n_1986),
.B(n_1684),
.Y(n_2397)
);

INVx3_ASAP7_75t_L g2398 ( 
.A(n_1839),
.Y(n_2398)
);

INVx2_ASAP7_75t_L g2399 ( 
.A(n_1940),
.Y(n_2399)
);

INVx1_ASAP7_75t_L g2400 ( 
.A(n_2048),
.Y(n_2400)
);

INVx2_ASAP7_75t_L g2401 ( 
.A(n_1944),
.Y(n_2401)
);

NAND2xp5_ASAP7_75t_SL g2402 ( 
.A(n_1813),
.B(n_1641),
.Y(n_2402)
);

NAND2xp5_ASAP7_75t_SL g2403 ( 
.A(n_1813),
.B(n_1656),
.Y(n_2403)
);

NOR2xp33_ASAP7_75t_L g2404 ( 
.A(n_2059),
.B(n_1332),
.Y(n_2404)
);

BUFx2_ASAP7_75t_L g2405 ( 
.A(n_1845),
.Y(n_2405)
);

OR2x2_ASAP7_75t_L g2406 ( 
.A(n_1845),
.B(n_1489),
.Y(n_2406)
);

INVx2_ASAP7_75t_L g2407 ( 
.A(n_1944),
.Y(n_2407)
);

INVx1_ASAP7_75t_L g2408 ( 
.A(n_2049),
.Y(n_2408)
);

INVx5_ASAP7_75t_L g2409 ( 
.A(n_2074),
.Y(n_2409)
);

BUFx6f_ASAP7_75t_L g2410 ( 
.A(n_1763),
.Y(n_2410)
);

INVx2_ASAP7_75t_L g2411 ( 
.A(n_1946),
.Y(n_2411)
);

NAND3xp33_ASAP7_75t_L g2412 ( 
.A(n_1927),
.B(n_1659),
.C(n_1637),
.Y(n_2412)
);

INVx2_ASAP7_75t_L g2413 ( 
.A(n_1946),
.Y(n_2413)
);

INVx1_ASAP7_75t_L g2414 ( 
.A(n_2052),
.Y(n_2414)
);

BUFx3_ASAP7_75t_L g2415 ( 
.A(n_1834),
.Y(n_2415)
);

BUFx10_ASAP7_75t_L g2416 ( 
.A(n_1814),
.Y(n_2416)
);

INVxp33_ASAP7_75t_L g2417 ( 
.A(n_1980),
.Y(n_2417)
);

HB1xp67_ASAP7_75t_L g2418 ( 
.A(n_1875),
.Y(n_2418)
);

INVx3_ASAP7_75t_L g2419 ( 
.A(n_1846),
.Y(n_2419)
);

INVx2_ASAP7_75t_L g2420 ( 
.A(n_1976),
.Y(n_2420)
);

NAND2xp5_ASAP7_75t_SL g2421 ( 
.A(n_1814),
.B(n_1656),
.Y(n_2421)
);

INVx2_ASAP7_75t_L g2422 ( 
.A(n_1976),
.Y(n_2422)
);

AND2x6_ASAP7_75t_L g2423 ( 
.A(n_1888),
.B(n_1132),
.Y(n_2423)
);

AO21x2_ASAP7_75t_L g2424 ( 
.A1(n_1978),
.A2(n_1698),
.B(n_1681),
.Y(n_2424)
);

INVx1_ASAP7_75t_L g2425 ( 
.A(n_2054),
.Y(n_2425)
);

NAND3xp33_ASAP7_75t_L g2426 ( 
.A(n_2027),
.B(n_1481),
.C(n_1452),
.Y(n_2426)
);

INVx2_ASAP7_75t_SL g2427 ( 
.A(n_1921),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_2056),
.Y(n_2428)
);

NAND2xp5_ASAP7_75t_L g2429 ( 
.A(n_1744),
.B(n_1332),
.Y(n_2429)
);

INVx1_ASAP7_75t_L g2430 ( 
.A(n_2058),
.Y(n_2430)
);

NAND2xp5_ASAP7_75t_L g2431 ( 
.A(n_1749),
.B(n_1217),
.Y(n_2431)
);

NAND2xp5_ASAP7_75t_SL g2432 ( 
.A(n_1814),
.B(n_1662),
.Y(n_2432)
);

INVx1_ASAP7_75t_L g2433 ( 
.A(n_2061),
.Y(n_2433)
);

INVx2_ASAP7_75t_L g2434 ( 
.A(n_1733),
.Y(n_2434)
);

INVx2_ASAP7_75t_L g2435 ( 
.A(n_1733),
.Y(n_2435)
);

CKINVDCx5p33_ASAP7_75t_R g2436 ( 
.A(n_1771),
.Y(n_2436)
);

INVx1_ASAP7_75t_L g2437 ( 
.A(n_2064),
.Y(n_2437)
);

NAND2xp5_ASAP7_75t_SL g2438 ( 
.A(n_1888),
.B(n_1662),
.Y(n_2438)
);

NAND2xp5_ASAP7_75t_L g2439 ( 
.A(n_1901),
.B(n_1220),
.Y(n_2439)
);

INVx1_ASAP7_75t_L g2440 ( 
.A(n_1738),
.Y(n_2440)
);

INVx4_ASAP7_75t_L g2441 ( 
.A(n_1846),
.Y(n_2441)
);

INVx2_ASAP7_75t_L g2442 ( 
.A(n_1738),
.Y(n_2442)
);

INVx2_ASAP7_75t_L g2443 ( 
.A(n_1739),
.Y(n_2443)
);

INVx2_ASAP7_75t_L g2444 ( 
.A(n_1739),
.Y(n_2444)
);

NAND2xp33_ASAP7_75t_L g2445 ( 
.A(n_2039),
.B(n_921),
.Y(n_2445)
);

NAND2xp5_ASAP7_75t_SL g2446 ( 
.A(n_1891),
.B(n_1670),
.Y(n_2446)
);

INVx2_ASAP7_75t_L g2447 ( 
.A(n_1747),
.Y(n_2447)
);

CKINVDCx5p33_ASAP7_75t_R g2448 ( 
.A(n_1771),
.Y(n_2448)
);

OR2x2_ASAP7_75t_L g2449 ( 
.A(n_1875),
.B(n_1545),
.Y(n_2449)
);

INVx1_ASAP7_75t_L g2450 ( 
.A(n_1747),
.Y(n_2450)
);

INVx3_ASAP7_75t_L g2451 ( 
.A(n_1846),
.Y(n_2451)
);

OAI22xp33_ASAP7_75t_L g2452 ( 
.A1(n_2024),
.A2(n_1670),
.B1(n_1708),
.B2(n_1693),
.Y(n_2452)
);

NAND2xp5_ASAP7_75t_SL g2453 ( 
.A(n_1891),
.B(n_1693),
.Y(n_2453)
);

INVx2_ASAP7_75t_L g2454 ( 
.A(n_1748),
.Y(n_2454)
);

INVx1_ASAP7_75t_L g2455 ( 
.A(n_1748),
.Y(n_2455)
);

INVx3_ASAP7_75t_L g2456 ( 
.A(n_1852),
.Y(n_2456)
);

INVx2_ASAP7_75t_L g2457 ( 
.A(n_1983),
.Y(n_2457)
);

INVx1_ASAP7_75t_SL g2458 ( 
.A(n_2042),
.Y(n_2458)
);

NAND2xp33_ASAP7_75t_L g2459 ( 
.A(n_2039),
.B(n_921),
.Y(n_2459)
);

INVx1_ASAP7_75t_L g2460 ( 
.A(n_1783),
.Y(n_2460)
);

NAND2xp5_ASAP7_75t_L g2461 ( 
.A(n_1901),
.B(n_1564),
.Y(n_2461)
);

INVx2_ASAP7_75t_L g2462 ( 
.A(n_1991),
.Y(n_2462)
);

INVx2_ASAP7_75t_L g2463 ( 
.A(n_1991),
.Y(n_2463)
);

INVx2_ASAP7_75t_L g2464 ( 
.A(n_1994),
.Y(n_2464)
);

NAND2xp5_ASAP7_75t_SL g2465 ( 
.A(n_1964),
.B(n_2025),
.Y(n_2465)
);

INVx4_ASAP7_75t_L g2466 ( 
.A(n_1852),
.Y(n_2466)
);

INVx2_ASAP7_75t_L g2467 ( 
.A(n_1994),
.Y(n_2467)
);

AND2x2_ASAP7_75t_L g2468 ( 
.A(n_2184),
.B(n_2230),
.Y(n_2468)
);

CKINVDCx5p33_ASAP7_75t_R g2469 ( 
.A(n_2277),
.Y(n_2469)
);

BUFx2_ASAP7_75t_L g2470 ( 
.A(n_2320),
.Y(n_2470)
);

OR2x2_ASAP7_75t_L g2471 ( 
.A(n_2458),
.B(n_1811),
.Y(n_2471)
);

INVx2_ASAP7_75t_L g2472 ( 
.A(n_2434),
.Y(n_2472)
);

NOR2xp33_ASAP7_75t_L g2473 ( 
.A(n_2162),
.B(n_2047),
.Y(n_2473)
);

INVx1_ASAP7_75t_L g2474 ( 
.A(n_2096),
.Y(n_2474)
);

INVx1_ASAP7_75t_L g2475 ( 
.A(n_2097),
.Y(n_2475)
);

INVx2_ASAP7_75t_L g2476 ( 
.A(n_2434),
.Y(n_2476)
);

NOR2xp33_ASAP7_75t_SL g2477 ( 
.A(n_2153),
.B(n_1847),
.Y(n_2477)
);

NAND2xp5_ASAP7_75t_L g2478 ( 
.A(n_2123),
.B(n_2039),
.Y(n_2478)
);

INVx1_ASAP7_75t_L g2479 ( 
.A(n_2101),
.Y(n_2479)
);

XNOR2xp5_ASAP7_75t_L g2480 ( 
.A(n_2385),
.B(n_1297),
.Y(n_2480)
);

INVxp33_ASAP7_75t_L g2481 ( 
.A(n_2316),
.Y(n_2481)
);

INVx2_ASAP7_75t_L g2482 ( 
.A(n_2435),
.Y(n_2482)
);

INVx1_ASAP7_75t_L g2483 ( 
.A(n_2103),
.Y(n_2483)
);

CKINVDCx5p33_ASAP7_75t_R g2484 ( 
.A(n_2277),
.Y(n_2484)
);

INVxp67_ASAP7_75t_L g2485 ( 
.A(n_2142),
.Y(n_2485)
);

CKINVDCx20_ASAP7_75t_R g2486 ( 
.A(n_2290),
.Y(n_2486)
);

INVx1_ASAP7_75t_L g2487 ( 
.A(n_2107),
.Y(n_2487)
);

INVx1_ASAP7_75t_L g2488 ( 
.A(n_2111),
.Y(n_2488)
);

INVx1_ASAP7_75t_L g2489 ( 
.A(n_2114),
.Y(n_2489)
);

INVx3_ASAP7_75t_L g2490 ( 
.A(n_2375),
.Y(n_2490)
);

INVx1_ASAP7_75t_L g2491 ( 
.A(n_2115),
.Y(n_2491)
);

CKINVDCx5p33_ASAP7_75t_R g2492 ( 
.A(n_2358),
.Y(n_2492)
);

INVx1_ASAP7_75t_L g2493 ( 
.A(n_2125),
.Y(n_2493)
);

INVx4_ASAP7_75t_SL g2494 ( 
.A(n_2109),
.Y(n_2494)
);

INVx1_ASAP7_75t_L g2495 ( 
.A(n_2129),
.Y(n_2495)
);

AND2x2_ASAP7_75t_SL g2496 ( 
.A(n_2312),
.B(n_1545),
.Y(n_2496)
);

BUFx6f_ASAP7_75t_L g2497 ( 
.A(n_2138),
.Y(n_2497)
);

XOR2xp5_ASAP7_75t_L g2498 ( 
.A(n_2436),
.B(n_1815),
.Y(n_2498)
);

INVx2_ASAP7_75t_L g2499 ( 
.A(n_2435),
.Y(n_2499)
);

INVx1_ASAP7_75t_L g2500 ( 
.A(n_2139),
.Y(n_2500)
);

INVxp33_ASAP7_75t_L g2501 ( 
.A(n_2316),
.Y(n_2501)
);

OR2x2_ASAP7_75t_L g2502 ( 
.A(n_2142),
.B(n_2320),
.Y(n_2502)
);

NAND2xp5_ASAP7_75t_SL g2503 ( 
.A(n_2127),
.B(n_2047),
.Y(n_2503)
);

INVx1_ASAP7_75t_L g2504 ( 
.A(n_2145),
.Y(n_2504)
);

INVx1_ASAP7_75t_L g2505 ( 
.A(n_2167),
.Y(n_2505)
);

XOR2xp5_ASAP7_75t_L g2506 ( 
.A(n_2436),
.B(n_2032),
.Y(n_2506)
);

INVx2_ASAP7_75t_SL g2507 ( 
.A(n_2339),
.Y(n_2507)
);

XNOR2x2_ASAP7_75t_L g2508 ( 
.A(n_2385),
.B(n_1385),
.Y(n_2508)
);

INVx1_ASAP7_75t_L g2509 ( 
.A(n_2174),
.Y(n_2509)
);

CKINVDCx20_ASAP7_75t_R g2510 ( 
.A(n_2290),
.Y(n_2510)
);

INVx1_ASAP7_75t_L g2511 ( 
.A(n_2177),
.Y(n_2511)
);

NOR2xp33_ASAP7_75t_L g2512 ( 
.A(n_2169),
.B(n_2084),
.Y(n_2512)
);

BUFx6f_ASAP7_75t_L g2513 ( 
.A(n_2138),
.Y(n_2513)
);

INVx1_ASAP7_75t_L g2514 ( 
.A(n_2186),
.Y(n_2514)
);

NAND2x1p5_ASAP7_75t_L g2515 ( 
.A(n_2336),
.B(n_2347),
.Y(n_2515)
);

INVx1_ASAP7_75t_L g2516 ( 
.A(n_2187),
.Y(n_2516)
);

INVx1_ASAP7_75t_L g2517 ( 
.A(n_2199),
.Y(n_2517)
);

CKINVDCx5p33_ASAP7_75t_R g2518 ( 
.A(n_2358),
.Y(n_2518)
);

INVx1_ASAP7_75t_L g2519 ( 
.A(n_2203),
.Y(n_2519)
);

OR2x2_ASAP7_75t_L g2520 ( 
.A(n_2339),
.B(n_2084),
.Y(n_2520)
);

AOI21x1_ASAP7_75t_L g2521 ( 
.A1(n_2280),
.A2(n_2010),
.B(n_1995),
.Y(n_2521)
);

OR2x6_ASAP7_75t_L g2522 ( 
.A(n_2153),
.B(n_1890),
.Y(n_2522)
);

CKINVDCx20_ASAP7_75t_R g2523 ( 
.A(n_2249),
.Y(n_2523)
);

OR2x2_ASAP7_75t_L g2524 ( 
.A(n_2405),
.B(n_2037),
.Y(n_2524)
);

AOI21xp5_ASAP7_75t_L g2525 ( 
.A1(n_2118),
.A2(n_2029),
.B(n_2020),
.Y(n_2525)
);

INVx1_ASAP7_75t_L g2526 ( 
.A(n_2216),
.Y(n_2526)
);

INVx1_ASAP7_75t_L g2527 ( 
.A(n_2218),
.Y(n_2527)
);

INVx1_ASAP7_75t_L g2528 ( 
.A(n_2220),
.Y(n_2528)
);

INVxp33_ASAP7_75t_L g2529 ( 
.A(n_2374),
.Y(n_2529)
);

NOR2xp33_ASAP7_75t_L g2530 ( 
.A(n_2156),
.B(n_1885),
.Y(n_2530)
);

INVx1_ASAP7_75t_L g2531 ( 
.A(n_2224),
.Y(n_2531)
);

NOR2xp67_ASAP7_75t_L g2532 ( 
.A(n_2249),
.B(n_1564),
.Y(n_2532)
);

INVx2_ASAP7_75t_L g2533 ( 
.A(n_2442),
.Y(n_2533)
);

INVx2_ASAP7_75t_L g2534 ( 
.A(n_2442),
.Y(n_2534)
);

NOR2xp33_ASAP7_75t_L g2535 ( 
.A(n_2143),
.B(n_2144),
.Y(n_2535)
);

INVx2_ASAP7_75t_L g2536 ( 
.A(n_2443),
.Y(n_2536)
);

INVx1_ASAP7_75t_L g2537 ( 
.A(n_2227),
.Y(n_2537)
);

INVxp67_ASAP7_75t_SL g2538 ( 
.A(n_2340),
.Y(n_2538)
);

CKINVDCx5p33_ASAP7_75t_R g2539 ( 
.A(n_2198),
.Y(n_2539)
);

INVx1_ASAP7_75t_L g2540 ( 
.A(n_2231),
.Y(n_2540)
);

NOR2xp33_ASAP7_75t_L g2541 ( 
.A(n_2106),
.B(n_1315),
.Y(n_2541)
);

INVx1_ASAP7_75t_L g2542 ( 
.A(n_2237),
.Y(n_2542)
);

NAND2xp5_ASAP7_75t_L g2543 ( 
.A(n_2324),
.B(n_2039),
.Y(n_2543)
);

INVx1_ASAP7_75t_L g2544 ( 
.A(n_2239),
.Y(n_2544)
);

INVx1_ASAP7_75t_L g2545 ( 
.A(n_2460),
.Y(n_2545)
);

NOR2xp33_ASAP7_75t_L g2546 ( 
.A(n_2182),
.B(n_1893),
.Y(n_2546)
);

INVx1_ASAP7_75t_L g2547 ( 
.A(n_2377),
.Y(n_2547)
);

AND2x4_ASAP7_75t_L g2548 ( 
.A(n_2289),
.B(n_2336),
.Y(n_2548)
);

INVxp33_ASAP7_75t_L g2549 ( 
.A(n_2374),
.Y(n_2549)
);

INVx2_ASAP7_75t_L g2550 ( 
.A(n_2443),
.Y(n_2550)
);

AND2x2_ASAP7_75t_L g2551 ( 
.A(n_2140),
.B(n_2037),
.Y(n_2551)
);

INVx1_ASAP7_75t_L g2552 ( 
.A(n_2377),
.Y(n_2552)
);

XOR2xp5_ASAP7_75t_L g2553 ( 
.A(n_2448),
.B(n_2032),
.Y(n_2553)
);

INVx1_ASAP7_75t_SL g2554 ( 
.A(n_2405),
.Y(n_2554)
);

NAND2xp5_ASAP7_75t_L g2555 ( 
.A(n_2397),
.B(n_2053),
.Y(n_2555)
);

INVx1_ASAP7_75t_L g2556 ( 
.A(n_2311),
.Y(n_2556)
);

AND2x2_ASAP7_75t_SL g2557 ( 
.A(n_2319),
.B(n_1804),
.Y(n_2557)
);

INVx2_ASAP7_75t_SL g2558 ( 
.A(n_2140),
.Y(n_2558)
);

INVx1_ASAP7_75t_L g2559 ( 
.A(n_2311),
.Y(n_2559)
);

INVx1_ASAP7_75t_L g2560 ( 
.A(n_2151),
.Y(n_2560)
);

INVx1_ASAP7_75t_L g2561 ( 
.A(n_2163),
.Y(n_2561)
);

NOR2xp33_ASAP7_75t_L g2562 ( 
.A(n_2189),
.B(n_1907),
.Y(n_2562)
);

INVx1_ASAP7_75t_L g2563 ( 
.A(n_2165),
.Y(n_2563)
);

INVx2_ASAP7_75t_L g2564 ( 
.A(n_2444),
.Y(n_2564)
);

CKINVDCx5p33_ASAP7_75t_R g2565 ( 
.A(n_2198),
.Y(n_2565)
);

OR2x2_ASAP7_75t_L g2566 ( 
.A(n_2309),
.B(n_2037),
.Y(n_2566)
);

NOR2xp33_ASAP7_75t_L g2567 ( 
.A(n_2197),
.B(n_1929),
.Y(n_2567)
);

INVx1_ASAP7_75t_L g2568 ( 
.A(n_2235),
.Y(n_2568)
);

AND2x4_ASAP7_75t_L g2569 ( 
.A(n_2289),
.B(n_1964),
.Y(n_2569)
);

XOR2xp5_ASAP7_75t_L g2570 ( 
.A(n_2448),
.B(n_1315),
.Y(n_2570)
);

NAND2xp5_ASAP7_75t_L g2571 ( 
.A(n_2210),
.B(n_2053),
.Y(n_2571)
);

NOR2xp33_ASAP7_75t_L g2572 ( 
.A(n_2160),
.B(n_2076),
.Y(n_2572)
);

INVx2_ASAP7_75t_L g2573 ( 
.A(n_2444),
.Y(n_2573)
);

XOR2x2_ASAP7_75t_L g2574 ( 
.A(n_2426),
.B(n_1879),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_2242),
.Y(n_2575)
);

NAND2xp5_ASAP7_75t_L g2576 ( 
.A(n_2217),
.B(n_2053),
.Y(n_2576)
);

XOR2xp5_ASAP7_75t_L g2577 ( 
.A(n_2342),
.B(n_1338),
.Y(n_2577)
);

NOR2xp33_ASAP7_75t_L g2578 ( 
.A(n_2108),
.B(n_2087),
.Y(n_2578)
);

INVx1_ASAP7_75t_L g2579 ( 
.A(n_2246),
.Y(n_2579)
);

INVx1_ASAP7_75t_L g2580 ( 
.A(n_2250),
.Y(n_2580)
);

INVx1_ASAP7_75t_L g2581 ( 
.A(n_2252),
.Y(n_2581)
);

INVx2_ASAP7_75t_L g2582 ( 
.A(n_2447),
.Y(n_2582)
);

INVx1_ASAP7_75t_L g2583 ( 
.A(n_2254),
.Y(n_2583)
);

XOR2xp5_ASAP7_75t_L g2584 ( 
.A(n_2342),
.B(n_1338),
.Y(n_2584)
);

CKINVDCx5p33_ASAP7_75t_R g2585 ( 
.A(n_2204),
.Y(n_2585)
);

NAND2x1p5_ASAP7_75t_L g2586 ( 
.A(n_2347),
.B(n_1852),
.Y(n_2586)
);

INVx2_ASAP7_75t_SL g2587 ( 
.A(n_2449),
.Y(n_2587)
);

NOR2xp33_ASAP7_75t_L g2588 ( 
.A(n_2155),
.B(n_2088),
.Y(n_2588)
);

INVx1_ASAP7_75t_L g2589 ( 
.A(n_2258),
.Y(n_2589)
);

INVx1_ASAP7_75t_L g2590 ( 
.A(n_2263),
.Y(n_2590)
);

INVx1_ASAP7_75t_L g2591 ( 
.A(n_2267),
.Y(n_2591)
);

OR2x6_ASAP7_75t_L g2592 ( 
.A(n_2153),
.B(n_1708),
.Y(n_2592)
);

NOR2xp67_ASAP7_75t_L g2593 ( 
.A(n_2309),
.B(n_1588),
.Y(n_2593)
);

INVx1_ASAP7_75t_L g2594 ( 
.A(n_2268),
.Y(n_2594)
);

INVx1_ASAP7_75t_L g2595 ( 
.A(n_2273),
.Y(n_2595)
);

INVx1_ASAP7_75t_L g2596 ( 
.A(n_2274),
.Y(n_2596)
);

INVx1_ASAP7_75t_L g2597 ( 
.A(n_2275),
.Y(n_2597)
);

NOR2xp33_ASAP7_75t_L g2598 ( 
.A(n_2429),
.B(n_2090),
.Y(n_2598)
);

NAND2x1p5_ASAP7_75t_L g2599 ( 
.A(n_2371),
.B(n_1895),
.Y(n_2599)
);

AND2x2_ASAP7_75t_L g2600 ( 
.A(n_2257),
.B(n_2041),
.Y(n_2600)
);

AND2x2_ASAP7_75t_L g2601 ( 
.A(n_2257),
.B(n_2041),
.Y(n_2601)
);

NOR2xp33_ASAP7_75t_L g2602 ( 
.A(n_2172),
.B(n_2091),
.Y(n_2602)
);

NOR2xp33_ASAP7_75t_L g2603 ( 
.A(n_2461),
.B(n_2093),
.Y(n_2603)
);

AND2x2_ASAP7_75t_L g2604 ( 
.A(n_2260),
.B(n_2041),
.Y(n_2604)
);

NAND2x1p5_ASAP7_75t_L g2605 ( 
.A(n_2371),
.B(n_1895),
.Y(n_2605)
);

NOR2xp33_ASAP7_75t_L g2606 ( 
.A(n_2209),
.B(n_2325),
.Y(n_2606)
);

INVx1_ASAP7_75t_L g2607 ( 
.A(n_2276),
.Y(n_2607)
);

INVx1_ASAP7_75t_L g2608 ( 
.A(n_2278),
.Y(n_2608)
);

INVx1_ASAP7_75t_L g2609 ( 
.A(n_2295),
.Y(n_2609)
);

AND2x6_ASAP7_75t_L g2610 ( 
.A(n_2153),
.B(n_2045),
.Y(n_2610)
);

AND2x4_ASAP7_75t_L g2611 ( 
.A(n_2289),
.B(n_1964),
.Y(n_2611)
);

INVx1_ASAP7_75t_L g2612 ( 
.A(n_2300),
.Y(n_2612)
);

NAND2xp5_ASAP7_75t_L g2613 ( 
.A(n_2222),
.B(n_2053),
.Y(n_2613)
);

INVx1_ASAP7_75t_L g2614 ( 
.A(n_2308),
.Y(n_2614)
);

CKINVDCx5p33_ASAP7_75t_R g2615 ( 
.A(n_2204),
.Y(n_2615)
);

INVx1_ASAP7_75t_L g2616 ( 
.A(n_2323),
.Y(n_2616)
);

CKINVDCx14_ASAP7_75t_R g2617 ( 
.A(n_2406),
.Y(n_2617)
);

CKINVDCx20_ASAP7_75t_R g2618 ( 
.A(n_2134),
.Y(n_2618)
);

INVx1_ASAP7_75t_L g2619 ( 
.A(n_2331),
.Y(n_2619)
);

INVx1_ASAP7_75t_L g2620 ( 
.A(n_2334),
.Y(n_2620)
);

INVx1_ASAP7_75t_L g2621 ( 
.A(n_2341),
.Y(n_2621)
);

INVx1_ASAP7_75t_L g2622 ( 
.A(n_2344),
.Y(n_2622)
);

INVx1_ASAP7_75t_L g2623 ( 
.A(n_2359),
.Y(n_2623)
);

BUFx3_ASAP7_75t_L g2624 ( 
.A(n_2134),
.Y(n_2624)
);

INVx1_ASAP7_75t_L g2625 ( 
.A(n_2368),
.Y(n_2625)
);

BUFx4f_ASAP7_75t_L g2626 ( 
.A(n_2449),
.Y(n_2626)
);

AND2x4_ASAP7_75t_L g2627 ( 
.A(n_2427),
.B(n_2025),
.Y(n_2627)
);

AND2x2_ASAP7_75t_L g2628 ( 
.A(n_2260),
.B(n_2045),
.Y(n_2628)
);

NOR2xp33_ASAP7_75t_L g2629 ( 
.A(n_2350),
.B(n_2094),
.Y(n_2629)
);

XOR2xp5_ASAP7_75t_L g2630 ( 
.A(n_2146),
.B(n_1386),
.Y(n_2630)
);

XNOR2xp5_ASAP7_75t_L g2631 ( 
.A(n_2351),
.B(n_1386),
.Y(n_2631)
);

INVx2_ASAP7_75t_L g2632 ( 
.A(n_2447),
.Y(n_2632)
);

INVx2_ASAP7_75t_L g2633 ( 
.A(n_2454),
.Y(n_2633)
);

INVx2_ASAP7_75t_SL g2634 ( 
.A(n_2418),
.Y(n_2634)
);

INVx1_ASAP7_75t_L g2635 ( 
.A(n_2379),
.Y(n_2635)
);

INVx4_ASAP7_75t_L g2636 ( 
.A(n_2375),
.Y(n_2636)
);

NAND2xp33_ASAP7_75t_SL g2637 ( 
.A(n_2360),
.B(n_2192),
.Y(n_2637)
);

NOR2xp33_ASAP7_75t_L g2638 ( 
.A(n_2200),
.B(n_2045),
.Y(n_2638)
);

XOR2xp5_ASAP7_75t_L g2639 ( 
.A(n_2146),
.B(n_1154),
.Y(n_2639)
);

OR2x2_ASAP7_75t_L g2640 ( 
.A(n_2439),
.B(n_2431),
.Y(n_2640)
);

INVx1_ASAP7_75t_L g2641 ( 
.A(n_2389),
.Y(n_2641)
);

INVx2_ASAP7_75t_L g2642 ( 
.A(n_2454),
.Y(n_2642)
);

INVx1_ASAP7_75t_L g2643 ( 
.A(n_2394),
.Y(n_2643)
);

INVx1_ASAP7_75t_L g2644 ( 
.A(n_2395),
.Y(n_2644)
);

CKINVDCx20_ASAP7_75t_R g2645 ( 
.A(n_2134),
.Y(n_2645)
);

NAND2x1p5_ASAP7_75t_L g2646 ( 
.A(n_2427),
.B(n_1895),
.Y(n_2646)
);

CKINVDCx20_ASAP7_75t_R g2647 ( 
.A(n_2164),
.Y(n_2647)
);

XOR2x2_ASAP7_75t_L g2648 ( 
.A(n_2266),
.B(n_2406),
.Y(n_2648)
);

INVx1_ASAP7_75t_L g2649 ( 
.A(n_2400),
.Y(n_2649)
);

CKINVDCx5p33_ASAP7_75t_R g2650 ( 
.A(n_2164),
.Y(n_2650)
);

INVx2_ASAP7_75t_L g2651 ( 
.A(n_2099),
.Y(n_2651)
);

CKINVDCx20_ASAP7_75t_R g2652 ( 
.A(n_2164),
.Y(n_2652)
);

INVxp33_ASAP7_75t_L g2653 ( 
.A(n_2253),
.Y(n_2653)
);

INVx1_ASAP7_75t_L g2654 ( 
.A(n_2408),
.Y(n_2654)
);

INVx1_ASAP7_75t_L g2655 ( 
.A(n_2414),
.Y(n_2655)
);

INVx1_ASAP7_75t_L g2656 ( 
.A(n_2425),
.Y(n_2656)
);

INVx1_ASAP7_75t_L g2657 ( 
.A(n_2428),
.Y(n_2657)
);

INVx1_ASAP7_75t_L g2658 ( 
.A(n_2430),
.Y(n_2658)
);

BUFx3_ASAP7_75t_L g2659 ( 
.A(n_2175),
.Y(n_2659)
);

INVx1_ASAP7_75t_L g2660 ( 
.A(n_2433),
.Y(n_2660)
);

INVxp67_ASAP7_75t_L g2661 ( 
.A(n_2181),
.Y(n_2661)
);

INVx1_ASAP7_75t_L g2662 ( 
.A(n_2437),
.Y(n_2662)
);

INVx1_ASAP7_75t_L g2663 ( 
.A(n_2181),
.Y(n_2663)
);

INVx1_ASAP7_75t_L g2664 ( 
.A(n_2191),
.Y(n_2664)
);

NOR2xp67_ASAP7_75t_L g2665 ( 
.A(n_2365),
.B(n_1588),
.Y(n_2665)
);

INVx2_ASAP7_75t_L g2666 ( 
.A(n_2099),
.Y(n_2666)
);

INVx1_ASAP7_75t_L g2667 ( 
.A(n_2191),
.Y(n_2667)
);

CKINVDCx16_ASAP7_75t_R g2668 ( 
.A(n_2175),
.Y(n_2668)
);

XNOR2xp5_ASAP7_75t_L g2669 ( 
.A(n_2351),
.B(n_1155),
.Y(n_2669)
);

INVx1_ASAP7_75t_L g2670 ( 
.A(n_2244),
.Y(n_2670)
);

INVx1_ASAP7_75t_L g2671 ( 
.A(n_2244),
.Y(n_2671)
);

INVx1_ASAP7_75t_L g2672 ( 
.A(n_2465),
.Y(n_2672)
);

INVx1_ASAP7_75t_L g2673 ( 
.A(n_2440),
.Y(n_2673)
);

AOI21xp5_ASAP7_75t_L g2674 ( 
.A1(n_2118),
.A2(n_2345),
.B(n_2340),
.Y(n_2674)
);

INVx1_ASAP7_75t_L g2675 ( 
.A(n_2450),
.Y(n_2675)
);

INVx1_ASAP7_75t_L g2676 ( 
.A(n_2455),
.Y(n_2676)
);

NOR2xp33_ASAP7_75t_L g2677 ( 
.A(n_2135),
.B(n_1876),
.Y(n_2677)
);

INVx1_ASAP7_75t_L g2678 ( 
.A(n_2116),
.Y(n_2678)
);

INVx4_ASAP7_75t_L g2679 ( 
.A(n_2375),
.Y(n_2679)
);

INVx2_ASAP7_75t_L g2680 ( 
.A(n_2116),
.Y(n_2680)
);

INVx1_ASAP7_75t_L g2681 ( 
.A(n_2117),
.Y(n_2681)
);

NOR2xp33_ASAP7_75t_SL g2682 ( 
.A(n_2185),
.B(n_1990),
.Y(n_2682)
);

INVx1_ASAP7_75t_L g2683 ( 
.A(n_2117),
.Y(n_2683)
);

INVx1_ASAP7_75t_L g2684 ( 
.A(n_2121),
.Y(n_2684)
);

INVx1_ASAP7_75t_L g2685 ( 
.A(n_2121),
.Y(n_2685)
);

NAND2xp33_ASAP7_75t_R g2686 ( 
.A(n_2387),
.B(n_1700),
.Y(n_2686)
);

CKINVDCx5p33_ASAP7_75t_R g2687 ( 
.A(n_2175),
.Y(n_2687)
);

INVx2_ASAP7_75t_SL g2688 ( 
.A(n_2416),
.Y(n_2688)
);

INVxp33_ASAP7_75t_L g2689 ( 
.A(n_2256),
.Y(n_2689)
);

INVx1_ASAP7_75t_L g2690 ( 
.A(n_2124),
.Y(n_2690)
);

CKINVDCx5p33_ASAP7_75t_R g2691 ( 
.A(n_2326),
.Y(n_2691)
);

NOR2xp33_ASAP7_75t_L g2692 ( 
.A(n_2098),
.B(n_1880),
.Y(n_2692)
);

INVx1_ASAP7_75t_L g2693 ( 
.A(n_2124),
.Y(n_2693)
);

NOR2xp33_ASAP7_75t_L g2694 ( 
.A(n_2119),
.B(n_1881),
.Y(n_2694)
);

INVx1_ASAP7_75t_L g2695 ( 
.A(n_2128),
.Y(n_2695)
);

NOR2xp67_ASAP7_75t_L g2696 ( 
.A(n_2391),
.B(n_1595),
.Y(n_2696)
);

AND2x2_ASAP7_75t_L g2697 ( 
.A(n_2314),
.B(n_1966),
.Y(n_2697)
);

INVx1_ASAP7_75t_L g2698 ( 
.A(n_2128),
.Y(n_2698)
);

INVx2_ASAP7_75t_L g2699 ( 
.A(n_2130),
.Y(n_2699)
);

AND2x2_ASAP7_75t_L g2700 ( 
.A(n_2314),
.B(n_1966),
.Y(n_2700)
);

NAND2xp5_ASAP7_75t_L g2701 ( 
.A(n_2166),
.B(n_2053),
.Y(n_2701)
);

INVx1_ASAP7_75t_L g2702 ( 
.A(n_2130),
.Y(n_2702)
);

BUFx6f_ASAP7_75t_L g2703 ( 
.A(n_2138),
.Y(n_2703)
);

AND2x2_ASAP7_75t_L g2704 ( 
.A(n_2265),
.B(n_1973),
.Y(n_2704)
);

NAND2xp33_ASAP7_75t_R g2705 ( 
.A(n_2361),
.B(n_1700),
.Y(n_2705)
);

INVx1_ASAP7_75t_L g2706 ( 
.A(n_2131),
.Y(n_2706)
);

INVx2_ASAP7_75t_SL g2707 ( 
.A(n_2416),
.Y(n_2707)
);

AND2x2_ASAP7_75t_L g2708 ( 
.A(n_2265),
.B(n_1973),
.Y(n_2708)
);

INVx2_ASAP7_75t_L g2709 ( 
.A(n_2131),
.Y(n_2709)
);

INVx1_ASAP7_75t_L g2710 ( 
.A(n_2132),
.Y(n_2710)
);

INVx1_ASAP7_75t_L g2711 ( 
.A(n_2132),
.Y(n_2711)
);

INVx3_ASAP7_75t_L g2712 ( 
.A(n_2375),
.Y(n_2712)
);

OR2x2_ASAP7_75t_SL g2713 ( 
.A(n_2269),
.B(n_1905),
.Y(n_2713)
);

INVx1_ASAP7_75t_L g2714 ( 
.A(n_2136),
.Y(n_2714)
);

INVx1_ASAP7_75t_L g2715 ( 
.A(n_2136),
.Y(n_2715)
);

NOR2xp33_ASAP7_75t_SL g2716 ( 
.A(n_2185),
.B(n_1990),
.Y(n_2716)
);

INVx1_ASAP7_75t_L g2717 ( 
.A(n_2137),
.Y(n_2717)
);

AOI21xp5_ASAP7_75t_L g2718 ( 
.A1(n_2345),
.A2(n_2029),
.B(n_2020),
.Y(n_2718)
);

OAI21xp5_ASAP7_75t_L g2719 ( 
.A1(n_2318),
.A2(n_2029),
.B(n_2020),
.Y(n_2719)
);

NOR2xp33_ASAP7_75t_L g2720 ( 
.A(n_2211),
.B(n_1882),
.Y(n_2720)
);

NOR2xp33_ASAP7_75t_L g2721 ( 
.A(n_2234),
.B(n_2337),
.Y(n_2721)
);

INVx1_ASAP7_75t_L g2722 ( 
.A(n_2137),
.Y(n_2722)
);

NOR2xp33_ASAP7_75t_L g2723 ( 
.A(n_2343),
.B(n_1883),
.Y(n_2723)
);

INVx2_ASAP7_75t_L g2724 ( 
.A(n_2147),
.Y(n_2724)
);

INVx2_ASAP7_75t_L g2725 ( 
.A(n_2147),
.Y(n_2725)
);

XOR2xp5_ASAP7_75t_L g2726 ( 
.A(n_2326),
.B(n_1189),
.Y(n_2726)
);

NOR2xp33_ASAP7_75t_SL g2727 ( 
.A(n_2185),
.B(n_2205),
.Y(n_2727)
);

INVx1_ASAP7_75t_L g2728 ( 
.A(n_2148),
.Y(n_2728)
);

AND2x4_ASAP7_75t_L g2729 ( 
.A(n_2361),
.B(n_2025),
.Y(n_2729)
);

INVxp67_ASAP7_75t_SL g2730 ( 
.A(n_2315),
.Y(n_2730)
);

NAND2xp33_ASAP7_75t_R g2731 ( 
.A(n_2361),
.B(n_2396),
.Y(n_2731)
);

INVx1_ASAP7_75t_L g2732 ( 
.A(n_2148),
.Y(n_2732)
);

BUFx3_ASAP7_75t_L g2733 ( 
.A(n_2208),
.Y(n_2733)
);

INVx1_ASAP7_75t_L g2734 ( 
.A(n_2149),
.Y(n_2734)
);

AND2x2_ASAP7_75t_L g2735 ( 
.A(n_2287),
.B(n_1982),
.Y(n_2735)
);

XOR2xp5_ASAP7_75t_L g2736 ( 
.A(n_2161),
.B(n_1189),
.Y(n_2736)
);

INVx1_ASAP7_75t_L g2737 ( 
.A(n_2149),
.Y(n_2737)
);

INVx1_ASAP7_75t_L g2738 ( 
.A(n_2152),
.Y(n_2738)
);

BUFx3_ASAP7_75t_L g2739 ( 
.A(n_2208),
.Y(n_2739)
);

INVx1_ASAP7_75t_L g2740 ( 
.A(n_2152),
.Y(n_2740)
);

AOI21x1_ASAP7_75t_L g2741 ( 
.A1(n_2280),
.A2(n_2226),
.B(n_2102),
.Y(n_2741)
);

INVx1_ASAP7_75t_L g2742 ( 
.A(n_2154),
.Y(n_2742)
);

INVx1_ASAP7_75t_L g2743 ( 
.A(n_2154),
.Y(n_2743)
);

INVx1_ASAP7_75t_L g2744 ( 
.A(n_2158),
.Y(n_2744)
);

AND2x6_ASAP7_75t_L g2745 ( 
.A(n_2185),
.B(n_1982),
.Y(n_2745)
);

AND2x6_ASAP7_75t_L g2746 ( 
.A(n_2205),
.B(n_1998),
.Y(n_2746)
);

AND2x2_ASAP7_75t_L g2747 ( 
.A(n_2287),
.B(n_1998),
.Y(n_2747)
);

XOR2xp5_ASAP7_75t_L g2748 ( 
.A(n_2161),
.B(n_1204),
.Y(n_2748)
);

AND2x2_ASAP7_75t_L g2749 ( 
.A(n_2404),
.B(n_2007),
.Y(n_2749)
);

INVx1_ASAP7_75t_L g2750 ( 
.A(n_2158),
.Y(n_2750)
);

INVx2_ASAP7_75t_L g2751 ( 
.A(n_2159),
.Y(n_2751)
);

CKINVDCx20_ASAP7_75t_R g2752 ( 
.A(n_2378),
.Y(n_2752)
);

AND2x6_ASAP7_75t_L g2753 ( 
.A(n_2205),
.B(n_2007),
.Y(n_2753)
);

INVxp67_ASAP7_75t_L g2754 ( 
.A(n_2214),
.Y(n_2754)
);

INVx1_ASAP7_75t_L g2755 ( 
.A(n_2159),
.Y(n_2755)
);

INVx1_ASAP7_75t_L g2756 ( 
.A(n_2171),
.Y(n_2756)
);

XNOR2xp5_ASAP7_75t_L g2757 ( 
.A(n_2452),
.B(n_1204),
.Y(n_2757)
);

AND2x2_ASAP7_75t_L g2758 ( 
.A(n_2100),
.B(n_2012),
.Y(n_2758)
);

BUFx6f_ASAP7_75t_L g2759 ( 
.A(n_2138),
.Y(n_2759)
);

CKINVDCx20_ASAP7_75t_R g2760 ( 
.A(n_2378),
.Y(n_2760)
);

OR2x2_ASAP7_75t_L g2761 ( 
.A(n_2417),
.B(n_1965),
.Y(n_2761)
);

CKINVDCx14_ASAP7_75t_R g2762 ( 
.A(n_2208),
.Y(n_2762)
);

NAND2xp5_ASAP7_75t_L g2763 ( 
.A(n_2100),
.B(n_2112),
.Y(n_2763)
);

CKINVDCx20_ASAP7_75t_R g2764 ( 
.A(n_2367),
.Y(n_2764)
);

AND2x2_ASAP7_75t_L g2765 ( 
.A(n_2112),
.B(n_2012),
.Y(n_2765)
);

INVx1_ASAP7_75t_L g2766 ( 
.A(n_2171),
.Y(n_2766)
);

INVx1_ASAP7_75t_L g2767 ( 
.A(n_2173),
.Y(n_2767)
);

NAND2xp5_ASAP7_75t_L g2768 ( 
.A(n_2183),
.B(n_2053),
.Y(n_2768)
);

INVxp33_ASAP7_75t_L g2769 ( 
.A(n_2417),
.Y(n_2769)
);

AND2x2_ASAP7_75t_L g2770 ( 
.A(n_2183),
.B(n_2303),
.Y(n_2770)
);

INVx2_ASAP7_75t_L g2771 ( 
.A(n_2173),
.Y(n_2771)
);

CKINVDCx5p33_ASAP7_75t_R g2772 ( 
.A(n_2367),
.Y(n_2772)
);

INVx1_ASAP7_75t_L g2773 ( 
.A(n_2176),
.Y(n_2773)
);

CKINVDCx20_ASAP7_75t_R g2774 ( 
.A(n_2233),
.Y(n_2774)
);

INVx1_ASAP7_75t_L g2775 ( 
.A(n_2176),
.Y(n_2775)
);

INVx1_ASAP7_75t_L g2776 ( 
.A(n_2179),
.Y(n_2776)
);

INVx1_ASAP7_75t_L g2777 ( 
.A(n_2179),
.Y(n_2777)
);

INVx1_ASAP7_75t_L g2778 ( 
.A(n_2188),
.Y(n_2778)
);

INVx1_ASAP7_75t_L g2779 ( 
.A(n_2188),
.Y(n_2779)
);

NOR2xp33_ASAP7_75t_L g2780 ( 
.A(n_2354),
.B(n_1894),
.Y(n_2780)
);

INVx1_ASAP7_75t_L g2781 ( 
.A(n_2190),
.Y(n_2781)
);

INVx1_ASAP7_75t_L g2782 ( 
.A(n_2190),
.Y(n_2782)
);

INVx1_ASAP7_75t_L g2783 ( 
.A(n_2194),
.Y(n_2783)
);

INVx2_ASAP7_75t_L g2784 ( 
.A(n_2194),
.Y(n_2784)
);

INVx1_ASAP7_75t_L g2785 ( 
.A(n_2201),
.Y(n_2785)
);

BUFx2_ASAP7_75t_L g2786 ( 
.A(n_2423),
.Y(n_2786)
);

INVx2_ASAP7_75t_L g2787 ( 
.A(n_2201),
.Y(n_2787)
);

NAND2xp5_ASAP7_75t_L g2788 ( 
.A(n_2303),
.B(n_1910),
.Y(n_2788)
);

INVx1_ASAP7_75t_L g2789 ( 
.A(n_2206),
.Y(n_2789)
);

INVx1_ASAP7_75t_L g2790 ( 
.A(n_2206),
.Y(n_2790)
);

XOR2x2_ASAP7_75t_L g2791 ( 
.A(n_2438),
.B(n_1469),
.Y(n_2791)
);

AND2x2_ASAP7_75t_L g2792 ( 
.A(n_2302),
.B(n_2033),
.Y(n_2792)
);

AOI21xp5_ASAP7_75t_L g2793 ( 
.A1(n_2315),
.A2(n_2034),
.B(n_1922),
.Y(n_2793)
);

INVx2_ASAP7_75t_L g2794 ( 
.A(n_2221),
.Y(n_2794)
);

INVxp67_ASAP7_75t_L g2795 ( 
.A(n_2215),
.Y(n_2795)
);

INVx1_ASAP7_75t_L g2796 ( 
.A(n_2221),
.Y(n_2796)
);

XOR2xp5_ASAP7_75t_L g2797 ( 
.A(n_2382),
.B(n_1223),
.Y(n_2797)
);

INVx1_ASAP7_75t_L g2798 ( 
.A(n_2223),
.Y(n_2798)
);

INVx1_ASAP7_75t_SL g2799 ( 
.A(n_2416),
.Y(n_2799)
);

NAND2xp5_ASAP7_75t_SL g2800 ( 
.A(n_2352),
.B(n_2033),
.Y(n_2800)
);

AND2x6_ASAP7_75t_L g2801 ( 
.A(n_2205),
.B(n_1910),
.Y(n_2801)
);

NOR2xp33_ASAP7_75t_L g2802 ( 
.A(n_2120),
.B(n_1898),
.Y(n_2802)
);

INVxp33_ASAP7_75t_L g2803 ( 
.A(n_2282),
.Y(n_2803)
);

INVx1_ASAP7_75t_L g2804 ( 
.A(n_2223),
.Y(n_2804)
);

INVx1_ASAP7_75t_L g2805 ( 
.A(n_2225),
.Y(n_2805)
);

INVx1_ASAP7_75t_L g2806 ( 
.A(n_2225),
.Y(n_2806)
);

INVx1_ASAP7_75t_L g2807 ( 
.A(n_2228),
.Y(n_2807)
);

INVx1_ASAP7_75t_L g2808 ( 
.A(n_2228),
.Y(n_2808)
);

NAND2xp5_ASAP7_75t_L g2809 ( 
.A(n_2241),
.B(n_1930),
.Y(n_2809)
);

INVx1_ASAP7_75t_L g2810 ( 
.A(n_2229),
.Y(n_2810)
);

INVx1_ASAP7_75t_L g2811 ( 
.A(n_2229),
.Y(n_2811)
);

INVx1_ASAP7_75t_L g2812 ( 
.A(n_2238),
.Y(n_2812)
);

INVxp67_ASAP7_75t_L g2813 ( 
.A(n_2288),
.Y(n_2813)
);

INVx1_ASAP7_75t_L g2814 ( 
.A(n_2238),
.Y(n_2814)
);

INVx1_ASAP7_75t_L g2815 ( 
.A(n_2240),
.Y(n_2815)
);

INVx1_ASAP7_75t_L g2816 ( 
.A(n_2240),
.Y(n_2816)
);

XNOR2xp5_ASAP7_75t_L g2817 ( 
.A(n_2446),
.B(n_1223),
.Y(n_2817)
);

INVx1_ASAP7_75t_L g2818 ( 
.A(n_2248),
.Y(n_2818)
);

INVx2_ASAP7_75t_L g2819 ( 
.A(n_2248),
.Y(n_2819)
);

INVx2_ASAP7_75t_L g2820 ( 
.A(n_2251),
.Y(n_2820)
);

AND2x2_ASAP7_75t_SL g2821 ( 
.A(n_2362),
.B(n_1971),
.Y(n_2821)
);

AND2x2_ASAP7_75t_L g2822 ( 
.A(n_2291),
.B(n_2033),
.Y(n_2822)
);

INVx1_ASAP7_75t_L g2823 ( 
.A(n_2251),
.Y(n_2823)
);

AND2x2_ASAP7_75t_L g2824 ( 
.A(n_2364),
.B(n_2035),
.Y(n_2824)
);

AND2x2_ASAP7_75t_L g2825 ( 
.A(n_2364),
.B(n_2035),
.Y(n_2825)
);

XNOR2x1_ASAP7_75t_L g2826 ( 
.A(n_2322),
.B(n_1246),
.Y(n_2826)
);

CKINVDCx5p33_ASAP7_75t_R g2827 ( 
.A(n_2233),
.Y(n_2827)
);

OAI22xp33_ASAP7_75t_L g2828 ( 
.A1(n_2535),
.A2(n_1716),
.B1(n_1609),
.B2(n_1610),
.Y(n_2828)
);

OAI22xp33_ASAP7_75t_L g2829 ( 
.A1(n_2535),
.A2(n_1716),
.B1(n_1609),
.B2(n_1620),
.Y(n_2829)
);

INVx1_ASAP7_75t_L g2830 ( 
.A(n_2474),
.Y(n_2830)
);

INVx1_ASAP7_75t_L g2831 ( 
.A(n_2475),
.Y(n_2831)
);

AOI22xp5_ASAP7_75t_L g2832 ( 
.A1(n_2541),
.A2(n_2245),
.B1(n_2168),
.B2(n_1620),
.Y(n_2832)
);

NOR2xp33_ASAP7_75t_L g2833 ( 
.A(n_2653),
.B(n_1246),
.Y(n_2833)
);

NAND2xp5_ASAP7_75t_L g2834 ( 
.A(n_2530),
.B(n_2299),
.Y(n_2834)
);

NAND2xp5_ASAP7_75t_L g2835 ( 
.A(n_2530),
.B(n_2299),
.Y(n_2835)
);

NAND2xp5_ASAP7_75t_L g2836 ( 
.A(n_2568),
.B(n_2299),
.Y(n_2836)
);

INVx2_ASAP7_75t_L g2837 ( 
.A(n_2472),
.Y(n_2837)
);

NAND2xp5_ASAP7_75t_L g2838 ( 
.A(n_2629),
.B(n_2353),
.Y(n_2838)
);

AND2x2_ASAP7_75t_L g2839 ( 
.A(n_2468),
.B(n_2035),
.Y(n_2839)
);

NAND2xp5_ASAP7_75t_L g2840 ( 
.A(n_2629),
.B(n_2353),
.Y(n_2840)
);

NAND2xp5_ASAP7_75t_L g2841 ( 
.A(n_2606),
.B(n_2353),
.Y(n_2841)
);

INVx1_ASAP7_75t_L g2842 ( 
.A(n_2479),
.Y(n_2842)
);

NAND2xp33_ASAP7_75t_L g2843 ( 
.A(n_2478),
.B(n_2168),
.Y(n_2843)
);

NAND2xp5_ASAP7_75t_L g2844 ( 
.A(n_2606),
.B(n_2473),
.Y(n_2844)
);

NAND2xp5_ASAP7_75t_SL g2845 ( 
.A(n_2512),
.B(n_2364),
.Y(n_2845)
);

INVx2_ASAP7_75t_L g2846 ( 
.A(n_2476),
.Y(n_2846)
);

NAND2xp5_ASAP7_75t_L g2847 ( 
.A(n_2473),
.B(n_2105),
.Y(n_2847)
);

INVx1_ASAP7_75t_L g2848 ( 
.A(n_2483),
.Y(n_2848)
);

AOI22xp5_ASAP7_75t_L g2849 ( 
.A1(n_2512),
.A2(n_2245),
.B1(n_1595),
.B2(n_2213),
.Y(n_2849)
);

NOR3xp33_ASAP7_75t_L g2850 ( 
.A(n_2602),
.B(n_2213),
.C(n_2412),
.Y(n_2850)
);

BUFx5_ASAP7_75t_L g2851 ( 
.A(n_2801),
.Y(n_2851)
);

INVx3_ASAP7_75t_L g2852 ( 
.A(n_2636),
.Y(n_2852)
);

INVx2_ASAP7_75t_L g2853 ( 
.A(n_2482),
.Y(n_2853)
);

INVx1_ASAP7_75t_L g2854 ( 
.A(n_2487),
.Y(n_2854)
);

BUFx3_ASAP7_75t_L g2855 ( 
.A(n_2469),
.Y(n_2855)
);

NAND2xp5_ASAP7_75t_L g2856 ( 
.A(n_2572),
.B(n_2105),
.Y(n_2856)
);

NAND2xp5_ASAP7_75t_L g2857 ( 
.A(n_2572),
.B(n_2105),
.Y(n_2857)
);

NAND2xp5_ASAP7_75t_SL g2858 ( 
.A(n_2689),
.B(n_2307),
.Y(n_2858)
);

INVx2_ASAP7_75t_L g2859 ( 
.A(n_2499),
.Y(n_2859)
);

NAND2xp5_ASAP7_75t_SL g2860 ( 
.A(n_2729),
.B(n_2307),
.Y(n_2860)
);

NAND2xp5_ASAP7_75t_L g2861 ( 
.A(n_2598),
.B(n_2602),
.Y(n_2861)
);

INVx1_ASAP7_75t_L g2862 ( 
.A(n_2488),
.Y(n_2862)
);

NOR2xp33_ASAP7_75t_L g2863 ( 
.A(n_2554),
.B(n_1469),
.Y(n_2863)
);

NOR2xp33_ASAP7_75t_L g2864 ( 
.A(n_2554),
.B(n_1531),
.Y(n_2864)
);

AOI22xp33_ASAP7_75t_L g2865 ( 
.A1(n_2508),
.A2(n_2423),
.B1(n_1633),
.B2(n_2357),
.Y(n_2865)
);

NAND2xp5_ASAP7_75t_L g2866 ( 
.A(n_2598),
.B(n_2133),
.Y(n_2866)
);

INVx2_ASAP7_75t_L g2867 ( 
.A(n_2533),
.Y(n_2867)
);

INVx2_ASAP7_75t_L g2868 ( 
.A(n_2534),
.Y(n_2868)
);

NAND2xp5_ASAP7_75t_L g2869 ( 
.A(n_2546),
.B(n_2133),
.Y(n_2869)
);

INVx2_ASAP7_75t_L g2870 ( 
.A(n_2536),
.Y(n_2870)
);

OAI22xp33_ASAP7_75t_L g2871 ( 
.A1(n_2484),
.A2(n_1473),
.B1(n_1475),
.B2(n_1453),
.Y(n_2871)
);

NAND2xp5_ASAP7_75t_L g2872 ( 
.A(n_2546),
.B(n_2133),
.Y(n_2872)
);

NAND2xp5_ASAP7_75t_L g2873 ( 
.A(n_2562),
.B(n_2150),
.Y(n_2873)
);

AOI22xp33_ASAP7_75t_L g2874 ( 
.A1(n_2826),
.A2(n_2423),
.B1(n_1633),
.B2(n_1475),
.Y(n_2874)
);

INVx2_ASAP7_75t_L g2875 ( 
.A(n_2550),
.Y(n_2875)
);

NAND2xp5_ASAP7_75t_L g2876 ( 
.A(n_2562),
.B(n_2150),
.Y(n_2876)
);

NAND2xp5_ASAP7_75t_L g2877 ( 
.A(n_2770),
.B(n_2150),
.Y(n_2877)
);

AO221x1_ASAP7_75t_L g2878 ( 
.A1(n_2786),
.A2(n_2485),
.B1(n_2731),
.B2(n_2661),
.C(n_2754),
.Y(n_2878)
);

INVx1_ASAP7_75t_L g2879 ( 
.A(n_2489),
.Y(n_2879)
);

NOR2x1p5_ASAP7_75t_L g2880 ( 
.A(n_2492),
.B(n_1473),
.Y(n_2880)
);

NOR2xp67_ASAP7_75t_L g2881 ( 
.A(n_2518),
.B(n_1486),
.Y(n_2881)
);

NAND2xp5_ASAP7_75t_L g2882 ( 
.A(n_2792),
.B(n_2697),
.Y(n_2882)
);

AOI22xp33_ASAP7_75t_L g2883 ( 
.A1(n_2797),
.A2(n_2821),
.B1(n_2557),
.B2(n_2566),
.Y(n_2883)
);

INVx1_ASAP7_75t_L g2884 ( 
.A(n_2491),
.Y(n_2884)
);

INVx1_ASAP7_75t_L g2885 ( 
.A(n_2493),
.Y(n_2885)
);

OAI21xp33_ASAP7_75t_L g2886 ( 
.A1(n_2603),
.A2(n_2313),
.B(n_2296),
.Y(n_2886)
);

NAND2xp5_ASAP7_75t_L g2887 ( 
.A(n_2700),
.B(n_2704),
.Y(n_2887)
);

INVx2_ASAP7_75t_L g2888 ( 
.A(n_2564),
.Y(n_2888)
);

NAND2xp5_ASAP7_75t_L g2889 ( 
.A(n_2708),
.B(n_1930),
.Y(n_2889)
);

NAND2xp33_ASAP7_75t_L g2890 ( 
.A(n_2478),
.B(n_2393),
.Y(n_2890)
);

NAND2xp5_ASAP7_75t_SL g2891 ( 
.A(n_2729),
.B(n_2307),
.Y(n_2891)
);

INVx2_ASAP7_75t_L g2892 ( 
.A(n_2573),
.Y(n_2892)
);

NOR2xp33_ASAP7_75t_L g2893 ( 
.A(n_2485),
.B(n_1531),
.Y(n_2893)
);

O2A1O1Ixp5_ASAP7_75t_L g2894 ( 
.A1(n_2578),
.A2(n_2270),
.B(n_2102),
.C(n_2126),
.Y(n_2894)
);

INVx2_ASAP7_75t_L g2895 ( 
.A(n_2582),
.Y(n_2895)
);

NAND2xp5_ASAP7_75t_L g2896 ( 
.A(n_2735),
.B(n_2423),
.Y(n_2896)
);

AOI22xp5_ASAP7_75t_L g2897 ( 
.A1(n_2749),
.A2(n_1486),
.B1(n_2423),
.B2(n_2346),
.Y(n_2897)
);

INVx1_ASAP7_75t_L g2898 ( 
.A(n_2495),
.Y(n_2898)
);

INVxp67_ASAP7_75t_L g2899 ( 
.A(n_2520),
.Y(n_2899)
);

AOI22xp5_ASAP7_75t_L g2900 ( 
.A1(n_2686),
.A2(n_2423),
.B1(n_2270),
.B2(n_2403),
.Y(n_2900)
);

NOR2xp33_ASAP7_75t_L g2901 ( 
.A(n_2640),
.B(n_1580),
.Y(n_2901)
);

INVx1_ASAP7_75t_L g2902 ( 
.A(n_2500),
.Y(n_2902)
);

INVx1_ASAP7_75t_L g2903 ( 
.A(n_2504),
.Y(n_2903)
);

NAND2xp5_ASAP7_75t_L g2904 ( 
.A(n_2763),
.B(n_2157),
.Y(n_2904)
);

AOI22xp33_ASAP7_75t_L g2905 ( 
.A1(n_2480),
.A2(n_1591),
.B1(n_1594),
.B2(n_1580),
.Y(n_2905)
);

NAND2xp5_ASAP7_75t_SL g2906 ( 
.A(n_2626),
.B(n_2627),
.Y(n_2906)
);

INVx8_ASAP7_75t_L g2907 ( 
.A(n_2610),
.Y(n_2907)
);

INVx8_ASAP7_75t_L g2908 ( 
.A(n_2610),
.Y(n_2908)
);

NAND2xp5_ASAP7_75t_L g2909 ( 
.A(n_2763),
.B(n_2157),
.Y(n_2909)
);

NAND2xp5_ASAP7_75t_SL g2910 ( 
.A(n_2626),
.B(n_2307),
.Y(n_2910)
);

AOI22xp5_ASAP7_75t_L g2911 ( 
.A1(n_2774),
.A2(n_2402),
.B1(n_2432),
.B2(n_2421),
.Y(n_2911)
);

NAND2xp5_ASAP7_75t_L g2912 ( 
.A(n_2747),
.B(n_1842),
.Y(n_2912)
);

INVx3_ASAP7_75t_L g2913 ( 
.A(n_2636),
.Y(n_2913)
);

NAND2xp5_ASAP7_75t_L g2914 ( 
.A(n_2758),
.B(n_1848),
.Y(n_2914)
);

NAND2xp5_ASAP7_75t_L g2915 ( 
.A(n_2765),
.B(n_1785),
.Y(n_2915)
);

NAND2xp5_ASAP7_75t_L g2916 ( 
.A(n_2603),
.B(n_1788),
.Y(n_2916)
);

NOR2xp33_ASAP7_75t_L g2917 ( 
.A(n_2502),
.B(n_1591),
.Y(n_2917)
);

INVx2_ASAP7_75t_SL g2918 ( 
.A(n_2733),
.Y(n_2918)
);

NAND2xp5_ASAP7_75t_L g2919 ( 
.A(n_2788),
.B(n_1793),
.Y(n_2919)
);

NOR2xp33_ASAP7_75t_L g2920 ( 
.A(n_2470),
.B(n_1594),
.Y(n_2920)
);

NAND2xp5_ASAP7_75t_L g2921 ( 
.A(n_2788),
.B(n_2122),
.Y(n_2921)
);

INVx2_ASAP7_75t_L g2922 ( 
.A(n_2632),
.Y(n_2922)
);

NAND2xp5_ASAP7_75t_L g2923 ( 
.A(n_2547),
.B(n_2321),
.Y(n_2923)
);

INVx1_ASAP7_75t_L g2924 ( 
.A(n_2505),
.Y(n_2924)
);

INVx5_ASAP7_75t_L g2925 ( 
.A(n_2610),
.Y(n_2925)
);

NAND2xp5_ASAP7_75t_L g2926 ( 
.A(n_2552),
.B(n_2330),
.Y(n_2926)
);

INVx2_ASAP7_75t_L g2927 ( 
.A(n_2633),
.Y(n_2927)
);

NAND2xp5_ASAP7_75t_L g2928 ( 
.A(n_2556),
.B(n_2335),
.Y(n_2928)
);

INVx2_ASAP7_75t_L g2929 ( 
.A(n_2642),
.Y(n_2929)
);

INVx2_ASAP7_75t_L g2930 ( 
.A(n_2651),
.Y(n_2930)
);

INVx2_ASAP7_75t_L g2931 ( 
.A(n_2666),
.Y(n_2931)
);

OR2x6_ASAP7_75t_L g2932 ( 
.A(n_2592),
.B(n_2393),
.Y(n_2932)
);

INVx1_ASAP7_75t_L g2933 ( 
.A(n_2509),
.Y(n_2933)
);

NAND2xp5_ASAP7_75t_SL g2934 ( 
.A(n_2627),
.B(n_2307),
.Y(n_2934)
);

INVx1_ASAP7_75t_L g2935 ( 
.A(n_2511),
.Y(n_2935)
);

CKINVDCx5p33_ASAP7_75t_R g2936 ( 
.A(n_2486),
.Y(n_2936)
);

INVx2_ASAP7_75t_L g2937 ( 
.A(n_2680),
.Y(n_2937)
);

BUFx3_ASAP7_75t_L g2938 ( 
.A(n_2523),
.Y(n_2938)
);

NAND2xp5_ASAP7_75t_SL g2939 ( 
.A(n_2507),
.B(n_2441),
.Y(n_2939)
);

AOI22xp5_ASAP7_75t_L g2940 ( 
.A1(n_2587),
.A2(n_2453),
.B1(n_1516),
.B2(n_1452),
.Y(n_2940)
);

OAI22xp5_ASAP7_75t_L g2941 ( 
.A1(n_2538),
.A2(n_2202),
.B1(n_2466),
.B2(n_2441),
.Y(n_2941)
);

NAND2xp5_ASAP7_75t_L g2942 ( 
.A(n_2559),
.B(n_2241),
.Y(n_2942)
);

BUFx6f_ASAP7_75t_L g2943 ( 
.A(n_2497),
.Y(n_2943)
);

AND2x4_ASAP7_75t_L g2944 ( 
.A(n_2569),
.B(n_2196),
.Y(n_2944)
);

INVx2_ASAP7_75t_L g2945 ( 
.A(n_2699),
.Y(n_2945)
);

INVx1_ASAP7_75t_L g2946 ( 
.A(n_2514),
.Y(n_2946)
);

AOI22xp5_ASAP7_75t_L g2947 ( 
.A1(n_2705),
.A2(n_1516),
.B1(n_1452),
.B2(n_1481),
.Y(n_2947)
);

OAI22xp5_ASAP7_75t_L g2948 ( 
.A1(n_2538),
.A2(n_2466),
.B1(n_2441),
.B2(n_2456),
.Y(n_2948)
);

NAND2xp5_ASAP7_75t_SL g2949 ( 
.A(n_2569),
.B(n_2466),
.Y(n_2949)
);

OR2x6_ASAP7_75t_L g2950 ( 
.A(n_2592),
.B(n_2393),
.Y(n_2950)
);

BUFx3_ASAP7_75t_L g2951 ( 
.A(n_2739),
.Y(n_2951)
);

NAND2xp5_ASAP7_75t_SL g2952 ( 
.A(n_2611),
.B(n_2451),
.Y(n_2952)
);

NOR2xp33_ASAP7_75t_L g2953 ( 
.A(n_2769),
.B(n_1614),
.Y(n_2953)
);

NAND2xp5_ASAP7_75t_SL g2954 ( 
.A(n_2611),
.B(n_2451),
.Y(n_2954)
);

NAND2xp5_ASAP7_75t_L g2955 ( 
.A(n_2578),
.B(n_2241),
.Y(n_2955)
);

INVx1_ASAP7_75t_L g2956 ( 
.A(n_2516),
.Y(n_2956)
);

BUFx6f_ASAP7_75t_SL g2957 ( 
.A(n_2496),
.Y(n_2957)
);

NAND2xp5_ASAP7_75t_SL g2958 ( 
.A(n_2682),
.B(n_2451),
.Y(n_2958)
);

OR2x6_ASAP7_75t_L g2959 ( 
.A(n_2592),
.B(n_2393),
.Y(n_2959)
);

AND2x2_ASAP7_75t_L g2960 ( 
.A(n_2600),
.B(n_2196),
.Y(n_2960)
);

NAND2xp5_ASAP7_75t_L g2961 ( 
.A(n_2588),
.B(n_2363),
.Y(n_2961)
);

INVx2_ASAP7_75t_L g2962 ( 
.A(n_2709),
.Y(n_2962)
);

INVx2_ASAP7_75t_L g2963 ( 
.A(n_2724),
.Y(n_2963)
);

INVx2_ASAP7_75t_L g2964 ( 
.A(n_2725),
.Y(n_2964)
);

AOI22xp33_ASAP7_75t_L g2965 ( 
.A1(n_2824),
.A2(n_1651),
.B1(n_1658),
.B2(n_1614),
.Y(n_2965)
);

NAND2xp5_ASAP7_75t_SL g2966 ( 
.A(n_2682),
.B(n_2157),
.Y(n_2966)
);

NAND2xp5_ASAP7_75t_L g2967 ( 
.A(n_2588),
.B(n_2381),
.Y(n_2967)
);

NAND2xp5_ASAP7_75t_SL g2968 ( 
.A(n_2716),
.B(n_2178),
.Y(n_2968)
);

AOI22xp33_ASAP7_75t_L g2969 ( 
.A1(n_2825),
.A2(n_1658),
.B1(n_1651),
.B2(n_1280),
.Y(n_2969)
);

INVx1_ASAP7_75t_L g2970 ( 
.A(n_2517),
.Y(n_2970)
);

INVx2_ASAP7_75t_L g2971 ( 
.A(n_2751),
.Y(n_2971)
);

AND2x2_ASAP7_75t_L g2972 ( 
.A(n_2601),
.B(n_2207),
.Y(n_2972)
);

NAND2xp5_ASAP7_75t_SL g2973 ( 
.A(n_2716),
.B(n_2178),
.Y(n_2973)
);

INVxp33_ASAP7_75t_L g2974 ( 
.A(n_2736),
.Y(n_2974)
);

INVx2_ASAP7_75t_L g2975 ( 
.A(n_2771),
.Y(n_2975)
);

INVx2_ASAP7_75t_L g2976 ( 
.A(n_2784),
.Y(n_2976)
);

NOR2x1p5_ASAP7_75t_L g2977 ( 
.A(n_2539),
.B(n_1817),
.Y(n_2977)
);

INVx2_ASAP7_75t_L g2978 ( 
.A(n_2787),
.Y(n_2978)
);

INVx4_ASAP7_75t_L g2979 ( 
.A(n_2522),
.Y(n_2979)
);

INVx2_ASAP7_75t_L g2980 ( 
.A(n_2794),
.Y(n_2980)
);

INVxp67_ASAP7_75t_L g2981 ( 
.A(n_2471),
.Y(n_2981)
);

A2O1A1Ixp33_ASAP7_75t_L g2982 ( 
.A1(n_2567),
.A2(n_2459),
.B(n_2445),
.C(n_2193),
.Y(n_2982)
);

NOR2xp33_ASAP7_75t_L g2983 ( 
.A(n_2803),
.B(n_1247),
.Y(n_2983)
);

INVx2_ASAP7_75t_L g2984 ( 
.A(n_2819),
.Y(n_2984)
);

NAND2xp5_ASAP7_75t_L g2985 ( 
.A(n_2567),
.B(n_2207),
.Y(n_2985)
);

NOR3xp33_ASAP7_75t_L g2986 ( 
.A(n_2637),
.B(n_2328),
.C(n_916),
.Y(n_2986)
);

O2A1O1Ixp33_ASAP7_75t_L g2987 ( 
.A1(n_2503),
.A2(n_2193),
.B(n_2195),
.C(n_2178),
.Y(n_2987)
);

AND2x4_ASAP7_75t_SL g2988 ( 
.A(n_2522),
.B(n_2180),
.Y(n_2988)
);

INVx8_ASAP7_75t_L g2989 ( 
.A(n_2610),
.Y(n_2989)
);

OR2x6_ASAP7_75t_L g2990 ( 
.A(n_2522),
.B(n_2219),
.Y(n_2990)
);

AND2x2_ASAP7_75t_L g2991 ( 
.A(n_2604),
.B(n_2219),
.Y(n_2991)
);

NAND2xp5_ASAP7_75t_L g2992 ( 
.A(n_2551),
.B(n_2243),
.Y(n_2992)
);

NAND2xp5_ASAP7_75t_SL g2993 ( 
.A(n_2696),
.B(n_2419),
.Y(n_2993)
);

INVx2_ASAP7_75t_L g2994 ( 
.A(n_2820),
.Y(n_2994)
);

NAND2xp5_ASAP7_75t_L g2995 ( 
.A(n_2822),
.B(n_2243),
.Y(n_2995)
);

INVx1_ASAP7_75t_L g2996 ( 
.A(n_2519),
.Y(n_2996)
);

NOR2xp33_ASAP7_75t_L g2997 ( 
.A(n_2481),
.B(n_1481),
.Y(n_2997)
);

NOR2xp33_ASAP7_75t_L g2998 ( 
.A(n_2501),
.B(n_1516),
.Y(n_2998)
);

NAND2xp33_ASAP7_75t_L g2999 ( 
.A(n_2801),
.B(n_2193),
.Y(n_2999)
);

NAND2xp5_ASAP7_75t_L g3000 ( 
.A(n_2543),
.B(n_2195),
.Y(n_3000)
);

NOR3xp33_ASAP7_75t_L g3001 ( 
.A(n_2827),
.B(n_916),
.C(n_889),
.Y(n_3001)
);

OAI22xp5_ASAP7_75t_L g3002 ( 
.A1(n_2730),
.A2(n_2555),
.B1(n_2543),
.B2(n_2768),
.Y(n_3002)
);

AND2x2_ASAP7_75t_L g3003 ( 
.A(n_2628),
.B(n_2356),
.Y(n_3003)
);

NAND2xp5_ASAP7_75t_L g3004 ( 
.A(n_2809),
.B(n_2195),
.Y(n_3004)
);

INVx2_ASAP7_75t_SL g3005 ( 
.A(n_2624),
.Y(n_3005)
);

NAND3xp33_ASAP7_75t_L g3006 ( 
.A(n_2721),
.B(n_1821),
.C(n_1817),
.Y(n_3006)
);

NAND2xp33_ASAP7_75t_L g3007 ( 
.A(n_2801),
.B(n_2236),
.Y(n_3007)
);

INVx2_ASAP7_75t_L g3008 ( 
.A(n_2678),
.Y(n_3008)
);

NOR2xp33_ASAP7_75t_L g3009 ( 
.A(n_2529),
.B(n_2356),
.Y(n_3009)
);

AND2x6_ASAP7_75t_L g3010 ( 
.A(n_2490),
.B(n_2109),
.Y(n_3010)
);

CKINVDCx5p33_ASAP7_75t_R g3011 ( 
.A(n_2510),
.Y(n_3011)
);

NOR2xp33_ASAP7_75t_L g3012 ( 
.A(n_2549),
.B(n_2415),
.Y(n_3012)
);

INVx2_ASAP7_75t_L g3013 ( 
.A(n_2681),
.Y(n_3013)
);

OAI22xp5_ASAP7_75t_L g3014 ( 
.A1(n_2730),
.A2(n_2255),
.B1(n_2272),
.B2(n_2236),
.Y(n_3014)
);

NOR2xp33_ASAP7_75t_L g3015 ( 
.A(n_2634),
.B(n_2415),
.Y(n_3015)
);

NAND2xp5_ASAP7_75t_L g3016 ( 
.A(n_2809),
.B(n_2236),
.Y(n_3016)
);

NAND2xp5_ASAP7_75t_L g3017 ( 
.A(n_2555),
.B(n_2255),
.Y(n_3017)
);

INVx1_ASAP7_75t_L g3018 ( 
.A(n_2526),
.Y(n_3018)
);

NAND2xp5_ASAP7_75t_SL g3019 ( 
.A(n_2558),
.B(n_2255),
.Y(n_3019)
);

NAND2xp5_ASAP7_75t_L g3020 ( 
.A(n_2801),
.B(n_2272),
.Y(n_3020)
);

INVx2_ASAP7_75t_L g3021 ( 
.A(n_2683),
.Y(n_3021)
);

AOI221xp5_ASAP7_75t_L g3022 ( 
.A1(n_2545),
.A2(n_1139),
.B1(n_1140),
.B2(n_1135),
.C(n_1134),
.Y(n_3022)
);

NAND2xp5_ASAP7_75t_SL g3023 ( 
.A(n_2548),
.B(n_2419),
.Y(n_3023)
);

AOI22xp33_ASAP7_75t_L g3024 ( 
.A1(n_2748),
.A2(n_1613),
.B1(n_1821),
.B2(n_1817),
.Y(n_3024)
);

NAND2xp5_ASAP7_75t_L g3025 ( 
.A(n_2801),
.B(n_2721),
.Y(n_3025)
);

AOI22xp33_ASAP7_75t_L g3026 ( 
.A1(n_2548),
.A2(n_1613),
.B1(n_1868),
.B2(n_1821),
.Y(n_3026)
);

NAND2xp5_ASAP7_75t_L g3027 ( 
.A(n_2571),
.B(n_2272),
.Y(n_3027)
);

NAND2xp5_ASAP7_75t_SL g3028 ( 
.A(n_2665),
.B(n_2456),
.Y(n_3028)
);

NAND2xp5_ASAP7_75t_SL g3029 ( 
.A(n_2524),
.B(n_2456),
.Y(n_3029)
);

NAND2xp5_ASAP7_75t_L g3030 ( 
.A(n_2571),
.B(n_2304),
.Y(n_3030)
);

BUFx6f_ASAP7_75t_L g3031 ( 
.A(n_2497),
.Y(n_3031)
);

AOI22xp33_ASAP7_75t_L g3032 ( 
.A1(n_2648),
.A2(n_1613),
.B1(n_1937),
.B2(n_1868),
.Y(n_3032)
);

INVx2_ASAP7_75t_SL g3033 ( 
.A(n_2659),
.Y(n_3033)
);

INVx2_ASAP7_75t_L g3034 ( 
.A(n_2684),
.Y(n_3034)
);

NAND2xp5_ASAP7_75t_L g3035 ( 
.A(n_2576),
.B(n_2304),
.Y(n_3035)
);

BUFx6f_ASAP7_75t_L g3036 ( 
.A(n_2497),
.Y(n_3036)
);

NAND2xp5_ASAP7_75t_L g3037 ( 
.A(n_2576),
.B(n_2304),
.Y(n_3037)
);

INVx1_ASAP7_75t_L g3038 ( 
.A(n_2527),
.Y(n_3038)
);

INVx2_ASAP7_75t_L g3039 ( 
.A(n_2685),
.Y(n_3039)
);

INVx3_ASAP7_75t_L g3040 ( 
.A(n_2679),
.Y(n_3040)
);

NAND2xp5_ASAP7_75t_L g3041 ( 
.A(n_2768),
.B(n_2613),
.Y(n_3041)
);

NAND2xp5_ASAP7_75t_L g3042 ( 
.A(n_2613),
.B(n_2388),
.Y(n_3042)
);

OR2x2_ASAP7_75t_L g3043 ( 
.A(n_2761),
.B(n_1903),
.Y(n_3043)
);

NAND2xp5_ASAP7_75t_SL g3044 ( 
.A(n_2532),
.B(n_2388),
.Y(n_3044)
);

NAND2xp5_ASAP7_75t_L g3045 ( 
.A(n_2745),
.B(n_2388),
.Y(n_3045)
);

NOR2xp33_ASAP7_75t_L g3046 ( 
.A(n_2754),
.B(n_1868),
.Y(n_3046)
);

BUFx6f_ASAP7_75t_L g3047 ( 
.A(n_2513),
.Y(n_3047)
);

NOR2xp33_ASAP7_75t_L g3048 ( 
.A(n_2795),
.B(n_1937),
.Y(n_3048)
);

NAND2xp5_ASAP7_75t_L g3049 ( 
.A(n_2745),
.B(n_2398),
.Y(n_3049)
);

INVx2_ASAP7_75t_L g3050 ( 
.A(n_2690),
.Y(n_3050)
);

NOR2xp33_ASAP7_75t_L g3051 ( 
.A(n_2795),
.B(n_1937),
.Y(n_3051)
);

NOR2xp33_ASAP7_75t_L g3052 ( 
.A(n_2813),
.B(n_1988),
.Y(n_3052)
);

NAND2xp5_ASAP7_75t_SL g3053 ( 
.A(n_2593),
.B(n_2398),
.Y(n_3053)
);

INVx2_ASAP7_75t_L g3054 ( 
.A(n_2693),
.Y(n_3054)
);

NAND2xp5_ASAP7_75t_SL g3055 ( 
.A(n_2668),
.B(n_2398),
.Y(n_3055)
);

INVx2_ASAP7_75t_L g3056 ( 
.A(n_2695),
.Y(n_3056)
);

INVx2_ASAP7_75t_L g3057 ( 
.A(n_2698),
.Y(n_3057)
);

NOR2xp33_ASAP7_75t_L g3058 ( 
.A(n_2813),
.B(n_1988),
.Y(n_3058)
);

NOR2xp33_ASAP7_75t_L g3059 ( 
.A(n_2661),
.B(n_1988),
.Y(n_3059)
);

NOR2xp33_ASAP7_75t_L g3060 ( 
.A(n_2672),
.B(n_2078),
.Y(n_3060)
);

NAND2xp5_ASAP7_75t_L g3061 ( 
.A(n_2745),
.B(n_2419),
.Y(n_3061)
);

INVxp67_ASAP7_75t_SL g3062 ( 
.A(n_2513),
.Y(n_3062)
);

NOR2xp67_ASAP7_75t_L g3063 ( 
.A(n_2650),
.B(n_2067),
.Y(n_3063)
);

NAND2xp5_ASAP7_75t_SL g3064 ( 
.A(n_2687),
.B(n_2138),
.Y(n_3064)
);

INVx1_ASAP7_75t_L g3065 ( 
.A(n_2528),
.Y(n_3065)
);

INVx2_ASAP7_75t_L g3066 ( 
.A(n_2702),
.Y(n_3066)
);

NAND2xp5_ASAP7_75t_L g3067 ( 
.A(n_2745),
.B(n_2259),
.Y(n_3067)
);

NAND2xp5_ASAP7_75t_L g3068 ( 
.A(n_2745),
.B(n_2746),
.Y(n_3068)
);

INVx2_ASAP7_75t_L g3069 ( 
.A(n_2706),
.Y(n_3069)
);

NOR2xp33_ASAP7_75t_L g3070 ( 
.A(n_2617),
.B(n_2078),
.Y(n_3070)
);

NAND2xp5_ASAP7_75t_L g3071 ( 
.A(n_2746),
.B(n_2259),
.Y(n_3071)
);

INVx2_ASAP7_75t_L g3072 ( 
.A(n_2710),
.Y(n_3072)
);

AND2x2_ASAP7_75t_L g3073 ( 
.A(n_2691),
.B(n_1144),
.Y(n_3073)
);

INVx1_ASAP7_75t_L g3074 ( 
.A(n_2531),
.Y(n_3074)
);

O2A1O1Ixp33_ASAP7_75t_L g3075 ( 
.A1(n_2692),
.A2(n_1912),
.B(n_1914),
.C(n_1904),
.Y(n_3075)
);

A2O1A1Ixp33_ASAP7_75t_L g3076 ( 
.A1(n_2638),
.A2(n_2459),
.B(n_2445),
.C(n_1922),
.Y(n_3076)
);

INVx1_ASAP7_75t_L g3077 ( 
.A(n_2537),
.Y(n_3077)
);

NAND2xp5_ASAP7_75t_L g3078 ( 
.A(n_2746),
.B(n_2261),
.Y(n_3078)
);

AOI22xp33_ASAP7_75t_L g3079 ( 
.A1(n_2630),
.A2(n_2078),
.B1(n_2110),
.B2(n_2109),
.Y(n_3079)
);

NAND2xp5_ASAP7_75t_SL g3080 ( 
.A(n_2799),
.B(n_2170),
.Y(n_3080)
);

NAND2xp5_ASAP7_75t_L g3081 ( 
.A(n_2746),
.B(n_2261),
.Y(n_3081)
);

NOR2xp33_ASAP7_75t_L g3082 ( 
.A(n_2799),
.B(n_2065),
.Y(n_3082)
);

NAND2xp5_ASAP7_75t_L g3083 ( 
.A(n_2746),
.B(n_2262),
.Y(n_3083)
);

AOI22xp5_ASAP7_75t_L g3084 ( 
.A1(n_2752),
.A2(n_2110),
.B1(n_2212),
.B2(n_2065),
.Y(n_3084)
);

NAND2xp5_ASAP7_75t_L g3085 ( 
.A(n_2753),
.B(n_2262),
.Y(n_3085)
);

INVx2_ASAP7_75t_L g3086 ( 
.A(n_2711),
.Y(n_3086)
);

OAI21xp33_ASAP7_75t_L g3087 ( 
.A1(n_2540),
.A2(n_2544),
.B(n_2542),
.Y(n_3087)
);

NAND2xp5_ASAP7_75t_L g3088 ( 
.A(n_2753),
.B(n_2264),
.Y(n_3088)
);

NAND2xp5_ASAP7_75t_L g3089 ( 
.A(n_2753),
.B(n_2264),
.Y(n_3089)
);

NAND2xp5_ASAP7_75t_L g3090 ( 
.A(n_2753),
.B(n_2271),
.Y(n_3090)
);

INVx1_ASAP7_75t_L g3091 ( 
.A(n_2575),
.Y(n_3091)
);

AND2x6_ASAP7_75t_SL g3092 ( 
.A(n_2498),
.B(n_1146),
.Y(n_3092)
);

NAND2xp5_ASAP7_75t_L g3093 ( 
.A(n_2753),
.B(n_2271),
.Y(n_3093)
);

INVx2_ASAP7_75t_L g3094 ( 
.A(n_2714),
.Y(n_3094)
);

INVx1_ASAP7_75t_L g3095 ( 
.A(n_2579),
.Y(n_3095)
);

NAND2xp5_ASAP7_75t_L g3096 ( 
.A(n_2638),
.B(n_2279),
.Y(n_3096)
);

INVx1_ASAP7_75t_L g3097 ( 
.A(n_2580),
.Y(n_3097)
);

INVx2_ASAP7_75t_L g3098 ( 
.A(n_2715),
.Y(n_3098)
);

BUFx6f_ASAP7_75t_SL g3099 ( 
.A(n_2610),
.Y(n_3099)
);

INVx2_ASAP7_75t_L g3100 ( 
.A(n_2717),
.Y(n_3100)
);

AOI22xp5_ASAP7_75t_L g3101 ( 
.A1(n_2760),
.A2(n_2110),
.B1(n_2212),
.B2(n_2065),
.Y(n_3101)
);

INVx2_ASAP7_75t_L g3102 ( 
.A(n_2722),
.Y(n_3102)
);

INVx2_ASAP7_75t_L g3103 ( 
.A(n_2728),
.Y(n_3103)
);

AOI22xp5_ASAP7_75t_L g3104 ( 
.A1(n_2800),
.A2(n_2212),
.B1(n_1919),
.B2(n_1923),
.Y(n_3104)
);

INVxp67_ASAP7_75t_L g3105 ( 
.A(n_2570),
.Y(n_3105)
);

INVx2_ASAP7_75t_L g3106 ( 
.A(n_2732),
.Y(n_3106)
);

INVxp67_ASAP7_75t_SL g3107 ( 
.A(n_2513),
.Y(n_3107)
);

HB1xp67_ASAP7_75t_L g3108 ( 
.A(n_2669),
.Y(n_3108)
);

HB1xp67_ASAP7_75t_L g3109 ( 
.A(n_2631),
.Y(n_3109)
);

NOR2xp67_ASAP7_75t_L g3110 ( 
.A(n_2565),
.B(n_2409),
.Y(n_3110)
);

INVx1_ASAP7_75t_L g3111 ( 
.A(n_2581),
.Y(n_3111)
);

NOR2xp33_ASAP7_75t_L g3112 ( 
.A(n_2577),
.B(n_1920),
.Y(n_3112)
);

AOI22xp5_ASAP7_75t_L g3113 ( 
.A1(n_2764),
.A2(n_1932),
.B1(n_1935),
.B2(n_1924),
.Y(n_3113)
);

NAND2xp5_ASAP7_75t_L g3114 ( 
.A(n_2560),
.B(n_2279),
.Y(n_3114)
);

BUFx3_ASAP7_75t_L g3115 ( 
.A(n_2618),
.Y(n_3115)
);

NAND2xp5_ASAP7_75t_L g3116 ( 
.A(n_2561),
.B(n_2283),
.Y(n_3116)
);

INVx2_ASAP7_75t_SL g3117 ( 
.A(n_2585),
.Y(n_3117)
);

NAND2xp5_ASAP7_75t_L g3118 ( 
.A(n_2563),
.B(n_2283),
.Y(n_3118)
);

INVx3_ASAP7_75t_L g3119 ( 
.A(n_2679),
.Y(n_3119)
);

NAND2xp5_ASAP7_75t_L g3120 ( 
.A(n_2673),
.B(n_2284),
.Y(n_3120)
);

NOR2xp33_ASAP7_75t_L g3121 ( 
.A(n_2584),
.B(n_1949),
.Y(n_3121)
);

NAND2xp5_ASAP7_75t_L g3122 ( 
.A(n_2675),
.B(n_2284),
.Y(n_3122)
);

NAND2xp5_ASAP7_75t_SL g3123 ( 
.A(n_2477),
.B(n_2141),
.Y(n_3123)
);

NOR2x1_ASAP7_75t_L g3124 ( 
.A(n_2645),
.B(n_1950),
.Y(n_3124)
);

NAND2xp33_ASAP7_75t_L g3125 ( 
.A(n_2772),
.B(n_2141),
.Y(n_3125)
);

AND2x2_ASAP7_75t_L g3126 ( 
.A(n_2762),
.B(n_2817),
.Y(n_3126)
);

INVx2_ASAP7_75t_L g3127 ( 
.A(n_2734),
.Y(n_3127)
);

INVx4_ASAP7_75t_L g3128 ( 
.A(n_2494),
.Y(n_3128)
);

BUFx6f_ASAP7_75t_SL g3129 ( 
.A(n_2506),
.Y(n_3129)
);

INVx1_ASAP7_75t_L g3130 ( 
.A(n_2583),
.Y(n_3130)
);

INVx2_ASAP7_75t_L g3131 ( 
.A(n_2737),
.Y(n_3131)
);

INVx2_ASAP7_75t_L g3132 ( 
.A(n_2738),
.Y(n_3132)
);

AND2x4_ASAP7_75t_L g3133 ( 
.A(n_2494),
.B(n_2380),
.Y(n_3133)
);

NAND2xp5_ASAP7_75t_L g3134 ( 
.A(n_2676),
.B(n_2285),
.Y(n_3134)
);

NOR2xp33_ASAP7_75t_L g3135 ( 
.A(n_2677),
.B(n_2457),
.Y(n_3135)
);

NOR2xp33_ASAP7_75t_L g3136 ( 
.A(n_2677),
.B(n_2457),
.Y(n_3136)
);

INVx1_ASAP7_75t_L g3137 ( 
.A(n_2589),
.Y(n_3137)
);

AOI22xp33_ASAP7_75t_L g3138 ( 
.A1(n_2757),
.A2(n_2294),
.B1(n_2286),
.B2(n_2292),
.Y(n_3138)
);

NOR2xp33_ASAP7_75t_L g3139 ( 
.A(n_2692),
.B(n_2462),
.Y(n_3139)
);

INVx1_ASAP7_75t_L g3140 ( 
.A(n_2590),
.Y(n_3140)
);

AOI22xp33_ASAP7_75t_L g3141 ( 
.A1(n_2639),
.A2(n_2294),
.B1(n_2286),
.B2(n_2292),
.Y(n_3141)
);

AOI21xp5_ASAP7_75t_L g3142 ( 
.A1(n_2674),
.A2(n_2424),
.B(n_2317),
.Y(n_3142)
);

NAND2xp5_ASAP7_75t_SL g3143 ( 
.A(n_2477),
.B(n_2141),
.Y(n_3143)
);

AND2x2_ASAP7_75t_L g3144 ( 
.A(n_2574),
.B(n_1147),
.Y(n_3144)
);

NAND2xp5_ASAP7_75t_L g3145 ( 
.A(n_2740),
.B(n_2285),
.Y(n_3145)
);

BUFx12f_ASAP7_75t_L g3146 ( 
.A(n_2936),
.Y(n_3146)
);

INVx2_ASAP7_75t_SL g3147 ( 
.A(n_2951),
.Y(n_3147)
);

AOI21xp5_ASAP7_75t_L g3148 ( 
.A1(n_2861),
.A2(n_2674),
.B(n_2701),
.Y(n_3148)
);

O2A1O1Ixp33_ASAP7_75t_L g3149 ( 
.A1(n_2861),
.A2(n_2694),
.B(n_2594),
.C(n_2595),
.Y(n_3149)
);

INVx2_ASAP7_75t_L g3150 ( 
.A(n_3008),
.Y(n_3150)
);

NOR2xp33_ASAP7_75t_L g3151 ( 
.A(n_2844),
.B(n_2553),
.Y(n_3151)
);

A2O1A1Ixp33_ASAP7_75t_L g3152 ( 
.A1(n_2850),
.A2(n_2723),
.B(n_2780),
.C(n_2720),
.Y(n_3152)
);

BUFx4f_ASAP7_75t_L g3153 ( 
.A(n_2932),
.Y(n_3153)
);

OAI21xp5_ASAP7_75t_L g3154 ( 
.A1(n_2844),
.A2(n_2701),
.B(n_2793),
.Y(n_3154)
);

AOI21xp5_ASAP7_75t_L g3155 ( 
.A1(n_2834),
.A2(n_2835),
.B(n_2838),
.Y(n_3155)
);

OAI21xp5_ASAP7_75t_L g3156 ( 
.A1(n_2838),
.A2(n_2793),
.B(n_2694),
.Y(n_3156)
);

AND2x6_ASAP7_75t_L g3157 ( 
.A(n_3133),
.B(n_2494),
.Y(n_3157)
);

AOI21xp5_ASAP7_75t_L g3158 ( 
.A1(n_2834),
.A2(n_2718),
.B(n_2525),
.Y(n_3158)
);

NAND2x2_ASAP7_75t_L g3159 ( 
.A(n_3117),
.B(n_2615),
.Y(n_3159)
);

NAND2xp5_ASAP7_75t_SL g3160 ( 
.A(n_2832),
.B(n_2688),
.Y(n_3160)
);

AOI21xp5_ASAP7_75t_L g3161 ( 
.A1(n_2835),
.A2(n_2718),
.B(n_2525),
.Y(n_3161)
);

INVx1_ASAP7_75t_L g3162 ( 
.A(n_2830),
.Y(n_3162)
);

INVx2_ASAP7_75t_L g3163 ( 
.A(n_3013),
.Y(n_3163)
);

INVx1_ASAP7_75t_L g3164 ( 
.A(n_2831),
.Y(n_3164)
);

NOR2xp33_ASAP7_75t_L g3165 ( 
.A(n_2833),
.B(n_2726),
.Y(n_3165)
);

A2O1A1Ixp33_ASAP7_75t_L g3166 ( 
.A1(n_2849),
.A2(n_2723),
.B(n_2780),
.C(n_2720),
.Y(n_3166)
);

AOI22xp5_ASAP7_75t_L g3167 ( 
.A1(n_2901),
.A2(n_2652),
.B1(n_2647),
.B2(n_2791),
.Y(n_3167)
);

INVx2_ASAP7_75t_L g3168 ( 
.A(n_3021),
.Y(n_3168)
);

OAI21xp5_ASAP7_75t_L g3169 ( 
.A1(n_2840),
.A2(n_2802),
.B(n_2719),
.Y(n_3169)
);

INVx3_ASAP7_75t_L g3170 ( 
.A(n_2907),
.Y(n_3170)
);

NAND2xp5_ASAP7_75t_SL g3171 ( 
.A(n_2897),
.B(n_2707),
.Y(n_3171)
);

NOR2xp33_ASAP7_75t_L g3172 ( 
.A(n_2845),
.B(n_2899),
.Y(n_3172)
);

NAND2xp5_ASAP7_75t_L g3173 ( 
.A(n_2916),
.B(n_2591),
.Y(n_3173)
);

NAND2xp5_ASAP7_75t_SL g3174 ( 
.A(n_2900),
.B(n_2515),
.Y(n_3174)
);

NAND2xp5_ASAP7_75t_L g3175 ( 
.A(n_2839),
.B(n_2596),
.Y(n_3175)
);

AOI21xp5_ASAP7_75t_L g3176 ( 
.A1(n_2840),
.A2(n_2727),
.B(n_2719),
.Y(n_3176)
);

OAI21xp33_ASAP7_75t_L g3177 ( 
.A1(n_2886),
.A2(n_894),
.B(n_889),
.Y(n_3177)
);

NOR2xp33_ASAP7_75t_L g3178 ( 
.A(n_2887),
.B(n_2713),
.Y(n_3178)
);

NAND2xp5_ASAP7_75t_L g3179 ( 
.A(n_2889),
.B(n_2597),
.Y(n_3179)
);

AND2x2_ASAP7_75t_L g3180 ( 
.A(n_3073),
.B(n_2607),
.Y(n_3180)
);

NAND2xp5_ASAP7_75t_L g3181 ( 
.A(n_2912),
.B(n_2914),
.Y(n_3181)
);

O2A1O1Ixp33_ASAP7_75t_L g3182 ( 
.A1(n_2828),
.A2(n_2609),
.B(n_2612),
.C(n_2608),
.Y(n_3182)
);

AOI21xp5_ASAP7_75t_L g3183 ( 
.A1(n_2999),
.A2(n_2727),
.B(n_2703),
.Y(n_3183)
);

OAI21xp5_ASAP7_75t_L g3184 ( 
.A1(n_2841),
.A2(n_2894),
.B(n_2982),
.Y(n_3184)
);

OAI21xp5_ASAP7_75t_L g3185 ( 
.A1(n_2841),
.A2(n_2802),
.B(n_1922),
.Y(n_3185)
);

AOI21xp5_ASAP7_75t_L g3186 ( 
.A1(n_3007),
.A2(n_2759),
.B(n_2703),
.Y(n_3186)
);

AOI21xp5_ASAP7_75t_L g3187 ( 
.A1(n_2843),
.A2(n_2759),
.B(n_2703),
.Y(n_3187)
);

INVx3_ASAP7_75t_L g3188 ( 
.A(n_2907),
.Y(n_3188)
);

AOI21x1_ASAP7_75t_L g3189 ( 
.A1(n_3142),
.A2(n_2741),
.B(n_2521),
.Y(n_3189)
);

A2O1A1Ixp33_ASAP7_75t_L g3190 ( 
.A1(n_3135),
.A2(n_2664),
.B(n_2667),
.C(n_2663),
.Y(n_3190)
);

OAI21xp33_ASAP7_75t_L g3191 ( 
.A1(n_2856),
.A2(n_896),
.B(n_894),
.Y(n_3191)
);

HB1xp67_ASAP7_75t_L g3192 ( 
.A(n_2981),
.Y(n_3192)
);

O2A1O1Ixp33_ASAP7_75t_L g3193 ( 
.A1(n_2829),
.A2(n_2616),
.B(n_2619),
.C(n_2614),
.Y(n_3193)
);

AOI21xp5_ASAP7_75t_L g3194 ( 
.A1(n_2941),
.A2(n_2759),
.B(n_2424),
.Y(n_3194)
);

AOI21xp5_ASAP7_75t_L g3195 ( 
.A1(n_2856),
.A2(n_2424),
.B(n_2170),
.Y(n_3195)
);

INVx1_ASAP7_75t_L g3196 ( 
.A(n_2842),
.Y(n_3196)
);

BUFx6f_ASAP7_75t_SL g3197 ( 
.A(n_2938),
.Y(n_3197)
);

INVx2_ASAP7_75t_SL g3198 ( 
.A(n_2977),
.Y(n_3198)
);

INVx1_ASAP7_75t_L g3199 ( 
.A(n_2848),
.Y(n_3199)
);

INVx5_ASAP7_75t_L g3200 ( 
.A(n_2932),
.Y(n_3200)
);

INVx1_ASAP7_75t_L g3201 ( 
.A(n_2854),
.Y(n_3201)
);

INVx1_ASAP7_75t_L g3202 ( 
.A(n_2862),
.Y(n_3202)
);

AOI21xp5_ASAP7_75t_L g3203 ( 
.A1(n_2857),
.A2(n_2170),
.B(n_2141),
.Y(n_3203)
);

AOI21xp5_ASAP7_75t_L g3204 ( 
.A1(n_2857),
.A2(n_2170),
.B(n_2141),
.Y(n_3204)
);

NOR2xp67_ASAP7_75t_L g3205 ( 
.A(n_2925),
.B(n_2490),
.Y(n_3205)
);

INVx1_ASAP7_75t_L g3206 ( 
.A(n_2879),
.Y(n_3206)
);

AOI21xp5_ASAP7_75t_L g3207 ( 
.A1(n_2866),
.A2(n_2180),
.B(n_2170),
.Y(n_3207)
);

CKINVDCx10_ASAP7_75t_R g3208 ( 
.A(n_3129),
.Y(n_3208)
);

NAND2xp5_ASAP7_75t_L g3209 ( 
.A(n_2915),
.B(n_2620),
.Y(n_3209)
);

AOI21xp5_ASAP7_75t_L g3210 ( 
.A1(n_2866),
.A2(n_2247),
.B(n_2180),
.Y(n_3210)
);

NAND2xp5_ASAP7_75t_L g3211 ( 
.A(n_2882),
.B(n_2621),
.Y(n_3211)
);

OR2x6_ASAP7_75t_L g3212 ( 
.A(n_2907),
.B(n_2515),
.Y(n_3212)
);

OAI22xp5_ASAP7_75t_L g3213 ( 
.A1(n_2847),
.A2(n_2623),
.B1(n_2625),
.B2(n_2622),
.Y(n_3213)
);

INVx2_ASAP7_75t_L g3214 ( 
.A(n_3034),
.Y(n_3214)
);

NOR2xp67_ASAP7_75t_SL g3215 ( 
.A(n_3011),
.B(n_2380),
.Y(n_3215)
);

BUFx6f_ASAP7_75t_L g3216 ( 
.A(n_2944),
.Y(n_3216)
);

AOI22xp33_ASAP7_75t_L g3217 ( 
.A1(n_2865),
.A2(n_2641),
.B1(n_2643),
.B2(n_2635),
.Y(n_3217)
);

OAI21xp5_ASAP7_75t_L g3218 ( 
.A1(n_3076),
.A2(n_1939),
.B(n_1899),
.Y(n_3218)
);

INVx1_ASAP7_75t_L g3219 ( 
.A(n_2884),
.Y(n_3219)
);

INVx1_ASAP7_75t_L g3220 ( 
.A(n_2885),
.Y(n_3220)
);

NOR2xp33_ASAP7_75t_SL g3221 ( 
.A(n_3070),
.B(n_2670),
.Y(n_3221)
);

NAND2xp5_ASAP7_75t_L g3222 ( 
.A(n_2919),
.B(n_2644),
.Y(n_3222)
);

NAND2xp5_ASAP7_75t_L g3223 ( 
.A(n_2985),
.B(n_2649),
.Y(n_3223)
);

NAND2xp5_ASAP7_75t_L g3224 ( 
.A(n_2961),
.B(n_2654),
.Y(n_3224)
);

INVx3_ASAP7_75t_L g3225 ( 
.A(n_2908),
.Y(n_3225)
);

AOI21xp5_ASAP7_75t_L g3226 ( 
.A1(n_2890),
.A2(n_2247),
.B(n_2180),
.Y(n_3226)
);

INVx1_ASAP7_75t_SL g3227 ( 
.A(n_2855),
.Y(n_3227)
);

INVx1_ASAP7_75t_L g3228 ( 
.A(n_2898),
.Y(n_3228)
);

AND2x2_ASAP7_75t_L g3229 ( 
.A(n_3144),
.B(n_3112),
.Y(n_3229)
);

INVx2_ASAP7_75t_L g3230 ( 
.A(n_3039),
.Y(n_3230)
);

O2A1O1Ixp33_ASAP7_75t_L g3231 ( 
.A1(n_2921),
.A2(n_2656),
.B(n_2657),
.C(n_2655),
.Y(n_3231)
);

NAND2xp33_ASAP7_75t_L g3232 ( 
.A(n_2847),
.B(n_2586),
.Y(n_3232)
);

AND2x4_ASAP7_75t_L g3233 ( 
.A(n_2932),
.B(n_2671),
.Y(n_3233)
);

AND2x2_ASAP7_75t_L g3234 ( 
.A(n_3121),
.B(n_2658),
.Y(n_3234)
);

INVx3_ASAP7_75t_L g3235 ( 
.A(n_2908),
.Y(n_3235)
);

INVx1_ASAP7_75t_L g3236 ( 
.A(n_2902),
.Y(n_3236)
);

AND2x2_ASAP7_75t_L g3237 ( 
.A(n_2960),
.B(n_2660),
.Y(n_3237)
);

NAND2x1p5_ASAP7_75t_L g3238 ( 
.A(n_3128),
.B(n_2712),
.Y(n_3238)
);

INVx2_ASAP7_75t_L g3239 ( 
.A(n_3050),
.Y(n_3239)
);

AOI21xp5_ASAP7_75t_L g3240 ( 
.A1(n_2948),
.A2(n_2247),
.B(n_2180),
.Y(n_3240)
);

AND2x4_ASAP7_75t_L g3241 ( 
.A(n_2950),
.B(n_2662),
.Y(n_3241)
);

NAND2xp5_ASAP7_75t_L g3242 ( 
.A(n_2967),
.B(n_2742),
.Y(n_3242)
);

NAND2xp5_ASAP7_75t_L g3243 ( 
.A(n_2972),
.B(n_2743),
.Y(n_3243)
);

NAND2xp5_ASAP7_75t_L g3244 ( 
.A(n_2991),
.B(n_2744),
.Y(n_3244)
);

NAND2xp5_ASAP7_75t_L g3245 ( 
.A(n_3003),
.B(n_2750),
.Y(n_3245)
);

AND2x2_ASAP7_75t_L g3246 ( 
.A(n_2983),
.B(n_896),
.Y(n_3246)
);

AND2x2_ASAP7_75t_L g3247 ( 
.A(n_3126),
.B(n_899),
.Y(n_3247)
);

AND2x2_ASAP7_75t_L g3248 ( 
.A(n_2944),
.B(n_899),
.Y(n_3248)
);

INVx1_ASAP7_75t_L g3249 ( 
.A(n_2903),
.Y(n_3249)
);

INVx1_ASAP7_75t_L g3250 ( 
.A(n_2924),
.Y(n_3250)
);

NAND2xp5_ASAP7_75t_L g3251 ( 
.A(n_3136),
.B(n_2755),
.Y(n_3251)
);

INVx2_ASAP7_75t_L g3252 ( 
.A(n_3054),
.Y(n_3252)
);

AOI21xp5_ASAP7_75t_L g3253 ( 
.A1(n_2836),
.A2(n_2298),
.B(n_2247),
.Y(n_3253)
);

AOI22xp33_ASAP7_75t_L g3254 ( 
.A1(n_2974),
.A2(n_2766),
.B1(n_2767),
.B2(n_2756),
.Y(n_3254)
);

NAND2xp5_ASAP7_75t_L g3255 ( 
.A(n_3139),
.B(n_2773),
.Y(n_3255)
);

AOI21xp5_ASAP7_75t_L g3256 ( 
.A1(n_2836),
.A2(n_2298),
.B(n_2247),
.Y(n_3256)
);

NAND2xp5_ASAP7_75t_L g3257 ( 
.A(n_2883),
.B(n_2775),
.Y(n_3257)
);

OR2x2_ASAP7_75t_L g3258 ( 
.A(n_3108),
.B(n_2776),
.Y(n_3258)
);

NAND2xp5_ASAP7_75t_L g3259 ( 
.A(n_3009),
.B(n_2777),
.Y(n_3259)
);

OAI22xp5_ASAP7_75t_L g3260 ( 
.A1(n_2869),
.A2(n_2599),
.B1(n_2605),
.B2(n_2586),
.Y(n_3260)
);

NAND2xp5_ASAP7_75t_L g3261 ( 
.A(n_3012),
.B(n_2778),
.Y(n_3261)
);

AND2x2_ASAP7_75t_L g3262 ( 
.A(n_2917),
.B(n_900),
.Y(n_3262)
);

AOI21xp5_ASAP7_75t_L g3263 ( 
.A1(n_3004),
.A2(n_2301),
.B(n_2298),
.Y(n_3263)
);

AND2x4_ASAP7_75t_L g3264 ( 
.A(n_2950),
.B(n_2712),
.Y(n_3264)
);

AOI21xp5_ASAP7_75t_L g3265 ( 
.A1(n_3004),
.A2(n_2301),
.B(n_2298),
.Y(n_3265)
);

NAND2xp5_ASAP7_75t_L g3266 ( 
.A(n_3015),
.B(n_2779),
.Y(n_3266)
);

INVx2_ASAP7_75t_L g3267 ( 
.A(n_3056),
.Y(n_3267)
);

BUFx3_ASAP7_75t_L g3268 ( 
.A(n_2918),
.Y(n_3268)
);

AOI21xp5_ASAP7_75t_L g3269 ( 
.A1(n_3016),
.A2(n_2301),
.B(n_2298),
.Y(n_3269)
);

OAI21xp5_ASAP7_75t_L g3270 ( 
.A1(n_2869),
.A2(n_1939),
.B(n_1899),
.Y(n_3270)
);

AOI22xp5_ASAP7_75t_L g3271 ( 
.A1(n_3060),
.A2(n_710),
.B1(n_729),
.B2(n_687),
.Y(n_3271)
);

OAI22xp5_ASAP7_75t_L g3272 ( 
.A1(n_2872),
.A2(n_2605),
.B1(n_2646),
.B2(n_2599),
.Y(n_3272)
);

AOI21xp5_ASAP7_75t_L g3273 ( 
.A1(n_3016),
.A2(n_2327),
.B(n_2301),
.Y(n_3273)
);

NOR2xp33_ASAP7_75t_SL g3274 ( 
.A(n_3129),
.B(n_2881),
.Y(n_3274)
);

AOI21xp5_ASAP7_75t_L g3275 ( 
.A1(n_2872),
.A2(n_2327),
.B(n_2301),
.Y(n_3275)
);

AOI21x1_ASAP7_75t_L g3276 ( 
.A1(n_2955),
.A2(n_2126),
.B(n_2113),
.Y(n_3276)
);

O2A1O1Ixp33_ASAP7_75t_SL g3277 ( 
.A1(n_2873),
.A2(n_2876),
.B(n_3049),
.C(n_3045),
.Y(n_3277)
);

INVx2_ASAP7_75t_L g3278 ( 
.A(n_3057),
.Y(n_3278)
);

NOR2xp33_ASAP7_75t_R g3279 ( 
.A(n_3115),
.B(n_2113),
.Y(n_3279)
);

AND2x2_ASAP7_75t_SL g3280 ( 
.A(n_3128),
.B(n_2781),
.Y(n_3280)
);

NOR2xp33_ASAP7_75t_L g3281 ( 
.A(n_2863),
.B(n_2646),
.Y(n_3281)
);

AND2x4_ASAP7_75t_L g3282 ( 
.A(n_2950),
.B(n_2380),
.Y(n_3282)
);

AOI21xp5_ASAP7_75t_L g3283 ( 
.A1(n_2873),
.A2(n_2369),
.B(n_2327),
.Y(n_3283)
);

AOI21xp5_ASAP7_75t_L g3284 ( 
.A1(n_2876),
.A2(n_2369),
.B(n_2327),
.Y(n_3284)
);

NOR2xp33_ASAP7_75t_L g3285 ( 
.A(n_2864),
.B(n_900),
.Y(n_3285)
);

INVx2_ASAP7_75t_SL g3286 ( 
.A(n_2880),
.Y(n_3286)
);

INVxp67_ASAP7_75t_L g3287 ( 
.A(n_3109),
.Y(n_3287)
);

AOI21xp5_ASAP7_75t_L g3288 ( 
.A1(n_3027),
.A2(n_2369),
.B(n_2327),
.Y(n_3288)
);

AOI21xp5_ASAP7_75t_L g3289 ( 
.A1(n_3027),
.A2(n_2390),
.B(n_2369),
.Y(n_3289)
);

BUFx6f_ASAP7_75t_L g3290 ( 
.A(n_2990),
.Y(n_3290)
);

NOR2xp33_ASAP7_75t_L g3291 ( 
.A(n_2893),
.B(n_906),
.Y(n_3291)
);

NAND2xp5_ASAP7_75t_SL g3292 ( 
.A(n_3025),
.B(n_2369),
.Y(n_3292)
);

INVx3_ASAP7_75t_L g3293 ( 
.A(n_2908),
.Y(n_3293)
);

AOI21xp5_ASAP7_75t_L g3294 ( 
.A1(n_3030),
.A2(n_2410),
.B(n_2390),
.Y(n_3294)
);

INVx2_ASAP7_75t_SL g3295 ( 
.A(n_3005),
.Y(n_3295)
);

NAND2xp33_ASAP7_75t_L g3296 ( 
.A(n_2851),
.B(n_2390),
.Y(n_3296)
);

INVx2_ASAP7_75t_L g3297 ( 
.A(n_3066),
.Y(n_3297)
);

NAND2xp5_ASAP7_75t_L g3298 ( 
.A(n_2933),
.B(n_2935),
.Y(n_3298)
);

O2A1O1Ixp33_ASAP7_75t_L g3299 ( 
.A1(n_3029),
.A2(n_1266),
.B(n_1259),
.C(n_1151),
.Y(n_3299)
);

NAND2xp5_ASAP7_75t_L g3300 ( 
.A(n_2946),
.B(n_2782),
.Y(n_3300)
);

OAI22xp5_ASAP7_75t_L g3301 ( 
.A1(n_2896),
.A2(n_1939),
.B1(n_1899),
.B2(n_998),
.Y(n_3301)
);

AO21x1_ASAP7_75t_L g3302 ( 
.A1(n_3096),
.A2(n_2785),
.B(n_2783),
.Y(n_3302)
);

AOI21xp5_ASAP7_75t_L g3303 ( 
.A1(n_3030),
.A2(n_2410),
.B(n_2390),
.Y(n_3303)
);

AOI21xp5_ASAP7_75t_L g3304 ( 
.A1(n_3035),
.A2(n_2410),
.B(n_2390),
.Y(n_3304)
);

BUFx3_ASAP7_75t_L g3305 ( 
.A(n_3033),
.Y(n_3305)
);

O2A1O1Ixp5_ASAP7_75t_L g3306 ( 
.A1(n_2958),
.A2(n_2463),
.B(n_2464),
.C(n_2462),
.Y(n_3306)
);

INVx1_ASAP7_75t_L g3307 ( 
.A(n_2956),
.Y(n_3307)
);

INVx1_ASAP7_75t_L g3308 ( 
.A(n_2970),
.Y(n_3308)
);

AOI21xp5_ASAP7_75t_L g3309 ( 
.A1(n_3035),
.A2(n_2410),
.B(n_2317),
.Y(n_3309)
);

AO21x1_ASAP7_75t_L g3310 ( 
.A1(n_3096),
.A2(n_2790),
.B(n_2789),
.Y(n_3310)
);

INVx2_ASAP7_75t_SL g3311 ( 
.A(n_3043),
.Y(n_3311)
);

AOI22xp5_ASAP7_75t_L g3312 ( 
.A1(n_3046),
.A2(n_712),
.B1(n_740),
.B2(n_690),
.Y(n_3312)
);

BUFx3_ASAP7_75t_L g3313 ( 
.A(n_2920),
.Y(n_3313)
);

NAND2xp5_ASAP7_75t_L g3314 ( 
.A(n_2996),
.B(n_2796),
.Y(n_3314)
);

O2A1O1Ixp33_ASAP7_75t_L g3315 ( 
.A1(n_3001),
.A2(n_1153),
.B(n_1156),
.C(n_1148),
.Y(n_3315)
);

OAI321xp33_ASAP7_75t_L g3316 ( 
.A1(n_2871),
.A2(n_1211),
.A3(n_1208),
.B1(n_1212),
.B2(n_1209),
.C(n_1202),
.Y(n_3316)
);

NAND2x1p5_ASAP7_75t_L g3317 ( 
.A(n_2925),
.B(n_3133),
.Y(n_3317)
);

INVx2_ASAP7_75t_L g3318 ( 
.A(n_3069),
.Y(n_3318)
);

NOR2xp67_ASAP7_75t_L g3319 ( 
.A(n_2925),
.B(n_2380),
.Y(n_3319)
);

OAI22xp33_ASAP7_75t_L g3320 ( 
.A1(n_2947),
.A2(n_910),
.B1(n_913),
.B2(n_906),
.Y(n_3320)
);

NAND2xp5_ASAP7_75t_L g3321 ( 
.A(n_3018),
.B(n_2798),
.Y(n_3321)
);

AOI21xp5_ASAP7_75t_L g3322 ( 
.A1(n_3037),
.A2(n_2410),
.B(n_2317),
.Y(n_3322)
);

OAI22xp5_ASAP7_75t_L g3323 ( 
.A1(n_2877),
.A2(n_1004),
.B1(n_924),
.B2(n_913),
.Y(n_3323)
);

AOI21xp5_ASAP7_75t_L g3324 ( 
.A1(n_3037),
.A2(n_2409),
.B(n_2380),
.Y(n_3324)
);

NOR2xp33_ASAP7_75t_L g3325 ( 
.A(n_3105),
.B(n_910),
.Y(n_3325)
);

INVx2_ASAP7_75t_L g3326 ( 
.A(n_3072),
.Y(n_3326)
);

NAND2xp5_ASAP7_75t_SL g3327 ( 
.A(n_3025),
.B(n_2409),
.Y(n_3327)
);

O2A1O1Ixp33_ASAP7_75t_L g3328 ( 
.A1(n_2952),
.A2(n_1158),
.B(n_1159),
.C(n_1157),
.Y(n_3328)
);

NAND2xp5_ASAP7_75t_L g3329 ( 
.A(n_3038),
.B(n_3065),
.Y(n_3329)
);

OAI22xp5_ASAP7_75t_L g3330 ( 
.A1(n_2877),
.A2(n_933),
.B1(n_918),
.B2(n_920),
.Y(n_3330)
);

INVx3_ASAP7_75t_L g3331 ( 
.A(n_2989),
.Y(n_3331)
);

INVx2_ASAP7_75t_L g3332 ( 
.A(n_3086),
.Y(n_3332)
);

NAND2xp5_ASAP7_75t_L g3333 ( 
.A(n_3074),
.B(n_2804),
.Y(n_3333)
);

INVx5_ASAP7_75t_L g3334 ( 
.A(n_2959),
.Y(n_3334)
);

CKINVDCx20_ASAP7_75t_R g3335 ( 
.A(n_2953),
.Y(n_3335)
);

AND2x2_ASAP7_75t_L g3336 ( 
.A(n_2874),
.B(n_917),
.Y(n_3336)
);

NAND2xp5_ASAP7_75t_SL g3337 ( 
.A(n_2911),
.B(n_3113),
.Y(n_3337)
);

OR2x2_ASAP7_75t_L g3338 ( 
.A(n_3077),
.B(n_2805),
.Y(n_3338)
);

NOR3xp33_ASAP7_75t_L g3339 ( 
.A(n_2986),
.B(n_918),
.C(n_917),
.Y(n_3339)
);

AOI21xp5_ASAP7_75t_L g3340 ( 
.A1(n_3017),
.A2(n_2409),
.B(n_2034),
.Y(n_3340)
);

AOI21xp33_ASAP7_75t_L g3341 ( 
.A1(n_2942),
.A2(n_2294),
.B(n_2806),
.Y(n_3341)
);

BUFx6f_ASAP7_75t_L g3342 ( 
.A(n_2990),
.Y(n_3342)
);

OAI21xp5_ASAP7_75t_L g3343 ( 
.A1(n_2987),
.A2(n_2034),
.B(n_1812),
.Y(n_3343)
);

O2A1O1Ixp33_ASAP7_75t_SL g3344 ( 
.A1(n_3045),
.A2(n_2808),
.B(n_2810),
.C(n_2807),
.Y(n_3344)
);

INVx1_ASAP7_75t_L g3345 ( 
.A(n_3091),
.Y(n_3345)
);

AOI21xp5_ASAP7_75t_L g3346 ( 
.A1(n_3017),
.A2(n_2409),
.B(n_2811),
.Y(n_3346)
);

NAND2xp5_ASAP7_75t_L g3347 ( 
.A(n_3095),
.B(n_2812),
.Y(n_3347)
);

AOI21x1_ASAP7_75t_L g3348 ( 
.A1(n_3002),
.A2(n_2226),
.B(n_2814),
.Y(n_3348)
);

INVx3_ASAP7_75t_L g3349 ( 
.A(n_2989),
.Y(n_3349)
);

A2O1A1Ixp33_ASAP7_75t_L g3350 ( 
.A1(n_3087),
.A2(n_2816),
.B(n_2818),
.C(n_2815),
.Y(n_3350)
);

NAND2xp5_ASAP7_75t_L g3351 ( 
.A(n_3097),
.B(n_2823),
.Y(n_3351)
);

INVx3_ASAP7_75t_SL g3352 ( 
.A(n_2990),
.Y(n_3352)
);

NOR3xp33_ASAP7_75t_L g3353 ( 
.A(n_2993),
.B(n_924),
.C(n_920),
.Y(n_3353)
);

NAND2xp5_ASAP7_75t_L g3354 ( 
.A(n_3111),
.B(n_930),
.Y(n_3354)
);

NAND2xp5_ASAP7_75t_L g3355 ( 
.A(n_3130),
.B(n_3137),
.Y(n_3355)
);

AOI21xp5_ASAP7_75t_L g3356 ( 
.A1(n_3000),
.A2(n_1812),
.B(n_1760),
.Y(n_3356)
);

NAND2xp33_ASAP7_75t_L g3357 ( 
.A(n_2851),
.B(n_2989),
.Y(n_3357)
);

AOI21xp5_ASAP7_75t_L g3358 ( 
.A1(n_3000),
.A2(n_1812),
.B(n_1760),
.Y(n_3358)
);

AOI22xp33_ASAP7_75t_L g3359 ( 
.A1(n_3337),
.A2(n_3138),
.B1(n_3141),
.B2(n_2878),
.Y(n_3359)
);

OR2x6_ASAP7_75t_SL g3360 ( 
.A(n_3258),
.B(n_3006),
.Y(n_3360)
);

NAND2xp5_ASAP7_75t_L g3361 ( 
.A(n_3181),
.B(n_3140),
.Y(n_3361)
);

AOI21xp5_ASAP7_75t_L g3362 ( 
.A1(n_3155),
.A2(n_3125),
.B(n_2968),
.Y(n_3362)
);

HB1xp67_ASAP7_75t_L g3363 ( 
.A(n_3311),
.Y(n_3363)
);

OAI22xp5_ASAP7_75t_SL g3364 ( 
.A1(n_3151),
.A2(n_3167),
.B1(n_3285),
.B2(n_3312),
.Y(n_3364)
);

AND2x4_ASAP7_75t_L g3365 ( 
.A(n_3200),
.B(n_2979),
.Y(n_3365)
);

NAND2xp5_ASAP7_75t_L g3366 ( 
.A(n_3180),
.B(n_3048),
.Y(n_3366)
);

AOI21xp5_ASAP7_75t_L g3367 ( 
.A1(n_3158),
.A2(n_3161),
.B(n_3232),
.Y(n_3367)
);

A2O1A1Ixp33_ASAP7_75t_L g3368 ( 
.A1(n_3166),
.A2(n_3075),
.B(n_3059),
.C(n_2940),
.Y(n_3368)
);

INVx1_ASAP7_75t_L g3369 ( 
.A(n_3298),
.Y(n_3369)
);

AND2x4_ASAP7_75t_L g3370 ( 
.A(n_3200),
.B(n_2979),
.Y(n_3370)
);

NAND2xp5_ASAP7_75t_L g3371 ( 
.A(n_3234),
.B(n_3051),
.Y(n_3371)
);

AOI21xp5_ASAP7_75t_L g3372 ( 
.A1(n_3156),
.A2(n_2973),
.B(n_2966),
.Y(n_3372)
);

AOI21xp5_ASAP7_75t_L g3373 ( 
.A1(n_3296),
.A2(n_3014),
.B(n_3020),
.Y(n_3373)
);

NAND2xp5_ASAP7_75t_SL g3374 ( 
.A(n_3280),
.B(n_3221),
.Y(n_3374)
);

NAND2xp5_ASAP7_75t_SL g3375 ( 
.A(n_3152),
.B(n_3052),
.Y(n_3375)
);

O2A1O1Ixp33_ASAP7_75t_L g3376 ( 
.A1(n_3291),
.A2(n_3053),
.B(n_2954),
.C(n_3028),
.Y(n_3376)
);

INVx1_ASAP7_75t_L g3377 ( 
.A(n_3329),
.Y(n_3377)
);

INVx1_ASAP7_75t_L g3378 ( 
.A(n_3355),
.Y(n_3378)
);

AND2x2_ASAP7_75t_L g3379 ( 
.A(n_3237),
.B(n_3058),
.Y(n_3379)
);

AND2x2_ASAP7_75t_L g3380 ( 
.A(n_3229),
.B(n_3124),
.Y(n_3380)
);

NAND2xp5_ASAP7_75t_L g3381 ( 
.A(n_3211),
.B(n_2904),
.Y(n_3381)
);

NAND2xp5_ASAP7_75t_L g3382 ( 
.A(n_3173),
.B(n_2904),
.Y(n_3382)
);

AOI21xp5_ASAP7_75t_L g3383 ( 
.A1(n_3176),
.A2(n_3020),
.B(n_3049),
.Y(n_3383)
);

O2A1O1Ixp33_ASAP7_75t_L g3384 ( 
.A1(n_3182),
.A2(n_3193),
.B(n_3320),
.C(n_3191),
.Y(n_3384)
);

AND2x2_ASAP7_75t_L g3385 ( 
.A(n_3248),
.B(n_3082),
.Y(n_3385)
);

BUFx8_ASAP7_75t_L g3386 ( 
.A(n_3197),
.Y(n_3386)
);

BUFx6f_ASAP7_75t_L g3387 ( 
.A(n_3216),
.Y(n_3387)
);

NOR2xp33_ASAP7_75t_L g3388 ( 
.A(n_3227),
.B(n_3092),
.Y(n_3388)
);

OAI22xp5_ASAP7_75t_L g3389 ( 
.A1(n_3312),
.A2(n_2926),
.B1(n_2928),
.B2(n_2923),
.Y(n_3389)
);

OAI22x1_ASAP7_75t_L g3390 ( 
.A1(n_3271),
.A2(n_2998),
.B1(n_2997),
.B2(n_3055),
.Y(n_3390)
);

AOI21xp5_ASAP7_75t_L g3391 ( 
.A1(n_3169),
.A2(n_3061),
.B(n_3042),
.Y(n_3391)
);

A2O1A1Ixp33_ASAP7_75t_L g3392 ( 
.A1(n_3191),
.A2(n_2995),
.B(n_3104),
.C(n_3063),
.Y(n_3392)
);

NAND3xp33_ASAP7_75t_L g3393 ( 
.A(n_3271),
.B(n_3022),
.C(n_3064),
.Y(n_3393)
);

INVx1_ASAP7_75t_L g3394 ( 
.A(n_3162),
.Y(n_3394)
);

NAND2xp5_ASAP7_75t_L g3395 ( 
.A(n_3209),
.B(n_2909),
.Y(n_3395)
);

NAND2xp5_ASAP7_75t_L g3396 ( 
.A(n_3175),
.B(n_2909),
.Y(n_3396)
);

INVx1_ASAP7_75t_L g3397 ( 
.A(n_3164),
.Y(n_3397)
);

NAND2xp5_ASAP7_75t_L g3398 ( 
.A(n_3224),
.B(n_3094),
.Y(n_3398)
);

INVx1_ASAP7_75t_L g3399 ( 
.A(n_3196),
.Y(n_3399)
);

AOI21xp5_ASAP7_75t_L g3400 ( 
.A1(n_3184),
.A2(n_3061),
.B(n_3042),
.Y(n_3400)
);

NOR2x1p5_ASAP7_75t_SL g3401 ( 
.A(n_3189),
.B(n_2851),
.Y(n_3401)
);

AOI21xp5_ASAP7_75t_L g3402 ( 
.A1(n_3240),
.A2(n_3143),
.B(n_3123),
.Y(n_3402)
);

NAND2xp5_ASAP7_75t_SL g3403 ( 
.A(n_3149),
.B(n_2925),
.Y(n_3403)
);

NAND2x1_ASAP7_75t_L g3404 ( 
.A(n_3170),
.B(n_2852),
.Y(n_3404)
);

OAI22xp5_ASAP7_75t_SL g3405 ( 
.A1(n_3167),
.A2(n_2905),
.B1(n_2969),
.B2(n_3032),
.Y(n_3405)
);

NOR2xp33_ASAP7_75t_L g3406 ( 
.A(n_3313),
.B(n_2965),
.Y(n_3406)
);

AND2x2_ASAP7_75t_L g3407 ( 
.A(n_3246),
.B(n_2992),
.Y(n_3407)
);

NAND2xp5_ASAP7_75t_L g3408 ( 
.A(n_3179),
.B(n_3098),
.Y(n_3408)
);

AOI21xp5_ASAP7_75t_L g3409 ( 
.A1(n_3277),
.A2(n_3068),
.B(n_3067),
.Y(n_3409)
);

BUFx6f_ASAP7_75t_L g3410 ( 
.A(n_3216),
.Y(n_3410)
);

OAI22xp5_ASAP7_75t_L g3411 ( 
.A1(n_3213),
.A2(n_3110),
.B1(n_2949),
.B2(n_3026),
.Y(n_3411)
);

OAI22xp5_ASAP7_75t_L g3412 ( 
.A1(n_3177),
.A2(n_3024),
.B1(n_3023),
.B2(n_3084),
.Y(n_3412)
);

OAI22xp5_ASAP7_75t_L g3413 ( 
.A1(n_3217),
.A2(n_3222),
.B1(n_3178),
.B2(n_3262),
.Y(n_3413)
);

AOI21xp5_ASAP7_75t_L g3414 ( 
.A1(n_3148),
.A2(n_3068),
.B(n_3067),
.Y(n_3414)
);

AOI21xp5_ASAP7_75t_L g3415 ( 
.A1(n_3218),
.A2(n_3078),
.B(n_3071),
.Y(n_3415)
);

OAI22xp5_ASAP7_75t_L g3416 ( 
.A1(n_3281),
.A2(n_3223),
.B1(n_3354),
.B2(n_3172),
.Y(n_3416)
);

BUFx2_ASAP7_75t_L g3417 ( 
.A(n_3192),
.Y(n_3417)
);

OAI22xp5_ASAP7_75t_L g3418 ( 
.A1(n_3336),
.A2(n_3190),
.B1(n_3287),
.B2(n_3286),
.Y(n_3418)
);

NAND2xp5_ASAP7_75t_L g3419 ( 
.A(n_3251),
.B(n_3100),
.Y(n_3419)
);

INVx2_ASAP7_75t_L g3420 ( 
.A(n_3150),
.Y(n_3420)
);

INVx2_ASAP7_75t_L g3421 ( 
.A(n_3163),
.Y(n_3421)
);

AOI21xp5_ASAP7_75t_L g3422 ( 
.A1(n_3183),
.A2(n_3078),
.B(n_3071),
.Y(n_3422)
);

INVx1_ASAP7_75t_L g3423 ( 
.A(n_3199),
.Y(n_3423)
);

NAND2xp5_ASAP7_75t_L g3424 ( 
.A(n_3255),
.B(n_3102),
.Y(n_3424)
);

NAND3xp33_ASAP7_75t_L g3425 ( 
.A(n_3339),
.B(n_2858),
.C(n_933),
.Y(n_3425)
);

AOI21xp5_ASAP7_75t_L g3426 ( 
.A1(n_3253),
.A2(n_3083),
.B(n_3081),
.Y(n_3426)
);

NAND2xp5_ASAP7_75t_SL g3427 ( 
.A(n_3316),
.B(n_2943),
.Y(n_3427)
);

AOI21xp5_ASAP7_75t_L g3428 ( 
.A1(n_3256),
.A2(n_3083),
.B(n_3081),
.Y(n_3428)
);

BUFx6f_ASAP7_75t_L g3429 ( 
.A(n_3216),
.Y(n_3429)
);

A2O1A1Ixp33_ASAP7_75t_L g3430 ( 
.A1(n_3231),
.A2(n_3101),
.B(n_3088),
.C(n_3089),
.Y(n_3430)
);

AOI21xp5_ASAP7_75t_L g3431 ( 
.A1(n_3226),
.A2(n_3289),
.B(n_3288),
.Y(n_3431)
);

OAI21xp5_ASAP7_75t_L g3432 ( 
.A1(n_3185),
.A2(n_3041),
.B(n_3085),
.Y(n_3432)
);

NAND2xp5_ASAP7_75t_SL g3433 ( 
.A(n_3241),
.B(n_2943),
.Y(n_3433)
);

OR2x2_ASAP7_75t_L g3434 ( 
.A(n_3201),
.B(n_3103),
.Y(n_3434)
);

OAI21xp5_ASAP7_75t_L g3435 ( 
.A1(n_3203),
.A2(n_3204),
.B(n_3275),
.Y(n_3435)
);

O2A1O1Ixp5_ASAP7_75t_L g3436 ( 
.A1(n_3160),
.A2(n_2934),
.B(n_2860),
.C(n_2891),
.Y(n_3436)
);

NAND2xp5_ASAP7_75t_SL g3437 ( 
.A(n_3241),
.B(n_2943),
.Y(n_3437)
);

AOI21xp5_ASAP7_75t_L g3438 ( 
.A1(n_3294),
.A2(n_3088),
.B(n_3085),
.Y(n_3438)
);

NAND2xp5_ASAP7_75t_SL g3439 ( 
.A(n_3233),
.B(n_3031),
.Y(n_3439)
);

AOI21xp5_ASAP7_75t_L g3440 ( 
.A1(n_3303),
.A2(n_3090),
.B(n_3089),
.Y(n_3440)
);

AOI21xp5_ASAP7_75t_L g3441 ( 
.A1(n_3304),
.A2(n_3093),
.B(n_3090),
.Y(n_3441)
);

AOI21xp5_ASAP7_75t_L g3442 ( 
.A1(n_3309),
.A2(n_3093),
.B(n_3041),
.Y(n_3442)
);

NAND3xp33_ASAP7_75t_L g3443 ( 
.A(n_3353),
.B(n_939),
.C(n_930),
.Y(n_3443)
);

AND2x2_ASAP7_75t_SL g3444 ( 
.A(n_3153),
.B(n_3079),
.Y(n_3444)
);

AOI21x1_ASAP7_75t_L g3445 ( 
.A1(n_3348),
.A2(n_3080),
.B(n_3145),
.Y(n_3445)
);

AOI22xp33_ASAP7_75t_L g3446 ( 
.A1(n_3165),
.A2(n_2957),
.B1(n_2846),
.B2(n_2853),
.Y(n_3446)
);

AOI21xp5_ASAP7_75t_L g3447 ( 
.A1(n_3322),
.A2(n_3116),
.B(n_3114),
.Y(n_3447)
);

OAI21x1_ASAP7_75t_L g3448 ( 
.A1(n_3340),
.A2(n_3145),
.B(n_3122),
.Y(n_3448)
);

NAND2xp5_ASAP7_75t_L g3449 ( 
.A(n_3266),
.B(n_3106),
.Y(n_3449)
);

NAND2xp5_ASAP7_75t_L g3450 ( 
.A(n_3259),
.B(n_3127),
.Y(n_3450)
);

BUFx3_ASAP7_75t_L g3451 ( 
.A(n_3147),
.Y(n_3451)
);

AOI21xp5_ASAP7_75t_L g3452 ( 
.A1(n_3194),
.A2(n_3116),
.B(n_3114),
.Y(n_3452)
);

NAND2xp5_ASAP7_75t_SL g3453 ( 
.A(n_3233),
.B(n_3031),
.Y(n_3453)
);

AOI21xp5_ASAP7_75t_L g3454 ( 
.A1(n_3207),
.A2(n_3118),
.B(n_3120),
.Y(n_3454)
);

OAI21xp33_ASAP7_75t_L g3455 ( 
.A1(n_3323),
.A2(n_992),
.B(n_939),
.Y(n_3455)
);

NOR2xp33_ASAP7_75t_L g3456 ( 
.A(n_3247),
.B(n_3044),
.Y(n_3456)
);

NAND2xp5_ASAP7_75t_L g3457 ( 
.A(n_3261),
.B(n_3131),
.Y(n_3457)
);

BUFx6f_ASAP7_75t_L g3458 ( 
.A(n_3153),
.Y(n_3458)
);

CKINVDCx20_ASAP7_75t_R g3459 ( 
.A(n_3335),
.Y(n_3459)
);

INVx2_ASAP7_75t_SL g3460 ( 
.A(n_3208),
.Y(n_3460)
);

BUFx6f_ASAP7_75t_L g3461 ( 
.A(n_3157),
.Y(n_3461)
);

NAND3xp33_ASAP7_75t_L g3462 ( 
.A(n_3154),
.B(n_3019),
.C(n_998),
.Y(n_3462)
);

OAI22xp5_ASAP7_75t_L g3463 ( 
.A1(n_3330),
.A2(n_3325),
.B1(n_3159),
.B2(n_3305),
.Y(n_3463)
);

AOI22x1_ASAP7_75t_L g3464 ( 
.A1(n_3187),
.A2(n_3210),
.B1(n_3283),
.B2(n_3284),
.Y(n_3464)
);

INVx2_ASAP7_75t_L g3465 ( 
.A(n_3168),
.Y(n_3465)
);

OAI22xp5_ASAP7_75t_L g3466 ( 
.A1(n_3268),
.A2(n_2959),
.B1(n_2957),
.B2(n_2939),
.Y(n_3466)
);

NOR2xp33_ASAP7_75t_L g3467 ( 
.A(n_3208),
.B(n_3197),
.Y(n_3467)
);

INVx3_ASAP7_75t_SL g3468 ( 
.A(n_3198),
.Y(n_3468)
);

BUFx12f_ASAP7_75t_L g3469 ( 
.A(n_3146),
.Y(n_3469)
);

A2O1A1Ixp33_ASAP7_75t_L g3470 ( 
.A1(n_3171),
.A2(n_2910),
.B(n_2906),
.C(n_3118),
.Y(n_3470)
);

AND2x2_ASAP7_75t_SL g3471 ( 
.A(n_3290),
.B(n_3342),
.Y(n_3471)
);

NAND2xp5_ASAP7_75t_SL g3472 ( 
.A(n_3264),
.B(n_3031),
.Y(n_3472)
);

NAND2xp5_ASAP7_75t_SL g3473 ( 
.A(n_3264),
.B(n_3036),
.Y(n_3473)
);

AOI22xp5_ASAP7_75t_L g3474 ( 
.A1(n_3274),
.A2(n_3099),
.B1(n_2959),
.B2(n_999),
.Y(n_3474)
);

OAI21xp5_ASAP7_75t_L g3475 ( 
.A1(n_3346),
.A2(n_3107),
.B(n_3062),
.Y(n_3475)
);

OAI22xp5_ASAP7_75t_L g3476 ( 
.A1(n_3254),
.A2(n_3099),
.B1(n_2988),
.B2(n_2913),
.Y(n_3476)
);

OA22x2_ASAP7_75t_L g3477 ( 
.A1(n_3257),
.A2(n_3132),
.B1(n_3122),
.B2(n_3120),
.Y(n_3477)
);

NAND2xp5_ASAP7_75t_L g3478 ( 
.A(n_3243),
.B(n_3134),
.Y(n_3478)
);

AOI22xp5_ASAP7_75t_L g3479 ( 
.A1(n_3174),
.A2(n_999),
.B1(n_1000),
.B2(n_992),
.Y(n_3479)
);

NOR2xp33_ASAP7_75t_L g3480 ( 
.A(n_3295),
.B(n_1000),
.Y(n_3480)
);

INVx2_ASAP7_75t_L g3481 ( 
.A(n_3214),
.Y(n_3481)
);

BUFx3_ASAP7_75t_L g3482 ( 
.A(n_3352),
.Y(n_3482)
);

NAND2xp5_ASAP7_75t_L g3483 ( 
.A(n_3244),
.B(n_3134),
.Y(n_3483)
);

AOI21xp5_ASAP7_75t_L g3484 ( 
.A1(n_3324),
.A2(n_2913),
.B(n_2852),
.Y(n_3484)
);

NOR2xp33_ASAP7_75t_L g3485 ( 
.A(n_3202),
.B(n_1003),
.Y(n_3485)
);

NAND2xp5_ASAP7_75t_L g3486 ( 
.A(n_3245),
.B(n_2837),
.Y(n_3486)
);

NAND2xp5_ASAP7_75t_L g3487 ( 
.A(n_3206),
.B(n_3219),
.Y(n_3487)
);

OAI22xp5_ASAP7_75t_L g3488 ( 
.A1(n_3260),
.A2(n_3119),
.B1(n_3040),
.B2(n_1004),
.Y(n_3488)
);

AND2x4_ASAP7_75t_L g3489 ( 
.A(n_3200),
.B(n_3036),
.Y(n_3489)
);

AO21x1_ASAP7_75t_L g3490 ( 
.A1(n_3272),
.A2(n_1219),
.B(n_1215),
.Y(n_3490)
);

HB1xp67_ASAP7_75t_L g3491 ( 
.A(n_3220),
.Y(n_3491)
);

NOR2xp33_ASAP7_75t_L g3492 ( 
.A(n_3228),
.B(n_1003),
.Y(n_3492)
);

AOI21xp5_ASAP7_75t_L g3493 ( 
.A1(n_3263),
.A2(n_3119),
.B(n_3040),
.Y(n_3493)
);

NOR2xp33_ASAP7_75t_L g3494 ( 
.A(n_3236),
.B(n_1008),
.Y(n_3494)
);

NOR2xp33_ASAP7_75t_L g3495 ( 
.A(n_3249),
.B(n_1008),
.Y(n_3495)
);

OAI22xp5_ASAP7_75t_L g3496 ( 
.A1(n_3301),
.A2(n_3047),
.B1(n_3036),
.B2(n_682),
.Y(n_3496)
);

AOI21xp5_ASAP7_75t_L g3497 ( 
.A1(n_3265),
.A2(n_3047),
.B(n_1760),
.Y(n_3497)
);

AOI22xp33_ASAP7_75t_L g3498 ( 
.A1(n_3230),
.A2(n_2867),
.B1(n_2868),
.B2(n_2859),
.Y(n_3498)
);

NAND2xp5_ASAP7_75t_L g3499 ( 
.A(n_3250),
.B(n_2870),
.Y(n_3499)
);

NAND2xp5_ASAP7_75t_L g3500 ( 
.A(n_3307),
.B(n_2875),
.Y(n_3500)
);

NAND2xp5_ASAP7_75t_L g3501 ( 
.A(n_3308),
.B(n_2888),
.Y(n_3501)
);

BUFx3_ASAP7_75t_L g3502 ( 
.A(n_3290),
.Y(n_3502)
);

A2O1A1Ixp33_ASAP7_75t_L g3503 ( 
.A1(n_3242),
.A2(n_1163),
.B(n_1166),
.C(n_1161),
.Y(n_3503)
);

INVx1_ASAP7_75t_L g3504 ( 
.A(n_3345),
.Y(n_3504)
);

O2A1O1Ixp5_ASAP7_75t_L g3505 ( 
.A1(n_3292),
.A2(n_2463),
.B(n_2467),
.C(n_2464),
.Y(n_3505)
);

AOI21xp5_ASAP7_75t_L g3506 ( 
.A1(n_3269),
.A2(n_3047),
.B(n_2232),
.Y(n_3506)
);

NAND2xp5_ASAP7_75t_L g3507 ( 
.A(n_3338),
.B(n_3300),
.Y(n_3507)
);

NAND2xp5_ASAP7_75t_L g3508 ( 
.A(n_3314),
.B(n_2892),
.Y(n_3508)
);

AOI21xp5_ASAP7_75t_L g3509 ( 
.A1(n_3273),
.A2(n_2232),
.B(n_2104),
.Y(n_3509)
);

NAND2xp5_ASAP7_75t_L g3510 ( 
.A(n_3321),
.B(n_2895),
.Y(n_3510)
);

AOI22x1_ASAP7_75t_L g3511 ( 
.A1(n_3186),
.A2(n_692),
.B1(n_699),
.B2(n_681),
.Y(n_3511)
);

AOI21xp5_ASAP7_75t_L g3512 ( 
.A1(n_3195),
.A2(n_2232),
.B(n_2104),
.Y(n_3512)
);

OAI22xp5_ASAP7_75t_L g3513 ( 
.A1(n_3270),
.A2(n_703),
.B1(n_704),
.B2(n_702),
.Y(n_3513)
);

AOI21xp5_ASAP7_75t_L g3514 ( 
.A1(n_3357),
.A2(n_2232),
.B(n_2104),
.Y(n_3514)
);

NAND2xp5_ASAP7_75t_SL g3515 ( 
.A(n_3279),
.B(n_2851),
.Y(n_3515)
);

AOI21x1_ASAP7_75t_L g3516 ( 
.A1(n_3276),
.A2(n_2467),
.B(n_2010),
.Y(n_3516)
);

OAI21x1_ASAP7_75t_L g3517 ( 
.A1(n_3356),
.A2(n_2297),
.B(n_2293),
.Y(n_3517)
);

OAI22xp5_ASAP7_75t_L g3518 ( 
.A1(n_3334),
.A2(n_711),
.B1(n_713),
.B2(n_706),
.Y(n_3518)
);

INVx2_ASAP7_75t_L g3519 ( 
.A(n_3239),
.Y(n_3519)
);

NAND2xp5_ASAP7_75t_L g3520 ( 
.A(n_3333),
.B(n_2922),
.Y(n_3520)
);

AND2x4_ASAP7_75t_L g3521 ( 
.A(n_3334),
.B(n_2927),
.Y(n_3521)
);

BUFx6f_ASAP7_75t_L g3522 ( 
.A(n_3157),
.Y(n_3522)
);

NAND2xp5_ASAP7_75t_L g3523 ( 
.A(n_3347),
.B(n_2929),
.Y(n_3523)
);

AOI21xp5_ASAP7_75t_L g3524 ( 
.A1(n_3344),
.A2(n_2232),
.B(n_2104),
.Y(n_3524)
);

AOI21xp5_ASAP7_75t_L g3525 ( 
.A1(n_3358),
.A2(n_2281),
.B(n_2104),
.Y(n_3525)
);

AOI21xp5_ASAP7_75t_L g3526 ( 
.A1(n_3343),
.A2(n_2281),
.B(n_2851),
.Y(n_3526)
);

INVx2_ASAP7_75t_L g3527 ( 
.A(n_3252),
.Y(n_3527)
);

AO21x1_ASAP7_75t_L g3528 ( 
.A1(n_3327),
.A2(n_1222),
.B(n_1221),
.Y(n_3528)
);

AOI21xp5_ASAP7_75t_L g3529 ( 
.A1(n_3302),
.A2(n_2281),
.B(n_2851),
.Y(n_3529)
);

INVx2_ASAP7_75t_L g3530 ( 
.A(n_3267),
.Y(n_3530)
);

OA22x2_ASAP7_75t_L g3531 ( 
.A1(n_3351),
.A2(n_2931),
.B1(n_2937),
.B2(n_2930),
.Y(n_3531)
);

AOI21xp5_ASAP7_75t_L g3532 ( 
.A1(n_3310),
.A2(n_3319),
.B(n_3350),
.Y(n_3532)
);

AOI21xp5_ASAP7_75t_L g3533 ( 
.A1(n_3319),
.A2(n_2281),
.B(n_2293),
.Y(n_3533)
);

NAND2xp5_ASAP7_75t_L g3534 ( 
.A(n_3278),
.B(n_2945),
.Y(n_3534)
);

AOI21xp5_ASAP7_75t_L g3535 ( 
.A1(n_3341),
.A2(n_2281),
.B(n_2297),
.Y(n_3535)
);

OAI21xp5_ASAP7_75t_L g3536 ( 
.A1(n_3315),
.A2(n_1958),
.B(n_1956),
.Y(n_3536)
);

NAND2xp5_ASAP7_75t_SL g3537 ( 
.A(n_3282),
.B(n_2962),
.Y(n_3537)
);

AOI22xp5_ASAP7_75t_L g3538 ( 
.A1(n_3212),
.A2(n_717),
.B1(n_719),
.B2(n_716),
.Y(n_3538)
);

NOR2xp33_ASAP7_75t_L g3539 ( 
.A(n_3290),
.B(n_724),
.Y(n_3539)
);

NAND2xp5_ASAP7_75t_L g3540 ( 
.A(n_3297),
.B(n_2963),
.Y(n_3540)
);

AND2x2_ASAP7_75t_L g3541 ( 
.A(n_3318),
.B(n_1168),
.Y(n_3541)
);

NAND2xp5_ASAP7_75t_L g3542 ( 
.A(n_3326),
.B(n_2964),
.Y(n_3542)
);

AND2x2_ASAP7_75t_L g3543 ( 
.A(n_3332),
.B(n_1170),
.Y(n_3543)
);

A2O1A1Ixp33_ASAP7_75t_L g3544 ( 
.A1(n_3299),
.A2(n_1173),
.B(n_1175),
.C(n_1171),
.Y(n_3544)
);

NOR2xp33_ASAP7_75t_R g3545 ( 
.A(n_3170),
.B(n_3010),
.Y(n_3545)
);

AOI22x1_ASAP7_75t_L g3546 ( 
.A1(n_3238),
.A2(n_737),
.B1(n_747),
.B2(n_730),
.Y(n_3546)
);

OAI22xp5_ASAP7_75t_L g3547 ( 
.A1(n_3334),
.A2(n_752),
.B1(n_753),
.B2(n_750),
.Y(n_3547)
);

OAI22xp5_ASAP7_75t_L g3548 ( 
.A1(n_3188),
.A2(n_758),
.B1(n_763),
.B2(n_756),
.Y(n_3548)
);

AOI21xp5_ASAP7_75t_L g3549 ( 
.A1(n_3205),
.A2(n_2306),
.B(n_2305),
.Y(n_3549)
);

OAI22xp5_ASAP7_75t_L g3550 ( 
.A1(n_3188),
.A2(n_3235),
.B1(n_3293),
.B2(n_3225),
.Y(n_3550)
);

NAND2xp5_ASAP7_75t_L g3551 ( 
.A(n_3342),
.B(n_2971),
.Y(n_3551)
);

OAI22xp5_ASAP7_75t_L g3552 ( 
.A1(n_3225),
.A2(n_766),
.B1(n_767),
.B2(n_765),
.Y(n_3552)
);

BUFx2_ASAP7_75t_L g3553 ( 
.A(n_3342),
.Y(n_3553)
);

A2O1A1Ixp33_ASAP7_75t_SL g3554 ( 
.A1(n_3215),
.A2(n_1178),
.B(n_1180),
.C(n_1176),
.Y(n_3554)
);

INVx3_ASAP7_75t_L g3555 ( 
.A(n_3282),
.Y(n_3555)
);

HB1xp67_ASAP7_75t_L g3556 ( 
.A(n_3212),
.Y(n_3556)
);

A2O1A1Ixp33_ASAP7_75t_L g3557 ( 
.A1(n_3328),
.A2(n_3306),
.B(n_3235),
.C(n_3293),
.Y(n_3557)
);

AOI21xp5_ASAP7_75t_L g3558 ( 
.A1(n_3205),
.A2(n_2306),
.B(n_2305),
.Y(n_3558)
);

OAI21xp5_ASAP7_75t_L g3559 ( 
.A1(n_3331),
.A2(n_1958),
.B(n_1956),
.Y(n_3559)
);

OAI22xp5_ASAP7_75t_L g3560 ( 
.A1(n_3331),
.A2(n_781),
.B1(n_784),
.B2(n_771),
.Y(n_3560)
);

NOR2xp33_ASAP7_75t_L g3561 ( 
.A(n_3349),
.B(n_792),
.Y(n_3561)
);

O2A1O1Ixp5_ASAP7_75t_L g3562 ( 
.A1(n_3349),
.A2(n_2077),
.B(n_1958),
.C(n_1977),
.Y(n_3562)
);

AOI22x1_ASAP7_75t_L g3563 ( 
.A1(n_3317),
.A2(n_797),
.B1(n_805),
.B2(n_796),
.Y(n_3563)
);

INVx1_ASAP7_75t_L g3564 ( 
.A(n_3212),
.Y(n_3564)
);

AOI21xp5_ASAP7_75t_L g3565 ( 
.A1(n_3157),
.A2(n_2329),
.B(n_2310),
.Y(n_3565)
);

AOI21x1_ASAP7_75t_SL g3566 ( 
.A1(n_3366),
.A2(n_3385),
.B(n_3379),
.Y(n_3566)
);

NAND2xp5_ASAP7_75t_L g3567 ( 
.A(n_3369),
.B(n_808),
.Y(n_3567)
);

OAI21xp5_ASAP7_75t_L g3568 ( 
.A1(n_3375),
.A2(n_1182),
.B(n_1181),
.Y(n_3568)
);

OAI21x1_ASAP7_75t_L g3569 ( 
.A1(n_3516),
.A2(n_2976),
.B(n_2975),
.Y(n_3569)
);

OAI21x1_ASAP7_75t_L g3570 ( 
.A1(n_3431),
.A2(n_2980),
.B(n_2978),
.Y(n_3570)
);

NAND2xp5_ASAP7_75t_L g3571 ( 
.A(n_3377),
.B(n_809),
.Y(n_3571)
);

OAI21x1_ASAP7_75t_L g3572 ( 
.A1(n_3464),
.A2(n_2994),
.B(n_2984),
.Y(n_3572)
);

NAND3x1_ASAP7_75t_L g3573 ( 
.A(n_3467),
.B(n_1227),
.C(n_1226),
.Y(n_3573)
);

NOR2xp33_ASAP7_75t_R g3574 ( 
.A(n_3459),
.B(n_3157),
.Y(n_3574)
);

OAI21xp5_ASAP7_75t_L g3575 ( 
.A1(n_3384),
.A2(n_1187),
.B(n_1186),
.Y(n_3575)
);

AO31x2_ASAP7_75t_L g3576 ( 
.A1(n_3532),
.A2(n_2329),
.A3(n_2332),
.B(n_2310),
.Y(n_3576)
);

INVx1_ASAP7_75t_L g3577 ( 
.A(n_3491),
.Y(n_3577)
);

AO21x1_ASAP7_75t_L g3578 ( 
.A1(n_3413),
.A2(n_1229),
.B(n_1228),
.Y(n_3578)
);

INVx1_ASAP7_75t_SL g3579 ( 
.A(n_3417),
.Y(n_3579)
);

OAI21x1_ASAP7_75t_L g3580 ( 
.A1(n_3529),
.A2(n_2333),
.B(n_2332),
.Y(n_3580)
);

NAND2xp5_ASAP7_75t_L g3581 ( 
.A(n_3378),
.B(n_813),
.Y(n_3581)
);

NAND2xp5_ASAP7_75t_L g3582 ( 
.A(n_3507),
.B(n_824),
.Y(n_3582)
);

OAI21x1_ASAP7_75t_L g3583 ( 
.A1(n_3435),
.A2(n_2338),
.B(n_2333),
.Y(n_3583)
);

AOI21xp5_ASAP7_75t_L g3584 ( 
.A1(n_3367),
.A2(n_2348),
.B(n_2338),
.Y(n_3584)
);

AOI21xp5_ASAP7_75t_L g3585 ( 
.A1(n_3362),
.A2(n_2349),
.B(n_2348),
.Y(n_3585)
);

NAND2xp5_ASAP7_75t_L g3586 ( 
.A(n_3396),
.B(n_826),
.Y(n_3586)
);

NAND2xp5_ASAP7_75t_L g3587 ( 
.A(n_3361),
.B(n_830),
.Y(n_3587)
);

OAI21x1_ASAP7_75t_L g3588 ( 
.A1(n_3526),
.A2(n_2355),
.B(n_2349),
.Y(n_3588)
);

INVxp67_ASAP7_75t_SL g3589 ( 
.A(n_3400),
.Y(n_3589)
);

BUFx2_ASAP7_75t_L g3590 ( 
.A(n_3363),
.Y(n_3590)
);

AOI21x1_ASAP7_75t_SL g3591 ( 
.A1(n_3371),
.A2(n_10),
.B(n_11),
.Y(n_3591)
);

AOI21xp5_ASAP7_75t_L g3592 ( 
.A1(n_3403),
.A2(n_2366),
.B(n_2355),
.Y(n_3592)
);

A2O1A1Ixp33_ASAP7_75t_L g3593 ( 
.A1(n_3368),
.A2(n_1191),
.B(n_1192),
.C(n_1190),
.Y(n_3593)
);

OAI21x1_ASAP7_75t_L g3594 ( 
.A1(n_3525),
.A2(n_2370),
.B(n_2366),
.Y(n_3594)
);

INVx2_ASAP7_75t_L g3595 ( 
.A(n_3420),
.Y(n_3595)
);

BUFx12f_ASAP7_75t_L g3596 ( 
.A(n_3386),
.Y(n_3596)
);

OAI21x1_ASAP7_75t_L g3597 ( 
.A1(n_3535),
.A2(n_2372),
.B(n_2370),
.Y(n_3597)
);

CKINVDCx20_ASAP7_75t_R g3598 ( 
.A(n_3386),
.Y(n_3598)
);

NAND2xp5_ASAP7_75t_L g3599 ( 
.A(n_3381),
.B(n_832),
.Y(n_3599)
);

OAI21x1_ASAP7_75t_L g3600 ( 
.A1(n_3517),
.A2(n_3497),
.B(n_3445),
.Y(n_3600)
);

AOI21x1_ASAP7_75t_L g3601 ( 
.A1(n_3374),
.A2(n_1195),
.B(n_1193),
.Y(n_3601)
);

NOR2x1_ASAP7_75t_SL g3602 ( 
.A(n_3461),
.B(n_1234),
.Y(n_3602)
);

INVx1_ASAP7_75t_L g3603 ( 
.A(n_3394),
.Y(n_3603)
);

AOI21xp5_ASAP7_75t_L g3604 ( 
.A1(n_3524),
.A2(n_2373),
.B(n_2372),
.Y(n_3604)
);

OAI21xp5_ASAP7_75t_L g3605 ( 
.A1(n_3393),
.A2(n_1201),
.B(n_1199),
.Y(n_3605)
);

NAND2xp5_ASAP7_75t_L g3606 ( 
.A(n_3395),
.B(n_3416),
.Y(n_3606)
);

NAND2xp5_ASAP7_75t_L g3607 ( 
.A(n_3382),
.B(n_833),
.Y(n_3607)
);

NAND2xp5_ASAP7_75t_L g3608 ( 
.A(n_3478),
.B(n_3483),
.Y(n_3608)
);

OAI21x1_ASAP7_75t_L g3609 ( 
.A1(n_3452),
.A2(n_2376),
.B(n_2373),
.Y(n_3609)
);

AND2x2_ASAP7_75t_L g3610 ( 
.A(n_3407),
.B(n_1236),
.Y(n_3610)
);

AND2x4_ASAP7_75t_L g3611 ( 
.A(n_3555),
.B(n_3482),
.Y(n_3611)
);

OAI21x1_ASAP7_75t_L g3612 ( 
.A1(n_3448),
.A2(n_2383),
.B(n_2376),
.Y(n_3612)
);

AND2x4_ASAP7_75t_L g3613 ( 
.A(n_3555),
.B(n_3010),
.Y(n_3613)
);

CKINVDCx5p33_ASAP7_75t_R g3614 ( 
.A(n_3469),
.Y(n_3614)
);

OAI21xp33_ASAP7_75t_L g3615 ( 
.A1(n_3455),
.A2(n_838),
.B(n_835),
.Y(n_3615)
);

OAI21x1_ASAP7_75t_SL g3616 ( 
.A1(n_3550),
.A2(n_3411),
.B(n_3484),
.Y(n_3616)
);

INVx3_ASAP7_75t_L g3617 ( 
.A(n_3489),
.Y(n_3617)
);

INVx1_ASAP7_75t_L g3618 ( 
.A(n_3397),
.Y(n_3618)
);

INVx3_ASAP7_75t_L g3619 ( 
.A(n_3489),
.Y(n_3619)
);

INVx4_ASAP7_75t_L g3620 ( 
.A(n_3451),
.Y(n_3620)
);

NAND2xp5_ASAP7_75t_L g3621 ( 
.A(n_3449),
.B(n_840),
.Y(n_3621)
);

CKINVDCx5p33_ASAP7_75t_R g3622 ( 
.A(n_3460),
.Y(n_3622)
);

OAI21x1_ASAP7_75t_L g3623 ( 
.A1(n_3512),
.A2(n_2384),
.B(n_2383),
.Y(n_3623)
);

NAND2xp5_ASAP7_75t_L g3624 ( 
.A(n_3398),
.B(n_847),
.Y(n_3624)
);

A2O1A1Ixp33_ASAP7_75t_L g3625 ( 
.A1(n_3538),
.A2(n_1238),
.B(n_1241),
.C(n_1237),
.Y(n_3625)
);

AOI21xp5_ASAP7_75t_L g3626 ( 
.A1(n_3373),
.A2(n_2386),
.B(n_2384),
.Y(n_3626)
);

BUFx5_ASAP7_75t_L g3627 ( 
.A(n_3365),
.Y(n_3627)
);

AOI31xp67_ASAP7_75t_L g3628 ( 
.A1(n_3477),
.A2(n_2015),
.A3(n_2051),
.B(n_1995),
.Y(n_3628)
);

INVx1_ASAP7_75t_L g3629 ( 
.A(n_3399),
.Y(n_3629)
);

NOR2xp67_ASAP7_75t_SL g3630 ( 
.A(n_3462),
.B(n_1245),
.Y(n_3630)
);

AND2x2_ASAP7_75t_L g3631 ( 
.A(n_3380),
.B(n_1248),
.Y(n_3631)
);

AO22x2_ASAP7_75t_L g3632 ( 
.A1(n_3418),
.A2(n_1251),
.B1(n_1253),
.B2(n_1249),
.Y(n_3632)
);

OAI21xp5_ASAP7_75t_L g3633 ( 
.A1(n_3462),
.A2(n_1256),
.B(n_1254),
.Y(n_3633)
);

AND2x2_ASAP7_75t_L g3634 ( 
.A(n_3423),
.B(n_1257),
.Y(n_3634)
);

OAI22x1_ASAP7_75t_L g3635 ( 
.A1(n_3474),
.A2(n_3388),
.B1(n_3504),
.B2(n_3406),
.Y(n_3635)
);

INVx1_ASAP7_75t_L g3636 ( 
.A(n_3487),
.Y(n_3636)
);

NAND2xp5_ASAP7_75t_L g3637 ( 
.A(n_3408),
.B(n_857),
.Y(n_3637)
);

NAND2xp5_ASAP7_75t_SL g3638 ( 
.A(n_3364),
.B(n_3444),
.Y(n_3638)
);

OAI21x1_ASAP7_75t_L g3639 ( 
.A1(n_3454),
.A2(n_2392),
.B(n_2386),
.Y(n_3639)
);

AOI21xp5_ASAP7_75t_L g3640 ( 
.A1(n_3514),
.A2(n_2399),
.B(n_2392),
.Y(n_3640)
);

OAI21x1_ASAP7_75t_L g3641 ( 
.A1(n_3447),
.A2(n_2401),
.B(n_2399),
.Y(n_3641)
);

AO31x2_ASAP7_75t_L g3642 ( 
.A1(n_3490),
.A2(n_2407),
.A3(n_2411),
.B(n_2401),
.Y(n_3642)
);

OAI21x1_ASAP7_75t_L g3643 ( 
.A1(n_3414),
.A2(n_3383),
.B(n_3402),
.Y(n_3643)
);

AOI21xp5_ASAP7_75t_L g3644 ( 
.A1(n_3509),
.A2(n_2411),
.B(n_2407),
.Y(n_3644)
);

NAND2xp5_ASAP7_75t_L g3645 ( 
.A(n_3450),
.B(n_859),
.Y(n_3645)
);

AOI21xp5_ASAP7_75t_L g3646 ( 
.A1(n_3391),
.A2(n_2420),
.B(n_2413),
.Y(n_3646)
);

OAI21x1_ASAP7_75t_L g3647 ( 
.A1(n_3493),
.A2(n_2420),
.B(n_2413),
.Y(n_3647)
);

INVxp67_ASAP7_75t_L g3648 ( 
.A(n_3456),
.Y(n_3648)
);

NAND2xp5_ASAP7_75t_SL g3649 ( 
.A(n_3364),
.B(n_1258),
.Y(n_3649)
);

OAI22xp5_ASAP7_75t_L g3650 ( 
.A1(n_3479),
.A2(n_861),
.B1(n_866),
.B2(n_860),
.Y(n_3650)
);

OAI21x1_ASAP7_75t_L g3651 ( 
.A1(n_3438),
.A2(n_2422),
.B(n_2051),
.Y(n_3651)
);

NOR2xp67_ASAP7_75t_L g3652 ( 
.A(n_3409),
.B(n_2422),
.Y(n_3652)
);

INVxp33_ASAP7_75t_L g3653 ( 
.A(n_3539),
.Y(n_3653)
);

OAI21x1_ASAP7_75t_L g3654 ( 
.A1(n_3440),
.A2(n_2060),
.B(n_2015),
.Y(n_3654)
);

NAND2xp5_ASAP7_75t_L g3655 ( 
.A(n_3457),
.B(n_3419),
.Y(n_3655)
);

OAI21x1_ASAP7_75t_L g3656 ( 
.A1(n_3441),
.A2(n_2069),
.B(n_2060),
.Y(n_3656)
);

NAND2xp5_ASAP7_75t_L g3657 ( 
.A(n_3424),
.B(n_868),
.Y(n_3657)
);

OAI21xp5_ASAP7_75t_L g3658 ( 
.A1(n_3455),
.A2(n_3470),
.B(n_3392),
.Y(n_3658)
);

OAI21x1_ASAP7_75t_L g3659 ( 
.A1(n_3426),
.A2(n_2069),
.B(n_1977),
.Y(n_3659)
);

OAI22xp5_ASAP7_75t_L g3660 ( 
.A1(n_3479),
.A2(n_870),
.B1(n_875),
.B2(n_869),
.Y(n_3660)
);

INVx2_ASAP7_75t_L g3661 ( 
.A(n_3421),
.Y(n_3661)
);

O2A1O1Ixp5_ASAP7_75t_L g3662 ( 
.A1(n_3372),
.A2(n_1977),
.B(n_2000),
.C(n_1956),
.Y(n_3662)
);

BUFx2_ASAP7_75t_L g3663 ( 
.A(n_3360),
.Y(n_3663)
);

NAND2xp5_ASAP7_75t_L g3664 ( 
.A(n_3434),
.B(n_879),
.Y(n_3664)
);

OAI21x1_ASAP7_75t_L g3665 ( 
.A1(n_3428),
.A2(n_2017),
.B(n_2000),
.Y(n_3665)
);

OR2x2_ASAP7_75t_L g3666 ( 
.A(n_3499),
.B(n_12),
.Y(n_3666)
);

NAND2xp5_ASAP7_75t_L g3667 ( 
.A(n_3486),
.B(n_942),
.Y(n_3667)
);

OAI21x1_ASAP7_75t_L g3668 ( 
.A1(n_3422),
.A2(n_2017),
.B(n_2000),
.Y(n_3668)
);

NAND2xp5_ASAP7_75t_L g3669 ( 
.A(n_3500),
.B(n_944),
.Y(n_3669)
);

INVx3_ASAP7_75t_L g3670 ( 
.A(n_3365),
.Y(n_3670)
);

AND2x2_ASAP7_75t_L g3671 ( 
.A(n_3553),
.B(n_13),
.Y(n_3671)
);

AOI21xp5_ASAP7_75t_L g3672 ( 
.A1(n_3442),
.A2(n_2081),
.B(n_2080),
.Y(n_3672)
);

AOI21x1_ASAP7_75t_L g3673 ( 
.A1(n_3390),
.A2(n_2081),
.B(n_2080),
.Y(n_3673)
);

INVx1_ASAP7_75t_L g3674 ( 
.A(n_3501),
.Y(n_3674)
);

NAND2xp5_ASAP7_75t_L g3675 ( 
.A(n_3508),
.B(n_946),
.Y(n_3675)
);

NAND2xp5_ASAP7_75t_L g3676 ( 
.A(n_3510),
.B(n_947),
.Y(n_3676)
);

OAI21x1_ASAP7_75t_L g3677 ( 
.A1(n_3505),
.A2(n_2031),
.B(n_2017),
.Y(n_3677)
);

HB1xp67_ASAP7_75t_L g3678 ( 
.A(n_3432),
.Y(n_3678)
);

OAI21x1_ASAP7_75t_L g3679 ( 
.A1(n_3506),
.A2(n_2040),
.B(n_2031),
.Y(n_3679)
);

NAND2xp5_ASAP7_75t_L g3680 ( 
.A(n_3520),
.B(n_948),
.Y(n_3680)
);

OAI21x1_ASAP7_75t_L g3681 ( 
.A1(n_3475),
.A2(n_2040),
.B(n_2031),
.Y(n_3681)
);

NAND2xp5_ASAP7_75t_L g3682 ( 
.A(n_3523),
.B(n_949),
.Y(n_3682)
);

AOI222xp33_ASAP7_75t_SL g3683 ( 
.A1(n_3463),
.A2(n_17),
.B1(n_20),
.B2(n_14),
.C1(n_15),
.C2(n_18),
.Y(n_3683)
);

A2O1A1Ixp33_ASAP7_75t_L g3684 ( 
.A1(n_3538),
.A2(n_959),
.B(n_960),
.C(n_954),
.Y(n_3684)
);

INVx1_ASAP7_75t_SL g3685 ( 
.A(n_3502),
.Y(n_3685)
);

BUFx3_ASAP7_75t_L g3686 ( 
.A(n_3468),
.Y(n_3686)
);

AO31x2_ASAP7_75t_L g3687 ( 
.A1(n_3430),
.A2(n_2092),
.A3(n_3010),
.B(n_1766),
.Y(n_3687)
);

BUFx4f_ASAP7_75t_L g3688 ( 
.A(n_3458),
.Y(n_3688)
);

NOR2xp33_ASAP7_75t_L g3689 ( 
.A(n_3480),
.B(n_961),
.Y(n_3689)
);

AO31x2_ASAP7_75t_L g3690 ( 
.A1(n_3415),
.A2(n_2092),
.A3(n_3010),
.B(n_1766),
.Y(n_3690)
);

INVx1_ASAP7_75t_L g3691 ( 
.A(n_3465),
.Y(n_3691)
);

NOR2xp67_ASAP7_75t_L g3692 ( 
.A(n_3564),
.B(n_2077),
.Y(n_3692)
);

OAI21x1_ASAP7_75t_L g3693 ( 
.A1(n_3562),
.A2(n_2070),
.B(n_2040),
.Y(n_3693)
);

AOI21x1_ASAP7_75t_L g3694 ( 
.A1(n_3515),
.A2(n_2077),
.B(n_2074),
.Y(n_3694)
);

OA22x2_ASAP7_75t_L g3695 ( 
.A1(n_3474),
.A2(n_966),
.B1(n_968),
.B2(n_964),
.Y(n_3695)
);

AO31x2_ASAP7_75t_L g3696 ( 
.A1(n_3528),
.A2(n_3010),
.A3(n_1766),
.B(n_1768),
.Y(n_3696)
);

AOI21xp5_ASAP7_75t_L g3697 ( 
.A1(n_3557),
.A2(n_2072),
.B(n_2070),
.Y(n_3697)
);

INVx2_ASAP7_75t_SL g3698 ( 
.A(n_3387),
.Y(n_3698)
);

BUFx10_ASAP7_75t_L g3699 ( 
.A(n_3561),
.Y(n_3699)
);

CKINVDCx5p33_ASAP7_75t_R g3700 ( 
.A(n_3387),
.Y(n_3700)
);

INVx2_ASAP7_75t_L g3701 ( 
.A(n_3481),
.Y(n_3701)
);

OAI21x1_ASAP7_75t_L g3702 ( 
.A1(n_3533),
.A2(n_2072),
.B(n_2070),
.Y(n_3702)
);

INVx1_ASAP7_75t_L g3703 ( 
.A(n_3519),
.Y(n_3703)
);

O2A1O1Ixp5_ASAP7_75t_L g3704 ( 
.A1(n_3427),
.A2(n_2072),
.B(n_21),
.C(n_18),
.Y(n_3704)
);

AOI21x1_ASAP7_75t_L g3705 ( 
.A1(n_3488),
.A2(n_2082),
.B(n_2074),
.Y(n_3705)
);

INVx3_ASAP7_75t_L g3706 ( 
.A(n_3370),
.Y(n_3706)
);

OAI21xp5_ASAP7_75t_L g3707 ( 
.A1(n_3389),
.A2(n_970),
.B(n_969),
.Y(n_3707)
);

NAND2xp5_ASAP7_75t_L g3708 ( 
.A(n_3527),
.B(n_973),
.Y(n_3708)
);

INVx5_ASAP7_75t_L g3709 ( 
.A(n_3461),
.Y(n_3709)
);

OAI22xp5_ASAP7_75t_L g3710 ( 
.A1(n_3405),
.A2(n_976),
.B1(n_979),
.B2(n_975),
.Y(n_3710)
);

INVx2_ASAP7_75t_L g3711 ( 
.A(n_3530),
.Y(n_3711)
);

NAND2xp5_ASAP7_75t_L g3712 ( 
.A(n_3485),
.B(n_981),
.Y(n_3712)
);

NAND2xp5_ASAP7_75t_L g3713 ( 
.A(n_3492),
.B(n_984),
.Y(n_3713)
);

OAI21xp5_ASAP7_75t_L g3714 ( 
.A1(n_3436),
.A2(n_3376),
.B(n_3359),
.Y(n_3714)
);

AOI21xp5_ASAP7_75t_SL g3715 ( 
.A1(n_3461),
.A2(n_853),
.B(n_842),
.Y(n_3715)
);

BUFx6f_ASAP7_75t_L g3716 ( 
.A(n_3458),
.Y(n_3716)
);

AOI21xp5_ASAP7_75t_L g3717 ( 
.A1(n_3404),
.A2(n_1766),
.B(n_1763),
.Y(n_3717)
);

NAND2xp5_ASAP7_75t_SL g3718 ( 
.A(n_3466),
.B(n_1768),
.Y(n_3718)
);

INVx2_ASAP7_75t_L g3719 ( 
.A(n_3534),
.Y(n_3719)
);

NAND2xp5_ASAP7_75t_L g3720 ( 
.A(n_3494),
.B(n_3495),
.Y(n_3720)
);

AND2x2_ASAP7_75t_L g3721 ( 
.A(n_3556),
.B(n_20),
.Y(n_3721)
);

OAI21x1_ASAP7_75t_L g3722 ( 
.A1(n_3549),
.A2(n_1784),
.B(n_1768),
.Y(n_3722)
);

NOR2xp33_ASAP7_75t_L g3723 ( 
.A(n_3405),
.B(n_988),
.Y(n_3723)
);

NAND2xp5_ASAP7_75t_L g3724 ( 
.A(n_3541),
.B(n_990),
.Y(n_3724)
);

AO31x2_ASAP7_75t_L g3725 ( 
.A1(n_3558),
.A2(n_1784),
.A3(n_1789),
.B(n_1768),
.Y(n_3725)
);

NOR2xp33_ASAP7_75t_L g3726 ( 
.A(n_3518),
.B(n_991),
.Y(n_3726)
);

NAND2xp5_ASAP7_75t_L g3727 ( 
.A(n_3543),
.B(n_22),
.Y(n_3727)
);

NAND2x1p5_ASAP7_75t_L g3728 ( 
.A(n_3522),
.B(n_1784),
.Y(n_3728)
);

NAND2xp5_ASAP7_75t_L g3729 ( 
.A(n_3387),
.B(n_3410),
.Y(n_3729)
);

AOI21x1_ASAP7_75t_L g3730 ( 
.A1(n_3412),
.A2(n_2089),
.B(n_2082),
.Y(n_3730)
);

AOI21xp5_ASAP7_75t_L g3731 ( 
.A1(n_3554),
.A2(n_1789),
.B(n_1784),
.Y(n_3731)
);

NAND2xp5_ASAP7_75t_L g3732 ( 
.A(n_3410),
.B(n_22),
.Y(n_3732)
);

NAND2x1p5_ASAP7_75t_L g3733 ( 
.A(n_3522),
.B(n_1789),
.Y(n_3733)
);

NAND2xp5_ASAP7_75t_L g3734 ( 
.A(n_3410),
.B(n_23),
.Y(n_3734)
);

INVx1_ASAP7_75t_L g3735 ( 
.A(n_3540),
.Y(n_3735)
);

OAI21x1_ASAP7_75t_L g3736 ( 
.A1(n_3565),
.A2(n_1800),
.B(n_1789),
.Y(n_3736)
);

OAI21xp5_ASAP7_75t_L g3737 ( 
.A1(n_3513),
.A2(n_3503),
.B(n_3425),
.Y(n_3737)
);

BUFx8_ASAP7_75t_L g3738 ( 
.A(n_3458),
.Y(n_3738)
);

NAND2xp5_ASAP7_75t_L g3739 ( 
.A(n_3429),
.B(n_23),
.Y(n_3739)
);

NAND2xp5_ASAP7_75t_L g3740 ( 
.A(n_3429),
.B(n_25),
.Y(n_3740)
);

BUFx12f_ASAP7_75t_L g3741 ( 
.A(n_3429),
.Y(n_3741)
);

AOI21xp5_ASAP7_75t_L g3742 ( 
.A1(n_3559),
.A2(n_1803),
.B(n_1800),
.Y(n_3742)
);

OAI21xp5_ASAP7_75t_L g3743 ( 
.A1(n_3547),
.A2(n_862),
.B(n_854),
.Y(n_3743)
);

O2A1O1Ixp5_ASAP7_75t_L g3744 ( 
.A1(n_3496),
.A2(n_29),
.B(n_25),
.C(n_27),
.Y(n_3744)
);

NOR2xp33_ASAP7_75t_L g3745 ( 
.A(n_3443),
.B(n_29),
.Y(n_3745)
);

O2A1O1Ixp5_ASAP7_75t_L g3746 ( 
.A1(n_3472),
.A2(n_35),
.B(n_30),
.C(n_34),
.Y(n_3746)
);

OAI21x1_ASAP7_75t_L g3747 ( 
.A1(n_3476),
.A2(n_3531),
.B(n_3536),
.Y(n_3747)
);

A2O1A1Ixp33_ASAP7_75t_L g3748 ( 
.A1(n_3446),
.A2(n_940),
.B(n_958),
.C(n_878),
.Y(n_3748)
);

INVxp67_ASAP7_75t_SL g3749 ( 
.A(n_3551),
.Y(n_3749)
);

AOI21xp33_ASAP7_75t_L g3750 ( 
.A1(n_3511),
.A2(n_1803),
.B(n_1800),
.Y(n_3750)
);

OAI21xp5_ASAP7_75t_L g3751 ( 
.A1(n_3548),
.A2(n_972),
.B(n_967),
.Y(n_3751)
);

INVx1_ASAP7_75t_L g3752 ( 
.A(n_3542),
.Y(n_3752)
);

OAI21x1_ASAP7_75t_L g3753 ( 
.A1(n_3439),
.A2(n_3453),
.B(n_3473),
.Y(n_3753)
);

AOI21xp33_ASAP7_75t_L g3754 ( 
.A1(n_3537),
.A2(n_1803),
.B(n_1800),
.Y(n_3754)
);

NAND2xp5_ASAP7_75t_L g3755 ( 
.A(n_3433),
.B(n_36),
.Y(n_3755)
);

AO31x2_ASAP7_75t_L g3756 ( 
.A1(n_3401),
.A2(n_3544),
.A3(n_3560),
.B(n_3552),
.Y(n_3756)
);

INVx1_ASAP7_75t_L g3757 ( 
.A(n_3521),
.Y(n_3757)
);

NOR2xp33_ASAP7_75t_L g3758 ( 
.A(n_3437),
.B(n_36),
.Y(n_3758)
);

INVx1_ASAP7_75t_L g3759 ( 
.A(n_3521),
.Y(n_3759)
);

NAND2xp5_ASAP7_75t_L g3760 ( 
.A(n_3471),
.B(n_37),
.Y(n_3760)
);

NOR4xp25_ASAP7_75t_L g3761 ( 
.A(n_3498),
.B(n_39),
.C(n_37),
.D(n_38),
.Y(n_3761)
);

INVx1_ASAP7_75t_L g3762 ( 
.A(n_3370),
.Y(n_3762)
);

AOI21x1_ASAP7_75t_L g3763 ( 
.A1(n_3545),
.A2(n_2089),
.B(n_2082),
.Y(n_3763)
);

AO21x2_ASAP7_75t_L g3764 ( 
.A1(n_3563),
.A2(n_1810),
.B(n_1803),
.Y(n_3764)
);

AOI21xp5_ASAP7_75t_L g3765 ( 
.A1(n_3522),
.A2(n_3546),
.B(n_1818),
.Y(n_3765)
);

INVx6_ASAP7_75t_L g3766 ( 
.A(n_3386),
.Y(n_3766)
);

OAI21x1_ASAP7_75t_L g3767 ( 
.A1(n_3516),
.A2(n_1818),
.B(n_1810),
.Y(n_3767)
);

OAI21x1_ASAP7_75t_L g3768 ( 
.A1(n_3516),
.A2(n_1818),
.B(n_1810),
.Y(n_3768)
);

OAI21xp5_ASAP7_75t_L g3769 ( 
.A1(n_3384),
.A2(n_987),
.B(n_983),
.Y(n_3769)
);

INVx1_ASAP7_75t_L g3770 ( 
.A(n_3491),
.Y(n_3770)
);

AOI221xp5_ASAP7_75t_SL g3771 ( 
.A1(n_3375),
.A2(n_41),
.B1(n_39),
.B2(n_40),
.C(n_42),
.Y(n_3771)
);

OA21x2_ASAP7_75t_L g3772 ( 
.A1(n_3367),
.A2(n_1818),
.B(n_1810),
.Y(n_3772)
);

NOR2xp67_ASAP7_75t_L g3773 ( 
.A(n_3532),
.B(n_353),
.Y(n_3773)
);

NAND2xp5_ASAP7_75t_L g3774 ( 
.A(n_3369),
.B(n_42),
.Y(n_3774)
);

AOI21x1_ASAP7_75t_L g3775 ( 
.A1(n_3375),
.A2(n_2089),
.B(n_2082),
.Y(n_3775)
);

AOI21x1_ASAP7_75t_L g3776 ( 
.A1(n_3375),
.A2(n_2095),
.B(n_2089),
.Y(n_3776)
);

OA21x2_ASAP7_75t_L g3777 ( 
.A1(n_3367),
.A2(n_1831),
.B(n_1825),
.Y(n_3777)
);

AOI21x1_ASAP7_75t_L g3778 ( 
.A1(n_3375),
.A2(n_2095),
.B(n_1831),
.Y(n_3778)
);

INVx3_ASAP7_75t_L g3779 ( 
.A(n_3555),
.Y(n_3779)
);

BUFx2_ASAP7_75t_L g3780 ( 
.A(n_3590),
.Y(n_3780)
);

AND2x2_ASAP7_75t_L g3781 ( 
.A(n_3579),
.B(n_43),
.Y(n_3781)
);

AOI22xp5_ASAP7_75t_L g3782 ( 
.A1(n_3683),
.A2(n_3638),
.B1(n_3723),
.B2(n_3658),
.Y(n_3782)
);

AND2x6_ASAP7_75t_L g3783 ( 
.A(n_3613),
.B(n_1825),
.Y(n_3783)
);

HB1xp67_ASAP7_75t_L g3784 ( 
.A(n_3577),
.Y(n_3784)
);

AND2x2_ASAP7_75t_L g3785 ( 
.A(n_3579),
.B(n_43),
.Y(n_3785)
);

INVx2_ASAP7_75t_SL g3786 ( 
.A(n_3766),
.Y(n_3786)
);

NAND2xp5_ASAP7_75t_L g3787 ( 
.A(n_3606),
.B(n_45),
.Y(n_3787)
);

INVx1_ASAP7_75t_L g3788 ( 
.A(n_3770),
.Y(n_3788)
);

INVx3_ASAP7_75t_L g3789 ( 
.A(n_3620),
.Y(n_3789)
);

HB1xp67_ASAP7_75t_L g3790 ( 
.A(n_3678),
.Y(n_3790)
);

OR2x2_ASAP7_75t_L g3791 ( 
.A(n_3603),
.B(n_45),
.Y(n_3791)
);

NOR2xp67_ASAP7_75t_L g3792 ( 
.A(n_3635),
.B(n_46),
.Y(n_3792)
);

HB1xp67_ASAP7_75t_L g3793 ( 
.A(n_3618),
.Y(n_3793)
);

BUFx3_ASAP7_75t_L g3794 ( 
.A(n_3686),
.Y(n_3794)
);

INVx1_ASAP7_75t_L g3795 ( 
.A(n_3629),
.Y(n_3795)
);

BUFx2_ASAP7_75t_L g3796 ( 
.A(n_3611),
.Y(n_3796)
);

CKINVDCx6p67_ASAP7_75t_R g3797 ( 
.A(n_3596),
.Y(n_3797)
);

NAND2xp5_ASAP7_75t_L g3798 ( 
.A(n_3608),
.B(n_46),
.Y(n_3798)
);

INVx2_ASAP7_75t_L g3799 ( 
.A(n_3595),
.Y(n_3799)
);

INVx4_ASAP7_75t_L g3800 ( 
.A(n_3620),
.Y(n_3800)
);

OAI22xp5_ASAP7_75t_L g3801 ( 
.A1(n_3720),
.A2(n_50),
.B1(n_48),
.B2(n_49),
.Y(n_3801)
);

NAND2xp5_ASAP7_75t_L g3802 ( 
.A(n_3636),
.B(n_49),
.Y(n_3802)
);

CKINVDCx5p33_ASAP7_75t_R g3803 ( 
.A(n_3614),
.Y(n_3803)
);

INVx2_ASAP7_75t_SL g3804 ( 
.A(n_3766),
.Y(n_3804)
);

AND2x2_ASAP7_75t_L g3805 ( 
.A(n_3663),
.B(n_51),
.Y(n_3805)
);

NAND2xp5_ASAP7_75t_L g3806 ( 
.A(n_3655),
.B(n_51),
.Y(n_3806)
);

INVx2_ASAP7_75t_SL g3807 ( 
.A(n_3700),
.Y(n_3807)
);

AOI21xp5_ASAP7_75t_L g3808 ( 
.A1(n_3589),
.A2(n_1831),
.B(n_1825),
.Y(n_3808)
);

INVx1_ASAP7_75t_L g3809 ( 
.A(n_3674),
.Y(n_3809)
);

INVx3_ASAP7_75t_L g3810 ( 
.A(n_3741),
.Y(n_3810)
);

AOI21xp5_ASAP7_75t_L g3811 ( 
.A1(n_3714),
.A2(n_1831),
.B(n_1825),
.Y(n_3811)
);

CKINVDCx20_ASAP7_75t_R g3812 ( 
.A(n_3598),
.Y(n_3812)
);

NOR2xp67_ASAP7_75t_SL g3813 ( 
.A(n_3715),
.B(n_2095),
.Y(n_3813)
);

NOR2xp33_ASAP7_75t_L g3814 ( 
.A(n_3699),
.B(n_52),
.Y(n_3814)
);

INVx2_ASAP7_75t_SL g3815 ( 
.A(n_3611),
.Y(n_3815)
);

O2A1O1Ixp33_ASAP7_75t_L g3816 ( 
.A1(n_3769),
.A2(n_56),
.B(n_54),
.C(n_55),
.Y(n_3816)
);

AOI22xp33_ASAP7_75t_L g3817 ( 
.A1(n_3769),
.A2(n_965),
.B1(n_921),
.B2(n_1832),
.Y(n_3817)
);

INVx2_ASAP7_75t_L g3818 ( 
.A(n_3661),
.Y(n_3818)
);

AND2x6_ASAP7_75t_L g3819 ( 
.A(n_3613),
.B(n_1832),
.Y(n_3819)
);

NAND3xp33_ASAP7_75t_L g3820 ( 
.A(n_3683),
.B(n_1418),
.C(n_1412),
.Y(n_3820)
);

AOI22xp33_ASAP7_75t_L g3821 ( 
.A1(n_3714),
.A2(n_965),
.B1(n_921),
.B2(n_1832),
.Y(n_3821)
);

AOI22xp33_ASAP7_75t_L g3822 ( 
.A1(n_3578),
.A2(n_965),
.B1(n_921),
.B2(n_1832),
.Y(n_3822)
);

AND2x4_ASAP7_75t_L g3823 ( 
.A(n_3670),
.B(n_54),
.Y(n_3823)
);

AOI22xp5_ASAP7_75t_L g3824 ( 
.A1(n_3649),
.A2(n_3615),
.B1(n_3632),
.B2(n_3573),
.Y(n_3824)
);

AOI22xp5_ASAP7_75t_L g3825 ( 
.A1(n_3615),
.A2(n_965),
.B1(n_921),
.B2(n_1861),
.Y(n_3825)
);

OR2x6_ASAP7_75t_L g3826 ( 
.A(n_3716),
.B(n_1412),
.Y(n_3826)
);

OA21x2_ASAP7_75t_L g3827 ( 
.A1(n_3643),
.A2(n_3600),
.B(n_3747),
.Y(n_3827)
);

AO31x2_ASAP7_75t_L g3828 ( 
.A1(n_3691),
.A2(n_1862),
.A3(n_1866),
.B(n_1861),
.Y(n_3828)
);

AOI22xp5_ASAP7_75t_L g3829 ( 
.A1(n_3632),
.A2(n_965),
.B1(n_921),
.B2(n_1861),
.Y(n_3829)
);

NOR2xp33_ASAP7_75t_L g3830 ( 
.A(n_3699),
.B(n_55),
.Y(n_3830)
);

NAND2xp5_ASAP7_75t_L g3831 ( 
.A(n_3610),
.B(n_57),
.Y(n_3831)
);

INVx1_ASAP7_75t_SL g3832 ( 
.A(n_3685),
.Y(n_3832)
);

A2O1A1Ixp33_ASAP7_75t_L g3833 ( 
.A1(n_3689),
.A2(n_59),
.B(n_57),
.C(n_58),
.Y(n_3833)
);

OAI22xp5_ASAP7_75t_L g3834 ( 
.A1(n_3737),
.A2(n_61),
.B1(n_58),
.B2(n_60),
.Y(n_3834)
);

INVx2_ASAP7_75t_L g3835 ( 
.A(n_3701),
.Y(n_3835)
);

INVx2_ASAP7_75t_SL g3836 ( 
.A(n_3685),
.Y(n_3836)
);

AND2x2_ASAP7_75t_L g3837 ( 
.A(n_3648),
.B(n_60),
.Y(n_3837)
);

AND2x2_ASAP7_75t_L g3838 ( 
.A(n_3779),
.B(n_3631),
.Y(n_3838)
);

O2A1O1Ixp33_ASAP7_75t_L g3839 ( 
.A1(n_3684),
.A2(n_64),
.B(n_62),
.C(n_63),
.Y(n_3839)
);

INVx2_ASAP7_75t_L g3840 ( 
.A(n_3711),
.Y(n_3840)
);

AND2x2_ASAP7_75t_L g3841 ( 
.A(n_3779),
.B(n_3670),
.Y(n_3841)
);

AND2x4_ASAP7_75t_L g3842 ( 
.A(n_3706),
.B(n_62),
.Y(n_3842)
);

INVx3_ASAP7_75t_SL g3843 ( 
.A(n_3622),
.Y(n_3843)
);

AOI21xp5_ASAP7_75t_L g3844 ( 
.A1(n_3616),
.A2(n_1862),
.B(n_1861),
.Y(n_3844)
);

BUFx10_ASAP7_75t_L g3845 ( 
.A(n_3758),
.Y(n_3845)
);

NAND2xp5_ASAP7_75t_L g3846 ( 
.A(n_3634),
.B(n_63),
.Y(n_3846)
);

NAND2xp5_ASAP7_75t_L g3847 ( 
.A(n_3749),
.B(n_3666),
.Y(n_3847)
);

INVx1_ASAP7_75t_L g3848 ( 
.A(n_3735),
.Y(n_3848)
);

AOI22xp5_ASAP7_75t_L g3849 ( 
.A1(n_3771),
.A2(n_965),
.B1(n_1866),
.B2(n_1862),
.Y(n_3849)
);

CKINVDCx20_ASAP7_75t_R g3850 ( 
.A(n_3738),
.Y(n_3850)
);

INVx2_ASAP7_75t_L g3851 ( 
.A(n_3703),
.Y(n_3851)
);

OAI22xp5_ASAP7_75t_L g3852 ( 
.A1(n_3737),
.A2(n_3707),
.B1(n_3745),
.B2(n_3726),
.Y(n_3852)
);

AND2x2_ASAP7_75t_L g3853 ( 
.A(n_3706),
.B(n_65),
.Y(n_3853)
);

INVx3_ASAP7_75t_L g3854 ( 
.A(n_3617),
.Y(n_3854)
);

INVx2_ASAP7_75t_L g3855 ( 
.A(n_3719),
.Y(n_3855)
);

INVx1_ASAP7_75t_L g3856 ( 
.A(n_3752),
.Y(n_3856)
);

AOI21xp5_ASAP7_75t_L g3857 ( 
.A1(n_3742),
.A2(n_1866),
.B(n_1862),
.Y(n_3857)
);

AOI21xp5_ASAP7_75t_L g3858 ( 
.A1(n_3662),
.A2(n_1867),
.B(n_1866),
.Y(n_3858)
);

BUFx6f_ASAP7_75t_L g3859 ( 
.A(n_3709),
.Y(n_3859)
);

NOR2xp33_ASAP7_75t_L g3860 ( 
.A(n_3653),
.B(n_66),
.Y(n_3860)
);

INVx1_ASAP7_75t_L g3861 ( 
.A(n_3757),
.Y(n_3861)
);

AOI221x1_ASAP7_75t_L g3862 ( 
.A1(n_3760),
.A2(n_1425),
.B1(n_1432),
.B2(n_1418),
.C(n_1412),
.Y(n_3862)
);

OR2x6_ASAP7_75t_L g3863 ( 
.A(n_3716),
.B(n_1418),
.Y(n_3863)
);

AND2x2_ASAP7_75t_SL g3864 ( 
.A(n_3761),
.B(n_66),
.Y(n_3864)
);

NAND2xp5_ASAP7_75t_L g3865 ( 
.A(n_3774),
.B(n_67),
.Y(n_3865)
);

INVx2_ASAP7_75t_L g3866 ( 
.A(n_3759),
.Y(n_3866)
);

NAND2xp5_ASAP7_75t_L g3867 ( 
.A(n_3599),
.B(n_67),
.Y(n_3867)
);

INVx1_ASAP7_75t_L g3868 ( 
.A(n_3570),
.Y(n_3868)
);

INVx2_ASAP7_75t_SL g3869 ( 
.A(n_3738),
.Y(n_3869)
);

AO32x1_ASAP7_75t_L g3870 ( 
.A1(n_3698),
.A2(n_70),
.A3(n_68),
.B1(n_69),
.B2(n_71),
.Y(n_3870)
);

NAND2x1_ASAP7_75t_L g3871 ( 
.A(n_3617),
.B(n_1418),
.Y(n_3871)
);

OAI21xp5_ASAP7_75t_L g3872 ( 
.A1(n_3761),
.A2(n_965),
.B(n_68),
.Y(n_3872)
);

NAND2xp5_ASAP7_75t_L g3873 ( 
.A(n_3607),
.B(n_69),
.Y(n_3873)
);

AOI22xp33_ASAP7_75t_L g3874 ( 
.A1(n_3695),
.A2(n_965),
.B1(n_1872),
.B2(n_1867),
.Y(n_3874)
);

OR2x2_ASAP7_75t_L g3875 ( 
.A(n_3727),
.B(n_3762),
.Y(n_3875)
);

INVx3_ASAP7_75t_L g3876 ( 
.A(n_3619),
.Y(n_3876)
);

INVx1_ASAP7_75t_L g3877 ( 
.A(n_3628),
.Y(n_3877)
);

AOI22xp5_ASAP7_75t_L g3878 ( 
.A1(n_3771),
.A2(n_1872),
.B1(n_1873),
.B2(n_1867),
.Y(n_3878)
);

AND2x2_ASAP7_75t_L g3879 ( 
.A(n_3671),
.B(n_71),
.Y(n_3879)
);

INVx2_ASAP7_75t_SL g3880 ( 
.A(n_3716),
.Y(n_3880)
);

NOR2xp33_ASAP7_75t_L g3881 ( 
.A(n_3712),
.B(n_3713),
.Y(n_3881)
);

BUFx10_ASAP7_75t_L g3882 ( 
.A(n_3574),
.Y(n_3882)
);

AND2x2_ASAP7_75t_L g3883 ( 
.A(n_3721),
.B(n_73),
.Y(n_3883)
);

OAI22xp5_ASAP7_75t_L g3884 ( 
.A1(n_3748),
.A2(n_3710),
.B1(n_3755),
.B2(n_3605),
.Y(n_3884)
);

INVx6_ASAP7_75t_L g3885 ( 
.A(n_3709),
.Y(n_3885)
);

INVx1_ASAP7_75t_L g3886 ( 
.A(n_3569),
.Y(n_3886)
);

INVx1_ASAP7_75t_L g3887 ( 
.A(n_3576),
.Y(n_3887)
);

INVx1_ASAP7_75t_L g3888 ( 
.A(n_3576),
.Y(n_3888)
);

INVx2_ASAP7_75t_L g3889 ( 
.A(n_3576),
.Y(n_3889)
);

OAI22xp5_ASAP7_75t_L g3890 ( 
.A1(n_3605),
.A2(n_77),
.B1(n_74),
.B2(n_76),
.Y(n_3890)
);

NAND2xp5_ASAP7_75t_L g3891 ( 
.A(n_3586),
.B(n_74),
.Y(n_3891)
);

AND2x4_ASAP7_75t_L g3892 ( 
.A(n_3619),
.B(n_76),
.Y(n_3892)
);

BUFx6f_ASAP7_75t_L g3893 ( 
.A(n_3709),
.Y(n_3893)
);

INVx3_ASAP7_75t_L g3894 ( 
.A(n_3627),
.Y(n_3894)
);

AOI22xp33_ASAP7_75t_L g3895 ( 
.A1(n_3724),
.A2(n_1872),
.B1(n_1873),
.B2(n_1867),
.Y(n_3895)
);

INVx1_ASAP7_75t_L g3896 ( 
.A(n_3572),
.Y(n_3896)
);

AOI22xp5_ASAP7_75t_L g3897 ( 
.A1(n_3630),
.A2(n_1873),
.B1(n_1886),
.B2(n_1872),
.Y(n_3897)
);

INVx1_ASAP7_75t_L g3898 ( 
.A(n_3732),
.Y(n_3898)
);

AOI21xp5_ASAP7_75t_L g3899 ( 
.A1(n_3773),
.A2(n_1886),
.B(n_1873),
.Y(n_3899)
);

NAND2xp5_ASAP7_75t_L g3900 ( 
.A(n_3621),
.B(n_78),
.Y(n_3900)
);

NAND2xp5_ASAP7_75t_L g3901 ( 
.A(n_3645),
.B(n_79),
.Y(n_3901)
);

AOI221x1_ASAP7_75t_L g3902 ( 
.A1(n_3734),
.A2(n_1472),
.B1(n_1477),
.B2(n_1432),
.C(n_1425),
.Y(n_3902)
);

NAND2xp5_ASAP7_75t_L g3903 ( 
.A(n_3657),
.B(n_79),
.Y(n_3903)
);

AOI21xp5_ASAP7_75t_L g3904 ( 
.A1(n_3773),
.A2(n_1887),
.B(n_1886),
.Y(n_3904)
);

INVx1_ASAP7_75t_L g3905 ( 
.A(n_3739),
.Y(n_3905)
);

INVx1_ASAP7_75t_L g3906 ( 
.A(n_3740),
.Y(n_3906)
);

HB1xp67_ASAP7_75t_L g3907 ( 
.A(n_3729),
.Y(n_3907)
);

AOI22xp5_ASAP7_75t_L g3908 ( 
.A1(n_3718),
.A2(n_3575),
.B1(n_3568),
.B2(n_3633),
.Y(n_3908)
);

NAND2xp5_ASAP7_75t_L g3909 ( 
.A(n_3587),
.B(n_80),
.Y(n_3909)
);

INVx1_ASAP7_75t_L g3910 ( 
.A(n_3753),
.Y(n_3910)
);

AO22x1_ASAP7_75t_L g3911 ( 
.A1(n_3575),
.A2(n_83),
.B1(n_81),
.B2(n_82),
.Y(n_3911)
);

AND2x4_ASAP7_75t_L g3912 ( 
.A(n_3692),
.B(n_81),
.Y(n_3912)
);

AOI21xp5_ASAP7_75t_L g3913 ( 
.A1(n_3584),
.A2(n_1887),
.B(n_1886),
.Y(n_3913)
);

INVx2_ASAP7_75t_L g3914 ( 
.A(n_3690),
.Y(n_3914)
);

HB1xp67_ASAP7_75t_L g3915 ( 
.A(n_3687),
.Y(n_3915)
);

BUFx4_ASAP7_75t_SL g3916 ( 
.A(n_3566),
.Y(n_3916)
);

INVx1_ASAP7_75t_L g3917 ( 
.A(n_3692),
.Y(n_3917)
);

INVx1_ASAP7_75t_L g3918 ( 
.A(n_3681),
.Y(n_3918)
);

INVx1_ASAP7_75t_L g3919 ( 
.A(n_3583),
.Y(n_3919)
);

NOR2xp67_ASAP7_75t_L g3920 ( 
.A(n_3664),
.B(n_84),
.Y(n_3920)
);

AND3x1_ASAP7_75t_SL g3921 ( 
.A(n_3591),
.B(n_85),
.C(n_86),
.Y(n_3921)
);

HB1xp67_ASAP7_75t_L g3922 ( 
.A(n_3687),
.Y(n_3922)
);

INVx4_ASAP7_75t_L g3923 ( 
.A(n_3688),
.Y(n_3923)
);

INVx2_ASAP7_75t_L g3924 ( 
.A(n_3690),
.Y(n_3924)
);

BUFx8_ASAP7_75t_L g3925 ( 
.A(n_3627),
.Y(n_3925)
);

AND2x4_ASAP7_75t_L g3926 ( 
.A(n_3602),
.B(n_85),
.Y(n_3926)
);

BUFx3_ASAP7_75t_L g3927 ( 
.A(n_3688),
.Y(n_3927)
);

INVx3_ASAP7_75t_L g3928 ( 
.A(n_3627),
.Y(n_3928)
);

NAND2xp5_ASAP7_75t_L g3929 ( 
.A(n_3624),
.B(n_87),
.Y(n_3929)
);

NAND2xp5_ASAP7_75t_L g3930 ( 
.A(n_3637),
.B(n_87),
.Y(n_3930)
);

NAND2xp5_ASAP7_75t_L g3931 ( 
.A(n_3675),
.B(n_88),
.Y(n_3931)
);

NAND2xp5_ASAP7_75t_L g3932 ( 
.A(n_3676),
.B(n_88),
.Y(n_3932)
);

AND2x4_ASAP7_75t_L g3933 ( 
.A(n_3673),
.B(n_90),
.Y(n_3933)
);

INVx1_ASAP7_75t_L g3934 ( 
.A(n_3687),
.Y(n_3934)
);

INVxp67_ASAP7_75t_L g3935 ( 
.A(n_3708),
.Y(n_3935)
);

INVx1_ASAP7_75t_L g3936 ( 
.A(n_3690),
.Y(n_3936)
);

INVx2_ASAP7_75t_L g3937 ( 
.A(n_3725),
.Y(n_3937)
);

AOI21xp5_ASAP7_75t_L g3938 ( 
.A1(n_3652),
.A2(n_1909),
.B(n_1887),
.Y(n_3938)
);

AND2x2_ASAP7_75t_L g3939 ( 
.A(n_3627),
.B(n_90),
.Y(n_3939)
);

AND2x2_ASAP7_75t_L g3940 ( 
.A(n_3627),
.B(n_91),
.Y(n_3940)
);

AND2x4_ASAP7_75t_L g3941 ( 
.A(n_3763),
.B(n_92),
.Y(n_3941)
);

OAI21xp5_ASAP7_75t_L g3942 ( 
.A1(n_3744),
.A2(n_93),
.B(n_95),
.Y(n_3942)
);

AND2x2_ASAP7_75t_L g3943 ( 
.A(n_3582),
.B(n_93),
.Y(n_3943)
);

AOI22xp5_ASAP7_75t_L g3944 ( 
.A1(n_3633),
.A2(n_1909),
.B1(n_1918),
.B2(n_1887),
.Y(n_3944)
);

NAND2xp5_ASAP7_75t_L g3945 ( 
.A(n_3680),
.B(n_96),
.Y(n_3945)
);

INVx2_ASAP7_75t_L g3946 ( 
.A(n_3725),
.Y(n_3946)
);

NAND2xp5_ASAP7_75t_L g3947 ( 
.A(n_3682),
.B(n_96),
.Y(n_3947)
);

NAND2xp5_ASAP7_75t_L g3948 ( 
.A(n_3667),
.B(n_97),
.Y(n_3948)
);

INVxp67_ASAP7_75t_L g3949 ( 
.A(n_3567),
.Y(n_3949)
);

NAND2xp5_ASAP7_75t_L g3950 ( 
.A(n_3669),
.B(n_97),
.Y(n_3950)
);

NAND2xp5_ASAP7_75t_L g3951 ( 
.A(n_3571),
.B(n_3581),
.Y(n_3951)
);

AOI21xp5_ASAP7_75t_L g3952 ( 
.A1(n_3652),
.A2(n_1918),
.B(n_1909),
.Y(n_3952)
);

HB1xp67_ASAP7_75t_L g3953 ( 
.A(n_3642),
.Y(n_3953)
);

CKINVDCx5p33_ASAP7_75t_R g3954 ( 
.A(n_3650),
.Y(n_3954)
);

NOR2xp33_ASAP7_75t_L g3955 ( 
.A(n_3660),
.B(n_98),
.Y(n_3955)
);

OAI22xp5_ASAP7_75t_L g3956 ( 
.A1(n_3593),
.A2(n_103),
.B1(n_99),
.B2(n_100),
.Y(n_3956)
);

BUFx2_ASAP7_75t_SL g3957 ( 
.A(n_3765),
.Y(n_3957)
);

INVx1_ASAP7_75t_L g3958 ( 
.A(n_3642),
.Y(n_3958)
);

OR2x6_ASAP7_75t_L g3959 ( 
.A(n_3601),
.B(n_1425),
.Y(n_3959)
);

AOI22xp33_ASAP7_75t_L g3960 ( 
.A1(n_3743),
.A2(n_1918),
.B1(n_1948),
.B2(n_1909),
.Y(n_3960)
);

AOI22xp5_ASAP7_75t_L g3961 ( 
.A1(n_3751),
.A2(n_1948),
.B1(n_1981),
.B2(n_1918),
.Y(n_3961)
);

AOI222xp33_ASAP7_75t_L g3962 ( 
.A1(n_3625),
.A2(n_104),
.B1(n_106),
.B2(n_100),
.C1(n_103),
.C2(n_105),
.Y(n_3962)
);

INVx3_ASAP7_75t_L g3963 ( 
.A(n_3694),
.Y(n_3963)
);

AOI21xp5_ASAP7_75t_L g3964 ( 
.A1(n_3626),
.A2(n_3585),
.B(n_3697),
.Y(n_3964)
);

AND2x2_ASAP7_75t_L g3965 ( 
.A(n_3772),
.B(n_104),
.Y(n_3965)
);

AND2x2_ASAP7_75t_SL g3966 ( 
.A(n_3772),
.B(n_3777),
.Y(n_3966)
);

OR2x2_ASAP7_75t_L g3967 ( 
.A(n_3777),
.B(n_107),
.Y(n_3967)
);

BUFx6f_ASAP7_75t_L g3968 ( 
.A(n_3728),
.Y(n_3968)
);

INVx2_ASAP7_75t_L g3969 ( 
.A(n_3725),
.Y(n_3969)
);

AOI22xp5_ASAP7_75t_L g3970 ( 
.A1(n_3764),
.A2(n_1981),
.B1(n_1992),
.B2(n_1948),
.Y(n_3970)
);

OAI22xp5_ASAP7_75t_L g3971 ( 
.A1(n_3731),
.A2(n_3705),
.B1(n_3733),
.B2(n_3717),
.Y(n_3971)
);

NAND2xp5_ASAP7_75t_L g3972 ( 
.A(n_3756),
.B(n_109),
.Y(n_3972)
);

INVx4_ASAP7_75t_L g3973 ( 
.A(n_3764),
.Y(n_3973)
);

INVx2_ASAP7_75t_L g3974 ( 
.A(n_3730),
.Y(n_3974)
);

INVx5_ASAP7_75t_L g3975 ( 
.A(n_3775),
.Y(n_3975)
);

INVx1_ASAP7_75t_L g3976 ( 
.A(n_3642),
.Y(n_3976)
);

HB1xp67_ASAP7_75t_L g3977 ( 
.A(n_3756),
.Y(n_3977)
);

NAND2xp5_ASAP7_75t_SL g3978 ( 
.A(n_3704),
.B(n_1425),
.Y(n_3978)
);

OR2x2_ASAP7_75t_L g3979 ( 
.A(n_3756),
.B(n_112),
.Y(n_3979)
);

OAI21xp33_ASAP7_75t_L g3980 ( 
.A1(n_3778),
.A2(n_3776),
.B(n_3672),
.Y(n_3980)
);

INVxp67_ASAP7_75t_L g3981 ( 
.A(n_3592),
.Y(n_3981)
);

BUFx3_ASAP7_75t_L g3982 ( 
.A(n_3679),
.Y(n_3982)
);

AOI22xp33_ASAP7_75t_L g3983 ( 
.A1(n_3754),
.A2(n_1981),
.B1(n_1992),
.B2(n_1948),
.Y(n_3983)
);

INVx2_ASAP7_75t_L g3984 ( 
.A(n_3597),
.Y(n_3984)
);

AOI21xp5_ASAP7_75t_L g3985 ( 
.A1(n_3646),
.A2(n_1992),
.B(n_1981),
.Y(n_3985)
);

NAND2xp5_ASAP7_75t_L g3986 ( 
.A(n_3665),
.B(n_112),
.Y(n_3986)
);

INVx1_ASAP7_75t_L g3987 ( 
.A(n_3612),
.Y(n_3987)
);

AOI21xp5_ASAP7_75t_L g3988 ( 
.A1(n_3604),
.A2(n_2005),
.B(n_1992),
.Y(n_3988)
);

OR2x6_ASAP7_75t_L g3989 ( 
.A(n_3644),
.B(n_1432),
.Y(n_3989)
);

AND2x2_ASAP7_75t_L g3990 ( 
.A(n_3696),
.B(n_113),
.Y(n_3990)
);

INVx4_ASAP7_75t_L g3991 ( 
.A(n_3746),
.Y(n_3991)
);

INVx1_ASAP7_75t_L g3992 ( 
.A(n_3609),
.Y(n_3992)
);

OAI22xp5_ASAP7_75t_L g3993 ( 
.A1(n_3750),
.A2(n_116),
.B1(n_114),
.B2(n_115),
.Y(n_3993)
);

AOI22xp5_ASAP7_75t_L g3994 ( 
.A1(n_3640),
.A2(n_2009),
.B1(n_2014),
.B2(n_2005),
.Y(n_3994)
);

AO21x2_ASAP7_75t_L g3995 ( 
.A1(n_3767),
.A2(n_2009),
.B(n_2005),
.Y(n_3995)
);

AOI22xp33_ASAP7_75t_L g3996 ( 
.A1(n_3580),
.A2(n_2009),
.B1(n_2014),
.B2(n_2005),
.Y(n_3996)
);

NAND2x1_ASAP7_75t_L g3997 ( 
.A(n_3668),
.B(n_1432),
.Y(n_3997)
);

NAND2xp5_ASAP7_75t_L g3998 ( 
.A(n_3639),
.B(n_114),
.Y(n_3998)
);

AOI22xp33_ASAP7_75t_L g3999 ( 
.A1(n_3864),
.A2(n_3641),
.B1(n_3588),
.B2(n_3647),
.Y(n_3999)
);

INVx2_ASAP7_75t_L g4000 ( 
.A(n_3851),
.Y(n_4000)
);

OAI22xp33_ASAP7_75t_L g4001 ( 
.A1(n_3782),
.A2(n_3696),
.B1(n_3702),
.B2(n_3722),
.Y(n_4001)
);

CKINVDCx5p33_ASAP7_75t_R g4002 ( 
.A(n_3803),
.Y(n_4002)
);

AOI21xp5_ASAP7_75t_L g4003 ( 
.A1(n_3852),
.A2(n_3736),
.B(n_3659),
.Y(n_4003)
);

OAI22xp5_ASAP7_75t_L g4004 ( 
.A1(n_3908),
.A2(n_120),
.B1(n_117),
.B2(n_118),
.Y(n_4004)
);

INVx3_ASAP7_75t_L g4005 ( 
.A(n_3800),
.Y(n_4005)
);

INVx2_ASAP7_75t_SL g4006 ( 
.A(n_3794),
.Y(n_4006)
);

INVx1_ASAP7_75t_L g4007 ( 
.A(n_3793),
.Y(n_4007)
);

OAI22xp33_ASAP7_75t_L g4008 ( 
.A1(n_3824),
.A2(n_3696),
.B1(n_2014),
.B2(n_2018),
.Y(n_4008)
);

INVx1_ASAP7_75t_L g4009 ( 
.A(n_3784),
.Y(n_4009)
);

BUFx3_ASAP7_75t_L g4010 ( 
.A(n_3850),
.Y(n_4010)
);

AO22x1_ASAP7_75t_L g4011 ( 
.A1(n_3805),
.A2(n_121),
.B1(n_117),
.B2(n_120),
.Y(n_4011)
);

INVx6_ASAP7_75t_L g4012 ( 
.A(n_3882),
.Y(n_4012)
);

NAND2xp5_ASAP7_75t_L g4013 ( 
.A(n_3790),
.B(n_3654),
.Y(n_4013)
);

CKINVDCx6p67_ASAP7_75t_R g4014 ( 
.A(n_3843),
.Y(n_4014)
);

HB1xp67_ASAP7_75t_L g4015 ( 
.A(n_3780),
.Y(n_4015)
);

AOI22xp33_ASAP7_75t_L g4016 ( 
.A1(n_3792),
.A2(n_3651),
.B1(n_3623),
.B2(n_3594),
.Y(n_4016)
);

NOR2x1_ASAP7_75t_L g4017 ( 
.A(n_3910),
.B(n_3768),
.Y(n_4017)
);

INVx1_ASAP7_75t_L g4018 ( 
.A(n_3795),
.Y(n_4018)
);

BUFx6f_ASAP7_75t_L g4019 ( 
.A(n_3859),
.Y(n_4019)
);

INVx2_ASAP7_75t_L g4020 ( 
.A(n_3799),
.Y(n_4020)
);

INVx6_ASAP7_75t_L g4021 ( 
.A(n_3882),
.Y(n_4021)
);

INVx1_ASAP7_75t_L g4022 ( 
.A(n_3809),
.Y(n_4022)
);

INVx1_ASAP7_75t_L g4023 ( 
.A(n_3848),
.Y(n_4023)
);

CKINVDCx11_ASAP7_75t_R g4024 ( 
.A(n_3812),
.Y(n_4024)
);

INVxp67_ASAP7_75t_SL g4025 ( 
.A(n_3977),
.Y(n_4025)
);

INVx1_ASAP7_75t_SL g4026 ( 
.A(n_3832),
.Y(n_4026)
);

BUFx2_ASAP7_75t_L g4027 ( 
.A(n_3796),
.Y(n_4027)
);

AOI22xp5_ASAP7_75t_SL g4028 ( 
.A1(n_3954),
.A2(n_123),
.B1(n_121),
.B2(n_122),
.Y(n_4028)
);

BUFx2_ASAP7_75t_L g4029 ( 
.A(n_3836),
.Y(n_4029)
);

INVx1_ASAP7_75t_L g4030 ( 
.A(n_3856),
.Y(n_4030)
);

INVx6_ASAP7_75t_L g4031 ( 
.A(n_3800),
.Y(n_4031)
);

AOI22xp33_ASAP7_75t_L g4032 ( 
.A1(n_3872),
.A2(n_3693),
.B1(n_3677),
.B2(n_3656),
.Y(n_4032)
);

AOI22xp5_ASAP7_75t_L g4033 ( 
.A1(n_3834),
.A2(n_2014),
.B1(n_2018),
.B2(n_2009),
.Y(n_4033)
);

INVx1_ASAP7_75t_L g4034 ( 
.A(n_3788),
.Y(n_4034)
);

BUFx2_ASAP7_75t_L g4035 ( 
.A(n_3815),
.Y(n_4035)
);

INVx1_ASAP7_75t_L g4036 ( 
.A(n_3861),
.Y(n_4036)
);

CKINVDCx11_ASAP7_75t_R g4037 ( 
.A(n_3797),
.Y(n_4037)
);

OAI21xp33_ASAP7_75t_L g4038 ( 
.A1(n_3955),
.A2(n_122),
.B(n_123),
.Y(n_4038)
);

INVx2_ASAP7_75t_L g4039 ( 
.A(n_3818),
.Y(n_4039)
);

INVx1_ASAP7_75t_SL g4040 ( 
.A(n_3807),
.Y(n_4040)
);

INVx3_ASAP7_75t_L g4041 ( 
.A(n_3854),
.Y(n_4041)
);

AOI22xp33_ASAP7_75t_L g4042 ( 
.A1(n_3979),
.A2(n_2026),
.B1(n_2028),
.B2(n_2018),
.Y(n_4042)
);

INVx1_ASAP7_75t_L g4043 ( 
.A(n_3847),
.Y(n_4043)
);

INVx1_ASAP7_75t_L g4044 ( 
.A(n_3907),
.Y(n_4044)
);

INVx3_ASAP7_75t_L g4045 ( 
.A(n_3854),
.Y(n_4045)
);

CKINVDCx20_ASAP7_75t_R g4046 ( 
.A(n_3786),
.Y(n_4046)
);

BUFx4_ASAP7_75t_SL g4047 ( 
.A(n_3927),
.Y(n_4047)
);

NAND2xp5_ASAP7_75t_L g4048 ( 
.A(n_3898),
.B(n_124),
.Y(n_4048)
);

CKINVDCx20_ASAP7_75t_R g4049 ( 
.A(n_3804),
.Y(n_4049)
);

INVx1_ASAP7_75t_L g4050 ( 
.A(n_3866),
.Y(n_4050)
);

INVx2_ASAP7_75t_L g4051 ( 
.A(n_3835),
.Y(n_4051)
);

INVx8_ASAP7_75t_L g4052 ( 
.A(n_3783),
.Y(n_4052)
);

CKINVDCx11_ASAP7_75t_R g4053 ( 
.A(n_3845),
.Y(n_4053)
);

OAI22xp33_ASAP7_75t_L g4054 ( 
.A1(n_3849),
.A2(n_2026),
.B1(n_2028),
.B2(n_2018),
.Y(n_4054)
);

BUFx6f_ASAP7_75t_L g4055 ( 
.A(n_3859),
.Y(n_4055)
);

OAI22xp5_ASAP7_75t_L g4056 ( 
.A1(n_3884),
.A2(n_128),
.B1(n_125),
.B2(n_126),
.Y(n_4056)
);

OAI22xp33_ASAP7_75t_L g4057 ( 
.A1(n_3972),
.A2(n_3991),
.B1(n_3890),
.B2(n_3878),
.Y(n_4057)
);

AOI22xp33_ASAP7_75t_L g4058 ( 
.A1(n_3991),
.A2(n_2028),
.B1(n_2050),
.B2(n_2026),
.Y(n_4058)
);

AND2x2_ASAP7_75t_L g4059 ( 
.A(n_3838),
.B(n_126),
.Y(n_4059)
);

INVx2_ASAP7_75t_L g4060 ( 
.A(n_3840),
.Y(n_4060)
);

CKINVDCx20_ASAP7_75t_R g4061 ( 
.A(n_3869),
.Y(n_4061)
);

AOI22xp33_ASAP7_75t_L g4062 ( 
.A1(n_3942),
.A2(n_2028),
.B1(n_2050),
.B2(n_2026),
.Y(n_4062)
);

BUFx3_ASAP7_75t_L g4063 ( 
.A(n_3789),
.Y(n_4063)
);

INVx1_ASAP7_75t_L g4064 ( 
.A(n_3905),
.Y(n_4064)
);

INVx2_ASAP7_75t_L g4065 ( 
.A(n_3855),
.Y(n_4065)
);

AOI22xp33_ASAP7_75t_L g4066 ( 
.A1(n_3935),
.A2(n_3949),
.B1(n_3951),
.B2(n_3881),
.Y(n_4066)
);

BUFx8_ASAP7_75t_SL g4067 ( 
.A(n_3810),
.Y(n_4067)
);

OAI21xp5_ASAP7_75t_SL g4068 ( 
.A1(n_3816),
.A2(n_129),
.B(n_131),
.Y(n_4068)
);

INVx4_ASAP7_75t_L g4069 ( 
.A(n_3923),
.Y(n_4069)
);

OAI22xp33_ASAP7_75t_L g4070 ( 
.A1(n_3829),
.A2(n_2062),
.B1(n_2066),
.B2(n_2050),
.Y(n_4070)
);

BUFx2_ASAP7_75t_SL g4071 ( 
.A(n_3920),
.Y(n_4071)
);

INVx2_ASAP7_75t_L g4072 ( 
.A(n_3917),
.Y(n_4072)
);

NAND2xp5_ASAP7_75t_L g4073 ( 
.A(n_3906),
.B(n_129),
.Y(n_4073)
);

INVx1_ASAP7_75t_L g4074 ( 
.A(n_3875),
.Y(n_4074)
);

INVx1_ASAP7_75t_L g4075 ( 
.A(n_3841),
.Y(n_4075)
);

INVx1_ASAP7_75t_L g4076 ( 
.A(n_3791),
.Y(n_4076)
);

INVx2_ASAP7_75t_L g4077 ( 
.A(n_3827),
.Y(n_4077)
);

INVx1_ASAP7_75t_L g4078 ( 
.A(n_3876),
.Y(n_4078)
);

INVx1_ASAP7_75t_SL g4079 ( 
.A(n_3837),
.Y(n_4079)
);

BUFx6f_ASAP7_75t_L g4080 ( 
.A(n_3859),
.Y(n_4080)
);

INVx2_ASAP7_75t_L g4081 ( 
.A(n_3827),
.Y(n_4081)
);

AOI22xp33_ASAP7_75t_L g4082 ( 
.A1(n_3962),
.A2(n_2062),
.B1(n_2066),
.B2(n_2050),
.Y(n_4082)
);

OAI21xp33_ASAP7_75t_L g4083 ( 
.A1(n_3833),
.A2(n_131),
.B(n_132),
.Y(n_4083)
);

INVx6_ASAP7_75t_L g4084 ( 
.A(n_3923),
.Y(n_4084)
);

CKINVDCx11_ASAP7_75t_R g4085 ( 
.A(n_3845),
.Y(n_4085)
);

AOI22xp5_ASAP7_75t_L g4086 ( 
.A1(n_3956),
.A2(n_2066),
.B1(n_2071),
.B2(n_2062),
.Y(n_4086)
);

INVxp67_ASAP7_75t_SL g4087 ( 
.A(n_3915),
.Y(n_4087)
);

BUFx12f_ASAP7_75t_L g4088 ( 
.A(n_3879),
.Y(n_4088)
);

INVx1_ASAP7_75t_SL g4089 ( 
.A(n_3781),
.Y(n_4089)
);

AOI22xp33_ASAP7_75t_SL g4090 ( 
.A1(n_3990),
.A2(n_134),
.B1(n_132),
.B2(n_133),
.Y(n_4090)
);

CKINVDCx11_ASAP7_75t_R g4091 ( 
.A(n_3893),
.Y(n_4091)
);

AOI22xp33_ASAP7_75t_L g4092 ( 
.A1(n_3817),
.A2(n_2066),
.B1(n_2071),
.B2(n_2062),
.Y(n_4092)
);

OAI22xp33_ASAP7_75t_L g4093 ( 
.A1(n_3787),
.A2(n_2071),
.B1(n_2095),
.B2(n_137),
.Y(n_4093)
);

HB1xp67_ASAP7_75t_L g4094 ( 
.A(n_3965),
.Y(n_4094)
);

OAI21xp5_ASAP7_75t_SL g4095 ( 
.A1(n_3801),
.A2(n_3830),
.B(n_3814),
.Y(n_4095)
);

OAI22xp5_ASAP7_75t_L g4096 ( 
.A1(n_3823),
.A2(n_140),
.B1(n_133),
.B2(n_136),
.Y(n_4096)
);

INVx1_ASAP7_75t_L g4097 ( 
.A(n_3876),
.Y(n_4097)
);

INVx6_ASAP7_75t_L g4098 ( 
.A(n_3925),
.Y(n_4098)
);

INVx1_ASAP7_75t_SL g4099 ( 
.A(n_3785),
.Y(n_4099)
);

BUFx3_ASAP7_75t_L g4100 ( 
.A(n_3892),
.Y(n_4100)
);

OAI22xp5_ASAP7_75t_L g4101 ( 
.A1(n_3823),
.A2(n_142),
.B1(n_136),
.B2(n_140),
.Y(n_4101)
);

INVx2_ASAP7_75t_SL g4102 ( 
.A(n_3885),
.Y(n_4102)
);

CKINVDCx11_ASAP7_75t_R g4103 ( 
.A(n_3893),
.Y(n_4103)
);

OR2x2_ASAP7_75t_L g4104 ( 
.A(n_3894),
.B(n_3928),
.Y(n_4104)
);

INVx2_ASAP7_75t_L g4105 ( 
.A(n_3967),
.Y(n_4105)
);

BUFx2_ASAP7_75t_L g4106 ( 
.A(n_3925),
.Y(n_4106)
);

AOI22xp33_ASAP7_75t_L g4107 ( 
.A1(n_3874),
.A2(n_2071),
.B1(n_1477),
.B2(n_1485),
.Y(n_4107)
);

INVx1_ASAP7_75t_L g4108 ( 
.A(n_3802),
.Y(n_4108)
);

AOI22xp33_ASAP7_75t_L g4109 ( 
.A1(n_3943),
.A2(n_1477),
.B1(n_1485),
.B2(n_1472),
.Y(n_4109)
);

OAI22xp5_ASAP7_75t_L g4110 ( 
.A1(n_3842),
.A2(n_145),
.B1(n_143),
.B2(n_144),
.Y(n_4110)
);

AOI22xp33_ASAP7_75t_L g4111 ( 
.A1(n_3821),
.A2(n_1477),
.B1(n_1485),
.B2(n_1472),
.Y(n_4111)
);

AOI22xp33_ASAP7_75t_SL g4112 ( 
.A1(n_3939),
.A2(n_147),
.B1(n_144),
.B2(n_146),
.Y(n_4112)
);

INVx1_ASAP7_75t_SL g4113 ( 
.A(n_3831),
.Y(n_4113)
);

INVx1_ASAP7_75t_L g4114 ( 
.A(n_3958),
.Y(n_4114)
);

INVx6_ASAP7_75t_L g4115 ( 
.A(n_3892),
.Y(n_4115)
);

OAI22xp5_ASAP7_75t_L g4116 ( 
.A1(n_3842),
.A2(n_3865),
.B1(n_3798),
.B2(n_3926),
.Y(n_4116)
);

INVx3_ASAP7_75t_L g4117 ( 
.A(n_3894),
.Y(n_4117)
);

INVx1_ASAP7_75t_L g4118 ( 
.A(n_3976),
.Y(n_4118)
);

OAI22xp33_ASAP7_75t_L g4119 ( 
.A1(n_3961),
.A2(n_150),
.B1(n_148),
.B2(n_149),
.Y(n_4119)
);

BUFx6f_ASAP7_75t_L g4120 ( 
.A(n_3893),
.Y(n_4120)
);

INVx1_ASAP7_75t_L g4121 ( 
.A(n_3828),
.Y(n_4121)
);

INVxp67_ASAP7_75t_SL g4122 ( 
.A(n_3922),
.Y(n_4122)
);

CKINVDCx5p33_ASAP7_75t_R g4123 ( 
.A(n_3880),
.Y(n_4123)
);

HB1xp67_ASAP7_75t_L g4124 ( 
.A(n_3981),
.Y(n_4124)
);

INVx1_ASAP7_75t_L g4125 ( 
.A(n_3828),
.Y(n_4125)
);

BUFx3_ASAP7_75t_L g4126 ( 
.A(n_3860),
.Y(n_4126)
);

INVx2_ASAP7_75t_L g4127 ( 
.A(n_3914),
.Y(n_4127)
);

INVx2_ASAP7_75t_L g4128 ( 
.A(n_3924),
.Y(n_4128)
);

OAI22xp5_ASAP7_75t_L g4129 ( 
.A1(n_3926),
.A2(n_153),
.B1(n_151),
.B2(n_152),
.Y(n_4129)
);

AOI22xp33_ASAP7_75t_L g4130 ( 
.A1(n_3825),
.A2(n_1485),
.B1(n_1487),
.B2(n_1472),
.Y(n_4130)
);

BUFx10_ASAP7_75t_L g4131 ( 
.A(n_3912),
.Y(n_4131)
);

INVx6_ASAP7_75t_L g4132 ( 
.A(n_3885),
.Y(n_4132)
);

CKINVDCx5p33_ASAP7_75t_R g4133 ( 
.A(n_3916),
.Y(n_4133)
);

CKINVDCx5p33_ASAP7_75t_R g4134 ( 
.A(n_3883),
.Y(n_4134)
);

BUFx2_ASAP7_75t_L g4135 ( 
.A(n_3928),
.Y(n_4135)
);

INVx2_ASAP7_75t_L g4136 ( 
.A(n_3886),
.Y(n_4136)
);

CKINVDCx5p33_ASAP7_75t_R g4137 ( 
.A(n_3867),
.Y(n_4137)
);

INVx2_ASAP7_75t_L g4138 ( 
.A(n_3828),
.Y(n_4138)
);

CKINVDCx11_ASAP7_75t_R g4139 ( 
.A(n_3968),
.Y(n_4139)
);

AOI22xp5_ASAP7_75t_L g4140 ( 
.A1(n_3911),
.A2(n_1499),
.B1(n_1507),
.B2(n_1487),
.Y(n_4140)
);

INVx1_ASAP7_75t_L g4141 ( 
.A(n_3953),
.Y(n_4141)
);

AOI22xp5_ASAP7_75t_SL g4142 ( 
.A1(n_3940),
.A2(n_156),
.B1(n_153),
.B2(n_154),
.Y(n_4142)
);

AOI21xp5_ASAP7_75t_L g4143 ( 
.A1(n_3811),
.A2(n_1499),
.B(n_1487),
.Y(n_4143)
);

INVx1_ASAP7_75t_L g4144 ( 
.A(n_3887),
.Y(n_4144)
);

AOI22xp33_ASAP7_75t_L g4145 ( 
.A1(n_3978),
.A2(n_3959),
.B1(n_3873),
.B2(n_3891),
.Y(n_4145)
);

BUFx2_ASAP7_75t_SL g4146 ( 
.A(n_3853),
.Y(n_4146)
);

BUFx6f_ASAP7_75t_L g4147 ( 
.A(n_3968),
.Y(n_4147)
);

AOI22xp5_ASAP7_75t_SL g4148 ( 
.A1(n_3806),
.A2(n_158),
.B1(n_156),
.B2(n_157),
.Y(n_4148)
);

BUFx6f_ASAP7_75t_L g4149 ( 
.A(n_3968),
.Y(n_4149)
);

OAI22xp33_ASAP7_75t_L g4150 ( 
.A1(n_3959),
.A2(n_162),
.B1(n_159),
.B2(n_160),
.Y(n_4150)
);

BUFx4_ASAP7_75t_R g4151 ( 
.A(n_3921),
.Y(n_4151)
);

INVx4_ASAP7_75t_L g4152 ( 
.A(n_3912),
.Y(n_4152)
);

INVx2_ASAP7_75t_L g4153 ( 
.A(n_3896),
.Y(n_4153)
);

OAI22xp5_ASAP7_75t_L g4154 ( 
.A1(n_3839),
.A2(n_163),
.B1(n_159),
.B2(n_160),
.Y(n_4154)
);

INVx1_ASAP7_75t_L g4155 ( 
.A(n_3888),
.Y(n_4155)
);

INVx4_ASAP7_75t_L g4156 ( 
.A(n_3941),
.Y(n_4156)
);

AOI22xp33_ASAP7_75t_L g4157 ( 
.A1(n_3822),
.A2(n_1499),
.B1(n_1507),
.B2(n_1487),
.Y(n_4157)
);

AOI22xp33_ASAP7_75t_L g4158 ( 
.A1(n_3909),
.A2(n_1507),
.B1(n_1513),
.B2(n_1499),
.Y(n_4158)
);

AOI22xp5_ASAP7_75t_L g4159 ( 
.A1(n_3993),
.A2(n_1513),
.B1(n_1507),
.B2(n_165),
.Y(n_4159)
);

INVx2_ASAP7_75t_L g4160 ( 
.A(n_3937),
.Y(n_4160)
);

CKINVDCx6p67_ASAP7_75t_R g4161 ( 
.A(n_3900),
.Y(n_4161)
);

BUFx6f_ASAP7_75t_L g4162 ( 
.A(n_3871),
.Y(n_4162)
);

OAI22xp5_ASAP7_75t_L g4163 ( 
.A1(n_3846),
.A2(n_166),
.B1(n_163),
.B2(n_164),
.Y(n_4163)
);

INVx3_ASAP7_75t_L g4164 ( 
.A(n_3982),
.Y(n_4164)
);

BUFx8_ASAP7_75t_SL g4165 ( 
.A(n_3901),
.Y(n_4165)
);

BUFx10_ASAP7_75t_L g4166 ( 
.A(n_3941),
.Y(n_4166)
);

OAI22xp5_ASAP7_75t_L g4167 ( 
.A1(n_3820),
.A2(n_168),
.B1(n_166),
.B2(n_167),
.Y(n_4167)
);

INVx1_ASAP7_75t_L g4168 ( 
.A(n_3998),
.Y(n_4168)
);

AOI22xp33_ASAP7_75t_L g4169 ( 
.A1(n_3933),
.A2(n_1513),
.B1(n_1520),
.B2(n_1514),
.Y(n_4169)
);

INVx2_ASAP7_75t_SL g4170 ( 
.A(n_3826),
.Y(n_4170)
);

CKINVDCx20_ASAP7_75t_R g4171 ( 
.A(n_3903),
.Y(n_4171)
);

AOI21x1_ASAP7_75t_SL g4172 ( 
.A1(n_4124),
.A2(n_3950),
.B(n_3930),
.Y(n_4172)
);

NAND2xp5_ASAP7_75t_L g4173 ( 
.A(n_4168),
.B(n_3877),
.Y(n_4173)
);

OAI22xp5_ASAP7_75t_L g4174 ( 
.A1(n_4068),
.A2(n_3986),
.B1(n_3929),
.B2(n_3932),
.Y(n_4174)
);

A2O1A1Ixp33_ASAP7_75t_L g4175 ( 
.A1(n_4038),
.A2(n_4083),
.B(n_4028),
.C(n_4095),
.Y(n_4175)
);

INVx1_ASAP7_75t_L g4176 ( 
.A(n_4007),
.Y(n_4176)
);

CKINVDCx20_ASAP7_75t_R g4177 ( 
.A(n_4024),
.Y(n_4177)
);

AND2x2_ASAP7_75t_L g4178 ( 
.A(n_4027),
.B(n_3918),
.Y(n_4178)
);

NAND2xp5_ASAP7_75t_L g4179 ( 
.A(n_4043),
.B(n_3931),
.Y(n_4179)
);

OR2x2_ASAP7_75t_L g4180 ( 
.A(n_4094),
.B(n_3934),
.Y(n_4180)
);

AND2x4_ASAP7_75t_L g4181 ( 
.A(n_4156),
.B(n_3868),
.Y(n_4181)
);

INVx2_ASAP7_75t_L g4182 ( 
.A(n_4072),
.Y(n_4182)
);

OR2x2_ASAP7_75t_L g4183 ( 
.A(n_4074),
.B(n_3936),
.Y(n_4183)
);

OA21x2_ASAP7_75t_L g4184 ( 
.A1(n_4077),
.A2(n_3969),
.B(n_3946),
.Y(n_4184)
);

OA21x2_ASAP7_75t_L g4185 ( 
.A1(n_4081),
.A2(n_3889),
.B(n_3844),
.Y(n_4185)
);

CKINVDCx8_ASAP7_75t_R g4186 ( 
.A(n_4071),
.Y(n_4186)
);

OR2x2_ASAP7_75t_L g4187 ( 
.A(n_4044),
.B(n_3919),
.Y(n_4187)
);

AOI21xp5_ASAP7_75t_L g4188 ( 
.A1(n_4057),
.A2(n_3808),
.B(n_3870),
.Y(n_4188)
);

O2A1O1Ixp5_ASAP7_75t_L g4189 ( 
.A1(n_4011),
.A2(n_3947),
.B(n_3948),
.C(n_3945),
.Y(n_4189)
);

AND2x2_ASAP7_75t_L g4190 ( 
.A(n_4035),
.B(n_3966),
.Y(n_4190)
);

AOI21xp5_ASAP7_75t_L g4191 ( 
.A1(n_4038),
.A2(n_3870),
.B(n_3964),
.Y(n_4191)
);

A2O1A1Ixp33_ASAP7_75t_L g4192 ( 
.A1(n_4083),
.A2(n_3813),
.B(n_3933),
.C(n_3960),
.Y(n_4192)
);

AOI21xp5_ASAP7_75t_L g4193 ( 
.A1(n_4003),
.A2(n_3971),
.B(n_3857),
.Y(n_4193)
);

AOI21xp5_ASAP7_75t_L g4194 ( 
.A1(n_4052),
.A2(n_3989),
.B(n_3862),
.Y(n_4194)
);

NAND2xp5_ASAP7_75t_L g4195 ( 
.A(n_4108),
.B(n_3963),
.Y(n_4195)
);

OA21x2_ASAP7_75t_L g4196 ( 
.A1(n_4141),
.A2(n_3980),
.B(n_3974),
.Y(n_4196)
);

OA21x2_ASAP7_75t_L g4197 ( 
.A1(n_4087),
.A2(n_4122),
.B(n_4025),
.Y(n_4197)
);

INVx3_ASAP7_75t_L g4198 ( 
.A(n_4132),
.Y(n_4198)
);

AOI221xp5_ASAP7_75t_L g4199 ( 
.A1(n_4056),
.A2(n_3895),
.B1(n_3973),
.B2(n_3957),
.C(n_3992),
.Y(n_4199)
);

AND2x2_ASAP7_75t_L g4200 ( 
.A(n_4015),
.B(n_3987),
.Y(n_4200)
);

NAND2xp5_ASAP7_75t_L g4201 ( 
.A(n_4009),
.B(n_3963),
.Y(n_4201)
);

NAND2xp5_ASAP7_75t_L g4202 ( 
.A(n_4026),
.B(n_3973),
.Y(n_4202)
);

OAI22xp5_ASAP7_75t_L g4203 ( 
.A1(n_4090),
.A2(n_3897),
.B1(n_3944),
.B2(n_3970),
.Y(n_4203)
);

AND2x2_ASAP7_75t_L g4204 ( 
.A(n_4029),
.B(n_3984),
.Y(n_4204)
);

NOR2xp67_ASAP7_75t_L g4205 ( 
.A(n_4164),
.B(n_3975),
.Y(n_4205)
);

BUFx3_ASAP7_75t_L g4206 ( 
.A(n_4010),
.Y(n_4206)
);

AND2x2_ASAP7_75t_L g4207 ( 
.A(n_4075),
.B(n_3989),
.Y(n_4207)
);

NOR2xp67_ASAP7_75t_L g4208 ( 
.A(n_4164),
.B(n_3975),
.Y(n_4208)
);

HB1xp67_ASAP7_75t_L g4209 ( 
.A(n_4034),
.Y(n_4209)
);

NAND2xp5_ASAP7_75t_L g4210 ( 
.A(n_4064),
.B(n_3975),
.Y(n_4210)
);

OAI22xp5_ASAP7_75t_L g4211 ( 
.A1(n_4161),
.A2(n_3994),
.B1(n_3863),
.B2(n_3826),
.Y(n_4211)
);

AND2x2_ASAP7_75t_L g4212 ( 
.A(n_4146),
.B(n_3783),
.Y(n_4212)
);

CKINVDCx5p33_ASAP7_75t_R g4213 ( 
.A(n_4002),
.Y(n_4213)
);

NOR2xp67_ASAP7_75t_L g4214 ( 
.A(n_4156),
.B(n_4069),
.Y(n_4214)
);

NOR2x1_ASAP7_75t_SL g4215 ( 
.A(n_4152),
.B(n_3863),
.Y(n_4215)
);

AND2x4_ASAP7_75t_L g4216 ( 
.A(n_4152),
.B(n_3783),
.Y(n_4216)
);

OAI22xp5_ASAP7_75t_L g4217 ( 
.A1(n_4066),
.A2(n_3996),
.B1(n_3997),
.B2(n_3983),
.Y(n_4217)
);

OAI22xp5_ASAP7_75t_L g4218 ( 
.A1(n_4145),
.A2(n_3899),
.B1(n_3904),
.B2(n_3858),
.Y(n_4218)
);

HB1xp67_ASAP7_75t_L g4219 ( 
.A(n_4036),
.Y(n_4219)
);

AOI21x1_ASAP7_75t_SL g4220 ( 
.A1(n_4013),
.A2(n_167),
.B(n_168),
.Y(n_4220)
);

O2A1O1Ixp5_ASAP7_75t_L g4221 ( 
.A1(n_4116),
.A2(n_3985),
.B(n_3988),
.C(n_3913),
.Y(n_4221)
);

OR2x2_ASAP7_75t_L g4222 ( 
.A(n_4105),
.B(n_3995),
.Y(n_4222)
);

AND2x4_ASAP7_75t_L g4223 ( 
.A(n_4102),
.B(n_3783),
.Y(n_4223)
);

AOI21x1_ASAP7_75t_SL g4224 ( 
.A1(n_4059),
.A2(n_170),
.B(n_171),
.Y(n_4224)
);

AOI21x1_ASAP7_75t_SL g4225 ( 
.A1(n_4048),
.A2(n_172),
.B(n_173),
.Y(n_4225)
);

INVx3_ASAP7_75t_L g4226 ( 
.A(n_4132),
.Y(n_4226)
);

OR2x2_ASAP7_75t_L g4227 ( 
.A(n_4076),
.B(n_3938),
.Y(n_4227)
);

NAND2xp5_ASAP7_75t_L g4228 ( 
.A(n_4022),
.B(n_3819),
.Y(n_4228)
);

AND2x2_ASAP7_75t_L g4229 ( 
.A(n_4041),
.B(n_3819),
.Y(n_4229)
);

AOI221x1_ASAP7_75t_SL g4230 ( 
.A1(n_4004),
.A2(n_175),
.B1(n_172),
.B2(n_174),
.C(n_176),
.Y(n_4230)
);

INVx1_ASAP7_75t_L g4231 ( 
.A(n_4018),
.Y(n_4231)
);

INVx1_ASAP7_75t_L g4232 ( 
.A(n_4023),
.Y(n_4232)
);

INVx1_ASAP7_75t_L g4233 ( 
.A(n_4030),
.Y(n_4233)
);

AOI21xp5_ASAP7_75t_SL g4234 ( 
.A1(n_4133),
.A2(n_3902),
.B(n_3952),
.Y(n_4234)
);

AND2x2_ASAP7_75t_L g4235 ( 
.A(n_4041),
.B(n_3819),
.Y(n_4235)
);

NAND2xp5_ASAP7_75t_L g4236 ( 
.A(n_4078),
.B(n_4097),
.Y(n_4236)
);

INVx2_ASAP7_75t_L g4237 ( 
.A(n_4000),
.Y(n_4237)
);

BUFx2_ASAP7_75t_L g4238 ( 
.A(n_4045),
.Y(n_4238)
);

NAND2xp5_ASAP7_75t_L g4239 ( 
.A(n_4113),
.B(n_4089),
.Y(n_4239)
);

CKINVDCx12_ASAP7_75t_R g4240 ( 
.A(n_4142),
.Y(n_4240)
);

AND2x4_ASAP7_75t_L g4241 ( 
.A(n_4100),
.B(n_3819),
.Y(n_4241)
);

OR2x2_ASAP7_75t_L g4242 ( 
.A(n_4099),
.B(n_4045),
.Y(n_4242)
);

AND2x2_ASAP7_75t_L g4243 ( 
.A(n_4079),
.B(n_174),
.Y(n_4243)
);

BUFx2_ASAP7_75t_L g4244 ( 
.A(n_4063),
.Y(n_4244)
);

OA21x2_ASAP7_75t_L g4245 ( 
.A1(n_4121),
.A2(n_177),
.B(n_178),
.Y(n_4245)
);

AOI21xp5_ASAP7_75t_L g4246 ( 
.A1(n_4052),
.A2(n_1513),
.B(n_1520),
.Y(n_4246)
);

O2A1O1Ixp33_ASAP7_75t_L g4247 ( 
.A1(n_4163),
.A2(n_181),
.B(n_177),
.C(n_180),
.Y(n_4247)
);

AND2x4_ASAP7_75t_L g4248 ( 
.A(n_4005),
.B(n_4117),
.Y(n_4248)
);

AOI221xp5_ASAP7_75t_L g4249 ( 
.A1(n_4154),
.A2(n_180),
.B1(n_184),
.B2(n_185),
.C(n_186),
.Y(n_4249)
);

INVx2_ASAP7_75t_L g4250 ( 
.A(n_4020),
.Y(n_4250)
);

NAND2xp5_ASAP7_75t_L g4251 ( 
.A(n_4136),
.B(n_184),
.Y(n_4251)
);

HB1xp67_ASAP7_75t_L g4252 ( 
.A(n_4135),
.Y(n_4252)
);

AND2x2_ASAP7_75t_L g4253 ( 
.A(n_4117),
.B(n_186),
.Y(n_4253)
);

AOI21xp5_ASAP7_75t_SL g4254 ( 
.A1(n_4140),
.A2(n_188),
.B(n_189),
.Y(n_4254)
);

INVx3_ASAP7_75t_SL g4255 ( 
.A(n_4014),
.Y(n_4255)
);

INVx1_ASAP7_75t_L g4256 ( 
.A(n_4050),
.Y(n_4256)
);

AOI21xp5_ASAP7_75t_SL g4257 ( 
.A1(n_4140),
.A2(n_188),
.B(n_189),
.Y(n_4257)
);

OAI22xp5_ASAP7_75t_L g4258 ( 
.A1(n_4112),
.A2(n_192),
.B1(n_190),
.B2(n_191),
.Y(n_4258)
);

HB1xp67_ASAP7_75t_L g4259 ( 
.A(n_4153),
.Y(n_4259)
);

AOI21x1_ASAP7_75t_SL g4260 ( 
.A1(n_4073),
.A2(n_190),
.B(n_191),
.Y(n_4260)
);

INVx2_ASAP7_75t_L g4261 ( 
.A(n_4039),
.Y(n_4261)
);

OAI22xp5_ASAP7_75t_L g4262 ( 
.A1(n_4159),
.A2(n_194),
.B1(n_192),
.B2(n_193),
.Y(n_4262)
);

A2O1A1Ixp33_ASAP7_75t_L g4263 ( 
.A1(n_4148),
.A2(n_196),
.B(n_194),
.C(n_195),
.Y(n_4263)
);

O2A1O1Ixp33_ASAP7_75t_L g4264 ( 
.A1(n_4167),
.A2(n_198),
.B(n_195),
.C(n_197),
.Y(n_4264)
);

AOI21xp5_ASAP7_75t_L g4265 ( 
.A1(n_4052),
.A2(n_1525),
.B(n_1520),
.Y(n_4265)
);

AOI21x1_ASAP7_75t_SL g4266 ( 
.A1(n_4151),
.A2(n_197),
.B(n_198),
.Y(n_4266)
);

A2O1A1Ixp33_ASAP7_75t_L g4267 ( 
.A1(n_4126),
.A2(n_203),
.B(n_200),
.C(n_202),
.Y(n_4267)
);

OR2x2_ASAP7_75t_L g4268 ( 
.A(n_4104),
.B(n_200),
.Y(n_4268)
);

AND2x2_ASAP7_75t_L g4269 ( 
.A(n_4006),
.B(n_203),
.Y(n_4269)
);

AOI21xp5_ASAP7_75t_L g4270 ( 
.A1(n_4001),
.A2(n_1525),
.B(n_1520),
.Y(n_4270)
);

AOI21x1_ASAP7_75t_SL g4271 ( 
.A1(n_4047),
.A2(n_204),
.B(n_207),
.Y(n_4271)
);

A2O1A1Ixp33_ASAP7_75t_L g4272 ( 
.A1(n_4082),
.A2(n_210),
.B(n_208),
.C(n_209),
.Y(n_4272)
);

HB1xp67_ASAP7_75t_L g4273 ( 
.A(n_4114),
.Y(n_4273)
);

NAND2xp5_ASAP7_75t_L g4274 ( 
.A(n_4005),
.B(n_208),
.Y(n_4274)
);

AOI21xp5_ASAP7_75t_L g4275 ( 
.A1(n_4119),
.A2(n_1542),
.B(n_1525),
.Y(n_4275)
);

CKINVDCx5p33_ASAP7_75t_R g4276 ( 
.A(n_4037),
.Y(n_4276)
);

OAI22xp5_ASAP7_75t_L g4277 ( 
.A1(n_4159),
.A2(n_4062),
.B1(n_4033),
.B2(n_4115),
.Y(n_4277)
);

OR2x2_ASAP7_75t_L g4278 ( 
.A(n_4118),
.B(n_209),
.Y(n_4278)
);

AND2x2_ASAP7_75t_L g4279 ( 
.A(n_4040),
.B(n_4106),
.Y(n_4279)
);

A2O1A1Ixp33_ASAP7_75t_L g4280 ( 
.A1(n_4137),
.A2(n_212),
.B(n_210),
.C(n_211),
.Y(n_4280)
);

AND2x2_ASAP7_75t_L g4281 ( 
.A(n_4053),
.B(n_213),
.Y(n_4281)
);

AND2x2_ASAP7_75t_L g4282 ( 
.A(n_4085),
.B(n_213),
.Y(n_4282)
);

NAND2xp5_ASAP7_75t_L g4283 ( 
.A(n_4166),
.B(n_214),
.Y(n_4283)
);

AOI21xp5_ASAP7_75t_L g4284 ( 
.A1(n_4143),
.A2(n_1542),
.B(n_1525),
.Y(n_4284)
);

INVx2_ASAP7_75t_L g4285 ( 
.A(n_4051),
.Y(n_4285)
);

A2O1A1Ixp33_ASAP7_75t_L g4286 ( 
.A1(n_4129),
.A2(n_216),
.B(n_214),
.C(n_215),
.Y(n_4286)
);

AND2x2_ASAP7_75t_L g4287 ( 
.A(n_4123),
.B(n_215),
.Y(n_4287)
);

AND2x2_ASAP7_75t_L g4288 ( 
.A(n_4166),
.B(n_218),
.Y(n_4288)
);

OR2x2_ASAP7_75t_L g4289 ( 
.A(n_4144),
.B(n_218),
.Y(n_4289)
);

HB1xp67_ASAP7_75t_L g4290 ( 
.A(n_4155),
.Y(n_4290)
);

AND2x2_ASAP7_75t_L g4291 ( 
.A(n_4012),
.B(n_219),
.Y(n_4291)
);

AOI21x1_ASAP7_75t_SL g4292 ( 
.A1(n_4067),
.A2(n_219),
.B(n_220),
.Y(n_4292)
);

NOR2xp67_ASAP7_75t_L g4293 ( 
.A(n_4069),
.B(n_222),
.Y(n_4293)
);

OAI22xp5_ASAP7_75t_L g4294 ( 
.A1(n_4033),
.A2(n_224),
.B1(n_222),
.B2(n_223),
.Y(n_4294)
);

AND2x2_ASAP7_75t_L g4295 ( 
.A(n_4012),
.B(n_223),
.Y(n_4295)
);

NOR2xp67_ASAP7_75t_L g4296 ( 
.A(n_4125),
.B(n_225),
.Y(n_4296)
);

HB1xp67_ASAP7_75t_L g4297 ( 
.A(n_4115),
.Y(n_4297)
);

OA21x2_ASAP7_75t_L g4298 ( 
.A1(n_4138),
.A2(n_226),
.B(n_227),
.Y(n_4298)
);

OR2x2_ASAP7_75t_L g4299 ( 
.A(n_4065),
.B(n_227),
.Y(n_4299)
);

AND2x4_ASAP7_75t_L g4300 ( 
.A(n_4019),
.B(n_228),
.Y(n_4300)
);

OAI22xp5_ASAP7_75t_L g4301 ( 
.A1(n_4171),
.A2(n_231),
.B1(n_228),
.B2(n_230),
.Y(n_4301)
);

AND2x2_ASAP7_75t_L g4302 ( 
.A(n_4021),
.B(n_230),
.Y(n_4302)
);

AND2x2_ASAP7_75t_L g4303 ( 
.A(n_4021),
.B(n_232),
.Y(n_4303)
);

O2A1O1Ixp5_ASAP7_75t_L g4304 ( 
.A1(n_4093),
.A2(n_234),
.B(n_232),
.C(n_233),
.Y(n_4304)
);

AOI21xp5_ASAP7_75t_SL g4305 ( 
.A1(n_4162),
.A2(n_236),
.B(n_238),
.Y(n_4305)
);

BUFx6f_ASAP7_75t_L g4306 ( 
.A(n_4091),
.Y(n_4306)
);

OAI22xp5_ASAP7_75t_L g4307 ( 
.A1(n_4150),
.A2(n_239),
.B1(n_236),
.B2(n_238),
.Y(n_4307)
);

O2A1O1Ixp33_ASAP7_75t_L g4308 ( 
.A1(n_4096),
.A2(n_241),
.B(n_239),
.C(n_240),
.Y(n_4308)
);

AND2x2_ASAP7_75t_L g4309 ( 
.A(n_4244),
.B(n_4103),
.Y(n_4309)
);

OR2x6_ASAP7_75t_L g4310 ( 
.A(n_4306),
.B(n_4098),
.Y(n_4310)
);

NAND2x1p5_ASAP7_75t_L g4311 ( 
.A(n_4306),
.B(n_4019),
.Y(n_4311)
);

NOR3xp33_ASAP7_75t_SL g4312 ( 
.A(n_4276),
.B(n_4134),
.C(n_4110),
.Y(n_4312)
);

INVx2_ASAP7_75t_SL g4313 ( 
.A(n_4306),
.Y(n_4313)
);

INVxp67_ASAP7_75t_L g4314 ( 
.A(n_4297),
.Y(n_4314)
);

BUFx3_ASAP7_75t_L g4315 ( 
.A(n_4177),
.Y(n_4315)
);

INVx2_ASAP7_75t_L g4316 ( 
.A(n_4182),
.Y(n_4316)
);

INVx1_ASAP7_75t_L g4317 ( 
.A(n_4209),
.Y(n_4317)
);

NAND2xp5_ASAP7_75t_L g4318 ( 
.A(n_4173),
.B(n_3999),
.Y(n_4318)
);

NOR2x1_ASAP7_75t_L g4319 ( 
.A(n_4198),
.B(n_4046),
.Y(n_4319)
);

AND2x2_ASAP7_75t_L g4320 ( 
.A(n_4190),
.B(n_4031),
.Y(n_4320)
);

BUFx6f_ASAP7_75t_L g4321 ( 
.A(n_4300),
.Y(n_4321)
);

INVx2_ASAP7_75t_L g4322 ( 
.A(n_4222),
.Y(n_4322)
);

CKINVDCx5p33_ASAP7_75t_R g4323 ( 
.A(n_4213),
.Y(n_4323)
);

INVx1_ASAP7_75t_L g4324 ( 
.A(n_4219),
.Y(n_4324)
);

OR2x6_ASAP7_75t_L g4325 ( 
.A(n_4293),
.B(n_4098),
.Y(n_4325)
);

AND2x2_ASAP7_75t_L g4326 ( 
.A(n_4248),
.B(n_4031),
.Y(n_4326)
);

OR2x2_ASAP7_75t_L g4327 ( 
.A(n_4179),
.B(n_4060),
.Y(n_4327)
);

OR2x2_ASAP7_75t_L g4328 ( 
.A(n_4242),
.B(n_4170),
.Y(n_4328)
);

INVx2_ASAP7_75t_L g4329 ( 
.A(n_4227),
.Y(n_4329)
);

NAND2xp33_ASAP7_75t_R g4330 ( 
.A(n_4197),
.B(n_241),
.Y(n_4330)
);

NOR3xp33_ASAP7_75t_SL g4331 ( 
.A(n_4175),
.B(n_4101),
.C(n_4008),
.Y(n_4331)
);

OR2x6_ASAP7_75t_L g4332 ( 
.A(n_4293),
.B(n_4084),
.Y(n_4332)
);

AND2x2_ASAP7_75t_SL g4333 ( 
.A(n_4216),
.B(n_4019),
.Y(n_4333)
);

NOR2xp33_ASAP7_75t_R g4334 ( 
.A(n_4186),
.B(n_4061),
.Y(n_4334)
);

NOR3xp33_ASAP7_75t_SL g4335 ( 
.A(n_4174),
.B(n_4301),
.C(n_4188),
.Y(n_4335)
);

NAND2xp33_ASAP7_75t_R g4336 ( 
.A(n_4197),
.B(n_242),
.Y(n_4336)
);

INVx3_ASAP7_75t_L g4337 ( 
.A(n_4181),
.Y(n_4337)
);

INVx8_ASAP7_75t_L g4338 ( 
.A(n_4300),
.Y(n_4338)
);

AND2x2_ASAP7_75t_L g4339 ( 
.A(n_4248),
.B(n_4055),
.Y(n_4339)
);

INVx1_ASAP7_75t_L g4340 ( 
.A(n_4273),
.Y(n_4340)
);

AO31x2_ASAP7_75t_L g4341 ( 
.A1(n_4174),
.A2(n_4160),
.A3(n_4128),
.B(n_4127),
.Y(n_4341)
);

CKINVDCx5p33_ASAP7_75t_R g4342 ( 
.A(n_4206),
.Y(n_4342)
);

NAND2x1_ASAP7_75t_L g4343 ( 
.A(n_4238),
.B(n_4181),
.Y(n_4343)
);

NOR2xp33_ASAP7_75t_R g4344 ( 
.A(n_4255),
.B(n_4049),
.Y(n_4344)
);

AND2x4_ASAP7_75t_SL g4345 ( 
.A(n_4198),
.B(n_4131),
.Y(n_4345)
);

NAND4xp25_ASAP7_75t_L g4346 ( 
.A(n_4230),
.B(n_4032),
.C(n_4058),
.D(n_4109),
.Y(n_4346)
);

AO31x2_ASAP7_75t_L g4347 ( 
.A1(n_4191),
.A2(n_4139),
.A3(n_4131),
.B(n_4165),
.Y(n_4347)
);

AOI22xp33_ASAP7_75t_SL g4348 ( 
.A1(n_4245),
.A2(n_4088),
.B1(n_4084),
.B2(n_4147),
.Y(n_4348)
);

AND2x2_ASAP7_75t_L g4349 ( 
.A(n_4252),
.B(n_4055),
.Y(n_4349)
);

INVx1_ASAP7_75t_L g4350 ( 
.A(n_4290),
.Y(n_4350)
);

NOR2xp33_ASAP7_75t_R g4351 ( 
.A(n_4240),
.B(n_4055),
.Y(n_4351)
);

INVx1_ASAP7_75t_L g4352 ( 
.A(n_4231),
.Y(n_4352)
);

NOR3xp33_ASAP7_75t_SL g4353 ( 
.A(n_4280),
.B(n_4195),
.C(n_4274),
.Y(n_4353)
);

INVx2_ASAP7_75t_L g4354 ( 
.A(n_4187),
.Y(n_4354)
);

AND2x2_ASAP7_75t_L g4355 ( 
.A(n_4226),
.B(n_4080),
.Y(n_4355)
);

NOR3xp33_ASAP7_75t_SL g4356 ( 
.A(n_4263),
.B(n_4283),
.C(n_4201),
.Y(n_4356)
);

INVx1_ASAP7_75t_L g4357 ( 
.A(n_4232),
.Y(n_4357)
);

OR2x2_ASAP7_75t_L g4358 ( 
.A(n_4180),
.B(n_4080),
.Y(n_4358)
);

INVx1_ASAP7_75t_L g4359 ( 
.A(n_4233),
.Y(n_4359)
);

OR2x2_ASAP7_75t_L g4360 ( 
.A(n_4176),
.B(n_4080),
.Y(n_4360)
);

AO31x2_ASAP7_75t_L g4361 ( 
.A1(n_4270),
.A2(n_4017),
.A3(n_4016),
.B(n_4042),
.Y(n_4361)
);

OAI22xp5_ASAP7_75t_L g4362 ( 
.A1(n_4277),
.A2(n_4192),
.B1(n_4216),
.B2(n_4267),
.Y(n_4362)
);

NOR2xp33_ASAP7_75t_L g4363 ( 
.A(n_4226),
.B(n_4279),
.Y(n_4363)
);

AOI22xp33_ASAP7_75t_SL g4364 ( 
.A1(n_4245),
.A2(n_4149),
.B1(n_4147),
.B2(n_4120),
.Y(n_4364)
);

INVx4_ASAP7_75t_L g4365 ( 
.A(n_4281),
.Y(n_4365)
);

INVx2_ASAP7_75t_L g4366 ( 
.A(n_4183),
.Y(n_4366)
);

INVx2_ASAP7_75t_L g4367 ( 
.A(n_4237),
.Y(n_4367)
);

AOI22xp33_ASAP7_75t_SL g4368 ( 
.A1(n_4196),
.A2(n_4149),
.B1(n_4147),
.B2(n_4120),
.Y(n_4368)
);

INVx2_ASAP7_75t_L g4369 ( 
.A(n_4250),
.Y(n_4369)
);

INVx2_ASAP7_75t_L g4370 ( 
.A(n_4261),
.Y(n_4370)
);

NOR2xp33_ASAP7_75t_R g4371 ( 
.A(n_4282),
.B(n_4120),
.Y(n_4371)
);

INVx2_ASAP7_75t_L g4372 ( 
.A(n_4285),
.Y(n_4372)
);

HB1xp67_ASAP7_75t_L g4373 ( 
.A(n_4200),
.Y(n_4373)
);

INVx2_ASAP7_75t_L g4374 ( 
.A(n_4204),
.Y(n_4374)
);

HB1xp67_ASAP7_75t_L g4375 ( 
.A(n_4210),
.Y(n_4375)
);

INVx2_ASAP7_75t_L g4376 ( 
.A(n_4178),
.Y(n_4376)
);

OR2x6_ASAP7_75t_L g4377 ( 
.A(n_4305),
.B(n_4149),
.Y(n_4377)
);

INVx1_ASAP7_75t_L g4378 ( 
.A(n_4256),
.Y(n_4378)
);

AOI22xp33_ASAP7_75t_SL g4379 ( 
.A1(n_4196),
.A2(n_4298),
.B1(n_4262),
.B2(n_4288),
.Y(n_4379)
);

BUFx4f_ASAP7_75t_SL g4380 ( 
.A(n_4287),
.Y(n_4380)
);

HB1xp67_ASAP7_75t_L g4381 ( 
.A(n_4236),
.Y(n_4381)
);

NAND2xp33_ASAP7_75t_R g4382 ( 
.A(n_4212),
.B(n_242),
.Y(n_4382)
);

CKINVDCx5p33_ASAP7_75t_R g4383 ( 
.A(n_4269),
.Y(n_4383)
);

AOI22xp33_ASAP7_75t_L g4384 ( 
.A1(n_4199),
.A2(n_4158),
.B1(n_4086),
.B2(n_4017),
.Y(n_4384)
);

INVx4_ASAP7_75t_SL g4385 ( 
.A(n_4291),
.Y(n_4385)
);

BUFx6f_ASAP7_75t_L g4386 ( 
.A(n_4298),
.Y(n_4386)
);

NAND2xp5_ASAP7_75t_L g4387 ( 
.A(n_4278),
.B(n_4289),
.Y(n_4387)
);

AND2x2_ASAP7_75t_L g4388 ( 
.A(n_4229),
.B(n_4162),
.Y(n_4388)
);

CKINVDCx5p33_ASAP7_75t_R g4389 ( 
.A(n_4295),
.Y(n_4389)
);

AND2x2_ASAP7_75t_L g4390 ( 
.A(n_4235),
.B(n_4162),
.Y(n_4390)
);

INVx2_ASAP7_75t_L g4391 ( 
.A(n_4259),
.Y(n_4391)
);

INVx1_ASAP7_75t_L g4392 ( 
.A(n_4251),
.Y(n_4392)
);

CKINVDCx5p33_ASAP7_75t_R g4393 ( 
.A(n_4302),
.Y(n_4393)
);

AO31x2_ASAP7_75t_L g4394 ( 
.A1(n_4218),
.A2(n_4169),
.A3(n_4086),
.B(n_4070),
.Y(n_4394)
);

OAI21x1_ASAP7_75t_L g4395 ( 
.A1(n_4172),
.A2(n_4202),
.B(n_4193),
.Y(n_4395)
);

HB1xp67_ASAP7_75t_L g4396 ( 
.A(n_4268),
.Y(n_4396)
);

AND2x2_ASAP7_75t_L g4397 ( 
.A(n_4214),
.B(n_4130),
.Y(n_4397)
);

CKINVDCx5p33_ASAP7_75t_R g4398 ( 
.A(n_4303),
.Y(n_4398)
);

CKINVDCx5p33_ASAP7_75t_R g4399 ( 
.A(n_4243),
.Y(n_4399)
);

BUFx3_ASAP7_75t_L g4400 ( 
.A(n_4239),
.Y(n_4400)
);

OR2x6_ASAP7_75t_L g4401 ( 
.A(n_4254),
.B(n_4054),
.Y(n_4401)
);

AND2x2_ASAP7_75t_L g4402 ( 
.A(n_4214),
.B(n_243),
.Y(n_4402)
);

NAND2xp5_ASAP7_75t_L g4403 ( 
.A(n_4253),
.B(n_243),
.Y(n_4403)
);

INVx2_ASAP7_75t_L g4404 ( 
.A(n_4228),
.Y(n_4404)
);

CKINVDCx16_ASAP7_75t_R g4405 ( 
.A(n_4241),
.Y(n_4405)
);

NOR2x1_ASAP7_75t_SL g4406 ( 
.A(n_4211),
.B(n_4215),
.Y(n_4406)
);

NAND2xp5_ASAP7_75t_L g4407 ( 
.A(n_4207),
.B(n_244),
.Y(n_4407)
);

OR2x2_ASAP7_75t_L g4408 ( 
.A(n_4299),
.B(n_245),
.Y(n_4408)
);

INVx1_ASAP7_75t_L g4409 ( 
.A(n_4296),
.Y(n_4409)
);

OR2x2_ASAP7_75t_L g4410 ( 
.A(n_4241),
.B(n_245),
.Y(n_4410)
);

OAI21xp5_ASAP7_75t_SL g4411 ( 
.A1(n_4247),
.A2(n_4264),
.B(n_4308),
.Y(n_4411)
);

CKINVDCx5p33_ASAP7_75t_R g4412 ( 
.A(n_4223),
.Y(n_4412)
);

BUFx3_ASAP7_75t_L g4413 ( 
.A(n_4223),
.Y(n_4413)
);

INVx2_ASAP7_75t_L g4414 ( 
.A(n_4184),
.Y(n_4414)
);

INVx1_ASAP7_75t_L g4415 ( 
.A(n_4296),
.Y(n_4415)
);

NOR2xp33_ASAP7_75t_R g4416 ( 
.A(n_4266),
.B(n_246),
.Y(n_4416)
);

NAND2xp5_ASAP7_75t_L g4417 ( 
.A(n_4230),
.B(n_246),
.Y(n_4417)
);

OR2x6_ASAP7_75t_L g4418 ( 
.A(n_4257),
.B(n_4107),
.Y(n_4418)
);

CKINVDCx11_ASAP7_75t_R g4419 ( 
.A(n_4258),
.Y(n_4419)
);

NOR2xp33_ASAP7_75t_R g4420 ( 
.A(n_4292),
.B(n_247),
.Y(n_4420)
);

INVxp67_ASAP7_75t_SL g4421 ( 
.A(n_4205),
.Y(n_4421)
);

OAI21xp5_ASAP7_75t_SL g4422 ( 
.A1(n_4249),
.A2(n_4111),
.B(n_4157),
.Y(n_4422)
);

AO32x1_ASAP7_75t_L g4423 ( 
.A1(n_4217),
.A2(n_4294),
.A3(n_4203),
.B1(n_4307),
.B2(n_4234),
.Y(n_4423)
);

INVx2_ASAP7_75t_L g4424 ( 
.A(n_4184),
.Y(n_4424)
);

HB1xp67_ASAP7_75t_L g4425 ( 
.A(n_4205),
.Y(n_4425)
);

AO31x2_ASAP7_75t_L g4426 ( 
.A1(n_4217),
.A2(n_4092),
.A3(n_250),
.B(n_247),
.Y(n_4426)
);

NAND3xp33_ASAP7_75t_SL g4427 ( 
.A(n_4189),
.B(n_249),
.C(n_250),
.Y(n_4427)
);

AND2x2_ASAP7_75t_L g4428 ( 
.A(n_4208),
.B(n_251),
.Y(n_4428)
);

NOR3xp33_ASAP7_75t_SL g4429 ( 
.A(n_4286),
.B(n_252),
.C(n_253),
.Y(n_4429)
);

NOR2xp33_ASAP7_75t_R g4430 ( 
.A(n_4271),
.B(n_252),
.Y(n_4430)
);

AND2x2_ASAP7_75t_L g4431 ( 
.A(n_4208),
.B(n_254),
.Y(n_4431)
);

BUFx4f_ASAP7_75t_SL g4432 ( 
.A(n_4225),
.Y(n_4432)
);

NAND2xp33_ASAP7_75t_R g4433 ( 
.A(n_4194),
.B(n_254),
.Y(n_4433)
);

AND2x4_ASAP7_75t_L g4434 ( 
.A(n_4265),
.B(n_4246),
.Y(n_4434)
);

INVx1_ASAP7_75t_L g4435 ( 
.A(n_4185),
.Y(n_4435)
);

INVx2_ASAP7_75t_L g4436 ( 
.A(n_4185),
.Y(n_4436)
);

AND2x2_ASAP7_75t_L g4437 ( 
.A(n_4221),
.B(n_255),
.Y(n_4437)
);

BUFx6f_ASAP7_75t_L g4438 ( 
.A(n_4310),
.Y(n_4438)
);

HB1xp67_ASAP7_75t_L g4439 ( 
.A(n_4381),
.Y(n_4439)
);

INVx3_ASAP7_75t_L g4440 ( 
.A(n_4405),
.Y(n_4440)
);

INVx1_ASAP7_75t_L g4441 ( 
.A(n_4352),
.Y(n_4441)
);

AOI33xp33_ASAP7_75t_L g4442 ( 
.A1(n_4379),
.A2(n_4260),
.A3(n_4224),
.B1(n_4220),
.B2(n_4304),
.B3(n_4307),
.Y(n_4442)
);

OR2x2_ASAP7_75t_L g4443 ( 
.A(n_4329),
.B(n_4294),
.Y(n_4443)
);

INVxp33_ASAP7_75t_L g4444 ( 
.A(n_4334),
.Y(n_4444)
);

OR2x2_ASAP7_75t_L g4445 ( 
.A(n_4391),
.B(n_4396),
.Y(n_4445)
);

AND2x2_ASAP7_75t_L g4446 ( 
.A(n_4333),
.B(n_4275),
.Y(n_4446)
);

NAND2xp5_ASAP7_75t_L g4447 ( 
.A(n_4437),
.B(n_4272),
.Y(n_4447)
);

INVx2_ASAP7_75t_L g4448 ( 
.A(n_4386),
.Y(n_4448)
);

AOI221xp5_ASAP7_75t_L g4449 ( 
.A1(n_4335),
.A2(n_4284),
.B1(n_258),
.B2(n_261),
.C(n_262),
.Y(n_4449)
);

INVx2_ASAP7_75t_L g4450 ( 
.A(n_4386),
.Y(n_4450)
);

AO21x2_ASAP7_75t_L g4451 ( 
.A1(n_4417),
.A2(n_256),
.B(n_258),
.Y(n_4451)
);

NAND2xp5_ASAP7_75t_L g4452 ( 
.A(n_4392),
.B(n_262),
.Y(n_4452)
);

AO21x2_ASAP7_75t_L g4453 ( 
.A1(n_4435),
.A2(n_4436),
.B(n_4318),
.Y(n_4453)
);

INVx1_ASAP7_75t_L g4454 ( 
.A(n_4352),
.Y(n_4454)
);

BUFx2_ASAP7_75t_L g4455 ( 
.A(n_4344),
.Y(n_4455)
);

INVx4_ASAP7_75t_L g4456 ( 
.A(n_4310),
.Y(n_4456)
);

INVx1_ASAP7_75t_L g4457 ( 
.A(n_4357),
.Y(n_4457)
);

INVx1_ASAP7_75t_L g4458 ( 
.A(n_4359),
.Y(n_4458)
);

AND2x2_ASAP7_75t_L g4459 ( 
.A(n_4337),
.B(n_263),
.Y(n_4459)
);

INVx3_ASAP7_75t_L g4460 ( 
.A(n_4343),
.Y(n_4460)
);

AND2x2_ASAP7_75t_L g4461 ( 
.A(n_4337),
.B(n_263),
.Y(n_4461)
);

INVx1_ASAP7_75t_L g4462 ( 
.A(n_4378),
.Y(n_4462)
);

INVx1_ASAP7_75t_L g4463 ( 
.A(n_4317),
.Y(n_4463)
);

OA21x2_ASAP7_75t_L g4464 ( 
.A1(n_4395),
.A2(n_265),
.B(n_266),
.Y(n_4464)
);

AO21x2_ASAP7_75t_L g4465 ( 
.A1(n_4427),
.A2(n_266),
.B(n_267),
.Y(n_4465)
);

NAND2xp5_ASAP7_75t_L g4466 ( 
.A(n_4350),
.B(n_268),
.Y(n_4466)
);

INVx1_ASAP7_75t_L g4467 ( 
.A(n_4324),
.Y(n_4467)
);

AND2x2_ASAP7_75t_L g4468 ( 
.A(n_4373),
.B(n_268),
.Y(n_4468)
);

NAND2xp5_ASAP7_75t_L g4469 ( 
.A(n_4324),
.B(n_269),
.Y(n_4469)
);

AND2x2_ASAP7_75t_L g4470 ( 
.A(n_4375),
.B(n_270),
.Y(n_4470)
);

BUFx6f_ASAP7_75t_L g4471 ( 
.A(n_4315),
.Y(n_4471)
);

INVxp67_ASAP7_75t_SL g4472 ( 
.A(n_4330),
.Y(n_4472)
);

INVx2_ASAP7_75t_L g4473 ( 
.A(n_4386),
.Y(n_4473)
);

INVx2_ASAP7_75t_L g4474 ( 
.A(n_4341),
.Y(n_4474)
);

INVx1_ASAP7_75t_L g4475 ( 
.A(n_4340),
.Y(n_4475)
);

INVxp33_ASAP7_75t_L g4476 ( 
.A(n_4351),
.Y(n_4476)
);

INVx1_ASAP7_75t_L g4477 ( 
.A(n_4340),
.Y(n_4477)
);

NAND2xp5_ASAP7_75t_L g4478 ( 
.A(n_4314),
.B(n_4353),
.Y(n_4478)
);

OR2x6_ASAP7_75t_L g4479 ( 
.A(n_4325),
.B(n_4332),
.Y(n_4479)
);

INVx2_ASAP7_75t_L g4480 ( 
.A(n_4341),
.Y(n_4480)
);

INVxp67_ASAP7_75t_SL g4481 ( 
.A(n_4336),
.Y(n_4481)
);

AND2x2_ASAP7_75t_L g4482 ( 
.A(n_4326),
.B(n_271),
.Y(n_4482)
);

INVx1_ASAP7_75t_L g4483 ( 
.A(n_4327),
.Y(n_4483)
);

OR2x2_ASAP7_75t_L g4484 ( 
.A(n_4354),
.B(n_272),
.Y(n_4484)
);

OAI21xp5_ASAP7_75t_L g4485 ( 
.A1(n_4331),
.A2(n_272),
.B(n_273),
.Y(n_4485)
);

AND2x2_ASAP7_75t_L g4486 ( 
.A(n_4339),
.B(n_273),
.Y(n_4486)
);

AND2x2_ASAP7_75t_L g4487 ( 
.A(n_4320),
.B(n_275),
.Y(n_4487)
);

AND2x2_ASAP7_75t_L g4488 ( 
.A(n_4347),
.B(n_276),
.Y(n_4488)
);

OAI221xp5_ASAP7_75t_L g4489 ( 
.A1(n_4433),
.A2(n_276),
.B1(n_277),
.B2(n_278),
.C(n_279),
.Y(n_4489)
);

INVx1_ASAP7_75t_L g4490 ( 
.A(n_4415),
.Y(n_4490)
);

INVx2_ASAP7_75t_SL g4491 ( 
.A(n_4319),
.Y(n_4491)
);

INVx1_ASAP7_75t_L g4492 ( 
.A(n_4366),
.Y(n_4492)
);

INVx2_ASAP7_75t_L g4493 ( 
.A(n_4341),
.Y(n_4493)
);

INVxp67_ASAP7_75t_SL g4494 ( 
.A(n_4382),
.Y(n_4494)
);

INVx1_ASAP7_75t_L g4495 ( 
.A(n_4409),
.Y(n_4495)
);

BUFx2_ASAP7_75t_L g4496 ( 
.A(n_4371),
.Y(n_4496)
);

INVx1_ASAP7_75t_L g4497 ( 
.A(n_4409),
.Y(n_4497)
);

AO21x2_ASAP7_75t_L g4498 ( 
.A1(n_4414),
.A2(n_277),
.B(n_279),
.Y(n_4498)
);

INVx1_ASAP7_75t_L g4499 ( 
.A(n_4387),
.Y(n_4499)
);

AO21x2_ASAP7_75t_L g4500 ( 
.A1(n_4424),
.A2(n_281),
.B(n_282),
.Y(n_4500)
);

INVx1_ASAP7_75t_L g4501 ( 
.A(n_4400),
.Y(n_4501)
);

INVx3_ASAP7_75t_L g4502 ( 
.A(n_4365),
.Y(n_4502)
);

AND2x2_ASAP7_75t_L g4503 ( 
.A(n_4347),
.B(n_283),
.Y(n_4503)
);

INVx2_ASAP7_75t_L g4504 ( 
.A(n_4316),
.Y(n_4504)
);

AOI21xp5_ASAP7_75t_SL g4505 ( 
.A1(n_4325),
.A2(n_284),
.B(n_285),
.Y(n_4505)
);

INVx1_ASAP7_75t_L g4506 ( 
.A(n_4328),
.Y(n_4506)
);

INVx1_ASAP7_75t_L g4507 ( 
.A(n_4404),
.Y(n_4507)
);

AND2x2_ASAP7_75t_L g4508 ( 
.A(n_4347),
.B(n_4388),
.Y(n_4508)
);

INVx1_ASAP7_75t_L g4509 ( 
.A(n_4408),
.Y(n_4509)
);

AO21x2_ASAP7_75t_L g4510 ( 
.A1(n_4407),
.A2(n_4431),
.B(n_4428),
.Y(n_4510)
);

A2O1A1Ixp33_ASAP7_75t_L g4511 ( 
.A1(n_4411),
.A2(n_4429),
.B(n_4356),
.C(n_4362),
.Y(n_4511)
);

CKINVDCx5p33_ASAP7_75t_R g4512 ( 
.A(n_4323),
.Y(n_4512)
);

OR2x2_ASAP7_75t_L g4513 ( 
.A(n_4376),
.B(n_4374),
.Y(n_4513)
);

BUFx2_ASAP7_75t_L g4514 ( 
.A(n_4365),
.Y(n_4514)
);

HB1xp67_ASAP7_75t_L g4515 ( 
.A(n_4360),
.Y(n_4515)
);

OAI21xp5_ASAP7_75t_L g4516 ( 
.A1(n_4364),
.A2(n_284),
.B(n_286),
.Y(n_4516)
);

AND2x2_ASAP7_75t_L g4517 ( 
.A(n_4390),
.B(n_4406),
.Y(n_4517)
);

NAND3xp33_ASAP7_75t_L g4518 ( 
.A(n_4368),
.B(n_286),
.C(n_288),
.Y(n_4518)
);

HB1xp67_ASAP7_75t_L g4519 ( 
.A(n_4358),
.Y(n_4519)
);

INVx2_ASAP7_75t_L g4520 ( 
.A(n_4322),
.Y(n_4520)
);

AO21x2_ASAP7_75t_L g4521 ( 
.A1(n_4403),
.A2(n_288),
.B(n_289),
.Y(n_4521)
);

HB1xp67_ASAP7_75t_L g4522 ( 
.A(n_4402),
.Y(n_4522)
);

INVx1_ASAP7_75t_L g4523 ( 
.A(n_4321),
.Y(n_4523)
);

OA21x2_ASAP7_75t_L g4524 ( 
.A1(n_4421),
.A2(n_290),
.B(n_291),
.Y(n_4524)
);

INVx1_ASAP7_75t_SL g4525 ( 
.A(n_4380),
.Y(n_4525)
);

OR2x2_ASAP7_75t_L g4526 ( 
.A(n_4413),
.B(n_4394),
.Y(n_4526)
);

INVx1_ASAP7_75t_L g4527 ( 
.A(n_4321),
.Y(n_4527)
);

AND2x2_ASAP7_75t_L g4528 ( 
.A(n_4406),
.B(n_291),
.Y(n_4528)
);

INVx1_ASAP7_75t_L g4529 ( 
.A(n_4321),
.Y(n_4529)
);

INVx1_ASAP7_75t_L g4530 ( 
.A(n_4410),
.Y(n_4530)
);

INVx1_ASAP7_75t_L g4531 ( 
.A(n_4363),
.Y(n_4531)
);

OA21x2_ASAP7_75t_L g4532 ( 
.A1(n_4425),
.A2(n_292),
.B(n_293),
.Y(n_4532)
);

INVx2_ASAP7_75t_L g4533 ( 
.A(n_4367),
.Y(n_4533)
);

INVx3_ASAP7_75t_L g4534 ( 
.A(n_4311),
.Y(n_4534)
);

BUFx2_ASAP7_75t_L g4535 ( 
.A(n_4309),
.Y(n_4535)
);

INVx3_ASAP7_75t_L g4536 ( 
.A(n_4332),
.Y(n_4536)
);

OAI21xp5_ASAP7_75t_L g4537 ( 
.A1(n_4348),
.A2(n_292),
.B(n_294),
.Y(n_4537)
);

AND2x2_ASAP7_75t_L g4538 ( 
.A(n_4349),
.B(n_294),
.Y(n_4538)
);

BUFx2_ASAP7_75t_L g4539 ( 
.A(n_4342),
.Y(n_4539)
);

AO21x2_ASAP7_75t_L g4540 ( 
.A1(n_4420),
.A2(n_296),
.B(n_297),
.Y(n_4540)
);

INVx1_ASAP7_75t_L g4541 ( 
.A(n_4441),
.Y(n_4541)
);

INVx4_ASAP7_75t_SL g4542 ( 
.A(n_4438),
.Y(n_4542)
);

INVx1_ASAP7_75t_L g4543 ( 
.A(n_4454),
.Y(n_4543)
);

INVx1_ASAP7_75t_L g4544 ( 
.A(n_4457),
.Y(n_4544)
);

AND2x4_ASAP7_75t_L g4545 ( 
.A(n_4440),
.B(n_4385),
.Y(n_4545)
);

NAND2xp5_ASAP7_75t_L g4546 ( 
.A(n_4451),
.B(n_4385),
.Y(n_4546)
);

HB1xp67_ASAP7_75t_L g4547 ( 
.A(n_4451),
.Y(n_4547)
);

BUFx2_ASAP7_75t_L g4548 ( 
.A(n_4455),
.Y(n_4548)
);

AND2x2_ASAP7_75t_L g4549 ( 
.A(n_4517),
.B(n_4345),
.Y(n_4549)
);

NAND2xp5_ASAP7_75t_L g4550 ( 
.A(n_4451),
.B(n_4338),
.Y(n_4550)
);

INVx1_ASAP7_75t_L g4551 ( 
.A(n_4458),
.Y(n_4551)
);

NAND2xp5_ASAP7_75t_L g4552 ( 
.A(n_4470),
.B(n_4338),
.Y(n_4552)
);

NAND2xp5_ASAP7_75t_L g4553 ( 
.A(n_4470),
.B(n_4432),
.Y(n_4553)
);

INVx2_ASAP7_75t_L g4554 ( 
.A(n_4532),
.Y(n_4554)
);

INVx1_ASAP7_75t_L g4555 ( 
.A(n_4462),
.Y(n_4555)
);

AND2x2_ASAP7_75t_L g4556 ( 
.A(n_4517),
.B(n_4355),
.Y(n_4556)
);

NAND2xp5_ASAP7_75t_L g4557 ( 
.A(n_4439),
.B(n_4399),
.Y(n_4557)
);

NAND2xp5_ASAP7_75t_L g4558 ( 
.A(n_4521),
.B(n_4312),
.Y(n_4558)
);

OAI22x1_ASAP7_75t_L g4559 ( 
.A1(n_4472),
.A2(n_4423),
.B1(n_4383),
.B2(n_4389),
.Y(n_4559)
);

OAI221xp5_ASAP7_75t_SL g4560 ( 
.A1(n_4511),
.A2(n_4423),
.B1(n_4401),
.B2(n_4418),
.C(n_4346),
.Y(n_4560)
);

AND2x2_ASAP7_75t_L g4561 ( 
.A(n_4440),
.B(n_4313),
.Y(n_4561)
);

INVx1_ASAP7_75t_L g4562 ( 
.A(n_4467),
.Y(n_4562)
);

INVx1_ASAP7_75t_L g4563 ( 
.A(n_4475),
.Y(n_4563)
);

AND2x2_ASAP7_75t_L g4564 ( 
.A(n_4440),
.B(n_4412),
.Y(n_4564)
);

CKINVDCx11_ASAP7_75t_R g4565 ( 
.A(n_4471),
.Y(n_4565)
);

OR2x2_ASAP7_75t_L g4566 ( 
.A(n_4499),
.B(n_4463),
.Y(n_4566)
);

AND2x2_ASAP7_75t_L g4567 ( 
.A(n_4535),
.B(n_4496),
.Y(n_4567)
);

INVx2_ASAP7_75t_SL g4568 ( 
.A(n_4471),
.Y(n_4568)
);

AND2x2_ASAP7_75t_L g4569 ( 
.A(n_4491),
.B(n_4502),
.Y(n_4569)
);

AND2x2_ASAP7_75t_L g4570 ( 
.A(n_4491),
.B(n_4397),
.Y(n_4570)
);

INVx2_ASAP7_75t_L g4571 ( 
.A(n_4532),
.Y(n_4571)
);

INVx1_ASAP7_75t_L g4572 ( 
.A(n_4477),
.Y(n_4572)
);

NOR2xp33_ASAP7_75t_L g4573 ( 
.A(n_4444),
.B(n_4476),
.Y(n_4573)
);

BUFx2_ASAP7_75t_L g4574 ( 
.A(n_4456),
.Y(n_4574)
);

HB1xp67_ASAP7_75t_L g4575 ( 
.A(n_4524),
.Y(n_4575)
);

INVx2_ASAP7_75t_L g4576 ( 
.A(n_4532),
.Y(n_4576)
);

NAND2xp5_ASAP7_75t_L g4577 ( 
.A(n_4521),
.B(n_4426),
.Y(n_4577)
);

INVx1_ASAP7_75t_L g4578 ( 
.A(n_4492),
.Y(n_4578)
);

INVx2_ASAP7_75t_L g4579 ( 
.A(n_4524),
.Y(n_4579)
);

NAND2xp5_ASAP7_75t_L g4580 ( 
.A(n_4521),
.B(n_4426),
.Y(n_4580)
);

OR2x2_ASAP7_75t_L g4581 ( 
.A(n_4443),
.B(n_4394),
.Y(n_4581)
);

NAND2xp5_ASAP7_75t_L g4582 ( 
.A(n_4468),
.B(n_4426),
.Y(n_4582)
);

INVxp67_ASAP7_75t_SL g4583 ( 
.A(n_4471),
.Y(n_4583)
);

INVx1_ASAP7_75t_L g4584 ( 
.A(n_4509),
.Y(n_4584)
);

INVx2_ASAP7_75t_L g4585 ( 
.A(n_4524),
.Y(n_4585)
);

AND2x2_ASAP7_75t_L g4586 ( 
.A(n_4502),
.B(n_4393),
.Y(n_4586)
);

INVx2_ASAP7_75t_L g4587 ( 
.A(n_4540),
.Y(n_4587)
);

INVx1_ASAP7_75t_L g4588 ( 
.A(n_4445),
.Y(n_4588)
);

BUFx2_ASAP7_75t_L g4589 ( 
.A(n_4456),
.Y(n_4589)
);

INVx1_ASAP7_75t_L g4590 ( 
.A(n_4483),
.Y(n_4590)
);

INVx1_ASAP7_75t_L g4591 ( 
.A(n_4468),
.Y(n_4591)
);

INVx1_ASAP7_75t_L g4592 ( 
.A(n_4484),
.Y(n_4592)
);

OR2x2_ASAP7_75t_L g4593 ( 
.A(n_4513),
.B(n_4394),
.Y(n_4593)
);

HB1xp67_ASAP7_75t_L g4594 ( 
.A(n_4522),
.Y(n_4594)
);

INVx1_ASAP7_75t_L g4595 ( 
.A(n_4498),
.Y(n_4595)
);

AOI222xp33_ASAP7_75t_L g4596 ( 
.A1(n_4481),
.A2(n_4419),
.B1(n_4422),
.B2(n_4384),
.C1(n_4369),
.C2(n_4370),
.Y(n_4596)
);

INVx1_ASAP7_75t_L g4597 ( 
.A(n_4498),
.Y(n_4597)
);

INVx2_ASAP7_75t_L g4598 ( 
.A(n_4540),
.Y(n_4598)
);

OR2x2_ASAP7_75t_L g4599 ( 
.A(n_4506),
.B(n_4361),
.Y(n_4599)
);

INVx1_ASAP7_75t_L g4600 ( 
.A(n_4498),
.Y(n_4600)
);

INVx1_ASAP7_75t_L g4601 ( 
.A(n_4500),
.Y(n_4601)
);

BUFx2_ASAP7_75t_L g4602 ( 
.A(n_4456),
.Y(n_4602)
);

AND2x2_ASAP7_75t_L g4603 ( 
.A(n_4502),
.B(n_4398),
.Y(n_4603)
);

AND2x2_ASAP7_75t_L g4604 ( 
.A(n_4514),
.B(n_4434),
.Y(n_4604)
);

OR2x2_ASAP7_75t_L g4605 ( 
.A(n_4495),
.B(n_4361),
.Y(n_4605)
);

CKINVDCx11_ASAP7_75t_R g4606 ( 
.A(n_4471),
.Y(n_4606)
);

INVx2_ASAP7_75t_L g4607 ( 
.A(n_4540),
.Y(n_4607)
);

INVx2_ASAP7_75t_L g4608 ( 
.A(n_4500),
.Y(n_4608)
);

AND2x2_ASAP7_75t_L g4609 ( 
.A(n_4508),
.B(n_4434),
.Y(n_4609)
);

INVxp67_ASAP7_75t_L g4610 ( 
.A(n_4573),
.Y(n_4610)
);

AND2x2_ASAP7_75t_L g4611 ( 
.A(n_4567),
.B(n_4508),
.Y(n_4611)
);

OR2x6_ASAP7_75t_L g4612 ( 
.A(n_4587),
.B(n_4505),
.Y(n_4612)
);

OAI22xp5_ASAP7_75t_L g4613 ( 
.A1(n_4560),
.A2(n_4511),
.B1(n_4478),
.B2(n_4518),
.Y(n_4613)
);

HB1xp67_ASAP7_75t_L g4614 ( 
.A(n_4548),
.Y(n_4614)
);

INVxp67_ASAP7_75t_L g4615 ( 
.A(n_4573),
.Y(n_4615)
);

AND2x2_ASAP7_75t_L g4616 ( 
.A(n_4567),
.B(n_4519),
.Y(n_4616)
);

NOR2xp33_ASAP7_75t_L g4617 ( 
.A(n_4565),
.B(n_4444),
.Y(n_4617)
);

AND2x2_ASAP7_75t_SL g4618 ( 
.A(n_4575),
.B(n_4528),
.Y(n_4618)
);

INVx2_ASAP7_75t_L g4619 ( 
.A(n_4554),
.Y(n_4619)
);

AND2x4_ASAP7_75t_L g4620 ( 
.A(n_4545),
.B(n_4438),
.Y(n_4620)
);

AOI222xp33_ASAP7_75t_L g4621 ( 
.A1(n_4559),
.A2(n_4494),
.B1(n_4489),
.B2(n_4485),
.C1(n_4503),
.C2(n_4488),
.Y(n_4621)
);

NAND3xp33_ASAP7_75t_L g4622 ( 
.A(n_4579),
.B(n_4449),
.C(n_4585),
.Y(n_4622)
);

BUFx2_ASAP7_75t_SL g4623 ( 
.A(n_4568),
.Y(n_4623)
);

AOI21xp5_ASAP7_75t_L g4624 ( 
.A1(n_4559),
.A2(n_4447),
.B(n_4528),
.Y(n_4624)
);

INVxp67_ASAP7_75t_L g4625 ( 
.A(n_4564),
.Y(n_4625)
);

HB1xp67_ASAP7_75t_L g4626 ( 
.A(n_4591),
.Y(n_4626)
);

AOI22xp33_ASAP7_75t_L g4627 ( 
.A1(n_4554),
.A2(n_4453),
.B1(n_4503),
.B2(n_4488),
.Y(n_4627)
);

AND2x2_ASAP7_75t_L g4628 ( 
.A(n_4545),
.B(n_4515),
.Y(n_4628)
);

BUFx2_ASAP7_75t_L g4629 ( 
.A(n_4545),
.Y(n_4629)
);

NAND2xp5_ASAP7_75t_L g4630 ( 
.A(n_4579),
.B(n_4510),
.Y(n_4630)
);

OR2x2_ASAP7_75t_L g4631 ( 
.A(n_4594),
.B(n_4490),
.Y(n_4631)
);

INVx2_ASAP7_75t_L g4632 ( 
.A(n_4571),
.Y(n_4632)
);

INVx2_ASAP7_75t_L g4633 ( 
.A(n_4571),
.Y(n_4633)
);

INVx1_ASAP7_75t_L g4634 ( 
.A(n_4566),
.Y(n_4634)
);

INVx2_ASAP7_75t_SL g4635 ( 
.A(n_4564),
.Y(n_4635)
);

AOI221xp5_ASAP7_75t_L g4636 ( 
.A1(n_4547),
.A2(n_4453),
.B1(n_4473),
.B2(n_4450),
.C(n_4448),
.Y(n_4636)
);

INVx2_ASAP7_75t_L g4637 ( 
.A(n_4576),
.Y(n_4637)
);

OAI222xp33_ASAP7_75t_L g4638 ( 
.A1(n_4581),
.A2(n_4526),
.B1(n_4479),
.B2(n_4450),
.C1(n_4473),
.C2(n_4448),
.Y(n_4638)
);

OAI33xp33_ASAP7_75t_L g4639 ( 
.A1(n_4588),
.A2(n_4581),
.A3(n_4590),
.B1(n_4584),
.B2(n_4599),
.B3(n_4566),
.Y(n_4639)
);

OR2x2_ASAP7_75t_L g4640 ( 
.A(n_4582),
.B(n_4497),
.Y(n_4640)
);

INVxp67_ASAP7_75t_SL g4641 ( 
.A(n_4553),
.Y(n_4641)
);

AOI21x1_ASAP7_75t_L g4642 ( 
.A1(n_4574),
.A2(n_4479),
.B(n_4461),
.Y(n_4642)
);

INVx2_ASAP7_75t_L g4643 ( 
.A(n_4576),
.Y(n_4643)
);

INVx2_ASAP7_75t_SL g4644 ( 
.A(n_4561),
.Y(n_4644)
);

AOI22xp33_ASAP7_75t_L g4645 ( 
.A1(n_4587),
.A2(n_4464),
.B1(n_4516),
.B2(n_4465),
.Y(n_4645)
);

INVxp67_ASAP7_75t_L g4646 ( 
.A(n_4561),
.Y(n_4646)
);

AO21x2_ASAP7_75t_L g4647 ( 
.A1(n_4598),
.A2(n_4469),
.B(n_4466),
.Y(n_4647)
);

AND2x2_ASAP7_75t_L g4648 ( 
.A(n_4556),
.B(n_4464),
.Y(n_4648)
);

NOR2xp33_ASAP7_75t_R g4649 ( 
.A(n_4565),
.B(n_4512),
.Y(n_4649)
);

CKINVDCx5p33_ASAP7_75t_R g4650 ( 
.A(n_4606),
.Y(n_4650)
);

OAI21x1_ASAP7_75t_L g4651 ( 
.A1(n_4585),
.A2(n_4536),
.B(n_4598),
.Y(n_4651)
);

AND2x2_ASAP7_75t_L g4652 ( 
.A(n_4556),
.B(n_4464),
.Y(n_4652)
);

INVx1_ASAP7_75t_L g4653 ( 
.A(n_4619),
.Y(n_4653)
);

AND2x4_ASAP7_75t_L g4654 ( 
.A(n_4620),
.B(n_4586),
.Y(n_4654)
);

INVx2_ASAP7_75t_L g4655 ( 
.A(n_4612),
.Y(n_4655)
);

INVx1_ASAP7_75t_L g4656 ( 
.A(n_4619),
.Y(n_4656)
);

NAND2x1p5_ASAP7_75t_L g4657 ( 
.A(n_4620),
.B(n_4438),
.Y(n_4657)
);

OR2x2_ASAP7_75t_L g4658 ( 
.A(n_4614),
.B(n_4583),
.Y(n_4658)
);

AND2x2_ASAP7_75t_L g4659 ( 
.A(n_4616),
.B(n_4606),
.Y(n_4659)
);

OR2x2_ASAP7_75t_L g4660 ( 
.A(n_4610),
.B(n_4615),
.Y(n_4660)
);

OR2x2_ASAP7_75t_L g4661 ( 
.A(n_4616),
.B(n_4568),
.Y(n_4661)
);

NAND2xp5_ASAP7_75t_L g4662 ( 
.A(n_4627),
.B(n_4541),
.Y(n_4662)
);

INVx2_ASAP7_75t_L g4663 ( 
.A(n_4612),
.Y(n_4663)
);

OR2x2_ASAP7_75t_L g4664 ( 
.A(n_4626),
.B(n_4644),
.Y(n_4664)
);

AND2x4_ASAP7_75t_L g4665 ( 
.A(n_4620),
.B(n_4542),
.Y(n_4665)
);

INVx4_ASAP7_75t_L g4666 ( 
.A(n_4650),
.Y(n_4666)
);

AND2x2_ASAP7_75t_L g4667 ( 
.A(n_4611),
.B(n_4586),
.Y(n_4667)
);

OR2x2_ASAP7_75t_L g4668 ( 
.A(n_4644),
.B(n_4589),
.Y(n_4668)
);

OR2x2_ASAP7_75t_L g4669 ( 
.A(n_4634),
.B(n_4602),
.Y(n_4669)
);

NAND2xp5_ASAP7_75t_L g4670 ( 
.A(n_4632),
.B(n_4543),
.Y(n_4670)
);

BUFx2_ASAP7_75t_L g4671 ( 
.A(n_4649),
.Y(n_4671)
);

INVx1_ASAP7_75t_L g4672 ( 
.A(n_4632),
.Y(n_4672)
);

AND2x2_ASAP7_75t_L g4673 ( 
.A(n_4611),
.B(n_4603),
.Y(n_4673)
);

INVx1_ASAP7_75t_L g4674 ( 
.A(n_4633),
.Y(n_4674)
);

INVxp67_ASAP7_75t_L g4675 ( 
.A(n_4623),
.Y(n_4675)
);

AND2x2_ASAP7_75t_L g4676 ( 
.A(n_4650),
.B(n_4603),
.Y(n_4676)
);

NAND2xp5_ASAP7_75t_L g4677 ( 
.A(n_4633),
.B(n_4544),
.Y(n_4677)
);

AND2x2_ASAP7_75t_L g4678 ( 
.A(n_4618),
.B(n_4549),
.Y(n_4678)
);

INVxp67_ASAP7_75t_SL g4679 ( 
.A(n_4613),
.Y(n_4679)
);

NAND2xp5_ASAP7_75t_L g4680 ( 
.A(n_4637),
.B(n_4551),
.Y(n_4680)
);

OR2x2_ASAP7_75t_L g4681 ( 
.A(n_4660),
.B(n_4635),
.Y(n_4681)
);

AND2x4_ASAP7_75t_L g4682 ( 
.A(n_4665),
.B(n_4635),
.Y(n_4682)
);

INVx1_ASAP7_75t_L g4683 ( 
.A(n_4658),
.Y(n_4683)
);

OR2x2_ASAP7_75t_L g4684 ( 
.A(n_4664),
.B(n_4631),
.Y(n_4684)
);

AND2x4_ASAP7_75t_L g4685 ( 
.A(n_4665),
.B(n_4629),
.Y(n_4685)
);

OR2x2_ASAP7_75t_L g4686 ( 
.A(n_4661),
.B(n_4640),
.Y(n_4686)
);

NAND2xp5_ASAP7_75t_L g4687 ( 
.A(n_4679),
.B(n_4618),
.Y(n_4687)
);

NAND2xp5_ASAP7_75t_L g4688 ( 
.A(n_4679),
.B(n_4622),
.Y(n_4688)
);

HB1xp67_ASAP7_75t_L g4689 ( 
.A(n_4662),
.Y(n_4689)
);

INVx1_ASAP7_75t_L g4690 ( 
.A(n_4653),
.Y(n_4690)
);

AND2x2_ASAP7_75t_L g4691 ( 
.A(n_4659),
.B(n_4649),
.Y(n_4691)
);

BUFx2_ASAP7_75t_L g4692 ( 
.A(n_4665),
.Y(n_4692)
);

INVx1_ASAP7_75t_L g4693 ( 
.A(n_4656),
.Y(n_4693)
);

NOR2xp33_ASAP7_75t_L g4694 ( 
.A(n_4666),
.B(n_4639),
.Y(n_4694)
);

INVx3_ASAP7_75t_L g4695 ( 
.A(n_4666),
.Y(n_4695)
);

AND2x2_ASAP7_75t_L g4696 ( 
.A(n_4671),
.B(n_4628),
.Y(n_4696)
);

AND2x4_ASAP7_75t_L g4697 ( 
.A(n_4654),
.B(n_4625),
.Y(n_4697)
);

INVx1_ASAP7_75t_L g4698 ( 
.A(n_4672),
.Y(n_4698)
);

INVx1_ASAP7_75t_L g4699 ( 
.A(n_4674),
.Y(n_4699)
);

AND2x2_ASAP7_75t_L g4700 ( 
.A(n_4676),
.B(n_4628),
.Y(n_4700)
);

NAND2xp5_ASAP7_75t_SL g4701 ( 
.A(n_4688),
.B(n_4687),
.Y(n_4701)
);

OAI21xp33_ASAP7_75t_L g4702 ( 
.A1(n_4694),
.A2(n_4678),
.B(n_4641),
.Y(n_4702)
);

AND2x2_ASAP7_75t_L g4703 ( 
.A(n_4696),
.B(n_4654),
.Y(n_4703)
);

INVx1_ASAP7_75t_L g4704 ( 
.A(n_4684),
.Y(n_4704)
);

INVx2_ASAP7_75t_L g4705 ( 
.A(n_4692),
.Y(n_4705)
);

AND2x2_ASAP7_75t_SL g4706 ( 
.A(n_4688),
.B(n_4617),
.Y(n_4706)
);

AND2x2_ASAP7_75t_L g4707 ( 
.A(n_4685),
.B(n_4667),
.Y(n_4707)
);

INVx1_ASAP7_75t_L g4708 ( 
.A(n_4683),
.Y(n_4708)
);

INVx1_ASAP7_75t_L g4709 ( 
.A(n_4681),
.Y(n_4709)
);

OR2x2_ASAP7_75t_L g4710 ( 
.A(n_4687),
.B(n_4686),
.Y(n_4710)
);

INVx1_ASAP7_75t_L g4711 ( 
.A(n_4689),
.Y(n_4711)
);

INVx1_ASAP7_75t_L g4712 ( 
.A(n_4689),
.Y(n_4712)
);

OR2x2_ASAP7_75t_L g4713 ( 
.A(n_4697),
.B(n_4669),
.Y(n_4713)
);

AND2x2_ASAP7_75t_L g4714 ( 
.A(n_4700),
.B(n_4673),
.Y(n_4714)
);

INVx2_ASAP7_75t_L g4715 ( 
.A(n_4685),
.Y(n_4715)
);

AND2x2_ASAP7_75t_L g4716 ( 
.A(n_4685),
.B(n_4675),
.Y(n_4716)
);

OR2x2_ASAP7_75t_L g4717 ( 
.A(n_4697),
.B(n_4668),
.Y(n_4717)
);

INVx2_ASAP7_75t_L g4718 ( 
.A(n_4682),
.Y(n_4718)
);

INVx1_ASAP7_75t_L g4719 ( 
.A(n_4690),
.Y(n_4719)
);

INVx1_ASAP7_75t_L g4720 ( 
.A(n_4705),
.Y(n_4720)
);

NAND2x1p5_ASAP7_75t_L g4721 ( 
.A(n_4716),
.B(n_4695),
.Y(n_4721)
);

O2A1O1Ixp33_ASAP7_75t_L g4722 ( 
.A1(n_4701),
.A2(n_4694),
.B(n_4662),
.C(n_4624),
.Y(n_4722)
);

BUFx2_ASAP7_75t_L g4723 ( 
.A(n_4703),
.Y(n_4723)
);

NAND2x1_ASAP7_75t_L g4724 ( 
.A(n_4707),
.B(n_4682),
.Y(n_4724)
);

INVx1_ASAP7_75t_L g4725 ( 
.A(n_4705),
.Y(n_4725)
);

INVx1_ASAP7_75t_L g4726 ( 
.A(n_4711),
.Y(n_4726)
);

AOI32xp33_ASAP7_75t_L g4727 ( 
.A1(n_4701),
.A2(n_4636),
.A3(n_4648),
.B1(n_4652),
.B2(n_4645),
.Y(n_4727)
);

OAI21xp33_ASAP7_75t_L g4728 ( 
.A1(n_4703),
.A2(n_4691),
.B(n_4646),
.Y(n_4728)
);

OR2x2_ASAP7_75t_L g4729 ( 
.A(n_4710),
.B(n_4695),
.Y(n_4729)
);

NAND2xp5_ASAP7_75t_L g4730 ( 
.A(n_4714),
.B(n_4675),
.Y(n_4730)
);

INVx1_ASAP7_75t_L g4731 ( 
.A(n_4712),
.Y(n_4731)
);

OAI22xp33_ASAP7_75t_L g4732 ( 
.A1(n_4704),
.A2(n_4612),
.B1(n_4546),
.B2(n_4558),
.Y(n_4732)
);

INVx2_ASAP7_75t_SL g4733 ( 
.A(n_4724),
.Y(n_4733)
);

AND2x2_ASAP7_75t_L g4734 ( 
.A(n_4723),
.B(n_4707),
.Y(n_4734)
);

AND2x2_ASAP7_75t_L g4735 ( 
.A(n_4721),
.B(n_4706),
.Y(n_4735)
);

HB1xp67_ASAP7_75t_L g4736 ( 
.A(n_4729),
.Y(n_4736)
);

INVx2_ASAP7_75t_L g4737 ( 
.A(n_4720),
.Y(n_4737)
);

INVx1_ASAP7_75t_SL g4738 ( 
.A(n_4730),
.Y(n_4738)
);

NAND2xp5_ASAP7_75t_L g4739 ( 
.A(n_4725),
.B(n_4706),
.Y(n_4739)
);

OR2x2_ASAP7_75t_L g4740 ( 
.A(n_4726),
.B(n_4718),
.Y(n_4740)
);

HB1xp67_ASAP7_75t_L g4741 ( 
.A(n_4731),
.Y(n_4741)
);

NAND2xp5_ASAP7_75t_L g4742 ( 
.A(n_4728),
.B(n_4716),
.Y(n_4742)
);

OAI22xp5_ASAP7_75t_L g4743 ( 
.A1(n_4738),
.A2(n_4739),
.B1(n_4736),
.B2(n_4722),
.Y(n_4743)
);

OAI21xp33_ASAP7_75t_L g4744 ( 
.A1(n_4734),
.A2(n_4702),
.B(n_4727),
.Y(n_4744)
);

OR2x2_ASAP7_75t_L g4745 ( 
.A(n_4738),
.B(n_4718),
.Y(n_4745)
);

NAND2xp5_ASAP7_75t_L g4746 ( 
.A(n_4735),
.B(n_4715),
.Y(n_4746)
);

INVx1_ASAP7_75t_L g4747 ( 
.A(n_4740),
.Y(n_4747)
);

INVx1_ASAP7_75t_L g4748 ( 
.A(n_4741),
.Y(n_4748)
);

NAND3xp33_ASAP7_75t_L g4749 ( 
.A(n_4733),
.B(n_4715),
.C(n_4709),
.Y(n_4749)
);

AOI222xp33_ASAP7_75t_L g4750 ( 
.A1(n_4737),
.A2(n_4643),
.B1(n_4637),
.B2(n_4630),
.C1(n_4607),
.C2(n_4680),
.Y(n_4750)
);

OAI21xp5_ASAP7_75t_SL g4751 ( 
.A1(n_4742),
.A2(n_4713),
.B(n_4717),
.Y(n_4751)
);

INVx1_ASAP7_75t_SL g4752 ( 
.A(n_4734),
.Y(n_4752)
);

OAI221xp5_ASAP7_75t_SL g4753 ( 
.A1(n_4738),
.A2(n_4732),
.B1(n_4708),
.B2(n_4643),
.C(n_4699),
.Y(n_4753)
);

INVx1_ASAP7_75t_L g4754 ( 
.A(n_4734),
.Y(n_4754)
);

INVxp67_ASAP7_75t_L g4755 ( 
.A(n_4734),
.Y(n_4755)
);

AND2x2_ASAP7_75t_L g4756 ( 
.A(n_4752),
.B(n_4609),
.Y(n_4756)
);

AND2x2_ASAP7_75t_L g4757 ( 
.A(n_4755),
.B(n_4609),
.Y(n_4757)
);

OAI21xp5_ASAP7_75t_L g4758 ( 
.A1(n_4749),
.A2(n_4657),
.B(n_4719),
.Y(n_4758)
);

INVx2_ASAP7_75t_L g4759 ( 
.A(n_4745),
.Y(n_4759)
);

NAND2xp5_ASAP7_75t_L g4760 ( 
.A(n_4747),
.B(n_4621),
.Y(n_4760)
);

INVx1_ASAP7_75t_L g4761 ( 
.A(n_4746),
.Y(n_4761)
);

NAND2xp5_ASAP7_75t_L g4762 ( 
.A(n_4751),
.B(n_4693),
.Y(n_4762)
);

INVx1_ASAP7_75t_L g4763 ( 
.A(n_4754),
.Y(n_4763)
);

AOI31xp33_ASAP7_75t_L g4764 ( 
.A1(n_4743),
.A2(n_4698),
.A3(n_4657),
.B(n_4525),
.Y(n_4764)
);

NAND2xp5_ASAP7_75t_L g4765 ( 
.A(n_4748),
.B(n_4647),
.Y(n_4765)
);

AND2x4_ASAP7_75t_L g4766 ( 
.A(n_4759),
.B(n_4756),
.Y(n_4766)
);

NAND2xp5_ASAP7_75t_L g4767 ( 
.A(n_4757),
.B(n_4744),
.Y(n_4767)
);

AND2x2_ASAP7_75t_L g4768 ( 
.A(n_4761),
.B(n_4570),
.Y(n_4768)
);

NOR2x1p5_ASAP7_75t_L g4769 ( 
.A(n_4762),
.B(n_4677),
.Y(n_4769)
);

INVx1_ASAP7_75t_SL g4770 ( 
.A(n_4760),
.Y(n_4770)
);

NAND2xp33_ASAP7_75t_SL g4771 ( 
.A(n_4763),
.B(n_4512),
.Y(n_4771)
);

OR2x2_ASAP7_75t_L g4772 ( 
.A(n_4764),
.B(n_4753),
.Y(n_4772)
);

INVx2_ASAP7_75t_L g4773 ( 
.A(n_4765),
.Y(n_4773)
);

INVx1_ASAP7_75t_L g4774 ( 
.A(n_4764),
.Y(n_4774)
);

OAI211xp5_ASAP7_75t_L g4775 ( 
.A1(n_4767),
.A2(n_4758),
.B(n_4750),
.C(n_4677),
.Y(n_4775)
);

NAND3xp33_ASAP7_75t_L g4776 ( 
.A(n_4774),
.B(n_4663),
.C(n_4655),
.Y(n_4776)
);

NAND3xp33_ASAP7_75t_SL g4777 ( 
.A(n_4770),
.B(n_4663),
.C(n_4655),
.Y(n_4777)
);

INVx1_ASAP7_75t_L g4778 ( 
.A(n_4768),
.Y(n_4778)
);

INVx1_ASAP7_75t_L g4779 ( 
.A(n_4766),
.Y(n_4779)
);

NAND2xp5_ASAP7_75t_L g4780 ( 
.A(n_4769),
.B(n_4647),
.Y(n_4780)
);

NAND4xp75_ASAP7_75t_L g4781 ( 
.A(n_4773),
.B(n_4680),
.C(n_4670),
.D(n_4648),
.Y(n_4781)
);

INVx2_ASAP7_75t_L g4782 ( 
.A(n_4772),
.Y(n_4782)
);

OAI21xp33_ASAP7_75t_L g4783 ( 
.A1(n_4771),
.A2(n_4670),
.B(n_4642),
.Y(n_4783)
);

OAI21xp33_ASAP7_75t_SL g4784 ( 
.A1(n_4767),
.A2(n_4569),
.B(n_4651),
.Y(n_4784)
);

INVx1_ASAP7_75t_L g4785 ( 
.A(n_4768),
.Y(n_4785)
);

NOR3xp33_ASAP7_75t_L g4786 ( 
.A(n_4770),
.B(n_4638),
.C(n_4651),
.Y(n_4786)
);

INVx1_ASAP7_75t_L g4787 ( 
.A(n_4768),
.Y(n_4787)
);

NAND4xp75_ASAP7_75t_L g4788 ( 
.A(n_4774),
.B(n_4652),
.C(n_4569),
.D(n_4550),
.Y(n_4788)
);

INVx1_ASAP7_75t_L g4789 ( 
.A(n_4779),
.Y(n_4789)
);

AND2x2_ASAP7_75t_L g4790 ( 
.A(n_4778),
.B(n_4570),
.Y(n_4790)
);

INVx1_ASAP7_75t_L g4791 ( 
.A(n_4781),
.Y(n_4791)
);

NOR2xp33_ASAP7_75t_L g4792 ( 
.A(n_4784),
.B(n_4647),
.Y(n_4792)
);

AOI21xp5_ASAP7_75t_L g4793 ( 
.A1(n_4775),
.A2(n_4557),
.B(n_4552),
.Y(n_4793)
);

INVxp67_ASAP7_75t_L g4794 ( 
.A(n_4777),
.Y(n_4794)
);

NAND2xp5_ASAP7_75t_SL g4795 ( 
.A(n_4783),
.B(n_4542),
.Y(n_4795)
);

INVxp67_ASAP7_75t_L g4796 ( 
.A(n_4785),
.Y(n_4796)
);

NOR2xp33_ASAP7_75t_L g4797 ( 
.A(n_4788),
.B(n_4476),
.Y(n_4797)
);

NAND4xp75_ASAP7_75t_L g4798 ( 
.A(n_4787),
.B(n_4607),
.C(n_4604),
.D(n_4537),
.Y(n_4798)
);

INVx1_ASAP7_75t_L g4799 ( 
.A(n_4780),
.Y(n_4799)
);

XOR2xp5_ASAP7_75t_L g4800 ( 
.A(n_4776),
.B(n_4539),
.Y(n_4800)
);

AND2x2_ASAP7_75t_SL g4801 ( 
.A(n_4782),
.B(n_4438),
.Y(n_4801)
);

INVx2_ASAP7_75t_L g4802 ( 
.A(n_4786),
.Y(n_4802)
);

NAND2xp5_ASAP7_75t_L g4803 ( 
.A(n_4781),
.B(n_4542),
.Y(n_4803)
);

NOR3xp33_ASAP7_75t_L g4804 ( 
.A(n_4777),
.B(n_4608),
.C(n_4580),
.Y(n_4804)
);

NAND2xp5_ASAP7_75t_SL g4805 ( 
.A(n_4779),
.B(n_4604),
.Y(n_4805)
);

NAND2xp5_ASAP7_75t_L g4806 ( 
.A(n_4781),
.B(n_4612),
.Y(n_4806)
);

INVx1_ASAP7_75t_L g4807 ( 
.A(n_4779),
.Y(n_4807)
);

NOR4xp25_ASAP7_75t_L g4808 ( 
.A(n_4779),
.B(n_4605),
.C(n_4599),
.D(n_4593),
.Y(n_4808)
);

AOI21xp5_ASAP7_75t_L g4809 ( 
.A1(n_4775),
.A2(n_4452),
.B(n_4605),
.Y(n_4809)
);

NOR3x1_ASAP7_75t_L g4810 ( 
.A(n_4775),
.B(n_4555),
.C(n_4562),
.Y(n_4810)
);

AND2x2_ASAP7_75t_L g4811 ( 
.A(n_4779),
.B(n_4549),
.Y(n_4811)
);

NOR3xp33_ASAP7_75t_L g4812 ( 
.A(n_4777),
.B(n_4608),
.C(n_4577),
.Y(n_4812)
);

OAI211xp5_ASAP7_75t_L g4813 ( 
.A1(n_4796),
.A2(n_4505),
.B(n_4596),
.C(n_4430),
.Y(n_4813)
);

AOI211xp5_ASAP7_75t_SL g4814 ( 
.A1(n_4791),
.A2(n_4460),
.B(n_4572),
.C(n_4563),
.Y(n_4814)
);

NOR3xp33_ASAP7_75t_L g4815 ( 
.A(n_4794),
.B(n_4597),
.C(n_4595),
.Y(n_4815)
);

AOI211xp5_ASAP7_75t_SL g4816 ( 
.A1(n_4797),
.A2(n_4460),
.B(n_4461),
.C(n_4459),
.Y(n_4816)
);

NAND4xp75_ASAP7_75t_L g4817 ( 
.A(n_4801),
.B(n_4459),
.C(n_4601),
.D(n_4600),
.Y(n_4817)
);

OAI211xp5_ASAP7_75t_L g4818 ( 
.A1(n_4803),
.A2(n_4416),
.B(n_4460),
.C(n_4501),
.Y(n_4818)
);

AOI211xp5_ASAP7_75t_L g4819 ( 
.A1(n_4795),
.A2(n_4593),
.B(n_4578),
.C(n_4487),
.Y(n_4819)
);

AOI22xp5_ASAP7_75t_L g4820 ( 
.A1(n_4802),
.A2(n_4792),
.B1(n_4790),
.B2(n_4800),
.Y(n_4820)
);

NOR4xp25_ASAP7_75t_L g4821 ( 
.A(n_4789),
.B(n_4536),
.C(n_4592),
.D(n_4487),
.Y(n_4821)
);

NAND5xp2_ASAP7_75t_L g4822 ( 
.A(n_4807),
.B(n_4482),
.C(n_4486),
.D(n_4446),
.E(n_4538),
.Y(n_4822)
);

AOI221xp5_ASAP7_75t_L g4823 ( 
.A1(n_4806),
.A2(n_4482),
.B1(n_4486),
.B2(n_4530),
.C(n_4538),
.Y(n_4823)
);

AOI211x1_ASAP7_75t_L g4824 ( 
.A1(n_4793),
.A2(n_4527),
.B(n_4529),
.C(n_4523),
.Y(n_4824)
);

INVx1_ASAP7_75t_L g4825 ( 
.A(n_4811),
.Y(n_4825)
);

NAND4xp25_ASAP7_75t_L g4826 ( 
.A(n_4805),
.B(n_4536),
.C(n_4442),
.D(n_4446),
.Y(n_4826)
);

NAND4xp75_ASAP7_75t_L g4827 ( 
.A(n_4810),
.B(n_4531),
.C(n_4479),
.D(n_4474),
.Y(n_4827)
);

NAND5xp2_ASAP7_75t_L g4828 ( 
.A(n_4804),
.B(n_4479),
.C(n_299),
.D(n_300),
.E(n_303),
.Y(n_4828)
);

NOR3xp33_ASAP7_75t_L g4829 ( 
.A(n_4799),
.B(n_4442),
.C(n_4474),
.Y(n_4829)
);

AND4x1_ASAP7_75t_L g4830 ( 
.A(n_4809),
.B(n_4808),
.C(n_4812),
.D(n_4798),
.Y(n_4830)
);

NOR2xp33_ASAP7_75t_SL g4831 ( 
.A(n_4808),
.B(n_4534),
.Y(n_4831)
);

NAND4xp25_ASAP7_75t_L g4832 ( 
.A(n_4797),
.B(n_4534),
.C(n_4493),
.D(n_4480),
.Y(n_4832)
);

AOI211xp5_ASAP7_75t_L g4833 ( 
.A1(n_4797),
.A2(n_4480),
.B(n_4493),
.C(n_4534),
.Y(n_4833)
);

NOR2xp33_ASAP7_75t_L g4834 ( 
.A(n_4794),
.B(n_4510),
.Y(n_4834)
);

NOR2xp67_ASAP7_75t_L g4835 ( 
.A(n_4803),
.B(n_298),
.Y(n_4835)
);

OAI221xp5_ASAP7_75t_L g4836 ( 
.A1(n_4800),
.A2(n_4377),
.B1(n_4507),
.B2(n_4520),
.C(n_4504),
.Y(n_4836)
);

NAND2xp5_ASAP7_75t_L g4837 ( 
.A(n_4801),
.B(n_4500),
.Y(n_4837)
);

INVx1_ASAP7_75t_L g4838 ( 
.A(n_4790),
.Y(n_4838)
);

AOI22x1_ASAP7_75t_L g4839 ( 
.A1(n_4800),
.A2(n_298),
.B1(n_304),
.B2(n_306),
.Y(n_4839)
);

NAND4xp25_ASAP7_75t_L g4840 ( 
.A(n_4820),
.B(n_306),
.C(n_307),
.D(n_308),
.Y(n_4840)
);

NAND3xp33_ASAP7_75t_SL g4841 ( 
.A(n_4830),
.B(n_4520),
.C(n_4504),
.Y(n_4841)
);

NAND2xp5_ASAP7_75t_SL g4842 ( 
.A(n_4825),
.B(n_4533),
.Y(n_4842)
);

OAI211xp5_ASAP7_75t_L g4843 ( 
.A1(n_4839),
.A2(n_308),
.B(n_309),
.C(n_310),
.Y(n_4843)
);

NOR3xp33_ASAP7_75t_L g4844 ( 
.A(n_4838),
.B(n_309),
.C(n_311),
.Y(n_4844)
);

AND2x2_ASAP7_75t_L g4845 ( 
.A(n_4821),
.B(n_4533),
.Y(n_4845)
);

AOI221xp5_ASAP7_75t_L g4846 ( 
.A1(n_4834),
.A2(n_4465),
.B1(n_314),
.B2(n_317),
.C(n_318),
.Y(n_4846)
);

NAND3xp33_ASAP7_75t_SL g4847 ( 
.A(n_4815),
.B(n_4465),
.C(n_313),
.Y(n_4847)
);

AND2x2_ASAP7_75t_L g4848 ( 
.A(n_4816),
.B(n_4377),
.Y(n_4848)
);

OAI211xp5_ASAP7_75t_SL g4849 ( 
.A1(n_4814),
.A2(n_4833),
.B(n_4837),
.C(n_4819),
.Y(n_4849)
);

INVx1_ASAP7_75t_L g4850 ( 
.A(n_4817),
.Y(n_4850)
);

INVxp33_ASAP7_75t_L g4851 ( 
.A(n_4835),
.Y(n_4851)
);

NAND2x1_ASAP7_75t_L g4852 ( 
.A(n_4824),
.B(n_4401),
.Y(n_4852)
);

NAND4xp25_ASAP7_75t_L g4853 ( 
.A(n_4828),
.B(n_317),
.C(n_319),
.D(n_320),
.Y(n_4853)
);

INVx2_ASAP7_75t_L g4854 ( 
.A(n_4827),
.Y(n_4854)
);

NAND4xp75_ASAP7_75t_L g4855 ( 
.A(n_4823),
.B(n_319),
.C(n_320),
.D(n_321),
.Y(n_4855)
);

OAI211xp5_ASAP7_75t_SL g4856 ( 
.A1(n_4829),
.A2(n_4836),
.B(n_4818),
.C(n_4831),
.Y(n_4856)
);

NOR2xp33_ASAP7_75t_L g4857 ( 
.A(n_4832),
.B(n_321),
.Y(n_4857)
);

NAND4xp25_ASAP7_75t_L g4858 ( 
.A(n_4826),
.B(n_4822),
.C(n_4813),
.D(n_326),
.Y(n_4858)
);

INVx1_ASAP7_75t_L g4859 ( 
.A(n_4825),
.Y(n_4859)
);

NAND4xp25_ASAP7_75t_L g4860 ( 
.A(n_4820),
.B(n_323),
.C(n_325),
.D(n_327),
.Y(n_4860)
);

NOR3x1_ASAP7_75t_L g4861 ( 
.A(n_4825),
.B(n_323),
.C(n_325),
.Y(n_4861)
);

INVx2_ASAP7_75t_L g4862 ( 
.A(n_4839),
.Y(n_4862)
);

OAI221xp5_ASAP7_75t_L g4863 ( 
.A1(n_4831),
.A2(n_4418),
.B1(n_330),
.B2(n_331),
.C(n_332),
.Y(n_4863)
);

AND2x2_ASAP7_75t_L g4864 ( 
.A(n_4848),
.B(n_4861),
.Y(n_4864)
);

NOR2x1_ASAP7_75t_L g4865 ( 
.A(n_4859),
.B(n_329),
.Y(n_4865)
);

AOI321xp33_ASAP7_75t_L g4866 ( 
.A1(n_4842),
.A2(n_329),
.A3(n_333),
.B1(n_334),
.B2(n_338),
.C(n_340),
.Y(n_4866)
);

OAI31xp33_ASAP7_75t_L g4867 ( 
.A1(n_4843),
.A2(n_4849),
.A3(n_4856),
.B(n_4863),
.Y(n_4867)
);

O2A1O1Ixp33_ASAP7_75t_L g4868 ( 
.A1(n_4854),
.A2(n_341),
.B(n_342),
.C(n_343),
.Y(n_4868)
);

INVx2_ASAP7_75t_L g4869 ( 
.A(n_4852),
.Y(n_4869)
);

INVx1_ASAP7_75t_SL g4870 ( 
.A(n_4855),
.Y(n_4870)
);

NAND3x1_ASAP7_75t_L g4871 ( 
.A(n_4850),
.B(n_341),
.C(n_345),
.Y(n_4871)
);

OAI21xp5_ASAP7_75t_SL g4872 ( 
.A1(n_4858),
.A2(n_346),
.B(n_347),
.Y(n_4872)
);

NOR2x1_ASAP7_75t_L g4873 ( 
.A(n_4840),
.B(n_348),
.Y(n_4873)
);

NAND2xp5_ASAP7_75t_SL g4874 ( 
.A(n_4862),
.B(n_349),
.Y(n_4874)
);

OAI22xp5_ASAP7_75t_L g4875 ( 
.A1(n_4857),
.A2(n_4372),
.B1(n_350),
.B2(n_349),
.Y(n_4875)
);

NAND2xp5_ASAP7_75t_L g4876 ( 
.A(n_4845),
.B(n_4851),
.Y(n_4876)
);

AOI22xp5_ASAP7_75t_L g4877 ( 
.A1(n_4847),
.A2(n_4841),
.B1(n_4853),
.B2(n_4846),
.Y(n_4877)
);

AO22x2_ASAP7_75t_L g4878 ( 
.A1(n_4844),
.A2(n_350),
.B1(n_4361),
.B2(n_357),
.Y(n_4878)
);

NOR2xp33_ASAP7_75t_L g4879 ( 
.A(n_4860),
.B(n_356),
.Y(n_4879)
);

OAI211xp5_ASAP7_75t_L g4880 ( 
.A1(n_4850),
.A2(n_1550),
.B(n_1542),
.C(n_1601),
.Y(n_4880)
);

AOI221xp5_ASAP7_75t_L g4881 ( 
.A1(n_4849),
.A2(n_1566),
.B1(n_1542),
.B2(n_1550),
.C(n_1551),
.Y(n_4881)
);

AOI22xp5_ASAP7_75t_L g4882 ( 
.A1(n_4864),
.A2(n_1566),
.B1(n_1550),
.B2(n_1551),
.Y(n_4882)
);

OAI22xp5_ASAP7_75t_L g4883 ( 
.A1(n_4876),
.A2(n_1566),
.B1(n_1550),
.B2(n_1551),
.Y(n_4883)
);

INVx2_ASAP7_75t_L g4884 ( 
.A(n_4865),
.Y(n_4884)
);

XOR2x1_ASAP7_75t_L g4885 ( 
.A(n_4869),
.B(n_364),
.Y(n_4885)
);

INVx2_ASAP7_75t_SL g4886 ( 
.A(n_4874),
.Y(n_4886)
);

NOR2x1_ASAP7_75t_L g4887 ( 
.A(n_4872),
.B(n_1551),
.Y(n_4887)
);

INVx1_ASAP7_75t_L g4888 ( 
.A(n_4871),
.Y(n_4888)
);

NOR2x1_ASAP7_75t_L g4889 ( 
.A(n_4868),
.B(n_1566),
.Y(n_4889)
);

OR2x2_ASAP7_75t_L g4890 ( 
.A(n_4870),
.B(n_368),
.Y(n_4890)
);

AND2x2_ASAP7_75t_L g4891 ( 
.A(n_4873),
.B(n_370),
.Y(n_4891)
);

OAI21xp5_ASAP7_75t_L g4892 ( 
.A1(n_4877),
.A2(n_1558),
.B(n_1406),
.Y(n_4892)
);

NOR2x1_ASAP7_75t_L g4893 ( 
.A(n_4880),
.B(n_4879),
.Y(n_4893)
);

NOR2x1_ASAP7_75t_L g4894 ( 
.A(n_4875),
.B(n_1573),
.Y(n_4894)
);

NAND3xp33_ASAP7_75t_L g4895 ( 
.A(n_4867),
.B(n_1574),
.C(n_1573),
.Y(n_4895)
);

HB1xp67_ASAP7_75t_L g4896 ( 
.A(n_4881),
.Y(n_4896)
);

INVx1_ASAP7_75t_L g4897 ( 
.A(n_4866),
.Y(n_4897)
);

AOI211xp5_ASAP7_75t_L g4898 ( 
.A1(n_4897),
.A2(n_4878),
.B(n_1601),
.C(n_1589),
.Y(n_4898)
);

A2O1A1Ixp33_ASAP7_75t_L g4899 ( 
.A1(n_4888),
.A2(n_4878),
.B(n_1573),
.C(n_1574),
.Y(n_4899)
);

OR2x2_ASAP7_75t_L g4900 ( 
.A(n_4884),
.B(n_375),
.Y(n_4900)
);

NAND4xp75_ASAP7_75t_L g4901 ( 
.A(n_4887),
.B(n_4893),
.C(n_4891),
.D(n_4886),
.Y(n_4901)
);

NOR3xp33_ASAP7_75t_SL g4902 ( 
.A(n_4892),
.B(n_380),
.C(n_386),
.Y(n_4902)
);

AOI211xp5_ASAP7_75t_L g4903 ( 
.A1(n_4896),
.A2(n_1601),
.B(n_1589),
.C(n_1586),
.Y(n_4903)
);

NAND3xp33_ASAP7_75t_L g4904 ( 
.A(n_4890),
.B(n_1574),
.C(n_1573),
.Y(n_4904)
);

NAND4xp25_ASAP7_75t_L g4905 ( 
.A(n_4889),
.B(n_4894),
.C(n_4895),
.D(n_4882),
.Y(n_4905)
);

NAND2xp5_ASAP7_75t_L g4906 ( 
.A(n_4885),
.B(n_390),
.Y(n_4906)
);

OR5x1_ASAP7_75t_L g4907 ( 
.A(n_4883),
.B(n_391),
.C(n_393),
.D(n_396),
.E(n_397),
.Y(n_4907)
);

NOR3xp33_ASAP7_75t_SL g4908 ( 
.A(n_4888),
.B(n_402),
.C(n_404),
.Y(n_4908)
);

NAND4xp25_ASAP7_75t_L g4909 ( 
.A(n_4888),
.B(n_406),
.C(n_407),
.D(n_408),
.Y(n_4909)
);

NOR3xp33_ASAP7_75t_L g4910 ( 
.A(n_4884),
.B(n_409),
.C(n_411),
.Y(n_4910)
);

OAI211xp5_ASAP7_75t_SL g4911 ( 
.A1(n_4888),
.A2(n_414),
.B(n_415),
.C(n_419),
.Y(n_4911)
);

INVx1_ASAP7_75t_L g4912 ( 
.A(n_4885),
.Y(n_4912)
);

INVx1_ASAP7_75t_L g4913 ( 
.A(n_4885),
.Y(n_4913)
);

NOR2x2_ASAP7_75t_L g4914 ( 
.A(n_4884),
.B(n_422),
.Y(n_4914)
);

NOR2x1p5_ASAP7_75t_L g4915 ( 
.A(n_4885),
.B(n_1574),
.Y(n_4915)
);

CKINVDCx16_ASAP7_75t_R g4916 ( 
.A(n_4912),
.Y(n_4916)
);

AOI22xp5_ASAP7_75t_L g4917 ( 
.A1(n_4913),
.A2(n_1581),
.B1(n_1586),
.B2(n_1589),
.Y(n_4917)
);

CKINVDCx5p33_ASAP7_75t_R g4918 ( 
.A(n_4915),
.Y(n_4918)
);

CKINVDCx5p33_ASAP7_75t_R g4919 ( 
.A(n_4906),
.Y(n_4919)
);

O2A1O1Ixp33_ASAP7_75t_L g4920 ( 
.A1(n_4899),
.A2(n_423),
.B(n_426),
.C(n_432),
.Y(n_4920)
);

CKINVDCx16_ASAP7_75t_R g4921 ( 
.A(n_4900),
.Y(n_4921)
);

BUFx2_ASAP7_75t_L g4922 ( 
.A(n_4914),
.Y(n_4922)
);

INVx1_ASAP7_75t_SL g4923 ( 
.A(n_4907),
.Y(n_4923)
);

CKINVDCx5p33_ASAP7_75t_R g4924 ( 
.A(n_4908),
.Y(n_4924)
);

INVx1_ASAP7_75t_L g4925 ( 
.A(n_4901),
.Y(n_4925)
);

INVx1_ASAP7_75t_L g4926 ( 
.A(n_4898),
.Y(n_4926)
);

INVxp67_ASAP7_75t_L g4927 ( 
.A(n_4904),
.Y(n_4927)
);

INVx2_ASAP7_75t_SL g4928 ( 
.A(n_4902),
.Y(n_4928)
);

OAI221xp5_ASAP7_75t_L g4929 ( 
.A1(n_4925),
.A2(n_4905),
.B1(n_4910),
.B2(n_4911),
.C(n_4909),
.Y(n_4929)
);

OAI22xp5_ASAP7_75t_SL g4930 ( 
.A1(n_4916),
.A2(n_4903),
.B1(n_439),
.B2(n_442),
.Y(n_4930)
);

OAI211xp5_ASAP7_75t_SL g4931 ( 
.A1(n_4926),
.A2(n_437),
.B(n_443),
.C(n_444),
.Y(n_4931)
);

OAI211xp5_ASAP7_75t_L g4932 ( 
.A1(n_4922),
.A2(n_1581),
.B(n_1586),
.C(n_1601),
.Y(n_4932)
);

INVx1_ASAP7_75t_L g4933 ( 
.A(n_4921),
.Y(n_4933)
);

INVx1_ASAP7_75t_L g4934 ( 
.A(n_4924),
.Y(n_4934)
);

INVx1_ASAP7_75t_L g4935 ( 
.A(n_4919),
.Y(n_4935)
);

AOI22xp5_ASAP7_75t_L g4936 ( 
.A1(n_4933),
.A2(n_4923),
.B1(n_4918),
.B2(n_4928),
.Y(n_4936)
);

OAI22xp5_ASAP7_75t_L g4937 ( 
.A1(n_4935),
.A2(n_4927),
.B1(n_4917),
.B2(n_4920),
.Y(n_4937)
);

INVx1_ASAP7_75t_L g4938 ( 
.A(n_4934),
.Y(n_4938)
);

AO22x2_ASAP7_75t_L g4939 ( 
.A1(n_4932),
.A2(n_446),
.B1(n_447),
.B2(n_448),
.Y(n_4939)
);

AND4x1_ASAP7_75t_L g4940 ( 
.A(n_4929),
.B(n_451),
.C(n_452),
.D(n_453),
.Y(n_4940)
);

CKINVDCx20_ASAP7_75t_R g4941 ( 
.A(n_4930),
.Y(n_4941)
);

AOI22xp5_ASAP7_75t_L g4942 ( 
.A1(n_4931),
.A2(n_1581),
.B1(n_1586),
.B2(n_1589),
.Y(n_4942)
);

AOI21xp5_ASAP7_75t_L g4943 ( 
.A1(n_4938),
.A2(n_1581),
.B(n_1606),
.Y(n_4943)
);

O2A1O1Ixp33_ASAP7_75t_L g4944 ( 
.A1(n_4937),
.A2(n_455),
.B(n_458),
.C(n_465),
.Y(n_4944)
);

NAND4xp75_ASAP7_75t_L g4945 ( 
.A(n_4936),
.B(n_466),
.C(n_468),
.D(n_469),
.Y(n_4945)
);

OAI211xp5_ASAP7_75t_SL g4946 ( 
.A1(n_4942),
.A2(n_471),
.B(n_479),
.C(n_482),
.Y(n_4946)
);

AOI221xp5_ASAP7_75t_L g4947 ( 
.A1(n_4941),
.A2(n_1607),
.B1(n_1606),
.B2(n_1596),
.C(n_1559),
.Y(n_4947)
);

OAI211xp5_ASAP7_75t_SL g4948 ( 
.A1(n_4939),
.A2(n_484),
.B(n_485),
.C(n_490),
.Y(n_4948)
);

AOI22xp5_ASAP7_75t_L g4949 ( 
.A1(n_4946),
.A2(n_4940),
.B1(n_1607),
.B2(n_1606),
.Y(n_4949)
);

NAND2xp5_ASAP7_75t_L g4950 ( 
.A(n_4945),
.B(n_4943),
.Y(n_4950)
);

HB1xp67_ASAP7_75t_L g4951 ( 
.A(n_4947),
.Y(n_4951)
);

INVx1_ASAP7_75t_L g4952 ( 
.A(n_4948),
.Y(n_4952)
);

HB1xp67_ASAP7_75t_L g4953 ( 
.A(n_4944),
.Y(n_4953)
);

OAI31xp33_ASAP7_75t_SL g4954 ( 
.A1(n_4952),
.A2(n_491),
.A3(n_492),
.B(n_493),
.Y(n_4954)
);

AOI21xp33_ASAP7_75t_L g4955 ( 
.A1(n_4953),
.A2(n_495),
.B(n_500),
.Y(n_4955)
);

AOI22xp5_ASAP7_75t_L g4956 ( 
.A1(n_4949),
.A2(n_1607),
.B1(n_1606),
.B2(n_1596),
.Y(n_4956)
);

XOR2xp5_ASAP7_75t_L g4957 ( 
.A(n_4950),
.B(n_503),
.Y(n_4957)
);

AOI22xp33_ASAP7_75t_L g4958 ( 
.A1(n_4957),
.A2(n_4951),
.B1(n_1401),
.B2(n_1406),
.Y(n_4958)
);

OR2x2_ASAP7_75t_L g4959 ( 
.A(n_4956),
.B(n_513),
.Y(n_4959)
);

NAND2x1p5_ASAP7_75t_L g4960 ( 
.A(n_4954),
.B(n_1401),
.Y(n_4960)
);

INVx1_ASAP7_75t_L g4961 ( 
.A(n_4955),
.Y(n_4961)
);

OAI22xp5_ASAP7_75t_SL g4962 ( 
.A1(n_4956),
.A2(n_1401),
.B1(n_1607),
.B2(n_1606),
.Y(n_4962)
);

XNOR2xp5_ASAP7_75t_L g4963 ( 
.A(n_4961),
.B(n_515),
.Y(n_4963)
);

OAI21xp5_ASAP7_75t_SL g4964 ( 
.A1(n_4960),
.A2(n_516),
.B(n_519),
.Y(n_4964)
);

OA22x2_ASAP7_75t_L g4965 ( 
.A1(n_4962),
.A2(n_524),
.B1(n_526),
.B2(n_528),
.Y(n_4965)
);

NAND2xp5_ASAP7_75t_L g4966 ( 
.A(n_4958),
.B(n_534),
.Y(n_4966)
);

NAND2xp5_ASAP7_75t_L g4967 ( 
.A(n_4959),
.B(n_535),
.Y(n_4967)
);

OAI21xp5_ASAP7_75t_L g4968 ( 
.A1(n_4961),
.A2(n_1435),
.B(n_1607),
.Y(n_4968)
);

NAND2xp5_ASAP7_75t_SL g4969 ( 
.A(n_4961),
.B(n_1435),
.Y(n_4969)
);

NAND2x1p5_ASAP7_75t_L g4970 ( 
.A(n_4961),
.B(n_1435),
.Y(n_4970)
);

INVxp67_ASAP7_75t_L g4971 ( 
.A(n_4961),
.Y(n_4971)
);

OAI21xp5_ASAP7_75t_L g4972 ( 
.A1(n_4961),
.A2(n_1435),
.B(n_1596),
.Y(n_4972)
);

OAI22xp5_ASAP7_75t_L g4973 ( 
.A1(n_4971),
.A2(n_1435),
.B1(n_1596),
.B2(n_1559),
.Y(n_4973)
);

OAI22xp5_ASAP7_75t_L g4974 ( 
.A1(n_4964),
.A2(n_1408),
.B1(n_1596),
.B2(n_1559),
.Y(n_4974)
);

AOI22xp5_ASAP7_75t_L g4975 ( 
.A1(n_4967),
.A2(n_4963),
.B1(n_4965),
.B2(n_4966),
.Y(n_4975)
);

OAI22xp5_ASAP7_75t_L g4976 ( 
.A1(n_4970),
.A2(n_1408),
.B1(n_1559),
.B2(n_1558),
.Y(n_4976)
);

OAI21xp5_ASAP7_75t_L g4977 ( 
.A1(n_4969),
.A2(n_1408),
.B(n_1559),
.Y(n_4977)
);

AOI22xp5_ASAP7_75t_L g4978 ( 
.A1(n_4968),
.A2(n_1406),
.B1(n_1558),
.B2(n_1519),
.Y(n_4978)
);

OAI22xp33_ASAP7_75t_L g4979 ( 
.A1(n_4972),
.A2(n_1406),
.B1(n_1558),
.B2(n_1519),
.Y(n_4979)
);

AOI22xp5_ASAP7_75t_L g4980 ( 
.A1(n_4971),
.A2(n_1406),
.B1(n_1558),
.B2(n_1519),
.Y(n_4980)
);

AOI22xp5_ASAP7_75t_L g4981 ( 
.A1(n_4971),
.A2(n_1401),
.B1(n_1519),
.B2(n_1500),
.Y(n_4981)
);

OAI22xp5_ASAP7_75t_L g4982 ( 
.A1(n_4971),
.A2(n_1401),
.B1(n_1519),
.B2(n_1500),
.Y(n_4982)
);

NAND2xp5_ASAP7_75t_L g4983 ( 
.A(n_4975),
.B(n_536),
.Y(n_4983)
);

BUFx3_ASAP7_75t_L g4984 ( 
.A(n_4978),
.Y(n_4984)
);

OAI22xp33_ASAP7_75t_L g4985 ( 
.A1(n_4974),
.A2(n_1408),
.B1(n_1500),
.B2(n_1494),
.Y(n_4985)
);

AOI21xp5_ASAP7_75t_L g4986 ( 
.A1(n_4976),
.A2(n_1408),
.B(n_1500),
.Y(n_4986)
);

NAND2xp5_ASAP7_75t_L g4987 ( 
.A(n_4977),
.B(n_541),
.Y(n_4987)
);

OAI221xp5_ASAP7_75t_L g4988 ( 
.A1(n_4980),
.A2(n_542),
.B1(n_543),
.B2(n_548),
.C(n_550),
.Y(n_4988)
);

NAND2xp5_ASAP7_75t_L g4989 ( 
.A(n_4979),
.B(n_553),
.Y(n_4989)
);

A2O1A1Ixp33_ASAP7_75t_L g4990 ( 
.A1(n_4981),
.A2(n_1468),
.B(n_1500),
.C(n_1494),
.Y(n_4990)
);

XNOR2xp5_ASAP7_75t_L g4991 ( 
.A(n_4984),
.B(n_4982),
.Y(n_4991)
);

OAI22xp33_ASAP7_75t_L g4992 ( 
.A1(n_4983),
.A2(n_4987),
.B1(n_4989),
.B2(n_4988),
.Y(n_4992)
);

OAI21xp5_ASAP7_75t_L g4993 ( 
.A1(n_4986),
.A2(n_4973),
.B(n_1468),
.Y(n_4993)
);

AOI22xp5_ASAP7_75t_L g4994 ( 
.A1(n_4985),
.A2(n_1468),
.B1(n_1494),
.B2(n_1492),
.Y(n_4994)
);

AOI221xp5_ASAP7_75t_L g4995 ( 
.A1(n_4992),
.A2(n_4990),
.B1(n_1468),
.B2(n_1484),
.C(n_1494),
.Y(n_4995)
);

AOI21xp33_ASAP7_75t_L g4996 ( 
.A1(n_4995),
.A2(n_4991),
.B(n_4993),
.Y(n_4996)
);

AOI211xp5_ASAP7_75t_L g4997 ( 
.A1(n_4996),
.A2(n_4994),
.B(n_555),
.C(n_556),
.Y(n_4997)
);


endmodule