module fake_jpeg_1287_n_150 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_150);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_150;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_7),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx2_ASAP7_75t_SL g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_1),
.B(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx2_ASAP7_75t_SL g30 ( 
.A(n_16),
.Y(n_30)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_31),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_2),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_32),
.B(n_35),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_14),
.B(n_6),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_8),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_36),
.B(n_41),
.Y(n_67)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

OR2x2_ASAP7_75t_SL g40 ( 
.A(n_21),
.B(n_3),
.Y(n_40)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_23),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_21),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_25),
.B(n_9),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_42),
.B(n_47),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

NAND2xp33_ASAP7_75t_SL g73 ( 
.A(n_44),
.B(n_11),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g45 ( 
.A1(n_22),
.A2(n_5),
.B(n_9),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_5),
.C(n_17),
.Y(n_62)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_28),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_45),
.A2(n_29),
.B1(n_16),
.B2(n_18),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_51),
.A2(n_55),
.B(n_60),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_31),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_52),
.B(n_50),
.Y(n_92)
);

CKINVDCx12_ASAP7_75t_R g54 ( 
.A(n_43),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_54),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_32),
.A2(n_29),
.B1(n_16),
.B2(n_18),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_62),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_30),
.A2(n_46),
.B1(n_20),
.B2(n_23),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_58),
.A2(n_59),
.B1(n_64),
.B2(n_39),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_49),
.A2(n_20),
.B1(n_19),
.B2(n_15),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_37),
.A2(n_19),
.B1(n_26),
.B2(n_17),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_33),
.A2(n_17),
.B1(n_10),
.B2(n_11),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_73),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_38),
.B(n_34),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_74),
.B(n_40),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_70),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_77),
.B(n_80),
.Y(n_98)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_81),
.B(n_83),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_57),
.B(n_44),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_82),
.Y(n_97)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_86),
.B(n_87),
.Y(n_107)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_88),
.A2(n_50),
.B1(n_69),
.B2(n_75),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_62),
.B(n_51),
.C(n_55),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_89),
.B(n_90),
.C(n_93),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_63),
.B(n_60),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_92),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_63),
.B(n_61),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_78),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_73),
.A2(n_67),
.B(n_75),
.Y(n_95)
);

O2A1O1Ixp33_ASAP7_75t_L g110 ( 
.A1(n_95),
.A2(n_82),
.B(n_84),
.C(n_90),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_100),
.A2(n_104),
.B1(n_90),
.B2(n_95),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_69),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_101),
.B(n_105),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_85),
.A2(n_56),
.B1(n_71),
.B2(n_88),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_76),
.B(n_71),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_76),
.B(n_71),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_106),
.B(n_111),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_108),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_110),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_76),
.B(n_82),
.C(n_93),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_101),
.A2(n_102),
.B(n_105),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_112),
.A2(n_114),
.B(n_117),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_102),
.A2(n_85),
.B(n_84),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_115),
.A2(n_100),
.B1(n_107),
.B2(n_96),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_93),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_116),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_110),
.A2(n_104),
.B(n_97),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_103),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_118),
.B(n_119),
.Y(n_127)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_99),
.Y(n_119)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_99),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_123),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_120),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_124),
.B(n_114),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_121),
.B(n_109),
.C(n_106),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_128),
.B(n_130),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_121),
.B(n_109),
.Y(n_130)
);

NOR4xp25_ASAP7_75t_L g131 ( 
.A(n_120),
.B(n_113),
.C(n_122),
.D(n_111),
.Y(n_131)
);

A2O1A1O1Ixp25_ASAP7_75t_L g137 ( 
.A1(n_131),
.A2(n_91),
.B(n_96),
.C(n_112),
.D(n_128),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_132),
.A2(n_115),
.B1(n_117),
.B2(n_122),
.Y(n_136)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_125),
.Y(n_133)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_133),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_135),
.B(n_136),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_137),
.A2(n_138),
.B(n_134),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_127),
.B(n_125),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_134),
.B(n_130),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_141),
.B(n_137),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_142),
.B(n_129),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_143),
.A2(n_144),
.B(n_129),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_140),
.B(n_126),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_145),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_146),
.B(n_139),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_147),
.C(n_141),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_136),
.Y(n_150)
);


endmodule