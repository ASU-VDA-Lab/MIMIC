module real_aes_6761_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_635;
wire n_503;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_555;
wire n_364;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_602;
wire n_552;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_713;
wire n_404;
wire n_288;
wire n_598;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_717;
wire n_359;
wire n_712;
wire n_183;
wire n_312;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_175;
wire n_168;
wire n_241;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g111 ( .A(n_0), .Y(n_111) );
INVx1_ASAP7_75t_L g490 ( .A(n_1), .Y(n_490) );
INVx1_ASAP7_75t_L g141 ( .A(n_2), .Y(n_141) );
AOI22xp33_ASAP7_75t_L g475 ( .A1(n_3), .A2(n_37), .B1(n_166), .B2(n_446), .Y(n_475) );
AOI21xp33_ASAP7_75t_L g185 ( .A1(n_4), .A2(n_157), .B(n_186), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_5), .B(n_155), .Y(n_501) );
AND2x6_ASAP7_75t_L g134 ( .A(n_6), .B(n_135), .Y(n_134) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_7), .A2(n_239), .B(n_240), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g112 ( .A(n_8), .B(n_38), .Y(n_112) );
INVx1_ASAP7_75t_L g191 ( .A(n_9), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_10), .B(n_220), .Y(n_219) );
INVx1_ASAP7_75t_L g126 ( .A(n_11), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_12), .B(n_147), .Y(n_454) );
INVx1_ASAP7_75t_L g245 ( .A(n_13), .Y(n_245) );
INVx1_ASAP7_75t_L g484 ( .A(n_14), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_15), .B(n_122), .Y(n_506) );
AO32x2_ASAP7_75t_L g473 ( .A1(n_16), .A2(n_121), .A3(n_155), .B1(n_448), .B2(n_474), .Y(n_473) );
NAND2xp5_ASAP7_75t_SL g457 ( .A(n_17), .B(n_166), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_18), .B(n_162), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_19), .B(n_122), .Y(n_492) );
AOI222xp33_ASAP7_75t_L g100 ( .A1(n_20), .A2(n_101), .B1(n_717), .B2(n_726), .C1(n_738), .C2(n_744), .Y(n_100) );
OAI22xp5_ASAP7_75t_SL g730 ( .A1(n_20), .A2(n_30), .B1(n_731), .B2(n_732), .Y(n_730) );
CKINVDCx20_ASAP7_75t_R g731 ( .A(n_20), .Y(n_731) );
AOI22xp33_ASAP7_75t_L g477 ( .A1(n_21), .A2(n_49), .B1(n_166), .B2(n_446), .Y(n_477) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_22), .B(n_157), .Y(n_202) );
AOI22xp33_ASAP7_75t_SL g447 ( .A1(n_23), .A2(n_76), .B1(n_147), .B2(n_166), .Y(n_447) );
NAND2xp5_ASAP7_75t_SL g469 ( .A(n_24), .B(n_166), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_25), .B(n_169), .Y(n_168) );
A2O1A1Ixp33_ASAP7_75t_L g242 ( .A1(n_26), .A2(n_243), .B(n_244), .C(n_246), .Y(n_242) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_27), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_28), .B(n_152), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_29), .B(n_145), .Y(n_144) );
CKINVDCx20_ASAP7_75t_R g732 ( .A(n_30), .Y(n_732) );
INVx1_ASAP7_75t_L g180 ( .A(n_31), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_32), .B(n_152), .Y(n_471) );
INVx2_ASAP7_75t_L g132 ( .A(n_33), .Y(n_132) );
NAND2xp5_ASAP7_75t_SL g520 ( .A(n_34), .B(n_166), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_35), .B(n_152), .Y(n_459) );
A2O1A1Ixp33_ASAP7_75t_L g203 ( .A1(n_36), .A2(n_134), .B(n_137), .C(n_204), .Y(n_203) );
INVx1_ASAP7_75t_L g178 ( .A(n_39), .Y(n_178) );
NAND2xp5_ASAP7_75t_SL g232 ( .A(n_40), .B(n_145), .Y(n_232) );
CKINVDCx20_ASAP7_75t_R g737 ( .A(n_41), .Y(n_737) );
NAND2xp5_ASAP7_75t_SL g496 ( .A(n_42), .B(n_166), .Y(n_496) );
AOI22xp33_ASAP7_75t_L g445 ( .A1(n_43), .A2(n_86), .B1(n_209), .B2(n_446), .Y(n_445) );
NAND2xp5_ASAP7_75t_SL g499 ( .A(n_44), .B(n_166), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_45), .B(n_166), .Y(n_485) );
CKINVDCx16_ASAP7_75t_R g181 ( .A(n_46), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_47), .B(n_489), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_48), .B(n_157), .Y(n_222) );
AOI22xp33_ASAP7_75t_SL g510 ( .A1(n_50), .A2(n_60), .B1(n_147), .B2(n_166), .Y(n_510) );
AOI222xp33_ASAP7_75t_SL g102 ( .A1(n_51), .A2(n_103), .B1(n_106), .B2(n_710), .C1(n_711), .C2(n_713), .Y(n_102) );
AOI22xp5_ASAP7_75t_L g175 ( .A1(n_52), .A2(n_137), .B1(n_147), .B2(n_176), .Y(n_175) );
CKINVDCx20_ASAP7_75t_R g212 ( .A(n_53), .Y(n_212) );
NAND2xp5_ASAP7_75t_SL g453 ( .A(n_54), .B(n_166), .Y(n_453) );
CKINVDCx16_ASAP7_75t_R g128 ( .A(n_55), .Y(n_128) );
NAND2xp5_ASAP7_75t_SL g524 ( .A(n_56), .B(n_166), .Y(n_524) );
A2O1A1Ixp33_ASAP7_75t_L g188 ( .A1(n_57), .A2(n_165), .B(n_189), .C(n_190), .Y(n_188) );
CKINVDCx20_ASAP7_75t_R g236 ( .A(n_58), .Y(n_236) );
INVx1_ASAP7_75t_L g187 ( .A(n_59), .Y(n_187) );
INVx1_ASAP7_75t_L g135 ( .A(n_61), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_62), .B(n_166), .Y(n_491) );
INVx1_ASAP7_75t_L g125 ( .A(n_63), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g722 ( .A(n_64), .Y(n_722) );
AO32x2_ASAP7_75t_L g443 ( .A1(n_65), .A2(n_155), .A3(n_214), .B1(n_444), .B2(n_448), .Y(n_443) );
INVx1_ASAP7_75t_L g523 ( .A(n_66), .Y(n_523) );
INVx1_ASAP7_75t_L g466 ( .A(n_67), .Y(n_466) );
OAI22xp5_ASAP7_75t_L g103 ( .A1(n_68), .A2(n_75), .B1(n_104), .B2(n_105), .Y(n_103) );
INVx1_ASAP7_75t_L g105 ( .A(n_68), .Y(n_105) );
A2O1A1Ixp33_ASAP7_75t_SL g161 ( .A1(n_69), .A2(n_162), .B(n_163), .C(n_165), .Y(n_161) );
INVxp67_ASAP7_75t_L g164 ( .A(n_70), .Y(n_164) );
NAND2xp5_ASAP7_75t_SL g467 ( .A(n_71), .B(n_147), .Y(n_467) );
INVx1_ASAP7_75t_L g721 ( .A(n_72), .Y(n_721) );
CKINVDCx20_ASAP7_75t_R g183 ( .A(n_73), .Y(n_183) );
INVx1_ASAP7_75t_L g229 ( .A(n_74), .Y(n_229) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_75), .Y(n_104) );
A2O1A1Ixp33_ASAP7_75t_L g230 ( .A1(n_77), .A2(n_134), .B(n_137), .C(n_231), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_78), .B(n_446), .Y(n_458) );
NAND2xp5_ASAP7_75t_SL g470 ( .A(n_79), .B(n_147), .Y(n_470) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_80), .B(n_142), .Y(n_205) );
INVx2_ASAP7_75t_L g123 ( .A(n_81), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_82), .B(n_162), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_83), .B(n_147), .Y(n_497) );
A2O1A1Ixp33_ASAP7_75t_L g136 ( .A1(n_84), .A2(n_134), .B(n_137), .C(n_140), .Y(n_136) );
OR2x2_ASAP7_75t_L g109 ( .A(n_85), .B(n_110), .Y(n_109) );
INVx2_ASAP7_75t_L g434 ( .A(n_85), .Y(n_434) );
OR2x2_ASAP7_75t_L g725 ( .A(n_85), .B(n_716), .Y(n_725) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_87), .A2(n_99), .B1(n_147), .B2(n_148), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_88), .B(n_152), .Y(n_192) );
CKINVDCx20_ASAP7_75t_R g150 ( .A(n_89), .Y(n_150) );
A2O1A1Ixp33_ASAP7_75t_L g216 ( .A1(n_90), .A2(n_134), .B(n_137), .C(n_217), .Y(n_216) );
CKINVDCx20_ASAP7_75t_R g224 ( .A(n_91), .Y(n_224) );
INVx1_ASAP7_75t_L g160 ( .A(n_92), .Y(n_160) );
CKINVDCx16_ASAP7_75t_R g241 ( .A(n_93), .Y(n_241) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_94), .B(n_142), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_95), .B(n_147), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_96), .B(n_155), .Y(n_247) );
AOI21xp5_ASAP7_75t_L g156 ( .A1(n_97), .A2(n_157), .B(n_158), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_98), .B(n_721), .Y(n_720) );
INVxp67_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
INVx1_ASAP7_75t_L g710 ( .A(n_103), .Y(n_710) );
OAI22xp5_ASAP7_75t_L g106 ( .A1(n_107), .A2(n_113), .B1(n_431), .B2(n_435), .Y(n_106) );
OAI22xp5_ASAP7_75t_SL g711 ( .A1(n_107), .A2(n_114), .B1(n_436), .B2(n_712), .Y(n_711) );
INVx2_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
OR2x2_ASAP7_75t_L g433 ( .A(n_110), .B(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g716 ( .A(n_110), .Y(n_716) );
AND2x2_ASAP7_75t_L g110 ( .A(n_111), .B(n_112), .Y(n_110) );
OAI22xp5_ASAP7_75t_SL g728 ( .A1(n_113), .A2(n_114), .B1(n_729), .B2(n_730), .Y(n_728) );
INVx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
OR4x1_ASAP7_75t_L g114 ( .A(n_115), .B(n_320), .C(n_380), .D(n_407), .Y(n_114) );
NAND4xp25_ASAP7_75t_SL g115 ( .A(n_116), .B(n_268), .C(n_299), .D(n_316), .Y(n_115) );
O2A1O1Ixp33_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_193), .B(n_195), .C(n_248), .Y(n_116) );
NOR2xp33_ASAP7_75t_L g117 ( .A(n_118), .B(n_171), .Y(n_117) );
INVx1_ASAP7_75t_L g310 ( .A(n_118), .Y(n_310) );
OAI22xp5_ASAP7_75t_L g428 ( .A1(n_118), .A2(n_351), .B1(n_399), .B2(n_429), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g118 ( .A(n_119), .B(n_153), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_119), .B(n_255), .Y(n_254) );
OR2x2_ASAP7_75t_L g261 ( .A(n_119), .B(n_173), .Y(n_261) );
AND2x2_ASAP7_75t_L g303 ( .A(n_119), .B(n_304), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_119), .B(n_194), .Y(n_315) );
INVx1_ASAP7_75t_L g355 ( .A(n_119), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_119), .B(n_409), .Y(n_408) );
INVx3_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
AND2x2_ASAP7_75t_L g283 ( .A(n_120), .B(n_173), .Y(n_283) );
INVx3_ASAP7_75t_L g287 ( .A(n_120), .Y(n_287) );
NAND2xp5_ASAP7_75t_SL g344 ( .A(n_120), .B(n_345), .Y(n_344) );
AO21x2_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_127), .B(n_149), .Y(n_120) );
AO21x2_ASAP7_75t_L g173 ( .A1(n_121), .A2(n_174), .B(n_182), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g182 ( .A(n_121), .B(n_183), .Y(n_182) );
INVx2_ASAP7_75t_L g210 ( .A(n_121), .Y(n_210) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_122), .Y(n_155) );
AND2x2_ASAP7_75t_L g122 ( .A(n_123), .B(n_124), .Y(n_122) );
AND2x2_ASAP7_75t_SL g152 ( .A(n_123), .B(n_124), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_125), .B(n_126), .Y(n_124) );
OAI21xp5_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_129), .B(n_136), .Y(n_127) );
OAI22xp33_ASAP7_75t_L g174 ( .A1(n_129), .A2(n_167), .B1(n_175), .B2(n_181), .Y(n_174) );
OAI21xp5_ASAP7_75t_L g228 ( .A1(n_129), .A2(n_229), .B(n_230), .Y(n_228) );
NAND2x1p5_ASAP7_75t_L g129 ( .A(n_130), .B(n_134), .Y(n_129) );
AND2x4_ASAP7_75t_L g157 ( .A(n_130), .B(n_134), .Y(n_157) );
AND2x2_ASAP7_75t_L g130 ( .A(n_131), .B(n_133), .Y(n_130) );
INVx1_ASAP7_75t_L g489 ( .A(n_131), .Y(n_489) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx2_ASAP7_75t_L g138 ( .A(n_132), .Y(n_138) );
INVx1_ASAP7_75t_L g148 ( .A(n_132), .Y(n_148) );
INVx1_ASAP7_75t_L g139 ( .A(n_133), .Y(n_139) );
INVx3_ASAP7_75t_L g143 ( .A(n_133), .Y(n_143) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_133), .Y(n_145) );
INVx1_ASAP7_75t_L g162 ( .A(n_133), .Y(n_162) );
BUFx6f_ASAP7_75t_L g177 ( .A(n_133), .Y(n_177) );
INVx4_ASAP7_75t_SL g167 ( .A(n_134), .Y(n_167) );
BUFx3_ASAP7_75t_L g448 ( .A(n_134), .Y(n_448) );
OAI21xp5_ASAP7_75t_L g451 ( .A1(n_134), .A2(n_452), .B(n_456), .Y(n_451) );
OAI21xp5_ASAP7_75t_L g464 ( .A1(n_134), .A2(n_465), .B(n_468), .Y(n_464) );
OAI21xp5_ASAP7_75t_L g482 ( .A1(n_134), .A2(n_483), .B(n_487), .Y(n_482) );
OAI21xp5_ASAP7_75t_L g494 ( .A1(n_134), .A2(n_495), .B(n_498), .Y(n_494) );
INVx5_ASAP7_75t_L g159 ( .A(n_137), .Y(n_159) );
AND2x6_ASAP7_75t_L g137 ( .A(n_138), .B(n_139), .Y(n_137) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_138), .Y(n_166) );
BUFx3_ASAP7_75t_L g209 ( .A(n_138), .Y(n_209) );
INVx1_ASAP7_75t_L g446 ( .A(n_138), .Y(n_446) );
O2A1O1Ixp33_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_142), .B(n_144), .C(n_146), .Y(n_140) );
O2A1O1Ixp5_ASAP7_75t_SL g465 ( .A1(n_142), .A2(n_165), .B(n_466), .C(n_467), .Y(n_465) );
INVx2_ASAP7_75t_L g476 ( .A(n_142), .Y(n_476) );
AOI21xp5_ASAP7_75t_L g495 ( .A1(n_142), .A2(n_496), .B(n_497), .Y(n_495) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_142), .A2(n_520), .B(n_521), .Y(n_519) );
INVx5_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
NOR2xp33_ASAP7_75t_L g163 ( .A(n_143), .B(n_164), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g190 ( .A(n_143), .B(n_191), .Y(n_190) );
OAI22xp5_ASAP7_75t_SL g444 ( .A1(n_143), .A2(n_145), .B1(n_445), .B2(n_447), .Y(n_444) );
INVx2_ASAP7_75t_L g189 ( .A(n_145), .Y(n_189) );
INVx4_ASAP7_75t_L g220 ( .A(n_145), .Y(n_220) );
OAI22xp5_ASAP7_75t_L g474 ( .A1(n_145), .A2(n_475), .B1(n_476), .B2(n_477), .Y(n_474) );
OAI22xp5_ASAP7_75t_L g508 ( .A1(n_145), .A2(n_476), .B1(n_509), .B2(n_510), .Y(n_508) );
O2A1O1Ixp33_ASAP7_75t_L g483 ( .A1(n_146), .A2(n_484), .B(n_485), .C(n_486), .Y(n_483) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx3_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
NOR2xp33_ASAP7_75t_L g149 ( .A(n_150), .B(n_151), .Y(n_149) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_151), .B(n_224), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_151), .B(n_236), .Y(n_235) );
INVx1_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g214 ( .A(n_152), .Y(n_214) );
OA21x2_ASAP7_75t_L g237 ( .A1(n_152), .A2(n_238), .B(n_247), .Y(n_237) );
OA21x2_ASAP7_75t_L g450 ( .A1(n_152), .A2(n_451), .B(n_459), .Y(n_450) );
OA21x2_ASAP7_75t_L g463 ( .A1(n_152), .A2(n_464), .B(n_471), .Y(n_463) );
AND2x2_ASAP7_75t_L g374 ( .A(n_153), .B(n_184), .Y(n_374) );
NOR2xp33_ASAP7_75t_L g393 ( .A(n_153), .B(n_287), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_153), .B(n_402), .Y(n_401) );
INVx3_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
AND2x2_ASAP7_75t_L g194 ( .A(n_154), .B(n_173), .Y(n_194) );
INVx1_ASAP7_75t_L g256 ( .A(n_154), .Y(n_256) );
BUFx2_ASAP7_75t_L g260 ( .A(n_154), .Y(n_260) );
AND2x2_ASAP7_75t_L g304 ( .A(n_154), .B(n_172), .Y(n_304) );
OR2x2_ASAP7_75t_L g343 ( .A(n_154), .B(n_172), .Y(n_343) );
AND2x2_ASAP7_75t_L g368 ( .A(n_154), .B(n_184), .Y(n_368) );
AND2x2_ASAP7_75t_L g427 ( .A(n_154), .B(n_257), .Y(n_427) );
OA21x2_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_156), .B(n_168), .Y(n_154) );
INVx4_ASAP7_75t_L g170 ( .A(n_155), .Y(n_170) );
OA21x2_ASAP7_75t_L g493 ( .A1(n_155), .A2(n_494), .B(n_501), .Y(n_493) );
BUFx2_ASAP7_75t_L g239 ( .A(n_157), .Y(n_239) );
O2A1O1Ixp33_ASAP7_75t_L g158 ( .A1(n_159), .A2(n_160), .B(n_161), .C(n_167), .Y(n_158) );
O2A1O1Ixp33_ASAP7_75t_L g186 ( .A1(n_159), .A2(n_167), .B(n_187), .C(n_188), .Y(n_186) );
O2A1O1Ixp33_ASAP7_75t_L g240 ( .A1(n_159), .A2(n_167), .B(n_241), .C(n_242), .Y(n_240) );
INVx1_ASAP7_75t_L g455 ( .A(n_162), .Y(n_455) );
INVx3_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
HB1xp67_ASAP7_75t_L g221 ( .A(n_166), .Y(n_221) );
OA21x2_ASAP7_75t_L g184 ( .A1(n_169), .A2(n_185), .B(n_192), .Y(n_184) );
INVx3_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
NOR2xp33_ASAP7_75t_SL g211 ( .A(n_170), .B(n_212), .Y(n_211) );
NAND3xp33_ASAP7_75t_L g507 ( .A(n_170), .B(n_448), .C(n_508), .Y(n_507) );
AO21x1_ASAP7_75t_L g554 ( .A1(n_170), .A2(n_508), .B(n_555), .Y(n_554) );
INVx1_ASAP7_75t_L g402 ( .A(n_171), .Y(n_402) );
OR2x2_ASAP7_75t_L g171 ( .A(n_172), .B(n_184), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_172), .B(n_184), .Y(n_288) );
AND2x2_ASAP7_75t_L g298 ( .A(n_172), .B(n_287), .Y(n_298) );
BUFx2_ASAP7_75t_L g309 ( .A(n_172), .Y(n_309) );
INVx3_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
AND2x2_ASAP7_75t_L g331 ( .A(n_173), .B(n_184), .Y(n_331) );
HB1xp67_ASAP7_75t_L g386 ( .A(n_173), .Y(n_386) );
OAI22xp5_ASAP7_75t_SL g176 ( .A1(n_177), .A2(n_178), .B1(n_179), .B2(n_180), .Y(n_176) );
INVx2_ASAP7_75t_L g179 ( .A(n_177), .Y(n_179) );
INVx4_ASAP7_75t_L g243 ( .A(n_177), .Y(n_243) );
AND2x2_ASAP7_75t_SL g193 ( .A(n_184), .B(n_194), .Y(n_193) );
INVx1_ASAP7_75t_SL g257 ( .A(n_184), .Y(n_257) );
BUFx2_ASAP7_75t_L g282 ( .A(n_184), .Y(n_282) );
INVx2_ASAP7_75t_L g301 ( .A(n_184), .Y(n_301) );
AND2x2_ASAP7_75t_L g363 ( .A(n_184), .B(n_287), .Y(n_363) );
AOI21xp5_ASAP7_75t_L g456 ( .A1(n_189), .A2(n_457), .B(n_458), .Y(n_456) );
O2A1O1Ixp5_ASAP7_75t_L g522 ( .A1(n_189), .A2(n_488), .B(n_523), .C(n_524), .Y(n_522) );
AOI321xp33_ASAP7_75t_L g382 ( .A1(n_193), .A2(n_383), .A3(n_384), .B1(n_385), .B2(n_387), .C(n_388), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_194), .B(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_194), .B(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_L g376 ( .A(n_194), .B(n_355), .Y(n_376) );
AND2x2_ASAP7_75t_L g409 ( .A(n_194), .B(n_301), .Y(n_409) );
INVx1_ASAP7_75t_SL g195 ( .A(n_196), .Y(n_195) );
OR2x2_ASAP7_75t_L g196 ( .A(n_197), .B(n_225), .Y(n_196) );
OR2x2_ASAP7_75t_L g311 ( .A(n_197), .B(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
AND2x2_ASAP7_75t_L g198 ( .A(n_199), .B(n_213), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
INVx3_ASAP7_75t_L g263 ( .A(n_200), .Y(n_263) );
AND2x2_ASAP7_75t_L g273 ( .A(n_200), .B(n_227), .Y(n_273) );
AND2x2_ASAP7_75t_L g278 ( .A(n_200), .B(n_253), .Y(n_278) );
INVx1_ASAP7_75t_L g295 ( .A(n_200), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_200), .B(n_276), .Y(n_314) );
AND2x2_ASAP7_75t_L g319 ( .A(n_200), .B(n_252), .Y(n_319) );
OR2x2_ASAP7_75t_L g351 ( .A(n_200), .B(n_340), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_200), .B(n_264), .Y(n_390) );
AND2x2_ASAP7_75t_L g424 ( .A(n_200), .B(n_250), .Y(n_424) );
OR2x6_ASAP7_75t_L g200 ( .A(n_201), .B(n_211), .Y(n_200) );
AOI21xp5_ASAP7_75t_SL g201 ( .A1(n_202), .A2(n_203), .B(n_210), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_206), .B(n_207), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_207), .A2(n_232), .B(n_233), .Y(n_231) );
INVx2_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx1_ASAP7_75t_L g246 ( .A(n_209), .Y(n_246) );
INVx1_ASAP7_75t_L g234 ( .A(n_210), .Y(n_234) );
OA21x2_ASAP7_75t_L g481 ( .A1(n_210), .A2(n_482), .B(n_492), .Y(n_481) );
OA21x2_ASAP7_75t_L g517 ( .A1(n_210), .A2(n_518), .B(n_525), .Y(n_517) );
INVx1_ASAP7_75t_L g251 ( .A(n_213), .Y(n_251) );
INVx2_ASAP7_75t_L g266 ( .A(n_213), .Y(n_266) );
AND2x2_ASAP7_75t_L g306 ( .A(n_213), .B(n_277), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_213), .B(n_253), .Y(n_328) );
AO21x2_ASAP7_75t_L g213 ( .A1(n_214), .A2(n_215), .B(n_223), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_216), .B(n_222), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_218), .A2(n_219), .B(n_221), .Y(n_217) );
INVx1_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
AND2x2_ASAP7_75t_L g412 ( .A(n_226), .B(n_263), .Y(n_412) );
AND2x2_ASAP7_75t_L g226 ( .A(n_227), .B(n_237), .Y(n_226) );
INVx2_ASAP7_75t_L g253 ( .A(n_227), .Y(n_253) );
AND2x2_ASAP7_75t_L g406 ( .A(n_227), .B(n_266), .Y(n_406) );
AO21x2_ASAP7_75t_L g227 ( .A1(n_228), .A2(n_234), .B(n_235), .Y(n_227) );
AND2x2_ASAP7_75t_L g252 ( .A(n_237), .B(n_253), .Y(n_252) );
INVx2_ASAP7_75t_L g267 ( .A(n_237), .Y(n_267) );
INVx1_ASAP7_75t_L g277 ( .A(n_237), .Y(n_277) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_243), .B(n_245), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g468 ( .A1(n_243), .A2(n_469), .B(n_470), .Y(n_468) );
INVx1_ASAP7_75t_L g486 ( .A(n_243), .Y(n_486) );
OAI22xp33_ASAP7_75t_L g248 ( .A1(n_249), .A2(n_254), .B1(n_258), .B2(n_262), .Y(n_248) );
OAI22xp33_ASAP7_75t_L g403 ( .A1(n_249), .A2(n_367), .B1(n_404), .B2(n_405), .Y(n_403) );
INVx1_ASAP7_75t_SL g249 ( .A(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_252), .Y(n_250) );
INVx1_ASAP7_75t_L g318 ( .A(n_251), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_252), .B(n_295), .Y(n_294) );
INVx2_ASAP7_75t_L g313 ( .A(n_253), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_253), .B(n_266), .Y(n_340) );
INVx1_ASAP7_75t_L g356 ( .A(n_253), .Y(n_356) );
AND2x2_ASAP7_75t_L g297 ( .A(n_255), .B(n_298), .Y(n_297) );
INVx3_ASAP7_75t_SL g336 ( .A(n_255), .Y(n_336) );
NOR2xp33_ASAP7_75t_L g413 ( .A(n_255), .B(n_261), .Y(n_413) );
AND2x4_ASAP7_75t_L g255 ( .A(n_256), .B(n_257), .Y(n_255) );
INVx1_ASAP7_75t_L g422 ( .A(n_258), .Y(n_422) );
OR2x2_ASAP7_75t_L g258 ( .A(n_259), .B(n_261), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_259), .B(n_355), .Y(n_397) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
INVx3_ASAP7_75t_SL g302 ( .A(n_261), .Y(n_302) );
NAND2x1_ASAP7_75t_SL g262 ( .A(n_263), .B(n_264), .Y(n_262) );
AND2x2_ASAP7_75t_L g323 ( .A(n_263), .B(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g330 ( .A(n_263), .B(n_267), .Y(n_330) );
AND2x2_ASAP7_75t_L g335 ( .A(n_263), .B(n_276), .Y(n_335) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_263), .Y(n_384) );
OAI311xp33_ASAP7_75t_L g407 ( .A1(n_264), .A2(n_408), .A3(n_410), .B1(n_411), .C1(n_421), .Y(n_407) );
INVx2_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
OR2x2_ASAP7_75t_L g420 ( .A(n_265), .B(n_293), .Y(n_420) );
OR2x2_ASAP7_75t_L g265 ( .A(n_266), .B(n_267), .Y(n_265) );
AND2x2_ASAP7_75t_L g276 ( .A(n_266), .B(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g324 ( .A(n_266), .B(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g379 ( .A(n_266), .Y(n_379) );
INVx1_ASAP7_75t_L g272 ( .A(n_267), .Y(n_272) );
INVx1_ASAP7_75t_L g292 ( .A(n_267), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_267), .B(n_313), .Y(n_312) );
INVx2_ASAP7_75t_L g325 ( .A(n_267), .Y(n_325) );
AOI221xp5_ASAP7_75t_SL g268 ( .A1(n_269), .A2(n_271), .B1(n_279), .B2(n_284), .C(n_289), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_270), .B(n_274), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g271 ( .A(n_272), .B(n_273), .Y(n_271) );
INVx4_ASAP7_75t_L g293 ( .A(n_273), .Y(n_293) );
AND2x2_ASAP7_75t_L g387 ( .A(n_273), .B(n_306), .Y(n_387) );
AND2x2_ASAP7_75t_L g394 ( .A(n_273), .B(n_276), .Y(n_394) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g275 ( .A(n_276), .B(n_278), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_276), .B(n_355), .Y(n_354) );
AND2x2_ASAP7_75t_L g305 ( .A(n_278), .B(n_306), .Y(n_305) );
INVx1_ASAP7_75t_SL g279 ( .A(n_280), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_281), .B(n_283), .Y(n_280) );
NOR2xp33_ASAP7_75t_L g353 ( .A(n_281), .B(n_354), .Y(n_353) );
INVx1_ASAP7_75t_SL g281 ( .A(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g430 ( .A(n_283), .B(n_374), .Y(n_430) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
OR2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_288), .Y(n_285) );
INVx1_ASAP7_75t_SL g286 ( .A(n_287), .Y(n_286) );
OR2x2_ASAP7_75t_L g415 ( .A(n_287), .B(n_343), .Y(n_415) );
OAI211xp5_ASAP7_75t_L g380 ( .A1(n_288), .A2(n_381), .B(n_382), .C(n_395), .Y(n_380) );
AOI21xp33_ASAP7_75t_SL g289 ( .A1(n_290), .A2(n_294), .B(n_296), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
NOR2xp67_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
INVx1_ASAP7_75t_L g359 ( .A(n_293), .Y(n_359) );
OAI221xp5_ASAP7_75t_L g388 ( .A1(n_294), .A2(n_389), .B1(n_390), .B2(n_391), .C(n_392), .Y(n_388) );
AND2x2_ASAP7_75t_L g365 ( .A(n_295), .B(n_306), .Y(n_365) );
AND2x2_ASAP7_75t_L g418 ( .A(n_295), .B(n_313), .Y(n_418) );
INVx2_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
NOR2xp33_ASAP7_75t_L g360 ( .A(n_298), .B(n_336), .Y(n_360) );
O2A1O1Ixp33_ASAP7_75t_L g299 ( .A1(n_300), .A2(n_303), .B(n_305), .C(n_307), .Y(n_299) );
AND2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
AND2x2_ASAP7_75t_L g346 ( .A(n_301), .B(n_304), .Y(n_346) );
OR2x2_ASAP7_75t_L g389 ( .A(n_301), .B(n_343), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_302), .B(n_368), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_302), .B(n_374), .Y(n_373) );
INVx1_ASAP7_75t_SL g333 ( .A(n_303), .Y(n_333) );
INVx1_ASAP7_75t_L g399 ( .A(n_306), .Y(n_399) );
OAI22xp5_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_311), .B1(n_314), .B2(n_315), .Y(n_307) );
INVx1_ASAP7_75t_L g322 ( .A(n_308), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_309), .B(n_310), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_309), .B(n_368), .Y(n_367) );
AND2x2_ASAP7_75t_L g385 ( .A(n_310), .B(n_386), .Y(n_385) );
INVxp67_ASAP7_75t_L g371 ( .A(n_312), .Y(n_371) );
NOR2xp33_ASAP7_75t_L g398 ( .A(n_313), .B(n_399), .Y(n_398) );
OAI22xp33_ASAP7_75t_L g372 ( .A1(n_314), .A2(n_373), .B1(n_375), .B2(n_377), .Y(n_372) );
INVx1_ASAP7_75t_L g381 ( .A(n_317), .Y(n_381) );
AND2x2_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
AND2x2_ASAP7_75t_L g423 ( .A(n_318), .B(n_418), .Y(n_423) );
AOI222xp33_ASAP7_75t_L g352 ( .A1(n_319), .A2(n_353), .B1(n_356), .B2(n_357), .C1(n_360), .C2(n_361), .Y(n_352) );
NAND4xp25_ASAP7_75t_SL g320 ( .A(n_321), .B(n_341), .C(n_352), .D(n_364), .Y(n_320) );
AOI221xp5_ASAP7_75t_L g321 ( .A1(n_322), .A2(n_323), .B1(n_326), .B2(n_331), .C(n_332), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_324), .B(n_359), .Y(n_358) );
INVxp67_ASAP7_75t_L g350 ( .A(n_325), .Y(n_350) );
AOI221xp5_ASAP7_75t_L g395 ( .A1(n_326), .A2(n_396), .B1(n_398), .B2(n_400), .C(n_403), .Y(n_395) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
OR2x2_ASAP7_75t_L g327 ( .A(n_328), .B(n_329), .Y(n_327) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g338 ( .A(n_330), .B(n_339), .Y(n_338) );
OAI21xp33_ASAP7_75t_L g392 ( .A1(n_331), .A2(n_393), .B(n_394), .Y(n_392) );
OAI22xp5_ASAP7_75t_L g332 ( .A1(n_333), .A2(n_334), .B1(n_336), .B2(n_337), .Y(n_332) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
OAI21xp5_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_344), .B(n_347), .Y(n_341) );
INVxp67_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
OR2x2_ASAP7_75t_L g348 ( .A(n_349), .B(n_351), .Y(n_348) );
HB1xp67_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g383 ( .A(n_354), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_355), .B(n_374), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_355), .B(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_359), .B(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_SL g391 ( .A(n_363), .Y(n_391) );
AOI221xp5_ASAP7_75t_L g364 ( .A1(n_365), .A2(n_366), .B1(n_369), .B2(n_371), .C(n_372), .Y(n_364) );
INVxp67_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
AOI222xp33_ASAP7_75t_L g411 ( .A1(n_374), .A2(n_412), .B1(n_413), .B2(n_414), .C1(n_416), .C2(n_419), .Y(n_411) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_378), .B(n_418), .Y(n_417) );
INVxp67_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g410 ( .A(n_384), .Y(n_410) );
INVxp67_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVxp33_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
AOI221xp5_ASAP7_75t_L g421 ( .A1(n_422), .A2(n_423), .B1(n_424), .B2(n_425), .C(n_428), .Y(n_421) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVxp67_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx2_ASAP7_75t_L g712 ( .A(n_432), .Y(n_712) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
NOR2x2_ASAP7_75t_L g715 ( .A(n_434), .B(n_716), .Y(n_715) );
INVx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
AND3x1_ASAP7_75t_L g437 ( .A(n_438), .B(n_630), .C(n_678), .Y(n_437) );
NOR4xp25_ASAP7_75t_L g438 ( .A(n_439), .B(n_558), .C(n_603), .D(n_617), .Y(n_438) );
OAI311xp33_ASAP7_75t_L g439 ( .A1(n_440), .A2(n_478), .A3(n_502), .B1(n_511), .C1(n_526), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_441), .B(n_449), .Y(n_440) );
OAI21xp33_ASAP7_75t_L g511 ( .A1(n_441), .A2(n_512), .B(n_514), .Y(n_511) );
AND2x2_ASAP7_75t_L g619 ( .A(n_441), .B(n_546), .Y(n_619) );
AND2x2_ASAP7_75t_L g676 ( .A(n_441), .B(n_562), .Y(n_676) );
BUFx2_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
AND2x2_ASAP7_75t_L g569 ( .A(n_442), .B(n_472), .Y(n_569) );
AND2x2_ASAP7_75t_L g626 ( .A(n_442), .B(n_574), .Y(n_626) );
INVx1_ASAP7_75t_L g667 ( .A(n_442), .Y(n_667) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
BUFx6f_ASAP7_75t_L g535 ( .A(n_443), .Y(n_535) );
AND2x2_ASAP7_75t_L g576 ( .A(n_443), .B(n_472), .Y(n_576) );
AND2x2_ASAP7_75t_L g580 ( .A(n_443), .B(n_473), .Y(n_580) );
INVx1_ASAP7_75t_L g592 ( .A(n_443), .Y(n_592) );
OAI21xp5_ASAP7_75t_L g518 ( .A1(n_448), .A2(n_519), .B(n_522), .Y(n_518) );
AND2x2_ASAP7_75t_L g449 ( .A(n_450), .B(n_460), .Y(n_449) );
AND2x2_ASAP7_75t_L g513 ( .A(n_450), .B(n_472), .Y(n_513) );
INVx2_ASAP7_75t_L g547 ( .A(n_450), .Y(n_547) );
AND2x2_ASAP7_75t_L g562 ( .A(n_450), .B(n_473), .Y(n_562) );
HB1xp67_ASAP7_75t_L g568 ( .A(n_450), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_450), .B(n_574), .Y(n_573) );
OR2x2_ASAP7_75t_L g582 ( .A(n_450), .B(n_545), .Y(n_582) );
INVx1_ASAP7_75t_L g594 ( .A(n_450), .Y(n_594) );
INVx1_ASAP7_75t_L g635 ( .A(n_450), .Y(n_635) );
NOR2xp33_ASAP7_75t_L g688 ( .A(n_450), .B(n_535), .Y(n_688) );
AOI21xp5_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_454), .B(n_455), .Y(n_452) );
NOR2xp67_ASAP7_75t_L g460 ( .A(n_461), .B(n_472), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
AND2x2_ASAP7_75t_L g512 ( .A(n_462), .B(n_513), .Y(n_512) );
HB1xp67_ASAP7_75t_L g540 ( .A(n_462), .Y(n_540) );
AND2x2_ASAP7_75t_SL g593 ( .A(n_462), .B(n_594), .Y(n_593) );
OR2x2_ASAP7_75t_L g597 ( .A(n_462), .B(n_472), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_462), .B(n_592), .Y(n_655) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx2_ASAP7_75t_L g545 ( .A(n_463), .Y(n_545) );
HB1xp67_ASAP7_75t_L g561 ( .A(n_463), .Y(n_561) );
OR2x2_ASAP7_75t_L g634 ( .A(n_463), .B(n_635), .Y(n_634) );
INVx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
BUFx2_ASAP7_75t_L g541 ( .A(n_473), .Y(n_541) );
AND2x2_ASAP7_75t_L g546 ( .A(n_473), .B(n_547), .Y(n_546) );
O2A1O1Ixp33_ASAP7_75t_L g487 ( .A1(n_476), .A2(n_488), .B(n_490), .C(n_491), .Y(n_487) );
AOI21xp5_ASAP7_75t_L g498 ( .A1(n_476), .A2(n_499), .B(n_500), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_478), .B(n_529), .Y(n_692) );
INVx1_ASAP7_75t_SL g478 ( .A(n_479), .Y(n_478) );
OR2x2_ASAP7_75t_L g662 ( .A(n_479), .B(n_504), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_480), .B(n_493), .Y(n_479) );
AND2x2_ASAP7_75t_L g538 ( .A(n_480), .B(n_529), .Y(n_538) );
INVx2_ASAP7_75t_L g550 ( .A(n_480), .Y(n_550) );
AND2x2_ASAP7_75t_L g584 ( .A(n_480), .B(n_532), .Y(n_584) );
AND2x2_ASAP7_75t_L g651 ( .A(n_480), .B(n_652), .Y(n_651) );
INVx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_481), .B(n_517), .Y(n_516) );
AND2x2_ASAP7_75t_L g531 ( .A(n_481), .B(n_532), .Y(n_531) );
AND2x2_ASAP7_75t_L g571 ( .A(n_481), .B(n_493), .Y(n_571) );
AND2x2_ASAP7_75t_L g588 ( .A(n_481), .B(n_589), .Y(n_588) );
INVx2_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
AND2x2_ASAP7_75t_L g514 ( .A(n_493), .B(n_515), .Y(n_514) );
INVx3_ASAP7_75t_L g532 ( .A(n_493), .Y(n_532) );
AND2x2_ASAP7_75t_L g537 ( .A(n_493), .B(n_517), .Y(n_537) );
AND2x2_ASAP7_75t_L g610 ( .A(n_493), .B(n_589), .Y(n_610) );
AND2x2_ASAP7_75t_L g675 ( .A(n_493), .B(n_665), .Y(n_675) );
OAI311xp33_ASAP7_75t_L g558 ( .A1(n_502), .A2(n_559), .A3(n_563), .B1(n_565), .C1(n_585), .Y(n_558) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
AND2x2_ASAP7_75t_L g570 ( .A(n_503), .B(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g629 ( .A(n_503), .B(n_537), .Y(n_629) );
AND2x2_ASAP7_75t_L g703 ( .A(n_503), .B(n_584), .Y(n_703) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
NOR2xp33_ASAP7_75t_L g515 ( .A(n_504), .B(n_516), .Y(n_515) );
INVx1_ASAP7_75t_L g638 ( .A(n_504), .Y(n_638) );
INVx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx3_ASAP7_75t_L g529 ( .A(n_505), .Y(n_529) );
NOR2x1_ASAP7_75t_L g601 ( .A(n_505), .B(n_602), .Y(n_601) );
AND2x2_ASAP7_75t_L g658 ( .A(n_505), .B(n_532), .Y(n_658) );
AND2x4_ASAP7_75t_L g505 ( .A(n_506), .B(n_507), .Y(n_505) );
INVx1_ASAP7_75t_L g555 ( .A(n_506), .Y(n_555) );
AND2x2_ASAP7_75t_L g533 ( .A(n_513), .B(n_534), .Y(n_533) );
AND2x2_ASAP7_75t_L g586 ( .A(n_513), .B(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g666 ( .A(n_513), .B(n_667), .Y(n_666) );
AOI221xp5_ASAP7_75t_L g565 ( .A1(n_514), .A2(n_546), .B1(n_566), .B2(n_570), .C(n_572), .Y(n_565) );
INVx1_ASAP7_75t_L g690 ( .A(n_515), .Y(n_690) );
OR2x2_ASAP7_75t_L g656 ( .A(n_516), .B(n_657), .Y(n_656) );
AND2x2_ASAP7_75t_L g551 ( .A(n_517), .B(n_532), .Y(n_551) );
OR2x2_ASAP7_75t_L g553 ( .A(n_517), .B(n_554), .Y(n_553) );
INVx1_ASAP7_75t_L g578 ( .A(n_517), .Y(n_578) );
INVx2_ASAP7_75t_L g589 ( .A(n_517), .Y(n_589) );
AND2x2_ASAP7_75t_L g616 ( .A(n_517), .B(n_554), .Y(n_616) );
HB1xp67_ASAP7_75t_L g645 ( .A(n_517), .Y(n_645) );
AOI221xp5_ASAP7_75t_L g526 ( .A1(n_527), .A2(n_533), .B1(n_536), .B2(n_539), .C(n_542), .Y(n_526) );
INVx1_ASAP7_75t_SL g527 ( .A(n_528), .Y(n_527) );
OR2x2_ASAP7_75t_L g528 ( .A(n_529), .B(n_530), .Y(n_528) );
AND2x2_ASAP7_75t_L g627 ( .A(n_529), .B(n_537), .Y(n_627) );
AND2x2_ASAP7_75t_L g677 ( .A(n_529), .B(n_531), .Y(n_677) );
INVx2_ASAP7_75t_SL g530 ( .A(n_531), .Y(n_530) );
AND2x2_ASAP7_75t_L g564 ( .A(n_531), .B(n_535), .Y(n_564) );
AND2x2_ASAP7_75t_L g643 ( .A(n_531), .B(n_616), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_532), .B(n_578), .Y(n_577) );
INVx2_ASAP7_75t_L g602 ( .A(n_532), .Y(n_602) );
OAI21xp33_ASAP7_75t_L g612 ( .A1(n_533), .A2(n_613), .B(n_615), .Y(n_612) );
OR2x2_ASAP7_75t_L g556 ( .A(n_534), .B(n_557), .Y(n_556) );
OR2x2_ASAP7_75t_L g622 ( .A(n_534), .B(n_582), .Y(n_622) );
NOR2xp33_ASAP7_75t_L g633 ( .A(n_534), .B(n_634), .Y(n_633) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
AND2x2_ASAP7_75t_L g599 ( .A(n_535), .B(n_568), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_535), .B(n_682), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_536), .B(n_562), .Y(n_672) );
AND2x2_ASAP7_75t_L g536 ( .A(n_537), .B(n_538), .Y(n_536) );
AND2x2_ASAP7_75t_L g595 ( .A(n_537), .B(n_550), .Y(n_595) );
INVx1_ASAP7_75t_L g611 ( .A(n_538), .Y(n_611) );
NOR2xp33_ASAP7_75t_L g539 ( .A(n_540), .B(n_541), .Y(n_539) );
OAI22xp5_ASAP7_75t_L g542 ( .A1(n_543), .A2(n_548), .B1(n_552), .B2(n_556), .Y(n_542) );
INVx2_ASAP7_75t_SL g543 ( .A(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_545), .B(n_546), .Y(n_544) );
INVx2_ASAP7_75t_L g574 ( .A(n_545), .Y(n_574) );
INVx1_ASAP7_75t_L g587 ( .A(n_545), .Y(n_587) );
INVx1_ASAP7_75t_L g557 ( .A(n_546), .Y(n_557) );
AND2x2_ASAP7_75t_L g628 ( .A(n_546), .B(n_574), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_546), .B(n_654), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_549), .B(n_551), .Y(n_548) );
OR2x2_ASAP7_75t_L g552 ( .A(n_549), .B(n_553), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_549), .B(n_665), .Y(n_664) );
NOR2xp67_ASAP7_75t_L g696 ( .A(n_549), .B(n_697), .Y(n_696) );
INVx3_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_L g699 ( .A(n_551), .B(n_651), .Y(n_699) );
INVx1_ASAP7_75t_SL g665 ( .A(n_553), .Y(n_665) );
AND2x2_ASAP7_75t_L g605 ( .A(n_554), .B(n_589), .Y(n_605) );
INVx1_ASAP7_75t_L g652 ( .A(n_554), .Y(n_652) );
OAI222xp33_ASAP7_75t_L g693 ( .A1(n_559), .A2(n_649), .B1(n_694), .B2(n_695), .C1(n_698), .C2(n_700), .Y(n_693) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_561), .B(n_562), .Y(n_560) );
INVx1_ASAP7_75t_L g614 ( .A(n_561), .Y(n_614) );
AND2x2_ASAP7_75t_L g625 ( .A(n_562), .B(n_626), .Y(n_625) );
NAND2xp5_ASAP7_75t_SL g694 ( .A(n_562), .B(n_667), .Y(n_694) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_564), .B(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g669 ( .A(n_566), .Y(n_669) );
AND2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_569), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx1_ASAP7_75t_SL g607 ( .A(n_569), .Y(n_607) );
AND2x2_ASAP7_75t_L g686 ( .A(n_569), .B(n_647), .Y(n_686) );
AND2x2_ASAP7_75t_L g709 ( .A(n_569), .B(n_593), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_571), .B(n_605), .Y(n_604) );
OAI32xp33_ASAP7_75t_L g572 ( .A1(n_573), .A2(n_575), .A3(n_577), .B1(n_579), .B2(n_583), .Y(n_572) );
BUFx2_ASAP7_75t_L g647 ( .A(n_574), .Y(n_647) );
NOR2xp33_ASAP7_75t_L g674 ( .A(n_575), .B(n_593), .Y(n_674) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g613 ( .A(n_576), .B(n_614), .Y(n_613) );
AND2x4_ASAP7_75t_L g681 ( .A(n_576), .B(n_682), .Y(n_681) );
OR2x2_ASAP7_75t_L g670 ( .A(n_577), .B(n_671), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_580), .B(n_581), .Y(n_579) );
AND2x2_ASAP7_75t_L g641 ( .A(n_580), .B(n_614), .Y(n_641) );
INVx2_ASAP7_75t_SL g581 ( .A(n_582), .Y(n_581) );
OAI221xp5_ASAP7_75t_SL g603 ( .A1(n_582), .A2(n_604), .B1(n_606), .B2(n_608), .C(n_612), .Y(n_603) );
INVx2_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g615 ( .A(n_584), .B(n_616), .Y(n_615) );
AND2x2_ASAP7_75t_L g621 ( .A(n_584), .B(n_605), .Y(n_621) );
AOI221xp5_ASAP7_75t_L g585 ( .A1(n_586), .A2(n_588), .B1(n_590), .B2(n_595), .C(n_596), .Y(n_585) );
INVx1_ASAP7_75t_L g704 ( .A(n_586), .Y(n_704) );
NAND2xp5_ASAP7_75t_SL g680 ( .A(n_587), .B(n_681), .Y(n_680) );
NAND2x1p5_ASAP7_75t_L g600 ( .A(n_588), .B(n_601), .Y(n_600) );
AND2x2_ASAP7_75t_L g590 ( .A(n_591), .B(n_593), .Y(n_590) );
HB1xp67_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_593), .B(n_607), .Y(n_606) );
INVx2_ASAP7_75t_L g659 ( .A(n_593), .Y(n_659) );
BUFx3_ASAP7_75t_L g682 ( .A(n_594), .Y(n_682) );
INVx1_ASAP7_75t_SL g623 ( .A(n_595), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_595), .B(n_637), .Y(n_636) );
AOI21xp33_ASAP7_75t_SL g596 ( .A1(n_597), .A2(n_598), .B(n_600), .Y(n_596) );
OAI221xp5_ASAP7_75t_L g701 ( .A1(n_597), .A2(n_698), .B1(n_702), .B2(n_704), .C(n_705), .Y(n_701) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g644 ( .A(n_602), .B(n_605), .Y(n_644) );
INVx1_ASAP7_75t_L g708 ( .A(n_602), .Y(n_708) );
INVx2_ASAP7_75t_L g697 ( .A(n_605), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_605), .B(n_708), .Y(n_707) );
OR2x2_ASAP7_75t_L g608 ( .A(n_609), .B(n_611), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g650 ( .A(n_610), .B(n_651), .Y(n_650) );
OAI221xp5_ASAP7_75t_SL g617 ( .A1(n_618), .A2(n_620), .B1(n_622), .B2(n_623), .C(n_624), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx1_ASAP7_75t_SL g620 ( .A(n_621), .Y(n_620) );
AOI22xp33_ASAP7_75t_L g624 ( .A1(n_625), .A2(n_627), .B1(n_628), .B2(n_629), .Y(n_624) );
AOI22xp5_ASAP7_75t_L g687 ( .A1(n_626), .A2(n_688), .B1(n_689), .B2(n_691), .Y(n_687) );
OAI21xp5_ASAP7_75t_L g705 ( .A1(n_629), .A2(n_706), .B(n_709), .Y(n_705) );
NOR4xp25_ASAP7_75t_SL g630 ( .A(n_631), .B(n_639), .C(n_648), .D(n_668), .Y(n_630) );
NOR2xp33_ASAP7_75t_L g631 ( .A(n_632), .B(n_636), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
OAI22xp5_ASAP7_75t_L g639 ( .A1(n_640), .A2(n_642), .B1(n_645), .B2(n_646), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
NOR2xp33_ASAP7_75t_L g642 ( .A(n_643), .B(n_644), .Y(n_642) );
INVx1_ASAP7_75t_L g684 ( .A(n_644), .Y(n_684) );
OAI221xp5_ASAP7_75t_L g648 ( .A1(n_649), .A2(n_653), .B1(n_656), .B2(n_659), .C(n_660), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g671 ( .A(n_651), .Y(n_671) );
INVx1_ASAP7_75t_SL g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
OAI21xp5_ASAP7_75t_SL g660 ( .A1(n_661), .A2(n_663), .B(n_666), .Y(n_660) );
INVx1_ASAP7_75t_SL g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
OAI211xp5_ASAP7_75t_L g668 ( .A1(n_669), .A2(n_670), .B(n_672), .C(n_673), .Y(n_668) );
AOI22xp5_ASAP7_75t_L g673 ( .A1(n_674), .A2(n_675), .B1(n_676), .B2(n_677), .Y(n_673) );
CKINVDCx14_ASAP7_75t_R g683 ( .A(n_677), .Y(n_683) );
NOR3xp33_ASAP7_75t_L g678 ( .A(n_679), .B(n_693), .C(n_701), .Y(n_678) );
OAI221xp5_ASAP7_75t_L g679 ( .A1(n_680), .A2(n_683), .B1(n_684), .B2(n_685), .C(n_687), .Y(n_679) );
INVxp67_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_SL g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
CKINVDCx16_ASAP7_75t_R g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_SL g713 ( .A(n_714), .Y(n_713) );
INVx3_ASAP7_75t_SL g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
NAND2xp33_ASAP7_75t_L g718 ( .A(n_719), .B(n_723), .Y(n_718) );
NOR2xp33_ASAP7_75t_SL g719 ( .A(n_720), .B(n_722), .Y(n_719) );
INVx1_ASAP7_75t_SL g743 ( .A(n_720), .Y(n_743) );
INVx1_ASAP7_75t_L g742 ( .A(n_722), .Y(n_742) );
OA21x2_ASAP7_75t_L g745 ( .A1(n_722), .A2(n_743), .B(n_746), .Y(n_745) );
INVx1_ASAP7_75t_SL g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_SL g724 ( .A(n_725), .Y(n_724) );
HB1xp67_ASAP7_75t_L g733 ( .A(n_725), .Y(n_733) );
INVx1_ASAP7_75t_SL g736 ( .A(n_725), .Y(n_736) );
BUFx2_ASAP7_75t_L g746 ( .A(n_725), .Y(n_746) );
INVxp67_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
AOI21xp5_ASAP7_75t_L g727 ( .A1(n_728), .A2(n_733), .B(n_734), .Y(n_727) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
NOR2xp33_ASAP7_75t_SL g734 ( .A(n_735), .B(n_737), .Y(n_734) );
INVx1_ASAP7_75t_SL g735 ( .A(n_736), .Y(n_735) );
CKINVDCx20_ASAP7_75t_R g738 ( .A(n_739), .Y(n_738) );
CKINVDCx6p67_ASAP7_75t_R g739 ( .A(n_740), .Y(n_739) );
AND2x2_ASAP7_75t_L g740 ( .A(n_741), .B(n_743), .Y(n_740) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx3_ASAP7_75t_SL g744 ( .A(n_745), .Y(n_744) );
endmodule