module fake_jpeg_3029_n_331 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_331);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_331;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx2_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_39),
.Y(n_91)
);

CKINVDCx5p33_ASAP7_75t_R g40 ( 
.A(n_25),
.Y(n_40)
);

INVx4_ASAP7_75t_SL g94 ( 
.A(n_40),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g76 ( 
.A(n_42),
.Y(n_76)
);

BUFx4f_ASAP7_75t_SL g43 ( 
.A(n_24),
.Y(n_43)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_43),
.Y(n_90)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

INVx2_ASAP7_75t_R g45 ( 
.A(n_36),
.Y(n_45)
);

BUFx2_ASAP7_75t_R g103 ( 
.A(n_45),
.Y(n_103)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_25),
.B(n_14),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_48),
.B(n_50),
.Y(n_84)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_24),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_28),
.B(n_0),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_51),
.B(n_54),
.Y(n_85)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_28),
.B(n_0),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

NAND2xp33_ASAP7_75t_SL g56 ( 
.A(n_36),
.B(n_0),
.Y(n_56)
);

A2O1A1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_56),
.A2(n_31),
.B(n_17),
.C(n_3),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

BUFx16f_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_32),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_60),
.B(n_71),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_54),
.A2(n_32),
.B1(n_37),
.B2(n_20),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_63),
.A2(n_83),
.B1(n_96),
.B2(n_104),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_45),
.A2(n_21),
.B1(n_19),
.B2(n_23),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_64),
.A2(n_66),
.B1(n_72),
.B2(n_97),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_45),
.A2(n_21),
.B1(n_23),
.B2(n_33),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_40),
.B(n_27),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_68),
.B(n_69),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_48),
.B(n_27),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_29),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_44),
.A2(n_20),
.B1(n_37),
.B2(n_33),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_50),
.B(n_39),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_73),
.B(n_80),
.Y(n_109)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_74),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_44),
.A2(n_37),
.B1(n_38),
.B2(n_35),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_75),
.A2(n_82),
.B1(n_106),
.B2(n_1),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_46),
.B(n_29),
.C(n_26),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_79),
.B(n_99),
.C(n_1),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_53),
.B(n_35),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_43),
.B(n_35),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_81),
.B(n_86),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_43),
.A2(n_38),
.B1(n_35),
.B2(n_26),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_52),
.A2(n_36),
.B1(n_38),
.B2(n_34),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_43),
.B(n_26),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_89),
.Y(n_110)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_42),
.Y(n_92)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_92),
.Y(n_118)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_93),
.Y(n_128)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_95),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_L g96 ( 
.A1(n_47),
.A2(n_30),
.B1(n_22),
.B2(n_34),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_49),
.A2(n_23),
.B1(n_26),
.B2(n_30),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_42),
.B(n_22),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_98),
.B(n_101),
.Y(n_140)
);

AOI21xp33_ASAP7_75t_SL g99 ( 
.A1(n_58),
.A2(n_23),
.B(n_17),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_100),
.B(n_2),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_58),
.B(n_15),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_58),
.A2(n_57),
.B1(n_55),
.B2(n_41),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_102),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_41),
.A2(n_57),
.B1(n_55),
.B2(n_31),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_40),
.B(n_15),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_105),
.B(n_12),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_51),
.A2(n_14),
.B1(n_12),
.B2(n_10),
.Y(n_106)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_78),
.Y(n_108)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_108),
.Y(n_164)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_90),
.Y(n_112)
);

BUFx4f_ASAP7_75t_SL g168 ( 
.A(n_112),
.Y(n_168)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_78),
.Y(n_113)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_113),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_114),
.A2(n_63),
.B1(n_82),
.B2(n_104),
.Y(n_159)
);

BUFx5_ASAP7_75t_L g115 ( 
.A(n_93),
.Y(n_115)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_115),
.Y(n_156)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_91),
.Y(n_116)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_116),
.Y(n_172)
);

BUFx5_ASAP7_75t_L g117 ( 
.A(n_76),
.Y(n_117)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_117),
.Y(n_158)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_90),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g153 ( 
.A(n_119),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_120),
.B(n_134),
.Y(n_141)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_91),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_122),
.Y(n_142)
);

AND2x2_ASAP7_75t_SL g149 ( 
.A(n_123),
.B(n_60),
.Y(n_149)
);

OA22x2_ASAP7_75t_L g124 ( 
.A1(n_83),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_124)
);

OA21x2_ASAP7_75t_L g166 ( 
.A1(n_124),
.A2(n_95),
.B(n_59),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_85),
.B(n_1),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_125),
.B(n_106),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_130),
.Y(n_174)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_59),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_131),
.Y(n_154)
);

INVxp67_ASAP7_75t_SL g132 ( 
.A(n_65),
.Y(n_132)
);

INVx13_ASAP7_75t_L g145 ( 
.A(n_132),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_133),
.A2(n_103),
.B1(n_100),
.B2(n_76),
.Y(n_157)
);

OR2x2_ASAP7_75t_L g134 ( 
.A(n_94),
.B(n_10),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_87),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_135),
.Y(n_173)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_87),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_136),
.B(n_139),
.Y(n_147)
);

BUFx12_ASAP7_75t_L g137 ( 
.A(n_65),
.Y(n_137)
);

INVx13_ASAP7_75t_L g177 ( 
.A(n_137),
.Y(n_177)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_88),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_107),
.B(n_94),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_143),
.B(n_151),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_110),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_144),
.B(n_148),
.Y(n_185)
);

OR2x2_ASAP7_75t_L g146 ( 
.A(n_116),
.B(n_71),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_146),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_149),
.B(n_161),
.Y(n_183)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_127),
.Y(n_150)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_150),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_109),
.B(n_84),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_140),
.B(n_79),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_152),
.B(n_160),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_111),
.B(n_77),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_155),
.B(n_144),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_157),
.A2(n_124),
.B(n_135),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_159),
.B(n_166),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_121),
.B(n_96),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_121),
.B(n_88),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_161),
.B(n_163),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_138),
.A2(n_72),
.B1(n_75),
.B2(n_99),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_162),
.A2(n_139),
.B1(n_118),
.B2(n_128),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_125),
.B(n_122),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_123),
.A2(n_62),
.B1(n_67),
.B2(n_70),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_165),
.A2(n_170),
.B1(n_171),
.B2(n_176),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_108),
.B(n_103),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_167),
.B(n_175),
.Y(n_190)
);

OAI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_126),
.A2(n_61),
.B1(n_77),
.B2(n_70),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_133),
.A2(n_67),
.B1(n_62),
.B2(n_61),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_133),
.B(n_10),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_138),
.A2(n_92),
.B1(n_74),
.B2(n_5),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_174),
.A2(n_119),
.B1(n_112),
.B2(n_113),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_178),
.Y(n_230)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_173),
.Y(n_181)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_181),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_SL g182 ( 
.A(n_149),
.B(n_134),
.C(n_120),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_182),
.B(n_189),
.C(n_199),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_183),
.B(n_156),
.Y(n_236)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_172),
.Y(n_186)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_186),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_167),
.B(n_146),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_187),
.A2(n_196),
.B(n_211),
.Y(n_234)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_172),
.Y(n_188)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_188),
.Y(n_238)
);

MAJx2_ASAP7_75t_L g189 ( 
.A(n_149),
.B(n_124),
.C(n_136),
.Y(n_189)
);

BUFx4f_ASAP7_75t_SL g191 ( 
.A(n_177),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_191),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_160),
.A2(n_110),
.B(n_131),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_192),
.A2(n_158),
.B(n_156),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g194 ( 
.A(n_173),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_194),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_163),
.B(n_128),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_197),
.B(n_212),
.Y(n_221)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_147),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_198),
.B(n_204),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_149),
.B(n_124),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_200),
.A2(n_202),
.B1(n_166),
.B2(n_176),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_162),
.A2(n_118),
.B1(n_127),
.B2(n_129),
.Y(n_202)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_147),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_152),
.B(n_115),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_205),
.B(n_209),
.Y(n_228)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_164),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_206),
.B(n_169),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_158),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_207),
.B(n_208),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_146),
.B(n_129),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_164),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_210),
.B(n_173),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_171),
.B(n_2),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_148),
.B(n_4),
.Y(n_212)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_213),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_179),
.A2(n_159),
.B1(n_166),
.B2(n_165),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_214),
.A2(n_216),
.B1(n_201),
.B2(n_192),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_179),
.A2(n_166),
.B1(n_142),
.B2(n_141),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_183),
.B(n_157),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_217),
.B(n_222),
.Y(n_240)
);

OR2x2_ASAP7_75t_L g244 ( 
.A(n_219),
.B(n_239),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_179),
.A2(n_141),
.B1(n_169),
.B2(n_150),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_220),
.A2(n_232),
.B1(n_211),
.B2(n_199),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_195),
.B(n_205),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_193),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_223),
.B(n_190),
.Y(n_245)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_231),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_201),
.A2(n_150),
.B1(n_175),
.B2(n_153),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_195),
.B(n_168),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_233),
.B(n_236),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_203),
.B(n_168),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_235),
.B(n_231),
.Y(n_247)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_237),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_184),
.A2(n_153),
.B(n_154),
.Y(n_239)
);

AO22x1_ASAP7_75t_L g242 ( 
.A1(n_220),
.A2(n_187),
.B1(n_202),
.B2(n_200),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_242),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_245),
.B(n_246),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_221),
.B(n_203),
.Y(n_246)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_247),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g248 ( 
.A(n_235),
.Y(n_248)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_248),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_225),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_250),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_215),
.B(n_185),
.Y(n_251)
);

INVxp33_ASAP7_75t_SL g268 ( 
.A(n_251),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_229),
.B(n_206),
.Y(n_252)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_252),
.Y(n_272)
);

OR2x2_ASAP7_75t_L g253 ( 
.A(n_216),
.B(n_187),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_253),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_254),
.A2(n_214),
.B1(n_213),
.B2(n_228),
.Y(n_276)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_229),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_256),
.A2(n_258),
.B1(n_259),
.B2(n_260),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_222),
.B(n_209),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_257),
.B(n_217),
.C(n_236),
.Y(n_270)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_238),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_233),
.B(n_189),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_238),
.B(n_180),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_261),
.A2(n_226),
.B1(n_218),
.B2(n_180),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_SL g262 ( 
.A(n_254),
.B(n_227),
.C(n_232),
.Y(n_262)
);

FAx1_ASAP7_75t_SL g283 ( 
.A(n_262),
.B(n_182),
.CI(n_243),
.CON(n_283),
.SN(n_283)
);

AOI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_241),
.A2(n_242),
.B1(n_230),
.B2(n_249),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_267),
.A2(n_276),
.B1(n_277),
.B2(n_196),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_240),
.B(n_227),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_269),
.B(n_270),
.C(n_257),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_274),
.A2(n_264),
.B1(n_266),
.B2(n_249),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_241),
.A2(n_219),
.B1(n_230),
.B2(n_234),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_240),
.B(n_228),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_278),
.B(n_218),
.C(n_207),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_273),
.B(n_250),
.Y(n_279)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_279),
.Y(n_294)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_280),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_268),
.B(n_255),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_281),
.B(n_285),
.Y(n_302)
);

OAI321xp33_ASAP7_75t_L g282 ( 
.A1(n_265),
.A2(n_253),
.A3(n_247),
.B1(n_259),
.B2(n_244),
.C(n_255),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_282),
.B(n_283),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_284),
.B(n_293),
.Y(n_298)
);

NAND3xp33_ASAP7_75t_L g285 ( 
.A(n_263),
.B(n_253),
.C(n_239),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_272),
.B(n_226),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_286),
.B(n_290),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_278),
.B(n_243),
.C(n_260),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_287),
.B(n_288),
.C(n_289),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_269),
.B(n_234),
.C(n_244),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_270),
.B(n_244),
.C(n_258),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_271),
.B(n_256),
.Y(n_290)
);

A2O1A1Ixp33_ASAP7_75t_SL g291 ( 
.A1(n_264),
.A2(n_242),
.B(n_211),
.C(n_224),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_291),
.A2(n_267),
.B(n_191),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_292),
.A2(n_277),
.B1(n_265),
.B2(n_262),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_289),
.A2(n_275),
.B(n_276),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_295),
.A2(n_291),
.B(n_154),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_299),
.Y(n_312)
);

XNOR2x1_ASAP7_75t_L g310 ( 
.A(n_300),
.B(n_168),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_291),
.A2(n_288),
.B(n_283),
.Y(n_304)
);

MAJx2_ASAP7_75t_L g307 ( 
.A(n_304),
.B(n_305),
.C(n_287),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_284),
.B(n_181),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_298),
.B(n_293),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_306),
.B(n_307),
.Y(n_315)
);

OAI21x1_ASAP7_75t_L g318 ( 
.A1(n_308),
.A2(n_300),
.B(n_294),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_303),
.A2(n_291),
.B(n_191),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_309),
.A2(n_299),
.B(n_296),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_310),
.B(n_314),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_298),
.B(n_177),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_311),
.B(n_313),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_302),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_296),
.B(n_168),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_312),
.A2(n_295),
.B(n_304),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_317),
.A2(n_310),
.B(n_301),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_318),
.B(n_319),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_312),
.B(n_297),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_321),
.B(n_320),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_323),
.A2(n_324),
.B(n_145),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_315),
.B(n_301),
.Y(n_324)
);

AOI322xp5_ASAP7_75t_L g326 ( 
.A1(n_325),
.A2(n_316),
.A3(n_305),
.B1(n_307),
.B2(n_177),
.C1(n_145),
.C2(n_137),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_326),
.B(n_327),
.C(n_322),
.Y(n_328)
);

OAI321xp33_ASAP7_75t_L g329 ( 
.A1(n_328),
.A2(n_145),
.A3(n_137),
.B1(n_117),
.B2(n_7),
.C(n_4),
.Y(n_329)
);

OAI311xp33_ASAP7_75t_L g330 ( 
.A1(n_329),
.A2(n_137),
.A3(n_5),
.B1(n_6),
.C1(n_8),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_4),
.Y(n_331)
);


endmodule