module fake_netlist_6_511_n_73 (n_7, n_6, n_12, n_4, n_2, n_15, n_16, n_3, n_5, n_1, n_14, n_13, n_0, n_9, n_11, n_8, n_17, n_10, n_73);

input n_7;
input n_6;
input n_12;
input n_4;
input n_2;
input n_15;
input n_16;
input n_3;
input n_5;
input n_1;
input n_14;
input n_13;
input n_0;
input n_9;
input n_11;
input n_8;
input n_17;
input n_10;

output n_73;

wire n_41;
wire n_52;
wire n_45;
wire n_46;
wire n_34;
wire n_42;
wire n_70;
wire n_21;
wire n_24;
wire n_18;
wire n_71;
wire n_37;
wire n_33;
wire n_54;
wire n_67;
wire n_27;
wire n_38;
wire n_72;
wire n_61;
wire n_39;
wire n_63;
wire n_60;
wire n_59;
wire n_32;
wire n_66;
wire n_36;
wire n_22;
wire n_26;
wire n_68;
wire n_55;
wire n_35;
wire n_28;
wire n_23;
wire n_58;
wire n_69;
wire n_20;
wire n_50;
wire n_49;
wire n_30;
wire n_64;
wire n_43;
wire n_19;
wire n_48;
wire n_62;
wire n_29;
wire n_47;
wire n_31;
wire n_65;
wire n_40;
wire n_25;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_17),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_L g19 ( 
.A1(n_1),
.A2(n_8),
.B1(n_4),
.B2(n_6),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_16),
.B(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_6),
.A2(n_2),
.B1(n_3),
.B2(n_14),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

AND2x6_ASAP7_75t_L g29 ( 
.A(n_7),
.B(n_5),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_10),
.B(n_5),
.Y(n_30)
);

AND2x4_ASAP7_75t_L g31 ( 
.A(n_0),
.B(n_12),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

CKINVDCx5p33_ASAP7_75t_R g33 ( 
.A(n_21),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_29),
.A2(n_0),
.B1(n_2),
.B2(n_31),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_36),
.B(n_31),
.Y(n_37)
);

NOR2xp67_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_20),
.Y(n_38)
);

A2O1A1Ixp33_ASAP7_75t_L g39 ( 
.A1(n_35),
.A2(n_30),
.B(n_23),
.C(n_26),
.Y(n_39)
);

CKINVDCx8_ASAP7_75t_R g40 ( 
.A(n_33),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_27),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_32),
.A2(n_28),
.B(n_22),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_37),
.A2(n_39),
.B1(n_40),
.B2(n_30),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_35),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_39),
.A2(n_19),
.B1(n_29),
.B2(n_23),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_25),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g53 ( 
.A(n_44),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_20),
.Y(n_54)
);

NAND4xp25_ASAP7_75t_L g55 ( 
.A(n_50),
.B(n_49),
.C(n_19),
.D(n_43),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g56 ( 
.A(n_50),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

NOR2xp67_ASAP7_75t_L g58 ( 
.A(n_53),
.B(n_45),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_57),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_56),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_57),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_60),
.B(n_53),
.Y(n_62)
);

NOR3x1_ASAP7_75t_L g63 ( 
.A(n_61),
.B(n_55),
.C(n_53),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g64 ( 
.A1(n_59),
.A2(n_54),
.B(n_52),
.Y(n_64)
);

OAI221xp5_ASAP7_75t_L g65 ( 
.A1(n_62),
.A2(n_58),
.B1(n_54),
.B2(n_51),
.C(n_52),
.Y(n_65)
);

AOI221x1_ASAP7_75t_L g66 ( 
.A1(n_64),
.A2(n_59),
.B1(n_48),
.B2(n_18),
.C(n_47),
.Y(n_66)
);

OAI221xp5_ASAP7_75t_L g67 ( 
.A1(n_65),
.A2(n_63),
.B1(n_48),
.B2(n_47),
.C(n_18),
.Y(n_67)
);

NOR3xp33_ASAP7_75t_L g68 ( 
.A(n_66),
.B(n_48),
.C(n_47),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_67),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_68),
.Y(n_70)
);

AOI22x1_ASAP7_75t_L g71 ( 
.A1(n_69),
.A2(n_18),
.B1(n_45),
.B2(n_29),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_71),
.A2(n_70),
.B(n_29),
.Y(n_72)
);

OR2x6_ASAP7_75t_L g73 ( 
.A(n_72),
.B(n_48),
.Y(n_73)
);


endmodule