module fake_netlist_5_58_n_1415 (n_137, n_294, n_318, n_82, n_194, n_316, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_61, n_127, n_75, n_235, n_226, n_74, n_57, n_351, n_111, n_155, n_43, n_116, n_22, n_284, n_46, n_245, n_21, n_139, n_38, n_105, n_280, n_4, n_17, n_254, n_33, n_23, n_302, n_265, n_293, n_244, n_47, n_173, n_198, n_247, n_314, n_8, n_321, n_292, n_100, n_212, n_119, n_275, n_252, n_26, n_295, n_133, n_330, n_2, n_6, n_39, n_147, n_67, n_307, n_87, n_150, n_106, n_209, n_259, n_301, n_68, n_93, n_186, n_134, n_191, n_51, n_63, n_171, n_153, n_341, n_204, n_250, n_260, n_298, n_320, n_286, n_122, n_282, n_331, n_10, n_24, n_325, n_132, n_90, n_101, n_281, n_240, n_189, n_220, n_291, n_231, n_257, n_31, n_13, n_152, n_317, n_9, n_323, n_195, n_42, n_227, n_45, n_271, n_94, n_335, n_123, n_167, n_234, n_343, n_308, n_267, n_297, n_156, n_5, n_225, n_219, n_157, n_131, n_192, n_223, n_158, n_138, n_264, n_109, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_347, n_169, n_59, n_255, n_215, n_350, n_196, n_211, n_218, n_181, n_3, n_290, n_221, n_178, n_287, n_344, n_72, n_104, n_41, n_56, n_141, n_15, n_336, n_145, n_48, n_50, n_337, n_313, n_88, n_216, n_168, n_164, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_296, n_241, n_184, n_65, n_78, n_144, n_114, n_96, n_165, n_213, n_129, n_342, n_98, n_197, n_107, n_69, n_236, n_1, n_249, n_304, n_329, n_203, n_274, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_333, n_309, n_30, n_14, n_84, n_130, n_322, n_258, n_29, n_79, n_151, n_25, n_306, n_288, n_188, n_190, n_201, n_263, n_44, n_224, n_40, n_34, n_228, n_283, n_112, n_85, n_239, n_55, n_49, n_310, n_54, n_12, n_76, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_312, n_345, n_210, n_91, n_176, n_182, n_143, n_83, n_237, n_180, n_340, n_207, n_37, n_346, n_229, n_108, n_66, n_177, n_60, n_16, n_0, n_58, n_18, n_117, n_326, n_233, n_205, n_113, n_246, n_179, n_125, n_269, n_128, n_285, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_193, n_251, n_352, n_53, n_160, n_154, n_62, n_148, n_71, n_300, n_159, n_334, n_175, n_262, n_238, n_99, n_319, n_20, n_121, n_242, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_115, n_324, n_199, n_187, n_32, n_103, n_348, n_97, n_166, n_11, n_7, n_256, n_305, n_52, n_278, n_110, n_1415);

input n_137;
input n_294;
input n_318;
input n_82;
input n_194;
input n_316;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_61;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_57;
input n_351;
input n_111;
input n_155;
input n_43;
input n_116;
input n_22;
input n_284;
input n_46;
input n_245;
input n_21;
input n_139;
input n_38;
input n_105;
input n_280;
input n_4;
input n_17;
input n_254;
input n_33;
input n_23;
input n_302;
input n_265;
input n_293;
input n_244;
input n_47;
input n_173;
input n_198;
input n_247;
input n_314;
input n_8;
input n_321;
input n_292;
input n_100;
input n_212;
input n_119;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_2;
input n_6;
input n_39;
input n_147;
input n_67;
input n_307;
input n_87;
input n_150;
input n_106;
input n_209;
input n_259;
input n_301;
input n_68;
input n_93;
input n_186;
input n_134;
input n_191;
input n_51;
input n_63;
input n_171;
input n_153;
input n_341;
input n_204;
input n_250;
input n_260;
input n_298;
input n_320;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_325;
input n_132;
input n_90;
input n_101;
input n_281;
input n_240;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_31;
input n_13;
input n_152;
input n_317;
input n_9;
input n_323;
input n_195;
input n_42;
input n_227;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_167;
input n_234;
input n_343;
input n_308;
input n_267;
input n_297;
input n_156;
input n_5;
input n_225;
input n_219;
input n_157;
input n_131;
input n_192;
input n_223;
input n_158;
input n_138;
input n_264;
input n_109;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_347;
input n_169;
input n_59;
input n_255;
input n_215;
input n_350;
input n_196;
input n_211;
input n_218;
input n_181;
input n_3;
input n_290;
input n_221;
input n_178;
input n_287;
input n_344;
input n_72;
input n_104;
input n_41;
input n_56;
input n_141;
input n_15;
input n_336;
input n_145;
input n_48;
input n_50;
input n_337;
input n_313;
input n_88;
input n_216;
input n_168;
input n_164;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_296;
input n_241;
input n_184;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_213;
input n_129;
input n_342;
input n_98;
input n_197;
input n_107;
input n_69;
input n_236;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_333;
input n_309;
input n_30;
input n_14;
input n_84;
input n_130;
input n_322;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_112;
input n_85;
input n_239;
input n_55;
input n_49;
input n_310;
input n_54;
input n_12;
input n_76;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_312;
input n_345;
input n_210;
input n_91;
input n_176;
input n_182;
input n_143;
input n_83;
input n_237;
input n_180;
input n_340;
input n_207;
input n_37;
input n_346;
input n_229;
input n_108;
input n_66;
input n_177;
input n_60;
input n_16;
input n_0;
input n_58;
input n_18;
input n_117;
input n_326;
input n_233;
input n_205;
input n_113;
input n_246;
input n_179;
input n_125;
input n_269;
input n_128;
input n_285;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_159;
input n_334;
input n_175;
input n_262;
input n_238;
input n_99;
input n_319;
input n_20;
input n_121;
input n_242;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_115;
input n_324;
input n_199;
input n_187;
input n_32;
input n_103;
input n_348;
input n_97;
input n_166;
input n_11;
input n_7;
input n_256;
input n_305;
input n_52;
input n_278;
input n_110;

output n_1415;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1166;
wire n_469;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_667;
wire n_790;
wire n_1055;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_688;
wire n_1353;
wire n_800;
wire n_1347;
wire n_671;
wire n_819;
wire n_1022;
wire n_915;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_625;
wire n_854;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_606;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_1285;
wire n_373;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_929;
wire n_1124;
wire n_902;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_731;
wire n_371;
wire n_1314;
wire n_709;
wire n_1236;
wire n_569;
wire n_920;
wire n_1289;
wire n_370;
wire n_976;
wire n_1078;
wire n_775;
wire n_600;
wire n_1374;
wire n_1328;
wire n_955;
wire n_1146;
wire n_882;
wire n_1036;
wire n_1097;
wire n_696;
wire n_550;
wire n_897;
wire n_798;
wire n_646;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_395;
wire n_901;
wire n_553;
wire n_813;
wire n_1284;
wire n_675;
wire n_888;
wire n_1167;
wire n_637;
wire n_1384;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_464;
wire n_363;
wire n_1069;
wire n_1075;
wire n_1322;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_461;
wire n_1211;
wire n_1197;
wire n_907;
wire n_1377;
wire n_989;
wire n_1039;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_838;
wire n_1053;
wire n_1224;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_534;
wire n_884;
wire n_944;
wire n_647;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_1162;
wire n_1199;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_887;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_434;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_759;
wire n_806;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_649;
wire n_547;
wire n_1191;
wire n_1128;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1233;
wire n_526;
wire n_372;
wire n_677;
wire n_1333;
wire n_1121;
wire n_368;
wire n_604;
wire n_433;
wire n_949;
wire n_1008;
wire n_946;
wire n_1001;
wire n_498;
wire n_689;
wire n_738;
wire n_640;
wire n_624;
wire n_1380;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_758;
wire n_999;
wire n_1158;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1306;
wire n_1068;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_592;
wire n_1169;
wire n_1017;
wire n_978;
wire n_1054;
wire n_1269;
wire n_1095;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_484;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_374;
wire n_396;
wire n_1383;
wire n_1073;
wire n_662;
wire n_459;
wire n_962;
wire n_1215;
wire n_1171;
wire n_723;
wire n_1065;
wire n_1336;
wire n_473;
wire n_1309;
wire n_1043;
wire n_355;
wire n_486;
wire n_614;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_743;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1006;
wire n_1270;
wire n_582;
wire n_1332;
wire n_1390;
wire n_512;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_1031;
wire n_609;
wire n_1041;
wire n_1265;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1304;
wire n_1324;
wire n_987;
wire n_767;
wire n_993;
wire n_1407;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_1209;
wire n_495;
wire n_602;
wire n_574;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_572;
wire n_366;
wire n_815;
wire n_1381;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1082;
wire n_589;
wire n_716;
wire n_562;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_960;
wire n_1290;
wire n_1123;
wire n_1047;
wire n_634;
wire n_1252;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_950;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_389;
wire n_418;
wire n_912;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_376;
wire n_967;
wire n_1139;
wire n_515;
wire n_885;
wire n_397;
wire n_1357;
wire n_483;
wire n_683;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_983;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_690;
wire n_583;
wire n_1343;
wire n_1203;
wire n_821;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_385;
wire n_507;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1329;
wire n_1312;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_943;
wire n_992;
wire n_543;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_883;
wire n_470;
wire n_449;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_1147;
wire n_1077;
wire n_540;
wire n_618;
wire n_896;
wire n_356;
wire n_894;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1096;
wire n_833;
wire n_1307;
wire n_988;
wire n_814;
wire n_1201;
wire n_1114;
wire n_655;
wire n_669;
wire n_472;
wire n_1176;
wire n_387;
wire n_1149;
wire n_398;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_1219;
wire n_1204;
wire n_1035;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_584;
wire n_681;
wire n_430;
wire n_510;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_875;
wire n_357;
wire n_1110;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_1338;
wire n_577;
wire n_693;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_778;
wire n_1122;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1187;
wire n_1392;
wire n_1164;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_876;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_1116;
wire n_1212;
wire n_726;
wire n_982;
wire n_818;
wire n_861;
wire n_1183;
wire n_899;
wire n_1253;
wire n_774;
wire n_1335;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_393;
wire n_487;
wire n_665;
wire n_421;
wire n_1356;
wire n_910;
wire n_768;
wire n_1302;
wire n_1136;
wire n_1313;
wire n_754;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_1109;
wire n_895;
wire n_1310;
wire n_427;
wire n_1399;
wire n_791;
wire n_732;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_766;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1352;
wire n_626;
wire n_1144;
wire n_1137;
wire n_1170;
wire n_676;
wire n_653;
wire n_642;
wire n_855;
wire n_1178;
wire n_850;
wire n_684;
wire n_664;
wire n_503;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_467;
wire n_1227;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_725;
wire n_1388;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_898;
wire n_1013;
wire n_718;
wire n_1120;
wire n_719;
wire n_443;
wire n_714;
wire n_909;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_733;
wire n_1376;
wire n_941;
wire n_981;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_518;
wire n_505;
wire n_752;
wire n_905;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_760;
wire n_381;
wire n_390;
wire n_1330;
wire n_481;
wire n_769;
wire n_1046;
wire n_934;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1361;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_1225;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1411;
wire n_622;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1247;
wire n_922;
wire n_816;
wire n_591;
wire n_1344;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_772;
wire n_499;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_740;
wire n_384;
wire n_1404;
wire n_1315;
wire n_1061;
wire n_1298;
wire n_462;
wire n_1193;
wire n_1255;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_471;
wire n_852;
wire n_1028;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_632;
wire n_699;
wire n_979;
wire n_1245;
wire n_846;
wire n_465;
wire n_362;
wire n_1321;
wire n_585;
wire n_616;
wire n_745;
wire n_1103;
wire n_648;
wire n_1379;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1220;
wire n_437;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_863;
wire n_805;
wire n_1275;
wire n_712;
wire n_1042;
wire n_1402;
wire n_412;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_566;
wire n_565;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1196;
wire n_651;
wire n_1340;
wire n_811;
wire n_807;
wire n_835;
wire n_666;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1251;

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_205),
.Y(n_353)
);

CKINVDCx16_ASAP7_75t_R g354 ( 
.A(n_56),
.Y(n_354)
);

INVx1_ASAP7_75t_SL g355 ( 
.A(n_231),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_124),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_352),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_137),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_49),
.Y(n_359)
);

INVx1_ASAP7_75t_SL g360 ( 
.A(n_202),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_79),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_134),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_149),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_42),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_155),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_327),
.Y(n_366)
);

HB1xp67_ASAP7_75t_L g367 ( 
.A(n_257),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_8),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_316),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_339),
.Y(n_370)
);

BUFx2_ASAP7_75t_SL g371 ( 
.A(n_210),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_76),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_342),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_35),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_263),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_92),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_307),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_203),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_338),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_314),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_261),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_187),
.Y(n_382)
);

INVx1_ASAP7_75t_SL g383 ( 
.A(n_174),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_168),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_196),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_115),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_65),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_68),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_209),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_304),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_3),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_200),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_157),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_260),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_350),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_71),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_349),
.Y(n_397)
);

INVx2_ASAP7_75t_SL g398 ( 
.A(n_332),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_252),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_35),
.Y(n_400)
);

BUFx2_ASAP7_75t_L g401 ( 
.A(n_222),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_132),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_170),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_54),
.Y(n_404)
);

CKINVDCx16_ASAP7_75t_R g405 ( 
.A(n_111),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_78),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_61),
.Y(n_407)
);

INVx1_ASAP7_75t_SL g408 ( 
.A(n_337),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_185),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_240),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_347),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_234),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_144),
.Y(n_413)
);

BUFx3_ASAP7_75t_L g414 ( 
.A(n_286),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_129),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_47),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_152),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_55),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_293),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_335),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_148),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_3),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_73),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_25),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_151),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_172),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_249),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_181),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_241),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_213),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_340),
.Y(n_431)
);

BUFx10_ASAP7_75t_L g432 ( 
.A(n_1),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_343),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_77),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_336),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_269),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_147),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_195),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_135),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_84),
.Y(n_440)
);

BUFx8_ASAP7_75t_SL g441 ( 
.A(n_331),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_284),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_289),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_321),
.Y(n_444)
);

INVx2_ASAP7_75t_SL g445 ( 
.A(n_82),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_180),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_160),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_186),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_232),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_258),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_216),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_219),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_298),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_292),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_16),
.Y(n_455)
);

BUFx2_ASAP7_75t_L g456 ( 
.A(n_320),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_117),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_43),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_50),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_72),
.Y(n_460)
);

INVx1_ASAP7_75t_SL g461 ( 
.A(n_60),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_344),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_58),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_334),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_11),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_282),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_341),
.Y(n_467)
);

BUFx2_ASAP7_75t_L g468 ( 
.A(n_17),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_207),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_14),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_175),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_291),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_52),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_333),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_167),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_218),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_211),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_318),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_44),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_109),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_7),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_204),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_235),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_212),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_215),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_281),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_217),
.Y(n_487)
);

BUFx3_ASAP7_75t_L g488 ( 
.A(n_279),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_50),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_165),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_297),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_221),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_262),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_52),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_346),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_206),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_345),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_237),
.Y(n_498)
);

BUFx6f_ASAP7_75t_L g499 ( 
.A(n_322),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_81),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_87),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_278),
.Y(n_502)
);

CKINVDCx16_ASAP7_75t_R g503 ( 
.A(n_190),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_351),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_19),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_315),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_296),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_191),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_53),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_164),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_171),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_176),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_308),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_254),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_326),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_146),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_184),
.Y(n_517)
);

CKINVDCx16_ASAP7_75t_R g518 ( 
.A(n_265),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_201),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_158),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_301),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_189),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_95),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_123),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_131),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_245),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_182),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_30),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_163),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_348),
.Y(n_530)
);

INVx2_ASAP7_75t_SL g531 ( 
.A(n_270),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_114),
.Y(n_532)
);

CKINVDCx16_ASAP7_75t_R g533 ( 
.A(n_251),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_121),
.Y(n_534)
);

INVx1_ASAP7_75t_SL g535 ( 
.A(n_27),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_283),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_69),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_310),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_47),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_16),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_274),
.Y(n_541)
);

INVx1_ASAP7_75t_SL g542 ( 
.A(n_119),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_330),
.Y(n_543)
);

CKINVDCx20_ASAP7_75t_R g544 ( 
.A(n_106),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_259),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_2),
.Y(n_546)
);

BUFx10_ASAP7_75t_L g547 ( 
.A(n_104),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_8),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_177),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_239),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_223),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_306),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_63),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_162),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_374),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_468),
.B(n_0),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_391),
.Y(n_557)
);

CKINVDCx20_ASAP7_75t_R g558 ( 
.A(n_478),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_400),
.Y(n_559)
);

INVxp67_ASAP7_75t_SL g560 ( 
.A(n_367),
.Y(n_560)
);

CKINVDCx20_ASAP7_75t_R g561 ( 
.A(n_386),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_422),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_353),
.Y(n_563)
);

INVxp67_ASAP7_75t_SL g564 ( 
.A(n_401),
.Y(n_564)
);

INVxp67_ASAP7_75t_SL g565 ( 
.A(n_456),
.Y(n_565)
);

CKINVDCx20_ASAP7_75t_R g566 ( 
.A(n_386),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_356),
.Y(n_567)
);

NOR2xp67_ASAP7_75t_L g568 ( 
.A(n_455),
.B(n_0),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_458),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_470),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_489),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_361),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_362),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_505),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g575 ( 
.A(n_395),
.Y(n_575)
);

INVxp67_ASAP7_75t_L g576 ( 
.A(n_432),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_366),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_398),
.B(n_1),
.Y(n_578)
);

CKINVDCx20_ASAP7_75t_R g579 ( 
.A(n_395),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_355),
.B(n_2),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_369),
.Y(n_581)
);

CKINVDCx20_ASAP7_75t_R g582 ( 
.A(n_469),
.Y(n_582)
);

CKINVDCx16_ASAP7_75t_R g583 ( 
.A(n_354),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_372),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_528),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_546),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_375),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_414),
.Y(n_588)
);

CKINVDCx20_ASAP7_75t_R g589 ( 
.A(n_469),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_414),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_376),
.Y(n_591)
);

INVxp67_ASAP7_75t_SL g592 ( 
.A(n_488),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_445),
.B(n_4),
.Y(n_593)
);

INVxp33_ASAP7_75t_L g594 ( 
.A(n_455),
.Y(n_594)
);

BUFx2_ASAP7_75t_SL g595 ( 
.A(n_544),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_488),
.Y(n_596)
);

NOR2xp67_ASAP7_75t_L g597 ( 
.A(n_378),
.B(n_4),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_377),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_358),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_379),
.Y(n_600)
);

CKINVDCx20_ASAP7_75t_R g601 ( 
.A(n_544),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_363),
.Y(n_602)
);

CKINVDCx16_ASAP7_75t_R g603 ( 
.A(n_405),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_365),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_380),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_370),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_382),
.Y(n_607)
);

CKINVDCx20_ASAP7_75t_R g608 ( 
.A(n_441),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_388),
.Y(n_609)
);

CKINVDCx20_ASAP7_75t_R g610 ( 
.A(n_441),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_531),
.B(n_5),
.Y(n_611)
);

CKINVDCx20_ASAP7_75t_R g612 ( 
.A(n_503),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_378),
.B(n_392),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_R g614 ( 
.A(n_518),
.B(n_5),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_373),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_389),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_381),
.Y(n_617)
);

CKINVDCx20_ASAP7_75t_R g618 ( 
.A(n_533),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_385),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_387),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_397),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_390),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_360),
.B(n_6),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_383),
.B(n_6),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_415),
.Y(n_625)
);

INVxp33_ASAP7_75t_SL g626 ( 
.A(n_359),
.Y(n_626)
);

BUFx2_ASAP7_75t_SL g627 ( 
.A(n_547),
.Y(n_627)
);

INVx3_ASAP7_75t_L g628 ( 
.A(n_432),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_429),
.Y(n_629)
);

INVxp67_ASAP7_75t_L g630 ( 
.A(n_432),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_393),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_430),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_434),
.Y(n_633)
);

NOR2xp67_ASAP7_75t_L g634 ( 
.A(n_392),
.B(n_7),
.Y(n_634)
);

BUFx6f_ASAP7_75t_L g635 ( 
.A(n_357),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_394),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_435),
.Y(n_637)
);

INVxp33_ASAP7_75t_SL g638 ( 
.A(n_364),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_444),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_396),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_450),
.Y(n_641)
);

INVxp67_ASAP7_75t_L g642 ( 
.A(n_535),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_452),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_399),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_453),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_454),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_457),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_466),
.Y(n_648)
);

CKINVDCx20_ASAP7_75t_R g649 ( 
.A(n_368),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_402),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_476),
.Y(n_651)
);

INVx2_ASAP7_75t_SL g652 ( 
.A(n_547),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_403),
.Y(n_653)
);

NOR2xp67_ASAP7_75t_L g654 ( 
.A(n_406),
.B(n_9),
.Y(n_654)
);

INVxp67_ASAP7_75t_SL g655 ( 
.A(n_477),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_599),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_563),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_602),
.Y(n_658)
);

AOI22xp5_ASAP7_75t_L g659 ( 
.A1(n_583),
.A2(n_416),
.B1(n_459),
.B2(n_424),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_635),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_604),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_655),
.B(n_404),
.Y(n_662)
);

CKINVDCx20_ASAP7_75t_R g663 ( 
.A(n_558),
.Y(n_663)
);

HB1xp67_ASAP7_75t_L g664 ( 
.A(n_642),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_606),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_615),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_635),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_617),
.B(n_407),
.Y(n_668)
);

INVx3_ASAP7_75t_L g669 ( 
.A(n_635),
.Y(n_669)
);

CKINVDCx20_ASAP7_75t_R g670 ( 
.A(n_566),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_567),
.Y(n_671)
);

NOR2x1_ASAP7_75t_L g672 ( 
.A(n_597),
.B(n_371),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_564),
.B(n_547),
.Y(n_673)
);

AND2x4_ASAP7_75t_L g674 ( 
.A(n_628),
.B(n_406),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_619),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_620),
.Y(n_676)
);

OA21x2_ASAP7_75t_L g677 ( 
.A1(n_613),
.A2(n_419),
.B(n_411),
.Y(n_677)
);

INVxp67_ASAP7_75t_L g678 ( 
.A(n_627),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_572),
.Y(n_679)
);

BUFx6f_ASAP7_75t_L g680 ( 
.A(n_635),
.Y(n_680)
);

INVx3_ASAP7_75t_L g681 ( 
.A(n_555),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_557),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_573),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_621),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_625),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_577),
.Y(n_686)
);

NAND2xp33_ASAP7_75t_R g687 ( 
.A(n_628),
.B(n_626),
.Y(n_687)
);

BUFx6f_ASAP7_75t_L g688 ( 
.A(n_559),
.Y(n_688)
);

INVxp67_ASAP7_75t_L g689 ( 
.A(n_592),
.Y(n_689)
);

INVx3_ASAP7_75t_L g690 ( 
.A(n_562),
.Y(n_690)
);

OA21x2_ASAP7_75t_L g691 ( 
.A1(n_578),
.A2(n_419),
.B(n_411),
.Y(n_691)
);

HB1xp67_ASAP7_75t_L g692 ( 
.A(n_576),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_629),
.Y(n_693)
);

INVx3_ASAP7_75t_L g694 ( 
.A(n_569),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_614),
.B(n_465),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_570),
.Y(n_696)
);

CKINVDCx20_ASAP7_75t_R g697 ( 
.A(n_575),
.Y(n_697)
);

BUFx6f_ASAP7_75t_L g698 ( 
.A(n_571),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_632),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_633),
.B(n_409),
.Y(n_700)
);

BUFx2_ASAP7_75t_L g701 ( 
.A(n_649),
.Y(n_701)
);

BUFx6f_ASAP7_75t_L g702 ( 
.A(n_574),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_637),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_565),
.B(n_408),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_639),
.Y(n_705)
);

OA21x2_ASAP7_75t_L g706 ( 
.A1(n_593),
.A2(n_426),
.B(n_423),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_581),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_641),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_584),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_585),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_587),
.Y(n_711)
);

INVx1_ASAP7_75t_SL g712 ( 
.A(n_595),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_586),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_643),
.Y(n_714)
);

NAND2xp33_ASAP7_75t_L g715 ( 
.A(n_614),
.B(n_473),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_591),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_645),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_646),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_647),
.B(n_410),
.Y(n_719)
);

BUFx6f_ASAP7_75t_L g720 ( 
.A(n_648),
.Y(n_720)
);

NAND2xp33_ASAP7_75t_SL g721 ( 
.A(n_556),
.B(n_479),
.Y(n_721)
);

BUFx10_ASAP7_75t_L g722 ( 
.A(n_598),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_651),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_588),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_590),
.Y(n_725)
);

BUFx6f_ASAP7_75t_L g726 ( 
.A(n_611),
.Y(n_726)
);

INVxp67_ASAP7_75t_SL g727 ( 
.A(n_594),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_596),
.Y(n_728)
);

CKINVDCx20_ASAP7_75t_R g729 ( 
.A(n_579),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_600),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_605),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_607),
.Y(n_732)
);

CKINVDCx6p67_ASAP7_75t_R g733 ( 
.A(n_608),
.Y(n_733)
);

XNOR2xp5_ASAP7_75t_L g734 ( 
.A(n_561),
.B(n_481),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_609),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_634),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_616),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_622),
.Y(n_738)
);

AND2x4_ASAP7_75t_L g739 ( 
.A(n_652),
.B(n_423),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_654),
.B(n_412),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_657),
.Y(n_741)
);

INVx5_ASAP7_75t_L g742 ( 
.A(n_680),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_727),
.B(n_603),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_727),
.B(n_631),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_656),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_664),
.B(n_636),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_669),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_671),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_669),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_678),
.B(n_640),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_678),
.B(n_644),
.Y(n_751)
);

BUFx6f_ASAP7_75t_L g752 ( 
.A(n_680),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_660),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_667),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_658),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_661),
.Y(n_756)
);

BUFx2_ASAP7_75t_L g757 ( 
.A(n_664),
.Y(n_757)
);

INVx5_ASAP7_75t_L g758 ( 
.A(n_680),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_704),
.B(n_650),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_689),
.B(n_638),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_712),
.B(n_653),
.Y(n_761)
);

AND2x4_ASAP7_75t_L g762 ( 
.A(n_674),
.B(n_560),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_712),
.B(n_612),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_714),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_665),
.Y(n_765)
);

AND2x2_ASAP7_75t_L g766 ( 
.A(n_689),
.B(n_594),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_666),
.Y(n_767)
);

AND2x2_ASAP7_75t_L g768 ( 
.A(n_673),
.B(n_692),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_677),
.B(n_426),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_675),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_676),
.Y(n_771)
);

INVx8_ASAP7_75t_L g772 ( 
.A(n_679),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_718),
.Y(n_773)
);

BUFx3_ASAP7_75t_L g774 ( 
.A(n_726),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_684),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_720),
.Y(n_776)
);

INVx4_ASAP7_75t_L g777 ( 
.A(n_726),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_685),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_726),
.B(n_618),
.Y(n_779)
);

INVx4_ASAP7_75t_L g780 ( 
.A(n_726),
.Y(n_780)
);

OAI22xp33_ASAP7_75t_SL g781 ( 
.A1(n_695),
.A2(n_728),
.B1(n_700),
.B2(n_719),
.Y(n_781)
);

AOI22xp33_ASAP7_75t_L g782 ( 
.A1(n_691),
.A2(n_568),
.B1(n_512),
.B2(n_431),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_693),
.Y(n_783)
);

BUFx3_ASAP7_75t_L g784 ( 
.A(n_699),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_692),
.B(n_630),
.Y(n_785)
);

OR2x2_ASAP7_75t_L g786 ( 
.A(n_662),
.B(n_580),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_720),
.Y(n_787)
);

BUFx6f_ASAP7_75t_L g788 ( 
.A(n_720),
.Y(n_788)
);

INVx4_ASAP7_75t_L g789 ( 
.A(n_720),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_703),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_683),
.B(n_580),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_686),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_682),
.Y(n_793)
);

INVx4_ASAP7_75t_L g794 ( 
.A(n_688),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_705),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_696),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_708),
.Y(n_797)
);

AND2x4_ASAP7_75t_L g798 ( 
.A(n_674),
.B(n_480),
.Y(n_798)
);

AOI22xp5_ASAP7_75t_SL g799 ( 
.A1(n_734),
.A2(n_601),
.B1(n_561),
.B2(n_589),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_710),
.Y(n_800)
);

BUFx2_ASAP7_75t_L g801 ( 
.A(n_721),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_707),
.B(n_623),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_677),
.B(n_431),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_709),
.Y(n_804)
);

BUFx6f_ASAP7_75t_L g805 ( 
.A(n_688),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_717),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_739),
.B(n_623),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_713),
.Y(n_808)
);

BUFx10_ASAP7_75t_L g809 ( 
.A(n_711),
.Y(n_809)
);

AND2x4_ASAP7_75t_L g810 ( 
.A(n_739),
.B(n_482),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_724),
.Y(n_811)
);

AND2x6_ASAP7_75t_L g812 ( 
.A(n_730),
.B(n_512),
.Y(n_812)
);

INVx1_ASAP7_75t_SL g813 ( 
.A(n_701),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_723),
.Y(n_814)
);

INVx1_ASAP7_75t_SL g815 ( 
.A(n_670),
.Y(n_815)
);

NAND2xp33_ASAP7_75t_L g816 ( 
.A(n_662),
.B(n_357),
.Y(n_816)
);

AND2x6_ASAP7_75t_L g817 ( 
.A(n_735),
.B(n_357),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_725),
.Y(n_818)
);

OR2x6_ASAP7_75t_L g819 ( 
.A(n_738),
.B(n_624),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_691),
.B(n_483),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_695),
.B(n_649),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_702),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_706),
.B(n_487),
.Y(n_823)
);

BUFx6f_ASAP7_75t_L g824 ( 
.A(n_688),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_716),
.B(n_624),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_688),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_668),
.B(n_582),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_731),
.B(n_413),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_706),
.B(n_492),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_SL g830 ( 
.A(n_732),
.B(n_461),
.Y(n_830)
);

AOI22xp33_ASAP7_75t_L g831 ( 
.A1(n_786),
.A2(n_782),
.B1(n_823),
.B2(n_820),
.Y(n_831)
);

AOI22xp33_ASAP7_75t_L g832 ( 
.A1(n_782),
.A2(n_721),
.B1(n_715),
.B2(n_498),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_781),
.B(n_668),
.Y(n_833)
);

INVx4_ASAP7_75t_L g834 ( 
.A(n_777),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_781),
.B(n_722),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_766),
.B(n_700),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_777),
.B(n_719),
.Y(n_837)
);

AOI22xp5_ASAP7_75t_L g838 ( 
.A1(n_827),
.A2(n_687),
.B1(n_737),
.B2(n_659),
.Y(n_838)
);

BUFx6f_ASAP7_75t_L g839 ( 
.A(n_774),
.Y(n_839)
);

INVx1_ASAP7_75t_SL g840 ( 
.A(n_757),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_780),
.B(n_740),
.Y(n_841)
);

AOI22xp5_ASAP7_75t_L g842 ( 
.A1(n_743),
.A2(n_687),
.B1(n_740),
.B2(n_672),
.Y(n_842)
);

BUFx3_ASAP7_75t_L g843 ( 
.A(n_772),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_741),
.Y(n_844)
);

NAND3xp33_ASAP7_75t_L g845 ( 
.A(n_760),
.B(n_736),
.C(n_509),
.Y(n_845)
);

AND2x4_ASAP7_75t_L g846 ( 
.A(n_784),
.B(n_681),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_780),
.B(n_698),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_807),
.B(n_698),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_762),
.B(n_698),
.Y(n_849)
);

AOI221xp5_ASAP7_75t_L g850 ( 
.A1(n_821),
.A2(n_540),
.B1(n_548),
.B2(n_539),
.C(n_494),
.Y(n_850)
);

INVx3_ASAP7_75t_L g851 ( 
.A(n_788),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_811),
.Y(n_852)
);

BUFx6f_ASAP7_75t_L g853 ( 
.A(n_752),
.Y(n_853)
);

OAI22xp5_ASAP7_75t_L g854 ( 
.A1(n_819),
.A2(n_542),
.B1(n_501),
.B2(n_502),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_762),
.B(n_745),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_755),
.B(n_698),
.Y(n_856)
);

OR2x6_ASAP7_75t_L g857 ( 
.A(n_772),
.B(n_681),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_756),
.B(n_690),
.Y(n_858)
);

BUFx3_ASAP7_75t_L g859 ( 
.A(n_772),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_765),
.B(n_690),
.Y(n_860)
);

HB1xp67_ASAP7_75t_L g861 ( 
.A(n_813),
.Y(n_861)
);

BUFx6f_ASAP7_75t_L g862 ( 
.A(n_752),
.Y(n_862)
);

OR2x2_ASAP7_75t_L g863 ( 
.A(n_785),
.B(n_733),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_767),
.B(n_770),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_771),
.B(n_694),
.Y(n_865)
);

INVx3_ASAP7_75t_L g866 ( 
.A(n_788),
.Y(n_866)
);

NAND2x1_ASAP7_75t_L g867 ( 
.A(n_789),
.B(n_357),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_818),
.Y(n_868)
);

AOI22xp33_ASAP7_75t_L g869 ( 
.A1(n_820),
.A2(n_497),
.B1(n_507),
.B2(n_506),
.Y(n_869)
);

AND2x2_ASAP7_75t_SL g870 ( 
.A(n_830),
.B(n_601),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_830),
.B(n_722),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_764),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_775),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_778),
.Y(n_874)
);

AOI22xp5_ASAP7_75t_L g875 ( 
.A1(n_768),
.A2(n_417),
.B1(n_420),
.B2(n_418),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_783),
.Y(n_876)
);

NAND2x1_ASAP7_75t_L g877 ( 
.A(n_789),
.B(n_384),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_746),
.B(n_744),
.Y(n_878)
);

NAND2xp33_ASAP7_75t_L g879 ( 
.A(n_812),
.B(n_421),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_773),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_793),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_759),
.B(n_702),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_790),
.B(n_694),
.Y(n_883)
);

AND2x4_ASAP7_75t_L g884 ( 
.A(n_795),
.B(n_702),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_797),
.B(n_513),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_806),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_814),
.B(n_516),
.Y(n_887)
);

AOI22xp33_ASAP7_75t_L g888 ( 
.A1(n_823),
.A2(n_525),
.B1(n_526),
.B2(n_520),
.Y(n_888)
);

INVxp67_ASAP7_75t_SL g889 ( 
.A(n_788),
.Y(n_889)
);

INVx2_ASAP7_75t_SL g890 ( 
.A(n_798),
.Y(n_890)
);

NAND3xp33_ASAP7_75t_L g891 ( 
.A(n_791),
.B(n_427),
.C(n_425),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_796),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_776),
.B(n_527),
.Y(n_893)
);

AOI22xp33_ASAP7_75t_L g894 ( 
.A1(n_829),
.A2(n_541),
.B1(n_549),
.B2(n_538),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_800),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_SL g896 ( 
.A(n_801),
.B(n_428),
.Y(n_896)
);

O2A1O1Ixp33_ASAP7_75t_L g897 ( 
.A1(n_829),
.A2(n_554),
.B(n_552),
.C(n_610),
.Y(n_897)
);

INVx2_ASAP7_75t_SL g898 ( 
.A(n_798),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_761),
.B(n_663),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_787),
.B(n_433),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_808),
.Y(n_901)
);

NOR2xp33_ASAP7_75t_L g902 ( 
.A(n_802),
.B(n_697),
.Y(n_902)
);

INVx4_ASAP7_75t_L g903 ( 
.A(n_805),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_753),
.Y(n_904)
);

BUFx3_ASAP7_75t_L g905 ( 
.A(n_809),
.Y(n_905)
);

AOI22xp33_ASAP7_75t_L g906 ( 
.A1(n_769),
.A2(n_803),
.B1(n_810),
.B2(n_812),
.Y(n_906)
);

NOR2xp33_ASAP7_75t_L g907 ( 
.A(n_825),
.B(n_729),
.Y(n_907)
);

A2O1A1Ixp33_ASAP7_75t_L g908 ( 
.A1(n_769),
.A2(n_436),
.B(n_438),
.C(n_437),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_826),
.B(n_439),
.Y(n_909)
);

AOI22xp33_ASAP7_75t_L g910 ( 
.A1(n_803),
.A2(n_499),
.B1(n_384),
.B2(n_442),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_794),
.B(n_440),
.Y(n_911)
);

INVx3_ASAP7_75t_L g912 ( 
.A(n_805),
.Y(n_912)
);

O2A1O1Ixp33_ASAP7_75t_L g913 ( 
.A1(n_816),
.A2(n_446),
.B(n_447),
.C(n_443),
.Y(n_913)
);

INVx3_ASAP7_75t_L g914 ( 
.A(n_805),
.Y(n_914)
);

NAND2x1p5_ASAP7_75t_L g915 ( 
.A(n_779),
.B(n_384),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_754),
.Y(n_916)
);

AND2x4_ASAP7_75t_L g917 ( 
.A(n_822),
.B(n_448),
.Y(n_917)
);

NOR2xp67_ASAP7_75t_L g918 ( 
.A(n_748),
.B(n_449),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_SL g919 ( 
.A(n_810),
.B(n_451),
.Y(n_919)
);

BUFx5_ASAP7_75t_L g920 ( 
.A(n_812),
.Y(n_920)
);

OR2x2_ASAP7_75t_L g921 ( 
.A(n_813),
.B(n_9),
.Y(n_921)
);

INVx4_ASAP7_75t_L g922 ( 
.A(n_824),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_747),
.Y(n_923)
);

NOR2xp33_ASAP7_75t_L g924 ( 
.A(n_750),
.B(n_460),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_794),
.B(n_462),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_749),
.Y(n_926)
);

CKINVDCx16_ASAP7_75t_R g927 ( 
.A(n_843),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_873),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_844),
.Y(n_929)
);

AOI22xp33_ASAP7_75t_SL g930 ( 
.A1(n_870),
.A2(n_799),
.B1(n_819),
.B2(n_804),
.Y(n_930)
);

BUFx3_ASAP7_75t_L g931 ( 
.A(n_859),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_874),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_916),
.Y(n_933)
);

OR2x4_ASAP7_75t_L g934 ( 
.A(n_921),
.B(n_799),
.Y(n_934)
);

INVxp67_ASAP7_75t_SL g935 ( 
.A(n_831),
.Y(n_935)
);

OR2x6_ASAP7_75t_L g936 ( 
.A(n_905),
.B(n_763),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_852),
.Y(n_937)
);

INVx2_ASAP7_75t_SL g938 ( 
.A(n_861),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_868),
.Y(n_939)
);

OR2x2_ASAP7_75t_L g940 ( 
.A(n_840),
.B(n_815),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_872),
.Y(n_941)
);

INVx4_ASAP7_75t_L g942 ( 
.A(n_839),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_836),
.B(n_819),
.Y(n_943)
);

BUFx2_ASAP7_75t_L g944 ( 
.A(n_846),
.Y(n_944)
);

BUFx4f_ASAP7_75t_L g945 ( 
.A(n_857),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_876),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_886),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_880),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_892),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_848),
.B(n_812),
.Y(n_950)
);

CKINVDCx20_ASAP7_75t_R g951 ( 
.A(n_838),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_881),
.Y(n_952)
);

NOR3xp33_ASAP7_75t_SL g953 ( 
.A(n_854),
.B(n_792),
.C(n_751),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_837),
.B(n_824),
.Y(n_954)
);

AND2x4_ASAP7_75t_L g955 ( 
.A(n_846),
.B(n_828),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_895),
.Y(n_956)
);

OAI22xp33_ASAP7_75t_L g957 ( 
.A1(n_833),
.A2(n_815),
.B1(n_499),
.B2(n_384),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_901),
.Y(n_958)
);

INVx3_ASAP7_75t_L g959 ( 
.A(n_851),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_904),
.Y(n_960)
);

INVx2_ASAP7_75t_SL g961 ( 
.A(n_917),
.Y(n_961)
);

BUFx3_ASAP7_75t_L g962 ( 
.A(n_839),
.Y(n_962)
);

HB1xp67_ASAP7_75t_L g963 ( 
.A(n_855),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_923),
.Y(n_964)
);

AND2x4_ASAP7_75t_L g965 ( 
.A(n_890),
.B(n_898),
.Y(n_965)
);

OAI22xp5_ASAP7_75t_L g966 ( 
.A1(n_906),
.A2(n_824),
.B1(n_464),
.B2(n_467),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_864),
.Y(n_967)
);

BUFx3_ASAP7_75t_L g968 ( 
.A(n_839),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_SL g969 ( 
.A(n_842),
.B(n_809),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_841),
.B(n_849),
.Y(n_970)
);

INVx2_ASAP7_75t_SL g971 ( 
.A(n_917),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_926),
.Y(n_972)
);

OR2x6_ASAP7_75t_L g973 ( 
.A(n_857),
.B(n_499),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_884),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_884),
.Y(n_975)
);

A2O1A1Ixp33_ASAP7_75t_L g976 ( 
.A1(n_897),
.A2(n_471),
.B(n_472),
.C(n_463),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_869),
.B(n_752),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_856),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_888),
.B(n_894),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_851),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_902),
.Y(n_981)
);

AND2x4_ASAP7_75t_L g982 ( 
.A(n_882),
.B(n_742),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_858),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_866),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_866),
.Y(n_985)
);

INVxp67_ASAP7_75t_L g986 ( 
.A(n_878),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_860),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_835),
.B(n_499),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_912),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_907),
.Y(n_990)
);

HB1xp67_ASAP7_75t_L g991 ( 
.A(n_853),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_912),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_914),
.Y(n_993)
);

INVx4_ASAP7_75t_L g994 ( 
.A(n_853),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_865),
.Y(n_995)
);

AOI22xp33_ASAP7_75t_L g996 ( 
.A1(n_832),
.A2(n_817),
.B1(n_475),
.B2(n_484),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_883),
.Y(n_997)
);

AND2x4_ASAP7_75t_L g998 ( 
.A(n_845),
.B(n_742),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_967),
.B(n_924),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_963),
.B(n_918),
.Y(n_1000)
);

BUFx4_ASAP7_75t_SL g1001 ( 
.A(n_931),
.Y(n_1001)
);

BUFx12f_ASAP7_75t_L g1002 ( 
.A(n_929),
.Y(n_1002)
);

INVx3_ASAP7_75t_L g1003 ( 
.A(n_959),
.Y(n_1003)
);

AND2x2_ASAP7_75t_L g1004 ( 
.A(n_943),
.B(n_899),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_928),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_SL g1006 ( 
.A1(n_935),
.A2(n_834),
.B(n_903),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_932),
.Y(n_1007)
);

INVx3_ASAP7_75t_L g1008 ( 
.A(n_959),
.Y(n_1008)
);

A2O1A1Ixp33_ASAP7_75t_L g1009 ( 
.A1(n_935),
.A2(n_850),
.B(n_891),
.C(n_871),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_963),
.B(n_834),
.Y(n_1010)
);

AND2x2_ASAP7_75t_L g1011 ( 
.A(n_981),
.B(n_990),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_970),
.A2(n_922),
.B(n_903),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_983),
.B(n_885),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_946),
.Y(n_1014)
);

AO31x2_ASAP7_75t_L g1015 ( 
.A1(n_976),
.A2(n_908),
.A3(n_950),
.B(n_954),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_987),
.B(n_887),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_933),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_995),
.B(n_896),
.Y(n_1018)
);

NOR2xp67_ASAP7_75t_L g1019 ( 
.A(n_938),
.B(n_940),
.Y(n_1019)
);

AOI21x1_ASAP7_75t_L g1020 ( 
.A1(n_988),
.A2(n_847),
.B(n_893),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_997),
.B(n_875),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_978),
.B(n_915),
.Y(n_1022)
);

AOI21x1_ASAP7_75t_L g1023 ( 
.A1(n_988),
.A2(n_925),
.B(n_911),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_986),
.B(n_910),
.Y(n_1024)
);

OAI21x1_ASAP7_75t_L g1025 ( 
.A1(n_980),
.A2(n_914),
.B(n_909),
.Y(n_1025)
);

NOR2xp33_ASAP7_75t_L g1026 ( 
.A(n_986),
.B(n_863),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_SL g1027 ( 
.A(n_955),
.B(n_853),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_947),
.B(n_889),
.Y(n_1028)
);

OAI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_979),
.A2(n_913),
.B(n_900),
.Y(n_1029)
);

OA21x2_ASAP7_75t_L g1030 ( 
.A1(n_980),
.A2(n_919),
.B(n_485),
.Y(n_1030)
);

BUFx6f_ASAP7_75t_L g1031 ( 
.A(n_962),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_960),
.B(n_922),
.Y(n_1032)
);

BUFx8_ASAP7_75t_L g1033 ( 
.A(n_931),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_977),
.A2(n_862),
.B(n_955),
.Y(n_1034)
);

AOI211x1_ASAP7_75t_L g1035 ( 
.A1(n_957),
.A2(n_12),
.B(n_10),
.C(n_11),
.Y(n_1035)
);

O2A1O1Ixp5_ASAP7_75t_SL g1036 ( 
.A1(n_969),
.A2(n_879),
.B(n_817),
.C(n_877),
.Y(n_1036)
);

OAI21x1_ASAP7_75t_L g1037 ( 
.A1(n_984),
.A2(n_867),
.B(n_920),
.Y(n_1037)
);

O2A1O1Ixp5_ASAP7_75t_L g1038 ( 
.A1(n_969),
.A2(n_920),
.B(n_817),
.C(n_862),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_966),
.A2(n_862),
.B(n_758),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_994),
.A2(n_758),
.B(n_742),
.Y(n_1040)
);

BUFx3_ASAP7_75t_L g1041 ( 
.A(n_962),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_960),
.B(n_920),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_933),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_937),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_972),
.B(n_920),
.Y(n_1045)
);

OAI22xp33_ASAP7_75t_L g1046 ( 
.A1(n_951),
.A2(n_486),
.B1(n_490),
.B2(n_474),
.Y(n_1046)
);

OAI22xp5_ASAP7_75t_L g1047 ( 
.A1(n_951),
.A2(n_493),
.B1(n_495),
.B2(n_491),
.Y(n_1047)
);

OAI21x1_ASAP7_75t_L g1048 ( 
.A1(n_984),
.A2(n_920),
.B(n_817),
.Y(n_1048)
);

OAI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_957),
.A2(n_500),
.B(n_496),
.Y(n_1049)
);

A2O1A1Ixp33_ASAP7_75t_L g1050 ( 
.A1(n_953),
.A2(n_508),
.B(n_510),
.C(n_504),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_SL g1051 ( 
.A(n_930),
.B(n_511),
.Y(n_1051)
);

INVx3_ASAP7_75t_L g1052 ( 
.A(n_994),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_974),
.A2(n_758),
.B(n_515),
.Y(n_1053)
);

OAI21x1_ASAP7_75t_L g1054 ( 
.A1(n_985),
.A2(n_59),
.B(n_57),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_975),
.A2(n_941),
.B(n_937),
.Y(n_1055)
);

NOR2xp33_ASAP7_75t_L g1056 ( 
.A(n_934),
.B(n_514),
.Y(n_1056)
);

A2O1A1Ixp33_ASAP7_75t_L g1057 ( 
.A1(n_953),
.A2(n_519),
.B(n_521),
.C(n_517),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_1017),
.Y(n_1058)
);

CKINVDCx6p67_ASAP7_75t_R g1059 ( 
.A(n_1002),
.Y(n_1059)
);

OAI21x1_ASAP7_75t_L g1060 ( 
.A1(n_1025),
.A2(n_992),
.B(n_985),
.Y(n_1060)
);

INVx6_ASAP7_75t_L g1061 ( 
.A(n_1033),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_1044),
.Y(n_1062)
);

AND2x2_ASAP7_75t_L g1063 ( 
.A(n_1004),
.B(n_930),
.Y(n_1063)
);

OAI21x1_ASAP7_75t_L g1064 ( 
.A1(n_1037),
.A2(n_992),
.B(n_972),
.Y(n_1064)
);

INVx3_ASAP7_75t_L g1065 ( 
.A(n_1052),
.Y(n_1065)
);

OAI21x1_ASAP7_75t_L g1066 ( 
.A1(n_1048),
.A2(n_948),
.B(n_941),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_999),
.A2(n_996),
.B(n_998),
.Y(n_1067)
);

NOR2xp33_ASAP7_75t_L g1068 ( 
.A(n_1021),
.B(n_934),
.Y(n_1068)
);

OA21x2_ASAP7_75t_L g1069 ( 
.A1(n_1038),
.A2(n_976),
.B(n_948),
.Y(n_1069)
);

OAI21x1_ASAP7_75t_L g1070 ( 
.A1(n_1054),
.A2(n_993),
.B(n_989),
.Y(n_1070)
);

AND2x2_ASAP7_75t_L g1071 ( 
.A(n_1011),
.B(n_944),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_1005),
.Y(n_1072)
);

NOR2xp67_ASAP7_75t_SL g1073 ( 
.A(n_1006),
.B(n_927),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_L g1074 ( 
.A(n_1018),
.B(n_956),
.Y(n_1074)
);

OA21x2_ASAP7_75t_L g1075 ( 
.A1(n_1029),
.A2(n_949),
.B(n_964),
.Y(n_1075)
);

OAI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_1029),
.A2(n_996),
.B(n_958),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_1013),
.B(n_991),
.Y(n_1077)
);

OAI21x1_ASAP7_75t_L g1078 ( 
.A1(n_1023),
.A2(n_952),
.B(n_939),
.Y(n_1078)
);

OR2x2_ASAP7_75t_L g1079 ( 
.A(n_1016),
.B(n_936),
.Y(n_1079)
);

AND2x2_ASAP7_75t_L g1080 ( 
.A(n_1026),
.B(n_965),
.Y(n_1080)
);

OAI21x1_ASAP7_75t_L g1081 ( 
.A1(n_1020),
.A2(n_991),
.B(n_998),
.Y(n_1081)
);

INVx1_ASAP7_75t_SL g1082 ( 
.A(n_1001),
.Y(n_1082)
);

AO21x2_ASAP7_75t_L g1083 ( 
.A1(n_1012),
.A2(n_982),
.B(n_965),
.Y(n_1083)
);

OA21x2_ASAP7_75t_L g1084 ( 
.A1(n_1055),
.A2(n_982),
.B(n_971),
.Y(n_1084)
);

NAND2xp33_ASAP7_75t_SL g1085 ( 
.A(n_1031),
.B(n_942),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_1007),
.Y(n_1086)
);

O2A1O1Ixp33_ASAP7_75t_SL g1087 ( 
.A1(n_1009),
.A2(n_961),
.B(n_973),
.C(n_13),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_1014),
.Y(n_1088)
);

AND2x4_ASAP7_75t_L g1089 ( 
.A(n_1041),
.B(n_968),
.Y(n_1089)
);

OAI21x1_ASAP7_75t_L g1090 ( 
.A1(n_1036),
.A2(n_945),
.B(n_942),
.Y(n_1090)
);

AO21x2_ASAP7_75t_L g1091 ( 
.A1(n_1039),
.A2(n_973),
.B(n_968),
.Y(n_1091)
);

CKINVDCx8_ASAP7_75t_R g1092 ( 
.A(n_1031),
.Y(n_1092)
);

OAI21x1_ASAP7_75t_L g1093 ( 
.A1(n_1034),
.A2(n_945),
.B(n_973),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_1043),
.Y(n_1094)
);

OR2x2_ASAP7_75t_L g1095 ( 
.A(n_1000),
.B(n_936),
.Y(n_1095)
);

NAND3xp33_ASAP7_75t_L g1096 ( 
.A(n_1047),
.B(n_936),
.C(n_523),
.Y(n_1096)
);

OAI21x1_ASAP7_75t_L g1097 ( 
.A1(n_1042),
.A2(n_64),
.B(n_62),
.Y(n_1097)
);

BUFx2_ASAP7_75t_L g1098 ( 
.A(n_1033),
.Y(n_1098)
);

OAI22xp5_ASAP7_75t_L g1099 ( 
.A1(n_1035),
.A2(n_524),
.B1(n_529),
.B2(n_522),
.Y(n_1099)
);

BUFx4f_ASAP7_75t_L g1100 ( 
.A(n_1031),
.Y(n_1100)
);

OAI21x1_ASAP7_75t_L g1101 ( 
.A1(n_1045),
.A2(n_67),
.B(n_66),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_1024),
.B(n_530),
.Y(n_1102)
);

NOR2x1_ASAP7_75t_SL g1103 ( 
.A(n_1022),
.B(n_70),
.Y(n_1103)
);

HB1xp67_ASAP7_75t_L g1104 ( 
.A(n_1019),
.Y(n_1104)
);

INVx8_ASAP7_75t_L g1105 ( 
.A(n_1052),
.Y(n_1105)
);

INVx2_ASAP7_75t_L g1106 ( 
.A(n_1003),
.Y(n_1106)
);

OAI21x1_ASAP7_75t_L g1107 ( 
.A1(n_1032),
.A2(n_75),
.B(n_74),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_1010),
.A2(n_553),
.B(n_534),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_SL g1109 ( 
.A(n_1050),
.B(n_532),
.Y(n_1109)
);

NOR2xp33_ASAP7_75t_L g1110 ( 
.A(n_1051),
.B(n_536),
.Y(n_1110)
);

AO31x2_ASAP7_75t_L g1111 ( 
.A1(n_1057),
.A2(n_10),
.A3(n_12),
.B(n_13),
.Y(n_1111)
);

A2O1A1Ixp33_ASAP7_75t_L g1112 ( 
.A1(n_1056),
.A2(n_551),
.B(n_550),
.C(n_545),
.Y(n_1112)
);

NOR3xp33_ASAP7_75t_SL g1113 ( 
.A(n_1096),
.B(n_1046),
.C(n_1047),
.Y(n_1113)
);

OAI21x1_ASAP7_75t_L g1114 ( 
.A1(n_1070),
.A2(n_1030),
.B(n_1053),
.Y(n_1114)
);

OR2x6_ASAP7_75t_L g1115 ( 
.A(n_1093),
.B(n_1028),
.Y(n_1115)
);

HB1xp67_ASAP7_75t_L g1116 ( 
.A(n_1080),
.Y(n_1116)
);

OAI22xp5_ASAP7_75t_SL g1117 ( 
.A1(n_1068),
.A2(n_1049),
.B1(n_1030),
.B2(n_1028),
.Y(n_1117)
);

OAI22xp5_ASAP7_75t_L g1118 ( 
.A1(n_1068),
.A2(n_1079),
.B1(n_1095),
.B2(n_1096),
.Y(n_1118)
);

AOI22xp33_ASAP7_75t_SL g1119 ( 
.A1(n_1110),
.A2(n_1049),
.B1(n_1008),
.B2(n_1003),
.Y(n_1119)
);

OR2x6_ASAP7_75t_L g1120 ( 
.A(n_1061),
.B(n_1027),
.Y(n_1120)
);

NAND2xp33_ASAP7_75t_SL g1121 ( 
.A(n_1104),
.B(n_1008),
.Y(n_1121)
);

BUFx3_ASAP7_75t_L g1122 ( 
.A(n_1092),
.Y(n_1122)
);

AND2x2_ASAP7_75t_L g1123 ( 
.A(n_1063),
.B(n_1071),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_1076),
.A2(n_1067),
.B(n_1084),
.Y(n_1124)
);

AND2x2_ASAP7_75t_L g1125 ( 
.A(n_1074),
.B(n_537),
.Y(n_1125)
);

AOI221x1_ASAP7_75t_L g1126 ( 
.A1(n_1099),
.A2(n_1040),
.B1(n_1015),
.B2(n_17),
.C(n_18),
.Y(n_1126)
);

BUFx2_ASAP7_75t_L g1127 ( 
.A(n_1089),
.Y(n_1127)
);

OAI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_1067),
.A2(n_543),
.B(n_1015),
.Y(n_1128)
);

NAND2xp33_ASAP7_75t_R g1129 ( 
.A(n_1098),
.B(n_80),
.Y(n_1129)
);

CKINVDCx16_ASAP7_75t_R g1130 ( 
.A(n_1082),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1086),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_1094),
.Y(n_1132)
);

AND2x2_ASAP7_75t_L g1133 ( 
.A(n_1074),
.B(n_1077),
.Y(n_1133)
);

CKINVDCx11_ASAP7_75t_R g1134 ( 
.A(n_1059),
.Y(n_1134)
);

AOI22xp33_ASAP7_75t_L g1135 ( 
.A1(n_1110),
.A2(n_1015),
.B1(n_15),
.B2(n_18),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_1058),
.Y(n_1136)
);

INVx1_ASAP7_75t_SL g1137 ( 
.A(n_1104),
.Y(n_1137)
);

CKINVDCx20_ASAP7_75t_R g1138 ( 
.A(n_1082),
.Y(n_1138)
);

OAI22xp33_ASAP7_75t_L g1139 ( 
.A1(n_1102),
.A2(n_14),
.B1(n_15),
.B2(n_19),
.Y(n_1139)
);

AND2x2_ASAP7_75t_L g1140 ( 
.A(n_1077),
.B(n_20),
.Y(n_1140)
);

CKINVDCx16_ASAP7_75t_R g1141 ( 
.A(n_1089),
.Y(n_1141)
);

OAI21x1_ASAP7_75t_L g1142 ( 
.A1(n_1060),
.A2(n_85),
.B(n_83),
.Y(n_1142)
);

OR2x2_ASAP7_75t_L g1143 ( 
.A(n_1102),
.B(n_20),
.Y(n_1143)
);

AOI22xp5_ASAP7_75t_L g1144 ( 
.A1(n_1087),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_1061),
.Y(n_1145)
);

NAND2xp33_ASAP7_75t_R g1146 ( 
.A(n_1075),
.B(n_86),
.Y(n_1146)
);

AOI222xp33_ASAP7_75t_L g1147 ( 
.A1(n_1099),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.C1(n_24),
.C2(n_25),
.Y(n_1147)
);

AO221x2_ASAP7_75t_L g1148 ( 
.A1(n_1076),
.A2(n_24),
.B1(n_26),
.B2(n_27),
.C(n_28),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_1062),
.Y(n_1149)
);

INVxp33_ASAP7_75t_L g1150 ( 
.A(n_1100),
.Y(n_1150)
);

OAI22xp33_ASAP7_75t_L g1151 ( 
.A1(n_1061),
.A2(n_26),
.B1(n_28),
.B2(n_29),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1072),
.Y(n_1152)
);

AND2x2_ASAP7_75t_L g1153 ( 
.A(n_1088),
.B(n_29),
.Y(n_1153)
);

OAI22xp33_ASAP7_75t_L g1154 ( 
.A1(n_1100),
.A2(n_1108),
.B1(n_1065),
.B2(n_1105),
.Y(n_1154)
);

OAI22xp5_ASAP7_75t_L g1155 ( 
.A1(n_1112),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1106),
.Y(n_1156)
);

AOI22xp33_ASAP7_75t_L g1157 ( 
.A1(n_1109),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_1157)
);

AND2x4_ASAP7_75t_L g1158 ( 
.A(n_1065),
.B(n_88),
.Y(n_1158)
);

OAI22xp5_ASAP7_75t_L g1159 ( 
.A1(n_1108),
.A2(n_1109),
.B1(n_1105),
.B2(n_1084),
.Y(n_1159)
);

CKINVDCx14_ASAP7_75t_R g1160 ( 
.A(n_1085),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1073),
.B(n_33),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_1105),
.Y(n_1162)
);

OAI21x1_ASAP7_75t_L g1163 ( 
.A1(n_1078),
.A2(n_90),
.B(n_89),
.Y(n_1163)
);

AOI22xp5_ASAP7_75t_L g1164 ( 
.A1(n_1087),
.A2(n_1075),
.B1(n_1091),
.B2(n_1083),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1081),
.Y(n_1165)
);

OR2x2_ASAP7_75t_L g1166 ( 
.A(n_1111),
.B(n_34),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_1103),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1111),
.Y(n_1168)
);

AND2x4_ASAP7_75t_L g1169 ( 
.A(n_1091),
.B(n_1083),
.Y(n_1169)
);

AOI221xp5_ASAP7_75t_L g1170 ( 
.A1(n_1139),
.A2(n_1111),
.B1(n_36),
.B2(n_37),
.C(n_38),
.Y(n_1170)
);

CKINVDCx14_ASAP7_75t_R g1171 ( 
.A(n_1134),
.Y(n_1171)
);

OAI22xp5_ASAP7_75t_L g1172 ( 
.A1(n_1113),
.A2(n_1069),
.B1(n_1090),
.B2(n_1107),
.Y(n_1172)
);

BUFx2_ASAP7_75t_L g1173 ( 
.A(n_1127),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_1124),
.A2(n_1069),
.B(n_1064),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_1130),
.Y(n_1175)
);

AOI22xp33_ASAP7_75t_L g1176 ( 
.A1(n_1148),
.A2(n_1101),
.B1(n_1097),
.B2(n_1066),
.Y(n_1176)
);

OAI21xp33_ASAP7_75t_L g1177 ( 
.A1(n_1147),
.A2(n_34),
.B(n_36),
.Y(n_1177)
);

AND2x2_ASAP7_75t_L g1178 ( 
.A(n_1123),
.B(n_91),
.Y(n_1178)
);

BUFx3_ASAP7_75t_L g1179 ( 
.A(n_1122),
.Y(n_1179)
);

INVx3_ASAP7_75t_L g1180 ( 
.A(n_1158),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1152),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1131),
.Y(n_1182)
);

OAI211xp5_ASAP7_75t_SL g1183 ( 
.A1(n_1143),
.A2(n_1137),
.B(n_1118),
.C(n_1144),
.Y(n_1183)
);

AND2x4_ASAP7_75t_L g1184 ( 
.A(n_1120),
.B(n_93),
.Y(n_1184)
);

AOI222xp33_ASAP7_75t_L g1185 ( 
.A1(n_1155),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.C1(n_40),
.C2(n_41),
.Y(n_1185)
);

OAI221xp5_ASAP7_75t_L g1186 ( 
.A1(n_1157),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.C(n_42),
.Y(n_1186)
);

OAI22xp5_ASAP7_75t_L g1187 ( 
.A1(n_1160),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_1187)
);

OAI22xp5_ASAP7_75t_L g1188 ( 
.A1(n_1133),
.A2(n_45),
.B1(n_46),
.B2(n_48),
.Y(n_1188)
);

AOI22xp33_ASAP7_75t_L g1189 ( 
.A1(n_1148),
.A2(n_46),
.B1(n_48),
.B2(n_49),
.Y(n_1189)
);

AND2x4_ASAP7_75t_L g1190 ( 
.A(n_1120),
.B(n_94),
.Y(n_1190)
);

OAI22xp33_ASAP7_75t_L g1191 ( 
.A1(n_1144),
.A2(n_51),
.B1(n_53),
.B2(n_96),
.Y(n_1191)
);

AOI22xp33_ASAP7_75t_L g1192 ( 
.A1(n_1117),
.A2(n_51),
.B1(n_97),
.B2(n_98),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1132),
.Y(n_1193)
);

AOI22xp33_ASAP7_75t_L g1194 ( 
.A1(n_1135),
.A2(n_99),
.B1(n_100),
.B2(n_101),
.Y(n_1194)
);

INVx3_ASAP7_75t_L g1195 ( 
.A(n_1158),
.Y(n_1195)
);

OAI22xp33_ASAP7_75t_L g1196 ( 
.A1(n_1129),
.A2(n_102),
.B1(n_103),
.B2(n_105),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1159),
.A2(n_1128),
.B(n_1115),
.Y(n_1197)
);

A2O1A1Ixp33_ASAP7_75t_L g1198 ( 
.A1(n_1161),
.A2(n_107),
.B(n_108),
.C(n_110),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_L g1199 ( 
.A(n_1116),
.B(n_112),
.Y(n_1199)
);

INVx2_ASAP7_75t_L g1200 ( 
.A(n_1136),
.Y(n_1200)
);

AOI33xp33_ASAP7_75t_L g1201 ( 
.A1(n_1151),
.A2(n_113),
.A3(n_116),
.B1(n_118),
.B2(n_120),
.B3(n_122),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1149),
.Y(n_1202)
);

OAI211xp5_ASAP7_75t_L g1203 ( 
.A1(n_1126),
.A2(n_125),
.B(n_126),
.C(n_127),
.Y(n_1203)
);

INVx1_ASAP7_75t_SL g1204 ( 
.A(n_1121),
.Y(n_1204)
);

NOR2xp33_ASAP7_75t_L g1205 ( 
.A(n_1141),
.B(n_128),
.Y(n_1205)
);

OAI22xp5_ASAP7_75t_L g1206 ( 
.A1(n_1120),
.A2(n_130),
.B1(n_133),
.B2(n_136),
.Y(n_1206)
);

NAND3xp33_ASAP7_75t_L g1207 ( 
.A(n_1119),
.B(n_138),
.C(n_139),
.Y(n_1207)
);

AND2x2_ASAP7_75t_L g1208 ( 
.A(n_1140),
.B(n_140),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_1138),
.Y(n_1209)
);

AOI222xp33_ASAP7_75t_L g1210 ( 
.A1(n_1125),
.A2(n_141),
.B1(n_142),
.B2(n_143),
.C1(n_145),
.C2(n_150),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_1156),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1168),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1167),
.B(n_153),
.Y(n_1213)
);

AOI22xp5_ASAP7_75t_L g1214 ( 
.A1(n_1154),
.A2(n_154),
.B1(n_156),
.B2(n_159),
.Y(n_1214)
);

OAI22xp33_ASAP7_75t_L g1215 ( 
.A1(n_1146),
.A2(n_1166),
.B1(n_1150),
.B2(n_1145),
.Y(n_1215)
);

A2O1A1Ixp33_ASAP7_75t_L g1216 ( 
.A1(n_1164),
.A2(n_1169),
.B(n_1114),
.C(n_1163),
.Y(n_1216)
);

AOI22xp33_ASAP7_75t_L g1217 ( 
.A1(n_1115),
.A2(n_161),
.B1(n_166),
.B2(n_169),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1115),
.Y(n_1218)
);

AOI22xp33_ASAP7_75t_L g1219 ( 
.A1(n_1153),
.A2(n_173),
.B1(n_178),
.B2(n_179),
.Y(n_1219)
);

HB1xp67_ASAP7_75t_L g1220 ( 
.A(n_1169),
.Y(n_1220)
);

AOI221xp5_ASAP7_75t_L g1221 ( 
.A1(n_1164),
.A2(n_183),
.B1(n_188),
.B2(n_192),
.C(n_193),
.Y(n_1221)
);

BUFx2_ASAP7_75t_L g1222 ( 
.A(n_1162),
.Y(n_1222)
);

AOI22xp33_ASAP7_75t_L g1223 ( 
.A1(n_1165),
.A2(n_194),
.B1(n_197),
.B2(n_198),
.Y(n_1223)
);

AOI222xp33_ASAP7_75t_L g1224 ( 
.A1(n_1142),
.A2(n_199),
.B1(n_208),
.B2(n_214),
.C1(n_220),
.C2(n_224),
.Y(n_1224)
);

AOI22xp33_ASAP7_75t_L g1225 ( 
.A1(n_1148),
.A2(n_225),
.B1(n_226),
.B2(n_227),
.Y(n_1225)
);

OR2x2_ASAP7_75t_L g1226 ( 
.A(n_1220),
.B(n_228),
.Y(n_1226)
);

BUFx3_ASAP7_75t_L g1227 ( 
.A(n_1173),
.Y(n_1227)
);

INVxp67_ASAP7_75t_L g1228 ( 
.A(n_1179),
.Y(n_1228)
);

AND2x2_ASAP7_75t_L g1229 ( 
.A(n_1181),
.B(n_229),
.Y(n_1229)
);

INVx3_ASAP7_75t_L g1230 ( 
.A(n_1218),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1182),
.B(n_230),
.Y(n_1231)
);

INVx2_ASAP7_75t_SL g1232 ( 
.A(n_1211),
.Y(n_1232)
);

AND2x2_ASAP7_75t_L g1233 ( 
.A(n_1212),
.B(n_233),
.Y(n_1233)
);

AND2x2_ASAP7_75t_L g1234 ( 
.A(n_1197),
.B(n_236),
.Y(n_1234)
);

AOI22xp33_ASAP7_75t_L g1235 ( 
.A1(n_1177),
.A2(n_238),
.B1(n_242),
.B2(n_243),
.Y(n_1235)
);

AND2x2_ASAP7_75t_L g1236 ( 
.A(n_1193),
.B(n_1202),
.Y(n_1236)
);

AND2x2_ASAP7_75t_L g1237 ( 
.A(n_1200),
.B(n_244),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1216),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_1172),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1204),
.Y(n_1240)
);

INVx3_ASAP7_75t_L g1241 ( 
.A(n_1180),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_1178),
.B(n_246),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1174),
.Y(n_1243)
);

BUFx6f_ASAP7_75t_L g1244 ( 
.A(n_1180),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1204),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1215),
.B(n_247),
.Y(n_1246)
);

INVx2_ASAP7_75t_L g1247 ( 
.A(n_1195),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1183),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1195),
.Y(n_1249)
);

OR2x2_ASAP7_75t_L g1250 ( 
.A(n_1176),
.B(n_1203),
.Y(n_1250)
);

INVx2_ASAP7_75t_L g1251 ( 
.A(n_1184),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1189),
.B(n_248),
.Y(n_1252)
);

INVx3_ASAP7_75t_L g1253 ( 
.A(n_1184),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1190),
.Y(n_1254)
);

BUFx2_ASAP7_75t_L g1255 ( 
.A(n_1190),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1199),
.B(n_250),
.Y(n_1256)
);

AND2x2_ASAP7_75t_L g1257 ( 
.A(n_1208),
.B(n_253),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_1207),
.Y(n_1258)
);

AND2x2_ASAP7_75t_L g1259 ( 
.A(n_1225),
.B(n_255),
.Y(n_1259)
);

AND2x2_ASAP7_75t_L g1260 ( 
.A(n_1192),
.B(n_256),
.Y(n_1260)
);

AO31x2_ASAP7_75t_L g1261 ( 
.A1(n_1198),
.A2(n_264),
.A3(n_266),
.B(n_267),
.Y(n_1261)
);

OR2x2_ASAP7_75t_L g1262 ( 
.A(n_1213),
.B(n_268),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1205),
.B(n_271),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1170),
.Y(n_1264)
);

NOR2x1_ASAP7_75t_L g1265 ( 
.A(n_1222),
.B(n_272),
.Y(n_1265)
);

INVx3_ASAP7_75t_L g1266 ( 
.A(n_1175),
.Y(n_1266)
);

OR2x2_ASAP7_75t_L g1267 ( 
.A(n_1188),
.B(n_273),
.Y(n_1267)
);

INVx2_ASAP7_75t_L g1268 ( 
.A(n_1214),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1201),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1232),
.Y(n_1270)
);

OAI22xp5_ASAP7_75t_L g1271 ( 
.A1(n_1235),
.A2(n_1186),
.B1(n_1191),
.B2(n_1194),
.Y(n_1271)
);

AND2x4_ASAP7_75t_L g1272 ( 
.A(n_1230),
.B(n_1217),
.Y(n_1272)
);

HB1xp67_ASAP7_75t_L g1273 ( 
.A(n_1232),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_1236),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_1236),
.Y(n_1275)
);

HB1xp67_ASAP7_75t_L g1276 ( 
.A(n_1240),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_1230),
.Y(n_1277)
);

AND2x2_ASAP7_75t_L g1278 ( 
.A(n_1230),
.B(n_1224),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1243),
.Y(n_1279)
);

HB1xp67_ASAP7_75t_L g1280 ( 
.A(n_1245),
.Y(n_1280)
);

OA21x2_ASAP7_75t_L g1281 ( 
.A1(n_1243),
.A2(n_1221),
.B(n_1223),
.Y(n_1281)
);

AO21x2_ASAP7_75t_L g1282 ( 
.A1(n_1238),
.A2(n_1239),
.B(n_1250),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1247),
.Y(n_1283)
);

BUFx2_ASAP7_75t_L g1284 ( 
.A(n_1227),
.Y(n_1284)
);

AND2x2_ASAP7_75t_L g1285 ( 
.A(n_1239),
.B(n_1224),
.Y(n_1285)
);

INVxp67_ASAP7_75t_SL g1286 ( 
.A(n_1227),
.Y(n_1286)
);

AO21x2_ASAP7_75t_L g1287 ( 
.A1(n_1238),
.A2(n_1196),
.B(n_1206),
.Y(n_1287)
);

OAI221xp5_ASAP7_75t_L g1288 ( 
.A1(n_1264),
.A2(n_1187),
.B1(n_1185),
.B2(n_1210),
.C(n_1219),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_1247),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_1249),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1241),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1241),
.Y(n_1292)
);

OR2x2_ASAP7_75t_L g1293 ( 
.A(n_1241),
.B(n_1209),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1274),
.Y(n_1294)
);

OR2x2_ASAP7_75t_L g1295 ( 
.A(n_1274),
.B(n_1255),
.Y(n_1295)
);

INVx2_ASAP7_75t_L g1296 ( 
.A(n_1283),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1275),
.Y(n_1297)
);

OR2x2_ASAP7_75t_L g1298 ( 
.A(n_1275),
.B(n_1255),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1282),
.B(n_1248),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_1279),
.Y(n_1300)
);

HB1xp67_ASAP7_75t_L g1301 ( 
.A(n_1279),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1290),
.Y(n_1302)
);

OR2x2_ASAP7_75t_L g1303 ( 
.A(n_1283),
.B(n_1251),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1290),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1276),
.Y(n_1305)
);

OR2x2_ASAP7_75t_L g1306 ( 
.A(n_1289),
.B(n_1251),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1280),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1284),
.B(n_1266),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1273),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1282),
.B(n_1234),
.Y(n_1310)
);

INVx2_ASAP7_75t_L g1311 ( 
.A(n_1289),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1302),
.Y(n_1312)
);

INVxp67_ASAP7_75t_L g1313 ( 
.A(n_1299),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1304),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1301),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1305),
.B(n_1282),
.Y(n_1316)
);

NAND3xp33_ASAP7_75t_SL g1317 ( 
.A(n_1310),
.B(n_1210),
.C(n_1234),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_SL g1318 ( 
.A(n_1310),
.B(n_1266),
.Y(n_1318)
);

OR2x2_ASAP7_75t_L g1319 ( 
.A(n_1295),
.B(n_1270),
.Y(n_1319)
);

OR2x2_ASAP7_75t_L g1320 ( 
.A(n_1298),
.B(n_1286),
.Y(n_1320)
);

AOI21xp33_ASAP7_75t_SL g1321 ( 
.A1(n_1299),
.A2(n_1288),
.B(n_1266),
.Y(n_1321)
);

NAND2x1p5_ASAP7_75t_L g1322 ( 
.A(n_1308),
.B(n_1253),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1322),
.B(n_1309),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1321),
.B(n_1307),
.Y(n_1324)
);

OAI211xp5_ASAP7_75t_SL g1325 ( 
.A1(n_1313),
.A2(n_1228),
.B(n_1269),
.C(n_1246),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_1320),
.B(n_1293),
.Y(n_1326)
);

BUFx2_ASAP7_75t_L g1327 ( 
.A(n_1319),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1321),
.B(n_1301),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1312),
.Y(n_1329)
);

NOR2xp33_ASAP7_75t_L g1330 ( 
.A(n_1317),
.B(n_1171),
.Y(n_1330)
);

AND2x2_ASAP7_75t_L g1331 ( 
.A(n_1318),
.B(n_1293),
.Y(n_1331)
);

OR2x2_ASAP7_75t_L g1332 ( 
.A(n_1316),
.B(n_1314),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1315),
.B(n_1294),
.Y(n_1333)
);

OR2x2_ASAP7_75t_L g1334 ( 
.A(n_1320),
.B(n_1303),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1322),
.B(n_1297),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1312),
.Y(n_1336)
);

OR2x2_ASAP7_75t_L g1337 ( 
.A(n_1320),
.B(n_1306),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1329),
.Y(n_1338)
);

OAI32xp33_ASAP7_75t_L g1339 ( 
.A1(n_1324),
.A2(n_1250),
.A3(n_1285),
.B1(n_1252),
.B2(n_1271),
.Y(n_1339)
);

AOI221xp5_ASAP7_75t_L g1340 ( 
.A1(n_1330),
.A2(n_1324),
.B1(n_1325),
.B2(n_1328),
.C(n_1327),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1326),
.B(n_1285),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1328),
.B(n_1296),
.Y(n_1342)
);

OR2x2_ASAP7_75t_L g1343 ( 
.A(n_1334),
.B(n_1311),
.Y(n_1343)
);

NAND3xp33_ASAP7_75t_L g1344 ( 
.A(n_1325),
.B(n_1258),
.C(n_1259),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1336),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1333),
.Y(n_1346)
);

INVx1_ASAP7_75t_SL g1347 ( 
.A(n_1341),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1340),
.B(n_1331),
.Y(n_1348)
);

OAI22xp5_ASAP7_75t_L g1349 ( 
.A1(n_1344),
.A2(n_1337),
.B1(n_1323),
.B2(n_1278),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1338),
.Y(n_1350)
);

NOR2xp33_ASAP7_75t_L g1351 ( 
.A(n_1339),
.B(n_1335),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1345),
.Y(n_1352)
);

INVxp67_ASAP7_75t_L g1353 ( 
.A(n_1342),
.Y(n_1353)
);

NAND3xp33_ASAP7_75t_L g1354 ( 
.A(n_1348),
.B(n_1346),
.C(n_1332),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1350),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_1352),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1347),
.B(n_1343),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1353),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_1351),
.B(n_1253),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1349),
.B(n_1291),
.Y(n_1360)
);

NOR3xp33_ASAP7_75t_L g1361 ( 
.A(n_1358),
.B(n_1263),
.C(n_1262),
.Y(n_1361)
);

INVxp67_ASAP7_75t_L g1362 ( 
.A(n_1357),
.Y(n_1362)
);

INVx1_ASAP7_75t_SL g1363 ( 
.A(n_1359),
.Y(n_1363)
);

NOR3xp33_ASAP7_75t_L g1364 ( 
.A(n_1354),
.B(n_1262),
.C(n_1256),
.Y(n_1364)
);

BUFx2_ASAP7_75t_L g1365 ( 
.A(n_1356),
.Y(n_1365)
);

NAND5xp2_ASAP7_75t_L g1366 ( 
.A(n_1355),
.B(n_1360),
.C(n_1259),
.D(n_1257),
.E(n_1242),
.Y(n_1366)
);

INVx2_ASAP7_75t_SL g1367 ( 
.A(n_1356),
.Y(n_1367)
);

NAND2xp33_ASAP7_75t_L g1368 ( 
.A(n_1357),
.B(n_1265),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1357),
.Y(n_1369)
);

AOI21xp5_ASAP7_75t_L g1370 ( 
.A1(n_1368),
.A2(n_1364),
.B(n_1362),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1363),
.B(n_1292),
.Y(n_1371)
);

AOI322xp5_ASAP7_75t_L g1372 ( 
.A1(n_1369),
.A2(n_1278),
.A3(n_1258),
.B1(n_1260),
.B2(n_1272),
.C1(n_1268),
.C2(n_1257),
.Y(n_1372)
);

NAND4xp75_ASAP7_75t_L g1373 ( 
.A(n_1367),
.B(n_1260),
.C(n_1242),
.D(n_1229),
.Y(n_1373)
);

BUFx2_ASAP7_75t_R g1374 ( 
.A(n_1365),
.Y(n_1374)
);

AOI21xp5_ASAP7_75t_L g1375 ( 
.A1(n_1366),
.A2(n_1231),
.B(n_1287),
.Y(n_1375)
);

AOI22xp5_ASAP7_75t_L g1376 ( 
.A1(n_1361),
.A2(n_1287),
.B1(n_1272),
.B2(n_1254),
.Y(n_1376)
);

HB1xp67_ASAP7_75t_L g1377 ( 
.A(n_1365),
.Y(n_1377)
);

OAI22xp33_ASAP7_75t_SL g1378 ( 
.A1(n_1377),
.A2(n_1371),
.B1(n_1370),
.B2(n_1376),
.Y(n_1378)
);

AND2x2_ASAP7_75t_SL g1379 ( 
.A(n_1374),
.B(n_1372),
.Y(n_1379)
);

NOR2xp33_ASAP7_75t_SL g1380 ( 
.A(n_1373),
.B(n_1375),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1377),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1377),
.Y(n_1382)
);

OAI211xp5_ASAP7_75t_SL g1383 ( 
.A1(n_1370),
.A2(n_1267),
.B(n_1226),
.C(n_1268),
.Y(n_1383)
);

NOR2xp33_ASAP7_75t_R g1384 ( 
.A(n_1377),
.B(n_1267),
.Y(n_1384)
);

NOR2xp33_ASAP7_75t_L g1385 ( 
.A(n_1374),
.B(n_1253),
.Y(n_1385)
);

AND2x4_ASAP7_75t_L g1386 ( 
.A(n_1381),
.B(n_1300),
.Y(n_1386)
);

INVx2_ASAP7_75t_L g1387 ( 
.A(n_1382),
.Y(n_1387)
);

OR5x1_ASAP7_75t_L g1388 ( 
.A(n_1383),
.B(n_1378),
.C(n_1379),
.D(n_1380),
.E(n_1385),
.Y(n_1388)
);

BUFx2_ASAP7_75t_L g1389 ( 
.A(n_1384),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1385),
.B(n_1300),
.Y(n_1390)
);

OA22x2_ASAP7_75t_SL g1391 ( 
.A1(n_1381),
.A2(n_1277),
.B1(n_1287),
.B2(n_1261),
.Y(n_1391)
);

AOI322xp5_ASAP7_75t_L g1392 ( 
.A1(n_1379),
.A2(n_1272),
.A3(n_1229),
.B1(n_1277),
.B2(n_1233),
.C1(n_1237),
.C2(n_1261),
.Y(n_1392)
);

XNOR2x1_ASAP7_75t_L g1393 ( 
.A(n_1387),
.B(n_1226),
.Y(n_1393)
);

AND4x1_ASAP7_75t_L g1394 ( 
.A(n_1388),
.B(n_1237),
.C(n_1233),
.D(n_277),
.Y(n_1394)
);

AOI211x1_ASAP7_75t_L g1395 ( 
.A1(n_1390),
.A2(n_1261),
.B(n_276),
.C(n_280),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1389),
.B(n_1386),
.Y(n_1396)
);

INVxp67_ASAP7_75t_L g1397 ( 
.A(n_1389),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1392),
.B(n_1261),
.Y(n_1398)
);

OAI322xp33_ASAP7_75t_L g1399 ( 
.A1(n_1391),
.A2(n_1261),
.A3(n_1244),
.B1(n_1281),
.B2(n_288),
.C1(n_290),
.C2(n_294),
.Y(n_1399)
);

OAI221xp5_ASAP7_75t_L g1400 ( 
.A1(n_1397),
.A2(n_1281),
.B1(n_1244),
.B2(n_287),
.C(n_295),
.Y(n_1400)
);

OAI22xp33_ASAP7_75t_SL g1401 ( 
.A1(n_1396),
.A2(n_1281),
.B1(n_285),
.B2(n_299),
.Y(n_1401)
);

O2A1O1Ixp33_ASAP7_75t_L g1402 ( 
.A1(n_1399),
.A2(n_275),
.B(n_300),
.C(n_302),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1400),
.Y(n_1403)
);

OAI21x1_ASAP7_75t_L g1404 ( 
.A1(n_1402),
.A2(n_1398),
.B(n_1394),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1401),
.Y(n_1405)
);

INVxp67_ASAP7_75t_L g1406 ( 
.A(n_1404),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1405),
.Y(n_1407)
);

OR2x6_ASAP7_75t_L g1408 ( 
.A(n_1407),
.B(n_1403),
.Y(n_1408)
);

BUFx2_ASAP7_75t_L g1409 ( 
.A(n_1406),
.Y(n_1409)
);

AOI21xp5_ASAP7_75t_L g1410 ( 
.A1(n_1409),
.A2(n_1408),
.B(n_1403),
.Y(n_1410)
);

AOI221xp5_ASAP7_75t_L g1411 ( 
.A1(n_1409),
.A2(n_1395),
.B1(n_1393),
.B2(n_1244),
.C(n_311),
.Y(n_1411)
);

AOI21xp33_ASAP7_75t_L g1412 ( 
.A1(n_1410),
.A2(n_303),
.B(n_305),
.Y(n_1412)
);

AOI322xp5_ASAP7_75t_L g1413 ( 
.A1(n_1412),
.A2(n_1411),
.A3(n_1244),
.B1(n_313),
.B2(n_317),
.C1(n_319),
.C2(n_323),
.Y(n_1413)
);

AOI221xp5_ASAP7_75t_L g1414 ( 
.A1(n_1413),
.A2(n_1244),
.B1(n_312),
.B2(n_324),
.C(n_325),
.Y(n_1414)
);

AOI211xp5_ASAP7_75t_L g1415 ( 
.A1(n_1414),
.A2(n_309),
.B(n_328),
.C(n_329),
.Y(n_1415)
);


endmodule