module fake_ibex_1734_n_6478 (n_151, n_1084, n_85, n_599, n_778, n_822, n_1042, n_507, n_743, n_1060, n_540, n_754, n_395, n_1104, n_1011, n_84, n_64, n_992, n_171, n_756, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_766, n_1041, n_688, n_130, n_1090, n_177, n_1110, n_946, n_707, n_76, n_273, n_309, n_330, n_926, n_1097, n_9, n_1079, n_1031, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_845, n_947, n_972, n_981, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_956, n_790, n_920, n_452, n_86, n_70, n_664, n_1067, n_255, n_175, n_586, n_773, n_994, n_638, n_398, n_59, n_28, n_125, n_304, n_821, n_191, n_873, n_962, n_593, n_5, n_62, n_71, n_153, n_862, n_545, n_909, n_583, n_887, n_1080, n_957, n_1015, n_678, n_663, n_969, n_194, n_249, n_334, n_634, n_733, n_961, n_991, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_1034, n_371, n_974, n_1036, n_403, n_872, n_423, n_608, n_864, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_930, n_336, n_959, n_258, n_861, n_1018, n_1044, n_1106, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_727, n_58, n_1077, n_43, n_216, n_996, n_915, n_911, n_33, n_652, n_781, n_421, n_828, n_738, n_475, n_802, n_166, n_163, n_1045, n_753, n_645, n_500, n_747, n_963, n_542, n_114, n_236, n_900, n_34, n_376, n_1098, n_377, n_584, n_531, n_647, n_15, n_761, n_556, n_748, n_24, n_189, n_498, n_698, n_280, n_317, n_340, n_375, n_708, n_901, n_1096, n_105, n_187, n_667, n_884, n_1061, n_1, n_154, n_682, n_850, n_182, n_196, n_326, n_327, n_879, n_89, n_1056, n_50, n_723, n_144, n_170, n_270, n_346, n_383, n_113, n_886, n_840, n_1010, n_561, n_883, n_117, n_417, n_471, n_846, n_739, n_755, n_265, n_853, n_504, n_948, n_158, n_1029, n_859, n_259, n_276, n_339, n_470, n_770, n_965, n_210, n_348, n_1109, n_220, n_875, n_941, n_674, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_671, n_228, n_711, n_876, n_147, n_552, n_251, n_384, n_632, n_989, n_373, n_1051, n_854, n_1008, n_458, n_244, n_73, n_1053, n_1112, n_343, n_310, n_714, n_1076, n_1032, n_936, n_703, n_426, n_323, n_469, n_829, n_1099, n_598, n_825, n_143, n_740, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_939, n_67, n_453, n_591, n_898, n_655, n_333, n_928, n_967, n_110, n_306, n_400, n_47, n_550, n_736, n_169, n_1055, n_10, n_673, n_21, n_732, n_798, n_832, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_641, n_7, n_109, n_127, n_1103, n_121, n_527, n_893, n_590, n_1025, n_465, n_1057, n_1068, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_690, n_914, n_120, n_1013, n_982, n_835, n_168, n_526, n_785, n_155, n_824, n_929, n_315, n_441, n_604, n_1024, n_13, n_637, n_122, n_523, n_116, n_694, n_787, n_977, n_1075, n_614, n_370, n_431, n_719, n_574, n_0, n_289, n_716, n_865, n_923, n_12, n_515, n_642, n_150, n_286, n_321, n_133, n_569, n_600, n_907, n_51, n_933, n_1081, n_215, n_279, n_49, n_1037, n_374, n_235, n_464, n_538, n_669, n_838, n_987, n_750, n_1021, n_746, n_22, n_136, n_261, n_742, n_521, n_665, n_459, n_30, n_1101, n_518, n_367, n_221, n_1052, n_852, n_789, n_880, n_654, n_1083, n_656, n_1014, n_724, n_437, n_731, n_602, n_904, n_842, n_938, n_355, n_767, n_474, n_878, n_758, n_594, n_636, n_710, n_720, n_407, n_102, n_490, n_1023, n_568, n_813, n_52, n_448, n_646, n_595, n_99, n_466, n_269, n_944, n_1001, n_156, n_570, n_126, n_623, n_585, n_1030, n_1094, n_715, n_791, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_769, n_1082, n_222, n_660, n_186, n_524, n_349, n_765, n_849, n_857, n_980, n_454, n_1070, n_1074, n_777, n_1017, n_295, n_730, n_331, n_576, n_230, n_96, n_759, n_917, n_185, n_388, n_953, n_625, n_968, n_619, n_1089, n_536, n_611, n_352, n_290, n_558, n_931, n_666, n_174, n_467, n_427, n_607, n_827, n_157, n_219, n_246, n_31, n_442, n_146, n_1064, n_1071, n_207, n_922, n_438, n_851, n_993, n_1012, n_1028, n_689, n_960, n_1022, n_793, n_167, n_676, n_128, n_937, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_973, n_358, n_771, n_205, n_618, n_488, n_139, n_514, n_705, n_999, n_1038, n_1092, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_659, n_267, n_662, n_910, n_1009, n_635, n_979, n_844, n_1066, n_245, n_589, n_571, n_229, n_209, n_472, n_648, n_783, n_347, n_1020, n_847, n_830, n_1062, n_1004, n_473, n_1027, n_445, n_629, n_335, n_413, n_1072, n_82, n_263, n_1069, n_27, n_573, n_353, n_966, n_359, n_826, n_299, n_87, n_262, n_433, n_75, n_439, n_704, n_949, n_1007, n_924, n_643, n_137, n_679, n_841, n_772, n_810, n_768, n_839, n_338, n_173, n_696, n_796, n_797, n_837, n_477, n_640, n_954, n_363, n_1006, n_402, n_725, n_180, n_369, n_976, n_596, n_201, n_699, n_14, n_1063, n_351, n_368, n_456, n_834, n_257, n_77, n_998, n_935, n_869, n_1115, n_925, n_718, n_801, n_918, n_1054, n_44, n_672, n_1100, n_1039, n_722, n_401, n_1046, n_553, n_554, n_1078, n_1043, n_66, n_735, n_305, n_882, n_942, n_713, n_307, n_192, n_804, n_140, n_484, n_566, n_480, n_416, n_581, n_651, n_365, n_721, n_4, n_814, n_955, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_630, n_516, n_548, n_567, n_943, n_1049, n_1086, n_763, n_745, n_329, n_447, n_940, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_868, n_546, n_199, n_788, n_795, n_1065, n_592, n_986, n_495, n_762, n_410, n_905, n_308, n_975, n_675, n_800, n_463, n_624, n_706, n_411, n_135, n_520, n_784, n_684, n_775, n_927, n_934, n_658, n_512, n_615, n_950, n_685, n_1026, n_283, n_366, n_397, n_111, n_803, n_894, n_1033, n_692, n_36, n_627, n_990, n_18, n_709, n_322, n_53, n_227, n_499, n_115, n_888, n_1087, n_757, n_11, n_248, n_92, n_702, n_451, n_712, n_971, n_101, n_190, n_906, n_138, n_650, n_776, n_1114, n_409, n_1093, n_582, n_978, n_818, n_653, n_214, n_238, n_579, n_843, n_899, n_1019, n_1059, n_902, n_332, n_799, n_517, n_211, n_744, n_817, n_218, n_314, n_691, n_563, n_132, n_277, n_555, n_337, n_522, n_700, n_479, n_534, n_225, n_360, n_881, n_272, n_951, n_511, n_23, n_734, n_468, n_1107, n_223, n_381, n_1073, n_1108, n_525, n_815, n_919, n_780, n_535, n_1002, n_382, n_502, n_681, n_633, n_1111, n_532, n_726, n_95, n_405, n_863, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_819, n_161, n_237, n_29, n_203, n_268, n_440, n_858, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_729, n_741, n_603, n_378, n_486, n_952, n_422, n_164, n_38, n_198, n_264, n_616, n_782, n_997, n_833, n_217, n_324, n_391, n_831, n_537, n_1113, n_728, n_78, n_805, n_670, n_820, n_20, n_69, n_892, n_390, n_544, n_891, n_913, n_39, n_178, n_509, n_695, n_786, n_639, n_303, n_362, n_717, n_93, n_505, n_162, n_482, n_240, n_1016, n_282, n_61, n_680, n_501, n_809, n_752, n_856, n_668, n_779, n_871, n_266, n_42, n_294, n_112, n_958, n_485, n_870, n_46, n_284, n_811, n_1047, n_808, n_80, n_172, n_250, n_945, n_493, n_460, n_609, n_1040, n_476, n_792, n_461, n_575, n_313, n_903, n_519, n_345, n_408, n_119, n_1085, n_361, n_1095, n_455, n_419, n_774, n_72, n_1048, n_319, n_1091, n_195, n_885, n_513, n_212, n_588, n_877, n_693, n_311, n_860, n_661, n_848, n_406, n_606, n_737, n_1088, n_896, n_97, n_197, n_528, n_181, n_1005, n_131, n_123, n_1102, n_631, n_683, n_260, n_620, n_794, n_836, n_462, n_302, n_450, n_443, n_686, n_985, n_572, n_867, n_983, n_1003, n_644, n_577, n_344, n_393, n_889, n_897, n_436, n_428, n_970, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_697, n_816, n_874, n_890, n_912, n_921, n_83, n_32, n_1058, n_1105, n_107, n_149, n_489, n_677, n_399, n_254, n_908, n_213, n_964, n_424, n_565, n_916, n_823, n_701, n_271, n_995, n_241, n_68, n_503, n_292, n_807, n_984, n_394, n_79, n_1000, n_81, n_35, n_364, n_687, n_895, n_988, n_159, n_202, n_231, n_298, n_587, n_1035, n_760, n_751, n_806, n_932, n_160, n_657, n_764, n_184, n_56, n_492, n_649, n_812, n_855, n_232, n_380, n_749, n_281, n_866, n_559, n_425, n_1050, n_6478);

input n_151;
input n_1084;
input n_85;
input n_599;
input n_778;
input n_822;
input n_1042;
input n_507;
input n_743;
input n_1060;
input n_540;
input n_754;
input n_395;
input n_1104;
input n_1011;
input n_84;
input n_64;
input n_992;
input n_171;
input n_756;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_766;
input n_1041;
input n_688;
input n_130;
input n_1090;
input n_177;
input n_1110;
input n_946;
input n_707;
input n_76;
input n_273;
input n_309;
input n_330;
input n_926;
input n_1097;
input n_9;
input n_1079;
input n_1031;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_845;
input n_947;
input n_972;
input n_981;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_956;
input n_790;
input n_920;
input n_452;
input n_86;
input n_70;
input n_664;
input n_1067;
input n_255;
input n_175;
input n_586;
input n_773;
input n_994;
input n_638;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_821;
input n_191;
input n_873;
input n_962;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_862;
input n_545;
input n_909;
input n_583;
input n_887;
input n_1080;
input n_957;
input n_1015;
input n_678;
input n_663;
input n_969;
input n_194;
input n_249;
input n_334;
input n_634;
input n_733;
input n_961;
input n_991;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_1034;
input n_371;
input n_974;
input n_1036;
input n_403;
input n_872;
input n_423;
input n_608;
input n_864;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_930;
input n_336;
input n_959;
input n_258;
input n_861;
input n_1018;
input n_1044;
input n_1106;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_727;
input n_58;
input n_1077;
input n_43;
input n_216;
input n_996;
input n_915;
input n_911;
input n_33;
input n_652;
input n_781;
input n_421;
input n_828;
input n_738;
input n_475;
input n_802;
input n_166;
input n_163;
input n_1045;
input n_753;
input n_645;
input n_500;
input n_747;
input n_963;
input n_542;
input n_114;
input n_236;
input n_900;
input n_34;
input n_376;
input n_1098;
input n_377;
input n_584;
input n_531;
input n_647;
input n_15;
input n_761;
input n_556;
input n_748;
input n_24;
input n_189;
input n_498;
input n_698;
input n_280;
input n_317;
input n_340;
input n_375;
input n_708;
input n_901;
input n_1096;
input n_105;
input n_187;
input n_667;
input n_884;
input n_1061;
input n_1;
input n_154;
input n_682;
input n_850;
input n_182;
input n_196;
input n_326;
input n_327;
input n_879;
input n_89;
input n_1056;
input n_50;
input n_723;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_886;
input n_840;
input n_1010;
input n_561;
input n_883;
input n_117;
input n_417;
input n_471;
input n_846;
input n_739;
input n_755;
input n_265;
input n_853;
input n_504;
input n_948;
input n_158;
input n_1029;
input n_859;
input n_259;
input n_276;
input n_339;
input n_470;
input n_770;
input n_965;
input n_210;
input n_348;
input n_1109;
input n_220;
input n_875;
input n_941;
input n_674;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_671;
input n_228;
input n_711;
input n_876;
input n_147;
input n_552;
input n_251;
input n_384;
input n_632;
input n_989;
input n_373;
input n_1051;
input n_854;
input n_1008;
input n_458;
input n_244;
input n_73;
input n_1053;
input n_1112;
input n_343;
input n_310;
input n_714;
input n_1076;
input n_1032;
input n_936;
input n_703;
input n_426;
input n_323;
input n_469;
input n_829;
input n_1099;
input n_598;
input n_825;
input n_143;
input n_740;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_939;
input n_67;
input n_453;
input n_591;
input n_898;
input n_655;
input n_333;
input n_928;
input n_967;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_736;
input n_169;
input n_1055;
input n_10;
input n_673;
input n_21;
input n_732;
input n_798;
input n_832;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_641;
input n_7;
input n_109;
input n_127;
input n_1103;
input n_121;
input n_527;
input n_893;
input n_590;
input n_1025;
input n_465;
input n_1057;
input n_1068;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_690;
input n_914;
input n_120;
input n_1013;
input n_982;
input n_835;
input n_168;
input n_526;
input n_785;
input n_155;
input n_824;
input n_929;
input n_315;
input n_441;
input n_604;
input n_1024;
input n_13;
input n_637;
input n_122;
input n_523;
input n_116;
input n_694;
input n_787;
input n_977;
input n_1075;
input n_614;
input n_370;
input n_431;
input n_719;
input n_574;
input n_0;
input n_289;
input n_716;
input n_865;
input n_923;
input n_12;
input n_515;
input n_642;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_907;
input n_51;
input n_933;
input n_1081;
input n_215;
input n_279;
input n_49;
input n_1037;
input n_374;
input n_235;
input n_464;
input n_538;
input n_669;
input n_838;
input n_987;
input n_750;
input n_1021;
input n_746;
input n_22;
input n_136;
input n_261;
input n_742;
input n_521;
input n_665;
input n_459;
input n_30;
input n_1101;
input n_518;
input n_367;
input n_221;
input n_1052;
input n_852;
input n_789;
input n_880;
input n_654;
input n_1083;
input n_656;
input n_1014;
input n_724;
input n_437;
input n_731;
input n_602;
input n_904;
input n_842;
input n_938;
input n_355;
input n_767;
input n_474;
input n_878;
input n_758;
input n_594;
input n_636;
input n_710;
input n_720;
input n_407;
input n_102;
input n_490;
input n_1023;
input n_568;
input n_813;
input n_52;
input n_448;
input n_646;
input n_595;
input n_99;
input n_466;
input n_269;
input n_944;
input n_1001;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_1030;
input n_1094;
input n_715;
input n_791;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_769;
input n_1082;
input n_222;
input n_660;
input n_186;
input n_524;
input n_349;
input n_765;
input n_849;
input n_857;
input n_980;
input n_454;
input n_1070;
input n_1074;
input n_777;
input n_1017;
input n_295;
input n_730;
input n_331;
input n_576;
input n_230;
input n_96;
input n_759;
input n_917;
input n_185;
input n_388;
input n_953;
input n_625;
input n_968;
input n_619;
input n_1089;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_931;
input n_666;
input n_174;
input n_467;
input n_427;
input n_607;
input n_827;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_1064;
input n_1071;
input n_207;
input n_922;
input n_438;
input n_851;
input n_993;
input n_1012;
input n_1028;
input n_689;
input n_960;
input n_1022;
input n_793;
input n_167;
input n_676;
input n_128;
input n_937;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_973;
input n_358;
input n_771;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_705;
input n_999;
input n_1038;
input n_1092;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_659;
input n_267;
input n_662;
input n_910;
input n_1009;
input n_635;
input n_979;
input n_844;
input n_1066;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_648;
input n_783;
input n_347;
input n_1020;
input n_847;
input n_830;
input n_1062;
input n_1004;
input n_473;
input n_1027;
input n_445;
input n_629;
input n_335;
input n_413;
input n_1072;
input n_82;
input n_263;
input n_1069;
input n_27;
input n_573;
input n_353;
input n_966;
input n_359;
input n_826;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_704;
input n_949;
input n_1007;
input n_924;
input n_643;
input n_137;
input n_679;
input n_841;
input n_772;
input n_810;
input n_768;
input n_839;
input n_338;
input n_173;
input n_696;
input n_796;
input n_797;
input n_837;
input n_477;
input n_640;
input n_954;
input n_363;
input n_1006;
input n_402;
input n_725;
input n_180;
input n_369;
input n_976;
input n_596;
input n_201;
input n_699;
input n_14;
input n_1063;
input n_351;
input n_368;
input n_456;
input n_834;
input n_257;
input n_77;
input n_998;
input n_935;
input n_869;
input n_1115;
input n_925;
input n_718;
input n_801;
input n_918;
input n_1054;
input n_44;
input n_672;
input n_1100;
input n_1039;
input n_722;
input n_401;
input n_1046;
input n_553;
input n_554;
input n_1078;
input n_1043;
input n_66;
input n_735;
input n_305;
input n_882;
input n_942;
input n_713;
input n_307;
input n_192;
input n_804;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_651;
input n_365;
input n_721;
input n_4;
input n_814;
input n_955;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_630;
input n_516;
input n_548;
input n_567;
input n_943;
input n_1049;
input n_1086;
input n_763;
input n_745;
input n_329;
input n_447;
input n_940;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_868;
input n_546;
input n_199;
input n_788;
input n_795;
input n_1065;
input n_592;
input n_986;
input n_495;
input n_762;
input n_410;
input n_905;
input n_308;
input n_975;
input n_675;
input n_800;
input n_463;
input n_624;
input n_706;
input n_411;
input n_135;
input n_520;
input n_784;
input n_684;
input n_775;
input n_927;
input n_934;
input n_658;
input n_512;
input n_615;
input n_950;
input n_685;
input n_1026;
input n_283;
input n_366;
input n_397;
input n_111;
input n_803;
input n_894;
input n_1033;
input n_692;
input n_36;
input n_627;
input n_990;
input n_18;
input n_709;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_888;
input n_1087;
input n_757;
input n_11;
input n_248;
input n_92;
input n_702;
input n_451;
input n_712;
input n_971;
input n_101;
input n_190;
input n_906;
input n_138;
input n_650;
input n_776;
input n_1114;
input n_409;
input n_1093;
input n_582;
input n_978;
input n_818;
input n_653;
input n_214;
input n_238;
input n_579;
input n_843;
input n_899;
input n_1019;
input n_1059;
input n_902;
input n_332;
input n_799;
input n_517;
input n_211;
input n_744;
input n_817;
input n_218;
input n_314;
input n_691;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_700;
input n_479;
input n_534;
input n_225;
input n_360;
input n_881;
input n_272;
input n_951;
input n_511;
input n_23;
input n_734;
input n_468;
input n_1107;
input n_223;
input n_381;
input n_1073;
input n_1108;
input n_525;
input n_815;
input n_919;
input n_780;
input n_535;
input n_1002;
input n_382;
input n_502;
input n_681;
input n_633;
input n_1111;
input n_532;
input n_726;
input n_95;
input n_405;
input n_863;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_819;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_858;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_729;
input n_741;
input n_603;
input n_378;
input n_486;
input n_952;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_782;
input n_997;
input n_833;
input n_217;
input n_324;
input n_391;
input n_831;
input n_537;
input n_1113;
input n_728;
input n_78;
input n_805;
input n_670;
input n_820;
input n_20;
input n_69;
input n_892;
input n_390;
input n_544;
input n_891;
input n_913;
input n_39;
input n_178;
input n_509;
input n_695;
input n_786;
input n_639;
input n_303;
input n_362;
input n_717;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_1016;
input n_282;
input n_61;
input n_680;
input n_501;
input n_809;
input n_752;
input n_856;
input n_668;
input n_779;
input n_871;
input n_266;
input n_42;
input n_294;
input n_112;
input n_958;
input n_485;
input n_870;
input n_46;
input n_284;
input n_811;
input n_1047;
input n_808;
input n_80;
input n_172;
input n_250;
input n_945;
input n_493;
input n_460;
input n_609;
input n_1040;
input n_476;
input n_792;
input n_461;
input n_575;
input n_313;
input n_903;
input n_519;
input n_345;
input n_408;
input n_119;
input n_1085;
input n_361;
input n_1095;
input n_455;
input n_419;
input n_774;
input n_72;
input n_1048;
input n_319;
input n_1091;
input n_195;
input n_885;
input n_513;
input n_212;
input n_588;
input n_877;
input n_693;
input n_311;
input n_860;
input n_661;
input n_848;
input n_406;
input n_606;
input n_737;
input n_1088;
input n_896;
input n_97;
input n_197;
input n_528;
input n_181;
input n_1005;
input n_131;
input n_123;
input n_1102;
input n_631;
input n_683;
input n_260;
input n_620;
input n_794;
input n_836;
input n_462;
input n_302;
input n_450;
input n_443;
input n_686;
input n_985;
input n_572;
input n_867;
input n_983;
input n_1003;
input n_644;
input n_577;
input n_344;
input n_393;
input n_889;
input n_897;
input n_436;
input n_428;
input n_970;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_697;
input n_816;
input n_874;
input n_890;
input n_912;
input n_921;
input n_83;
input n_32;
input n_1058;
input n_1105;
input n_107;
input n_149;
input n_489;
input n_677;
input n_399;
input n_254;
input n_908;
input n_213;
input n_964;
input n_424;
input n_565;
input n_916;
input n_823;
input n_701;
input n_271;
input n_995;
input n_241;
input n_68;
input n_503;
input n_292;
input n_807;
input n_984;
input n_394;
input n_79;
input n_1000;
input n_81;
input n_35;
input n_364;
input n_687;
input n_895;
input n_988;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_1035;
input n_760;
input n_751;
input n_806;
input n_932;
input n_160;
input n_657;
input n_764;
input n_184;
input n_56;
input n_492;
input n_649;
input n_812;
input n_855;
input n_232;
input n_380;
input n_749;
input n_281;
input n_866;
input n_559;
input n_425;
input n_1050;

output n_6478;

wire n_4557;
wire n_6210;
wire n_5285;
wire n_3590;
wire n_4056;
wire n_2960;
wire n_4983;
wire n_3548;
wire n_5647;
wire n_1382;
wire n_2949;
wire n_2840;
wire n_3319;
wire n_3915;
wire n_5002;
wire n_5155;
wire n_5130;
wire n_4204;
wire n_5899;
wire n_6259;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_1802;
wire n_3817;
wire n_2038;
wire n_2504;
wire n_4607;
wire n_4514;
wire n_3674;
wire n_4249;
wire n_4931;
wire n_1859;
wire n_5827;
wire n_4805;
wire n_1765;
wire n_2392;
wire n_5008;
wire n_6183;
wire n_3280;
wire n_4371;
wire n_4601;
wire n_6035;
wire n_5858;
wire n_5879;
wire n_3458;
wire n_3519;
wire n_2276;
wire n_1782;
wire n_2889;
wire n_2391;
wire n_4585;
wire n_1391;
wire n_3338;
wire n_3168;
wire n_2396;
wire n_3440;
wire n_4169;
wire n_3570;
wire n_5760;
wire n_4875;
wire n_1957;
wire n_4197;
wire n_2188;
wire n_1144;
wire n_2506;
wire n_6229;
wire n_3598;
wire n_1752;
wire n_4172;
wire n_1730;
wire n_5243;
wire n_3479;
wire n_5587;
wire n_3751;
wire n_3262;
wire n_4673;
wire n_3537;
wire n_5667;
wire n_2343;
wire n_5615;
wire n_1480;
wire n_6327;
wire n_1463;
wire n_1823;
wire n_4781;
wire n_6256;
wire n_4423;
wire n_5517;
wire n_1766;
wire n_4065;
wire n_3469;
wire n_3170;
wire n_1922;
wire n_5962;
wire n_3347;
wire n_3395;
wire n_4808;
wire n_4507;
wire n_3577;
wire n_2995;
wire n_4526;
wire n_6286;
wire n_3472;
wire n_5922;
wire n_1981;
wire n_3976;
wire n_4348;
wire n_5931;
wire n_3807;
wire n_2998;
wire n_3845;
wire n_2163;
wire n_4450;
wire n_4467;
wire n_6159;
wire n_4801;
wire n_6005;
wire n_3639;
wire n_5809;
wire n_1664;
wire n_4144;
wire n_3298;
wire n_1427;
wire n_4447;
wire n_4955;
wire n_3208;
wire n_5588;
wire n_4569;
wire n_5404;
wire n_3671;
wire n_1778;
wire n_2839;
wire n_4998;
wire n_1698;
wire n_1496;
wire n_2333;
wire n_2705;
wire n_5505;
wire n_1214;
wire n_1274;
wire n_1595;
wire n_4510;
wire n_5658;
wire n_4567;
wire n_5151;
wire n_2362;
wire n_5478;
wire n_2822;
wire n_1306;
wire n_5994;
wire n_1493;
wire n_2597;
wire n_2774;
wire n_3681;
wire n_2753;
wire n_3603;
wire n_5037;
wire n_5878;
wire n_5716;
wire n_1960;
wire n_3979;
wire n_3714;
wire n_2844;
wire n_6192;
wire n_3565;
wire n_5304;
wire n_3883;
wire n_5866;
wire n_5941;
wire n_3943;
wire n_4563;
wire n_1309;
wire n_5882;
wire n_1316;
wire n_1562;
wire n_6102;
wire n_4854;
wire n_3769;
wire n_6456;
wire n_1445;
wire n_6026;
wire n_2147;
wire n_5591;
wire n_6083;
wire n_2253;
wire n_4479;
wire n_5381;
wire n_3858;
wire n_4173;
wire n_5261;
wire n_5895;
wire n_5944;
wire n_6328;
wire n_5673;
wire n_4422;
wire n_5743;
wire n_1865;
wire n_5033;
wire n_4842;
wire n_4786;
wire n_1170;
wire n_3842;
wire n_2980;
wire n_6219;
wire n_5075;
wire n_1322;
wire n_4457;
wire n_4060;
wire n_6241;
wire n_1305;
wire n_2088;
wire n_1248;
wire n_2171;
wire n_3307;
wire n_1388;
wire n_3780;
wire n_5571;
wire n_1653;
wire n_1375;
wire n_6254;
wire n_1118;
wire n_6066;
wire n_1881;
wire n_3798;
wire n_4809;
wire n_5241;
wire n_3060;
wire n_5129;
wire n_4124;
wire n_4499;
wire n_1350;
wire n_3627;
wire n_5191;
wire n_2957;
wire n_2586;
wire n_3958;
wire n_2412;
wire n_2783;
wire n_5259;
wire n_3293;
wire n_2550;
wire n_5913;
wire n_6302;
wire n_5266;
wire n_3381;
wire n_2750;
wire n_1650;
wire n_1453;
wire n_5580;
wire n_6078;
wire n_1423;
wire n_3836;
wire n_1239;
wire n_4714;
wire n_5660;
wire n_5955;
wire n_1209;
wire n_5419;
wire n_3732;
wire n_6070;
wire n_3295;
wire n_3199;
wire n_1616;
wire n_2389;
wire n_5612;
wire n_6408;
wire n_2107;
wire n_3435;
wire n_4828;
wire n_4480;
wire n_1613;
wire n_3874;
wire n_2782;
wire n_4258;
wire n_1549;
wire n_4290;
wire n_1531;
wire n_2919;
wire n_6019;
wire n_4577;
wire n_1424;
wire n_2625;
wire n_2444;
wire n_3652;
wire n_4913;
wire n_2199;
wire n_1610;
wire n_4398;
wire n_1298;
wire n_1844;
wire n_4055;
wire n_3194;
wire n_4692;
wire n_5987;
wire n_6421;
wire n_6009;
wire n_2431;
wire n_2084;
wire n_1243;
wire n_3572;
wire n_6114;
wire n_1121;
wire n_4823;
wire n_5195;
wire n_5541;
wire n_6081;
wire n_3951;
wire n_4927;
wire n_3355;
wire n_2019;
wire n_1407;
wire n_4680;
wire n_1821;
wire n_5609;
wire n_5904;
wire n_4757;
wire n_5254;
wire n_6334;
wire n_3698;
wire n_2731;
wire n_4451;
wire n_5423;
wire n_4653;
wire n_3466;
wire n_3370;
wire n_1504;
wire n_1781;
wire n_4331;
wire n_2028;
wire n_3678;
wire n_4216;
wire n_2856;
wire n_1921;
wire n_5732;
wire n_5141;
wire n_1293;
wire n_3968;
wire n_4825;
wire n_6178;
wire n_3950;
wire n_5252;
wire n_6209;
wire n_1319;
wire n_4376;
wire n_4050;
wire n_4623;
wire n_4523;
wire n_4411;
wire n_3811;
wire n_1271;
wire n_6011;
wire n_3416;
wire n_3147;
wire n_3983;
wire n_3628;
wire n_2425;
wire n_2800;
wire n_4225;
wire n_5238;
wire n_3859;
wire n_4489;
wire n_3455;
wire n_1591;
wire n_2289;
wire n_2841;
wire n_4271;
wire n_1409;
wire n_2744;
wire n_3524;
wire n_6085;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_4404;
wire n_1521;
wire n_5502;
wire n_3054;
wire n_2456;
wire n_2924;
wire n_5288;
wire n_2264;
wire n_1987;
wire n_5749;
wire n_1129;
wire n_1244;
wire n_3365;
wire n_4974;
wire n_4725;
wire n_6431;
wire n_1932;
wire n_3775;
wire n_6196;
wire n_3741;
wire n_3854;
wire n_1217;
wire n_4658;
wire n_2655;
wire n_3487;
wire n_1715;
wire n_6377;
wire n_3300;
wire n_5920;
wire n_5969;
wire n_1713;
wire n_3621;
wire n_2036;
wire n_1255;
wire n_2740;
wire n_2622;
wire n_4250;
wire n_1218;
wire n_4572;
wire n_5705;
wire n_4374;
wire n_6146;
wire n_3708;
wire n_2626;
wire n_1446;
wire n_3218;
wire n_2880;
wire n_5887;
wire n_5948;
wire n_2423;
wire n_3849;
wire n_3490;
wire n_3055;
wire n_1633;
wire n_4469;
wire n_2580;
wire n_3222;
wire n_3529;
wire n_6124;
wire n_3352;
wire n_4180;
wire n_2964;
wire n_4062;
wire n_1498;
wire n_5199;
wire n_1207;
wire n_1735;
wire n_3813;
wire n_1825;
wire n_4232;
wire n_4199;
wire n_6061;
wire n_5099;
wire n_1210;
wire n_6136;
wire n_4033;
wire n_2522;
wire n_4608;
wire n_1201;
wire n_5859;
wire n_1246;
wire n_5258;
wire n_4231;
wire n_6187;
wire n_1724;
wire n_2838;
wire n_1540;
wire n_3243;
wire n_3214;
wire n_1890;
wire n_3128;
wire n_4073;
wire n_6402;
wire n_2549;
wire n_4325;
wire n_2440;
wire n_4113;
wire n_1440;
wire n_4646;
wire n_6305;
wire n_1751;
wire n_2146;
wire n_2341;
wire n_1737;
wire n_4819;
wire n_4261;
wire n_4884;
wire n_3205;
wire n_4490;
wire n_2358;
wire n_6128;
wire n_2361;
wire n_4128;
wire n_5213;
wire n_6469;
wire n_5354;
wire n_2062;
wire n_3932;
wire n_2339;
wire n_1963;
wire n_1418;
wire n_1137;
wire n_2552;
wire n_2590;
wire n_3119;
wire n_1977;
wire n_3345;
wire n_4114;
wire n_1776;
wire n_6113;
wire n_3544;
wire n_5049;
wire n_1279;
wire n_4209;
wire n_3692;
wire n_5163;
wire n_1408;
wire n_5707;
wire n_3913;
wire n_3535;
wire n_2287;
wire n_3597;
wire n_4190;
wire n_2954;
wire n_6379;
wire n_2046;
wire n_6454;
wire n_4443;
wire n_4151;
wire n_4625;
wire n_4170;
wire n_4424;
wire n_1465;
wire n_6071;
wire n_4674;
wire n_6450;
wire n_1232;
wire n_2715;
wire n_6270;
wire n_4679;
wire n_6065;
wire n_1345;
wire n_4456;
wire n_5574;
wire n_1590;
wire n_2133;
wire n_3553;
wire n_5081;
wire n_6332;
wire n_6345;
wire n_1471;
wire n_3441;
wire n_5385;
wire n_4559;
wire n_5336;
wire n_2551;
wire n_4641;
wire n_4064;
wire n_5668;
wire n_4110;
wire n_4379;
wire n_3397;
wire n_5310;
wire n_4145;
wire n_1627;
wire n_3880;
wire n_5192;
wire n_4664;
wire n_3829;
wire n_1864;
wire n_5206;
wire n_2010;
wire n_2733;
wire n_6120;
wire n_3796;
wire n_5719;
wire n_5157;
wire n_1836;
wire n_6384;
wire n_4753;
wire n_1420;
wire n_2651;
wire n_1699;
wire n_4894;
wire n_5892;
wire n_5216;
wire n_4115;
wire n_2905;
wire n_3460;
wire n_3978;
wire n_3954;
wire n_4321;
wire n_5375;
wire n_2418;
wire n_1599;
wire n_3070;
wire n_3477;
wire n_1575;
wire n_4416;
wire n_5998;
wire n_4024;
wire n_5521;
wire n_3975;
wire n_3164;
wire n_6314;
wire n_1448;
wire n_3034;
wire n_5433;
wire n_2628;
wire n_4361;
wire n_1705;
wire n_4237;
wire n_2263;
wire n_3495;
wire n_3169;
wire n_6349;
wire n_3759;
wire n_4777;
wire n_4800;
wire n_3629;
wire n_5573;
wire n_5620;
wire n_4117;
wire n_2884;
wire n_3383;
wire n_3687;
wire n_4154;
wire n_3459;
wire n_6105;
wire n_2691;
wire n_2243;
wire n_3092;
wire n_5330;
wire n_4385;
wire n_2759;
wire n_3434;
wire n_2654;
wire n_5729;
wire n_2975;
wire n_2503;
wire n_4072;
wire n_1512;
wire n_4908;
wire n_3885;
wire n_1426;
wire n_2365;
wire n_2245;
wire n_3877;
wire n_5083;
wire n_3260;
wire n_6463;
wire n_2776;
wire n_2630;
wire n_6348;
wire n_1967;
wire n_5801;
wire n_3834;
wire n_5579;
wire n_1378;
wire n_3257;
wire n_2459;
wire n_2439;
wire n_1430;
wire n_5365;
wire n_2450;
wire n_6459;
wire n_4195;
wire n_1475;
wire n_3337;
wire n_5263;
wire n_4851;
wire n_4963;
wire n_1122;
wire n_3387;
wire n_6126;
wire n_4495;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_1514;
wire n_2728;
wire n_4685;
wire n_6115;
wire n_3428;
wire n_5959;
wire n_6282;
wire n_2427;
wire n_5017;
wire n_1127;
wire n_5938;
wire n_1845;
wire n_3835;
wire n_3723;
wire n_3389;
wire n_5292;
wire n_2422;
wire n_6277;
wire n_5190;
wire n_1679;
wire n_2342;
wire n_5926;
wire n_2755;
wire n_2301;
wire n_1578;
wire n_2712;
wire n_5316;
wire n_4314;
wire n_2788;
wire n_2089;
wire n_1857;
wire n_1997;
wire n_3314;
wire n_5135;
wire n_1349;
wire n_3891;
wire n_4704;
wire n_1777;
wire n_3409;
wire n_1546;
wire n_6394;
wire n_4003;
wire n_4775;
wire n_3420;
wire n_5840;
wire n_4192;
wire n_4633;
wire n_1950;
wire n_6439;
wire n_6084;
wire n_4593;
wire n_3914;
wire n_3289;
wire n_1834;
wire n_3372;
wire n_4121;
wire n_2862;
wire n_3850;
wire n_4488;
wire n_3405;
wire n_1657;
wire n_1741;
wire n_4264;
wire n_4183;
wire n_4118;
wire n_4302;
wire n_2138;
wire n_4916;
wire n_4858;
wire n_1914;
wire n_3833;
wire n_5833;
wire n_3339;
wire n_3673;
wire n_5792;
wire n_2620;
wire n_1826;
wire n_1855;
wire n_4241;
wire n_3556;
wire n_5617;
wire n_1340;
wire n_2562;
wire n_6191;
wire n_3269;
wire n_5491;
wire n_2223;
wire n_5024;
wire n_3876;
wire n_4971;
wire n_1267;
wire n_2683;
wire n_3432;
wire n_5696;
wire n_1816;
wire n_4645;
wire n_4619;
wire n_2318;
wire n_2141;
wire n_1422;
wire n_6044;
wire n_4339;
wire n_5493;
wire n_4085;
wire n_3190;
wire n_3878;
wire n_4661;
wire n_2947;
wire n_4080;
wire n_5406;
wire n_1754;
wire n_3686;
wire n_2679;
wire n_4028;
wire n_5704;
wire n_1517;
wire n_5973;
wire n_3670;
wire n_3002;
wire n_2087;
wire n_2920;
wire n_4289;
wire n_5555;
wire n_1895;
wire n_1860;
wire n_5727;
wire n_5770;
wire n_1763;
wire n_3912;
wire n_5169;
wire n_1607;
wire n_2959;
wire n_2380;
wire n_2420;
wire n_3265;
wire n_2221;
wire n_1774;
wire n_5274;
wire n_2516;
wire n_2031;
wire n_1348;
wire n_1191;
wire n_4099;
wire n_3899;
wire n_6153;
wire n_4729;
wire n_5957;
wire n_1617;
wire n_2639;
wire n_5323;
wire n_3099;
wire n_6412;
wire n_4745;
wire n_4057;
wire n_2410;
wire n_3206;
wire n_2633;
wire n_2049;
wire n_6245;
wire n_2113;
wire n_1690;
wire n_4466;
wire n_4132;
wire n_3361;
wire n_5566;
wire n_6185;
wire n_5342;
wire n_4603;
wire n_1135;
wire n_4300;
wire n_3277;
wire n_2758;
wire n_5787;
wire n_4417;
wire n_5967;
wire n_1550;
wire n_1169;
wire n_6224;
wire n_1938;
wire n_3452;
wire n_4022;
wire n_5843;
wire n_2194;
wire n_6072;
wire n_4320;
wire n_1173;
wire n_2736;
wire n_2845;
wire n_3886;
wire n_1901;
wire n_5332;
wire n_6073;
wire n_3096;
wire n_6097;
wire n_2059;
wire n_1278;
wire n_5553;
wire n_4730;
wire n_5763;
wire n_4616;
wire n_4760;
wire n_1710;
wire n_3021;
wire n_1603;
wire n_5864;
wire n_5227;
wire n_3404;
wire n_2072;
wire n_2963;
wire n_1489;
wire n_1993;
wire n_4859;
wire n_1455;
wire n_2182;
wire n_3115;
wire n_5352;
wire n_4583;
wire n_1502;
wire n_4923;
wire n_3920;
wire n_5370;
wire n_4082;
wire n_3273;
wire n_4367;
wire n_4282;
wire n_5600;
wire n_4475;
wire n_2286;
wire n_2563;
wire n_4893;
wire n_3650;
wire n_5014;
wire n_3513;
wire n_2677;
wire n_2531;
wire n_4029;
wire n_3212;
wire n_1321;
wire n_1779;
wire n_2489;
wire n_2950;
wire n_2272;
wire n_3574;
wire n_2608;
wire n_5824;
wire n_6280;
wire n_5472;
wire n_5950;
wire n_3739;
wire n_2825;
wire n_4338;
wire n_5546;
wire n_6222;
wire n_5972;
wire n_4985;
wire n_2742;
wire n_3604;
wire n_1740;
wire n_3540;
wire n_2680;
wire n_1343;
wire n_1371;
wire n_4198;
wire n_5924;
wire n_4529;
wire n_2861;
wire n_2976;
wire n_2366;
wire n_6318;
wire n_6200;
wire n_4919;
wire n_4111;
wire n_4200;
wire n_1659;
wire n_4575;
wire n_4847;
wire n_1878;
wire n_4803;
wire n_1374;
wire n_2851;
wire n_2973;
wire n_3651;
wire n_4666;
wire n_5752;
wire n_1242;
wire n_2810;
wire n_1119;
wire n_3027;
wire n_4189;
wire n_4076;
wire n_5233;
wire n_3438;
wire n_4835;
wire n_3464;
wire n_4390;
wire n_5977;
wire n_4722;
wire n_1530;
wire n_3215;
wire n_5968;
wire n_2871;
wire n_2764;
wire n_5713;
wire n_3648;
wire n_3234;
wire n_4058;
wire n_6268;
wire n_5403;
wire n_4611;
wire n_5527;
wire n_2714;
wire n_2669;
wire n_4081;
wire n_4391;
wire n_5831;
wire n_1459;
wire n_4032;
wire n_6032;
wire n_2232;
wire n_4541;
wire n_4530;
wire n_1570;
wire n_5048;
wire n_5671;
wire n_6129;
wire n_1303;
wire n_1994;
wire n_6058;
wire n_1526;
wire n_4268;
wire n_2367;
wire n_3236;
wire n_1961;
wire n_3013;
wire n_4265;
wire n_3062;
wire n_3806;
wire n_3256;
wire n_3126;
wire n_5834;
wire n_1257;
wire n_2864;
wire n_1632;
wire n_3104;
wire n_5951;
wire n_4895;
wire n_5480;
wire n_3354;
wire n_4069;
wire n_5289;
wire n_3373;
wire n_2784;
wire n_4140;
wire n_1909;
wire n_4125;
wire n_2495;
wire n_4531;
wire n_4789;
wire n_4778;
wire n_2703;
wire n_6152;
wire n_2574;
wire n_5492;
wire n_1887;
wire n_6106;
wire n_3504;
wire n_3511;
wire n_2428;
wire n_3159;
wire n_1768;
wire n_3697;
wire n_2068;
wire n_2636;
wire n_3101;
wire n_5260;
wire n_6416;
wire n_5069;
wire n_2364;
wire n_2641;
wire n_4751;
wire n_5930;
wire n_5309;
wire n_3774;
wire n_2494;
wire n_3863;
wire n_5782;
wire n_2228;
wire n_4474;
wire n_5646;
wire n_1518;
wire n_4350;
wire n_5327;
wire n_4478;
wire n_2872;
wire n_2411;
wire n_3539;
wire n_2266;
wire n_4473;
wire n_3761;
wire n_2830;
wire n_4675;
wire n_3083;
wire n_5927;
wire n_3844;
wire n_4049;
wire n_2044;
wire n_2091;
wire n_4945;
wire n_3362;
wire n_3035;
wire n_4165;
wire n_5019;
wire n_4891;
wire n_2394;
wire n_1572;
wire n_1245;
wire n_4867;
wire n_2929;
wire n_6346;
wire n_4911;
wire n_5414;
wire n_1329;
wire n_2409;
wire n_6403;
wire n_2405;
wire n_2601;
wire n_4405;
wire n_3118;
wire n_6172;
wire n_3742;
wire n_6004;
wire n_3532;
wire n_6347;
wire n_5280;
wire n_5466;
wire n_5469;
wire n_4686;
wire n_6358;
wire n_4682;
wire n_5750;
wire n_5305;
wire n_2914;
wire n_1833;
wire n_5186;
wire n_1986;
wire n_2882;
wire n_4301;
wire n_2493;
wire n_6215;
wire n_2115;
wire n_2013;
wire n_1556;
wire n_3547;
wire n_4898;
wire n_3700;
wire n_5180;
wire n_6233;
wire n_4733;
wire n_5368;
wire n_6338;
wire n_5757;
wire n_3947;
wire n_4684;
wire n_3663;
wire n_2129;
wire n_3230;
wire n_2532;
wire n_3782;
wire n_1720;
wire n_3831;
wire n_2293;
wire n_3068;
wire n_3071;
wire n_3919;
wire n_3683;
wire n_6053;
wire n_2734;
wire n_1166;
wire n_5267;
wire n_6020;
wire n_2310;
wire n_2674;
wire n_1284;
wire n_6432;
wire n_6426;
wire n_2689;
wire n_1992;
wire n_4493;
wire n_4797;
wire n_4962;
wire n_5397;
wire n_2596;
wire n_1488;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_3606;
wire n_5232;
wire n_1866;
wire n_2169;
wire n_2111;
wire n_1262;
wire n_5890;
wire n_4644;
wire n_4412;
wire n_6068;
wire n_5802;
wire n_4266;
wire n_5815;
wire n_5605;
wire n_3124;
wire n_2634;
wire n_2982;
wire n_5384;
wire n_3015;
wire n_3321;
wire n_3081;
wire n_4639;
wire n_2291;
wire n_5664;
wire n_4102;
wire n_3612;
wire n_2172;
wire n_1728;
wire n_5863;
wire n_1230;
wire n_3622;
wire n_5276;
wire n_3857;
wire n_6042;
wire n_2357;
wire n_5197;
wire n_4354;
wire n_5320;
wire n_2937;
wire n_3728;
wire n_5265;
wire n_5087;
wire n_4401;
wire n_4727;
wire n_6265;
wire n_4296;
wire n_5312;
wire n_5534;
wire n_2967;
wire n_3005;
wire n_4627;
wire n_5107;
wire n_4309;
wire n_4027;
wire n_2056;
wire n_2054;
wire n_2226;
wire n_1402;
wire n_3267;
wire n_3008;
wire n_6452;
wire n_2802;
wire n_4728;
wire n_2279;
wire n_1536;
wire n_1719;
wire n_5281;
wire n_4046;
wire n_2961;
wire n_6458;
wire n_3689;
wire n_4631;
wire n_3283;
wire n_1736;
wire n_6176;
wire n_2907;
wire n_1948;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_6092;
wire n_3675;
wire n_2378;
wire n_2749;
wire n_3658;
wire n_4901;
wire n_3133;
wire n_3527;
wire n_2014;
wire n_3901;
wire n_5025;
wire n_4539;
wire n_1205;
wire n_5575;
wire n_2969;
wire n_6052;
wire n_5753;
wire n_3550;
wire n_5401;
wire n_5509;
wire n_3287;
wire n_3534;
wire n_1837;
wire n_6468;
wire n_1414;
wire n_5506;
wire n_6063;
wire n_2195;
wire n_2940;
wire n_4150;
wire n_3275;
wire n_2645;
wire n_5417;
wire n_1714;
wire n_1958;
wire n_1611;
wire n_5015;
wire n_5372;
wire n_1675;
wire n_1551;
wire n_1533;
wire n_3792;
wire n_2515;
wire n_3089;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_3406;
wire n_3988;
wire n_3758;
wire n_6418;
wire n_2353;
wire n_4251;
wire n_4106;
wire n_3662;
wire n_6344;
wire n_1354;
wire n_3329;
wire n_1277;
wire n_5995;
wire n_3233;
wire n_3193;
wire n_2582;
wire n_5253;
wire n_3789;
wire n_6308;
wire n_2174;
wire n_2510;
wire n_2435;
wire n_3934;
wire n_2583;
wire n_1678;
wire n_4606;
wire n_1287;
wire n_1525;
wire n_6461;
wire n_1150;
wire n_1674;
wire n_6304;
wire n_3980;
wire n_2912;
wire n_2710;
wire n_2970;
wire n_1393;
wire n_4691;
wire n_5937;
wire n_2978;
wire n_5291;
wire n_3502;
wire n_5460;
wire n_3935;
wire n_5379;
wire n_1854;
wire n_2804;
wire n_5390;
wire n_5691;
wire n_4926;
wire n_5043;
wire n_4688;
wire n_5097;
wire n_5675;
wire n_3144;
wire n_4234;
wire n_4146;
wire n_2835;
wire n_4656;
wire n_4932;
wire n_6179;
wire n_1930;
wire n_5577;
wire n_1234;
wire n_4881;
wire n_3755;
wire n_1469;
wire n_4632;
wire n_3255;
wire n_1652;
wire n_2183;
wire n_1883;
wire n_2037;
wire n_4550;
wire n_1226;
wire n_4651;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2682;
wire n_3605;
wire n_5181;
wire n_3105;
wire n_3146;
wire n_4892;
wire n_4343;
wire n_3931;
wire n_5745;
wire n_4421;
wire n_2322;
wire n_3025;
wire n_3411;
wire n_2955;
wire n_3235;
wire n_2989;
wire n_1856;
wire n_5893;
wire n_3843;
wire n_2847;
wire n_4399;
wire n_1308;
wire n_5067;
wire n_3904;
wire n_4378;
wire n_6455;
wire n_3729;
wire n_5637;
wire n_3484;
wire n_2485;
wire n_5614;
wire n_4477;
wire n_5177;
wire n_5643;
wire n_2179;
wire n_4654;
wire n_3984;
wire n_4233;
wire n_4765;
wire n_3086;
wire n_2475;
wire n_3721;
wire n_5695;
wire n_3726;
wire n_5438;
wire n_4277;
wire n_4431;
wire n_4771;
wire n_4652;
wire n_4970;
wire n_5179;
wire n_3804;
wire n_1908;
wire n_6457;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_4285;
wire n_4928;
wire n_3251;
wire n_2921;
wire n_3724;
wire n_3192;
wire n_3753;
wire n_5683;
wire n_3566;
wire n_2820;
wire n_2311;
wire n_5701;
wire n_4403;
wire n_3242;
wire n_1654;
wire n_6428;
wire n_5774;
wire n_3330;
wire n_2707;
wire n_4746;
wire n_4382;
wire n_4002;
wire n_3631;
wire n_2537;
wire n_1130;
wire n_4246;
wire n_2643;
wire n_4545;
wire n_2336;
wire n_3987;
wire n_3969;
wire n_4437;
wire n_3856;
wire n_1155;
wire n_5394;
wire n_1292;
wire n_5462;
wire n_2432;
wire n_3043;
wire n_2273;
wire n_5428;
wire n_4491;
wire n_4672;
wire n_5001;
wire n_2421;
wire n_3237;
wire n_6095;
wire n_1970;
wire n_3946;
wire n_2953;
wire n_3949;
wire n_3507;
wire n_6150;
wire n_3926;
wire n_3688;
wire n_2462;
wire n_2436;
wire n_1663;
wire n_4267;
wire n_5933;
wire n_4723;
wire n_2269;
wire n_2472;
wire n_2846;
wire n_3699;
wire n_4312;
wire n_5874;
wire n_5104;
wire n_2249;
wire n_3022;
wire n_4014;
wire n_3766;
wire n_3707;
wire n_4217;
wire n_3973;
wire n_5964;
wire n_5551;
wire n_4769;
wire n_4724;
wire n_2260;
wire n_5319;
wire n_5543;
wire n_4721;
wire n_2663;
wire n_3882;
wire n_2595;
wire n_5723;
wire n_5621;
wire n_5386;
wire n_4433;
wire n_5133;
wire n_5056;
wire n_3030;
wire n_5631;
wire n_5983;
wire n_5796;
wire n_4503;
wire n_6232;
wire n_3917;
wire n_3679;
wire n_4517;
wire n_6021;
wire n_3210;
wire n_3221;
wire n_4511;
wire n_1672;
wire n_4171;
wire n_3764;
wire n_5405;
wire n_6389;
wire n_3795;
wire n_6055;
wire n_4788;
wire n_4754;
wire n_1817;
wire n_5848;
wire n_5221;
wire n_1301;
wire n_5997;
wire n_4166;
wire n_2242;
wire n_4845;
wire n_1561;
wire n_5122;
wire n_2247;
wire n_3177;
wire n_3399;
wire n_5439;
wire n_4850;
wire n_1869;
wire n_2189;
wire n_2482;
wire n_3799;
wire n_3676;
wire n_1753;
wire n_6351;
wire n_4610;
wire n_6441;
wire n_5854;
wire n_4067;
wire n_4997;
wire n_5906;
wire n_4393;
wire n_5205;
wire n_3777;
wire n_5916;
wire n_5993;
wire n_4553;
wire n_5240;
wire n_3961;
wire n_1520;
wire n_2509;
wire n_5714;
wire n_4283;
wire n_4174;
wire n_4870;
wire n_2399;
wire n_1370;
wire n_1708;
wire n_3038;
wire n_6476;
wire n_5828;
wire n_6276;
wire n_5907;
wire n_5284;
wire n_4804;
wire n_3716;
wire n_1649;
wire n_3450;
wire n_5357;
wire n_4994;
wire n_4518;
wire n_4732;
wire n_1936;
wire n_1717;
wire n_6040;
wire n_2257;
wire n_4856;
wire n_5088;
wire n_5250;
wire n_1467;
wire n_6388;
wire n_3217;
wire n_2511;
wire n_5461;
wire n_6298;
wire n_3909;
wire n_3971;
wire n_1332;
wire n_2661;
wire n_4079;
wire n_3573;
wire n_3563;
wire n_4993;
wire n_3510;
wire n_4248;
wire n_2334;
wire n_2350;
wire n_5958;
wire n_5619;
wire n_1709;
wire n_2649;
wire n_3607;
wire n_4476;
wire n_6460;
wire n_3241;
wire n_2746;
wire n_5471;
wire n_2256;
wire n_5210;
wire n_2445;
wire n_1980;
wire n_3583;
wire n_4987;
wire n_3832;
wire n_4649;
wire n_3508;
wire n_6295;
wire n_1862;
wire n_4693;
wire n_3415;
wire n_2355;
wire n_4992;
wire n_1543;
wire n_3386;
wire n_4568;
wire n_4359;
wire n_3814;
wire n_1441;
wire n_4573;
wire n_4105;
wire n_4206;
wire n_5273;
wire n_4177;
wire n_1888;
wire n_3320;
wire n_1786;
wire n_2033;
wire n_5877;
wire n_5457;
wire n_5482;
wire n_4700;
wire n_2828;
wire n_1964;
wire n_6090;
wire n_3720;
wire n_1196;
wire n_1182;
wire n_4074;
wire n_5237;
wire n_5360;
wire n_3633;
wire n_1731;
wire n_5596;
wire n_2879;
wire n_3514;
wire n_3091;
wire n_5625;
wire n_4037;
wire n_4582;
wire n_5539;
wire n_3426;
wire n_4308;
wire n_2288;
wire n_3075;
wire n_1671;
wire n_3448;
wire n_3788;
wire n_6164;
wire n_6211;
wire n_2076;
wire n_3733;
wire n_1831;
wire n_4853;
wire n_6117;
wire n_1312;
wire n_5844;
wire n_6470;
wire n_6448;
wire n_3684;
wire n_1318;
wire n_4006;
wire n_1508;
wire n_6018;
wire n_6094;
wire n_3970;
wire n_3291;
wire n_2454;
wire n_4008;
wire n_4973;
wire n_2829;
wire n_4966;
wire n_2968;
wire n_4494;
wire n_3473;
wire n_5362;
wire n_6236;
wire n_6208;
wire n_5294;
wire n_6197;
wire n_3263;
wire n_4501;
wire n_1772;
wire n_2858;
wire n_1283;
wire n_1421;
wire n_4922;
wire n_6237;
wire n_5089;
wire n_2424;
wire n_1793;
wire n_2573;
wire n_2390;
wire n_4402;
wire n_2793;
wire n_4813;
wire n_3098;
wire n_6449;
wire n_1711;
wire n_3069;
wire n_5488;
wire n_3107;
wire n_5465;
wire n_4134;
wire n_4131;
wire n_4330;
wire n_5832;
wire n_2176;
wire n_2805;
wire n_5165;
wire n_2319;
wire n_5678;
wire n_3757;
wire n_5811;
wire n_1933;
wire n_1842;
wire n_3364;
wire n_3429;
wire n_3306;
wire n_5234;
wire n_3787;
wire n_5140;
wire n_3445;
wire n_2080;
wire n_5655;
wire n_5514;
wire n_2554;
wire n_6130;
wire n_1676;
wire n_5020;
wire n_5225;
wire n_1136;
wire n_1918;
wire n_3642;
wire n_2461;
wire n_1229;
wire n_1490;
wire n_1179;
wire n_4818;
wire n_4462;
wire n_1153;
wire n_2787;
wire n_4540;
wire n_4187;
wire n_1273;
wire n_3821;
wire n_2930;
wire n_2616;
wire n_4979;
wire n_3503;
wire n_2441;
wire n_4063;
wire n_4362;
wire n_5318;
wire n_3312;
wire n_1848;
wire n_4009;
wire n_2650;
wire n_2888;
wire n_3614;
wire n_5946;
wire n_6131;
wire n_3394;
wire n_6207;
wire n_5942;
wire n_2530;
wire n_2792;
wire n_2372;
wire n_4191;
wire n_4965;
wire n_1522;
wire n_2523;
wire n_6326;
wire n_3488;
wire n_6365;
wire n_2832;
wire n_4991;
wire n_4525;
wire n_4011;
wire n_3526;
wire n_5242;
wire n_2142;
wire n_3703;
wire n_5116;
wire n_4554;
wire n_1260;
wire n_4097;
wire n_4861;
wire n_3239;
wire n_6155;
wire n_5953;
wire n_2600;
wire n_3952;
wire n_1171;
wire n_1126;
wire n_6151;
wire n_6074;
wire n_4596;
wire n_2434;
wire n_3578;
wire n_4734;
wire n_5947;
wire n_4492;
wire n_3470;
wire n_1738;
wire n_6370;
wire n_1729;
wire n_5563;
wire n_2094;
wire n_1479;
wire n_2306;
wire n_5194;
wire n_4579;
wire n_5628;
wire n_2568;
wire n_2629;
wire n_3587;
wire n_4936;
wire n_2097;
wire n_2109;
wire n_2648;
wire n_6262;
wire n_2398;
wire n_1593;
wire n_1775;
wire n_6361;
wire n_2570;
wire n_4025;
wire n_2184;
wire n_3948;
wire n_2842;
wire n_1400;
wire n_2469;
wire n_6024;
wire n_3074;
wire n_4640;
wire n_5790;
wire n_5746;
wire n_5883;
wire n_5630;
wire n_3136;
wire n_3108;
wire n_2395;
wire n_6062;
wire n_4059;
wire n_4130;
wire n_2752;
wire n_2124;
wire n_3991;
wire n_3974;
wire n_4642;
wire n_3625;
wire n_1746;
wire n_2716;
wire n_2212;
wire n_4878;
wire n_3718;
wire n_1832;
wire n_1128;
wire n_2376;
wire n_3398;
wire n_6252;
wire n_5193;
wire n_2170;
wire n_6407;
wire n_4904;
wire n_1785;
wire n_3999;
wire n_1405;
wire n_4087;
wire n_5153;
wire n_6235;
wire n_5369;
wire n_3238;
wire n_4318;
wire n_3731;
wire n_3555;
wire n_3254;
wire n_5007;
wire n_4717;
wire n_4052;
wire n_6447;
wire n_2463;
wire n_6434;
wire n_2478;
wire n_3178;
wire n_4245;
wire n_3378;
wire n_5689;
wire n_3350;
wire n_6391;
wire n_5399;
wire n_4873;
wire n_3936;
wire n_1560;
wire n_5513;
wire n_3166;
wire n_3953;
wire n_3385;
wire n_1265;
wire n_2488;
wire n_2042;
wire n_5891;
wire n_1925;
wire n_1251;
wire n_3090;
wire n_1247;
wire n_5030;
wire n_3816;
wire n_5755;
wire n_5098;
wire n_4636;
wire n_5408;
wire n_4256;
wire n_1185;
wire n_3575;
wire n_2765;
wire n_4278;
wire n_6165;
wire n_6263;
wire n_4609;
wire n_5148;
wire n_4822;
wire n_2936;
wire n_2985;
wire n_3106;
wire n_4030;
wire n_4276;
wire n_6238;
wire n_4612;
wire n_1148;
wire n_1667;
wire n_6272;
wire n_5454;
wire n_3902;
wire n_1707;
wire n_4203;
wire n_5650;
wire n_2055;
wire n_4866;
wire n_2385;
wire n_3864;
wire n_3026;
wire n_3294;
wire n_4831;
wire n_5656;
wire n_1143;
wire n_2584;
wire n_4381;
wire n_5183;
wire n_2442;
wire n_5072;
wire n_4441;
wire n_2000;
wire n_4083;
wire n_2696;
wire n_4960;
wire n_5146;
wire n_5131;
wire n_1894;
wire n_2904;
wire n_3064;
wire n_2896;
wire n_4228;
wire n_4699;
wire n_5803;
wire n_1331;
wire n_1223;
wire n_5754;
wire n_1739;
wire n_3130;
wire n_1353;
wire n_5018;
wire n_2386;
wire n_3324;
wire n_3073;
wire n_2029;
wire n_4254;
wire n_4536;
wire n_1320;
wire n_4247;
wire n_4071;
wire n_2238;
wire n_4924;
wire n_6398;
wire n_5786;
wire n_4138;
wire n_3100;
wire n_1727;
wire n_6366;
wire n_1294;
wire n_1351;
wire n_5035;
wire n_5425;
wire n_1380;
wire n_6036;
wire n_3336;
wire n_6104;
wire n_1291;
wire n_5742;
wire n_5901;
wire n_3763;
wire n_4284;
wire n_5943;
wire n_4370;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_6253;
wire n_1830;
wire n_3476;
wire n_3990;
wire n_2011;
wire n_4044;
wire n_5499;
wire n_1662;
wire n_3443;
wire n_5143;
wire n_3029;
wire n_4135;
wire n_1626;
wire n_3995;
wire n_4104;
wire n_5302;
wire n_1660;
wire n_5640;
wire n_4000;
wire n_5841;
wire n_5011;
wire n_2556;
wire n_1537;
wire n_3908;
wire n_3696;
wire n_2902;
wire n_6242;
wire n_3608;
wire n_4269;
wire n_4016;
wire n_4915;
wire n_4286;
wire n_3048;
wire n_6414;
wire n_1962;
wire n_5296;
wire n_5159;
wire n_1624;
wire n_1952;
wire n_4795;
wire n_1598;
wire n_2952;
wire n_2250;
wire n_1491;
wire n_3778;
wire n_2075;
wire n_4816;
wire n_3335;
wire n_4846;
wire n_3669;
wire n_1899;
wire n_4001;
wire n_6029;
wire n_2892;
wire n_3356;
wire n_4377;
wire n_3220;
wire n_3422;
wire n_5798;
wire n_2309;
wire n_2274;
wire n_6278;
wire n_5096;
wire n_6443;
wire n_3712;
wire n_5805;
wire n_5171;
wire n_2143;
wire n_4637;
wire n_4976;
wire n_4021;
wire n_5351;
wire n_2739;
wire n_2528;
wire n_2548;
wire n_3216;
wire n_6157;
wire n_6453;
wire n_3061;
wire n_3717;
wire n_3424;
wire n_3745;
wire n_3245;
wire n_4855;
wire n_5851;
wire n_4643;
wire n_5217;
wire n_6030;
wire n_4736;
wire n_2817;
wire n_1790;
wire n_4202;
wire n_3196;
wire n_5767;
wire n_4287;
wire n_2809;
wire n_3921;
wire n_3480;
wire n_1494;
wire n_2060;
wire n_2214;
wire n_1726;
wire n_5751;
wire n_1241;
wire n_5929;
wire n_2589;
wire n_5928;
wire n_1231;
wire n_1208;
wire n_1604;
wire n_4947;
wire n_3506;
wire n_1976;
wire n_1337;
wire n_2984;
wire n_4890;
wire n_4538;
wire n_4023;
wire n_3031;
wire n_4920;
wire n_5862;
wire n_5869;
wire n_1238;
wire n_3959;
wire n_4288;
wire n_2452;
wire n_6274;
wire n_2144;
wire n_4763;
wire n_2592;
wire n_2251;
wire n_5201;
wire n_1644;
wire n_4586;
wire n_6190;
wire n_3860;
wire n_5353;
wire n_1871;
wire n_2868;
wire n_3044;
wire n_3493;
wire n_2818;
wire n_3486;
wire n_2426;
wire n_1403;
wire n_2181;
wire n_3253;
wire n_4034;
wire n_5444;
wire n_1149;
wire n_4905;
wire n_6100;
wire n_1457;
wire n_3172;
wire n_2159;
wire n_2700;
wire n_1222;
wire n_1630;
wire n_1959;
wire n_1198;
wire n_3637;
wire n_3393;
wire n_5772;
wire n_1261;
wire n_5520;
wire n_3327;
wire n_5277;
wire n_5900;
wire n_3647;
wire n_6240;
wire n_3619;
wire n_3928;
wire n_4043;
wire n_1846;
wire n_1573;
wire n_1956;
wire n_5569;
wire n_5779;
wire n_4270;
wire n_2983;
wire n_4273;
wire n_1669;
wire n_6247;
wire n_5109;
wire n_1885;
wire n_1989;
wire n_5837;
wire n_5402;
wire n_1801;
wire n_3740;
wire n_3001;
wire n_4181;
wire n_2161;
wire n_2191;
wire n_2329;
wire n_2576;
wire n_4344;
wire n_1342;
wire n_2756;
wire n_4408;
wire n_1175;
wire n_5473;
wire n_1221;
wire n_3875;
wire n_5113;
wire n_4341;
wire n_4759;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_2567;
wire n_5645;
wire n_2981;
wire n_2222;
wire n_4439;
wire n_5102;
wire n_6258;
wire n_6139;
wire n_5167;
wire n_4565;
wire n_5562;
wire n_1451;
wire n_4663;
wire n_2471;
wire n_5666;
wire n_1288;
wire n_1275;
wire n_4519;
wire n_2757;
wire n_1622;
wire n_3121;
wire n_2121;
wire n_4515;
wire n_1893;
wire n_5639;
wire n_5607;
wire n_2278;
wire n_2433;
wire n_2798;
wire n_3425;
wire n_1771;
wire n_3308;
wire n_6169;
wire n_1507;
wire n_5914;
wire n_1206;
wire n_3576;
wire n_5275;
wire n_3109;
wire n_4838;
wire n_2553;
wire n_4524;
wire n_2218;
wire n_2130;
wire n_4862;
wire n_5114;
wire n_4260;
wire n_4628;
wire n_4696;
wire n_3122;
wire n_3012;
wire n_5005;
wire n_5004;
wire n_3368;
wire n_3586;
wire n_2381;
wire n_2313;
wire n_4597;
wire n_1812;
wire n_5090;
wire n_4574;
wire n_4242;
wire n_4949;
wire n_4748;
wire n_4959;
wire n_1747;
wire n_3400;
wire n_2508;
wire n_4243;
wire n_2540;
wire n_3820;
wire n_5395;
wire n_2672;
wire n_3360;
wire n_1585;
wire n_5649;
wire n_2316;
wire n_5489;
wire n_1995;
wire n_4677;
wire n_1631;
wire n_2911;
wire n_1828;
wire n_1389;
wire n_6380;
wire n_5791;
wire n_1798;
wire n_5559;
wire n_4562;
wire n_1584;
wire n_5009;
wire n_6034;
wire n_1438;
wire n_1973;
wire n_2156;
wire n_4986;
wire n_4453;
wire n_1366;
wire n_1187;
wire n_3173;
wire n_6212;
wire n_4281;
wire n_4332;
wire n_3433;
wire n_3998;
wire n_1686;
wire n_4464;
wire n_3017;
wire n_4605;
wire n_4737;
wire n_6111;
wire n_2542;
wire n_2843;
wire n_3305;
wire n_1635;
wire n_5295;
wire n_6427;
wire n_4310;
wire n_3752;
wire n_2637;
wire n_5047;
wire n_5504;
wire n_5076;
wire n_3543;
wire n_5693;
wire n_3655;
wire n_3791;
wire n_2666;
wire n_3050;
wire n_4091;
wire n_4906;
wire n_4257;
wire n_5712;
wire n_4516;
wire n_2913;
wire n_5028;
wire n_1381;
wire n_2254;
wire n_1597;
wire n_1486;
wire n_6444;
wire n_5622;
wire n_4196;
wire n_5255;
wire n_2371;
wire n_6362;
wire n_3898;
wire n_3366;
wire n_3453;
wire n_4107;
wire n_1949;
wire n_1197;
wire n_2408;
wire n_4961;
wire n_6330;
wire n_5013;
wire n_2140;
wire n_2134;
wire n_2483;
wire n_2466;
wire n_3661;
wire n_5348;
wire n_6405;
wire n_2048;
wire n_2760;
wire n_1299;
wire n_2942;
wire n_4420;
wire n_4964;
wire n_5251;
wire n_5036;
wire n_3665;
wire n_2079;
wire n_4807;
wire n_4886;
wire n_4342;
wire n_5554;
wire n_2671;
wire n_3296;
wire n_5919;
wire n_5978;
wire n_6220;
wire n_1390;
wire n_2775;
wire n_3223;
wire n_2005;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_2848;
wire n_6087;
wire n_1784;
wire n_3200;
wire n_1213;
wire n_3483;
wire n_5702;
wire n_3207;
wire n_5450;
wire n_5806;
wire n_1180;
wire n_4657;
wire n_3869;
wire n_3852;
wire n_1220;
wire n_5071;
wire n_5308;
wire n_5982;
wire n_3036;
wire n_5012;
wire n_5376;
wire n_5778;
wire n_4207;
wire n_1760;
wire n_5208;
wire n_6396;
wire n_2173;
wire n_2824;
wire n_4038;
wire n_5503;
wire n_4793;
wire n_4472;
wire n_2588;
wire n_3046;
wire n_1142;
wire n_1385;
wire n_4395;
wire n_4274;
wire n_5644;
wire n_6368;
wire n_2533;
wire n_1500;
wire n_2706;
wire n_1868;
wire n_2303;
wire n_4532;
wire n_5235;
wire n_5062;
wire n_6309;
wire n_3332;
wire n_5161;
wire n_4413;
wire n_4743;
wire n_2403;
wire n_5016;
wire n_2702;
wire n_3922;
wire n_2791;
wire n_1450;
wire n_2092;
wire n_6248;
wire n_5996;
wire n_3189;
wire n_2797;
wire n_4275;
wire n_2988;
wire n_3945;
wire n_1882;
wire n_2996;
wire n_2836;
wire n_1404;
wire n_3582;
wire n_4830;
wire n_4442;
wire n_5700;
wire n_1442;
wire n_2168;
wire n_4689;
wire n_2886;
wire n_5699;
wire n_6287;
wire n_6022;
wire n_1968;
wire n_4018;
wire n_2609;
wire n_4613;
wire n_5940;
wire n_1483;
wire n_1703;
wire n_1953;
wire n_3715;
wire n_3261;
wire n_5324;
wire n_5421;
wire n_3861;
wire n_5175;
wire n_3161;
wire n_3313;
wire n_1807;
wire n_1310;
wire n_3198;
wire n_5820;
wire n_3463;
wire n_2559;
wire n_4188;
wire n_2619;
wire n_2726;
wire n_2917;
wire n_5340;
wire n_3738;
wire n_1640;
wire n_5694;
wire n_5022;
wire n_1145;
wire n_2307;
wire n_3546;
wire n_1511;
wire n_1651;
wire n_6297;
wire n_5245;
wire n_5651;
wire n_3944;
wire n_3595;
wire n_1732;
wire n_2167;
wire n_3079;
wire n_1696;
wire n_6367;
wire n_6198;
wire n_1355;
wire n_5364;
wire n_5459;
wire n_4534;
wire n_3635;
wire n_3270;
wire n_5168;
wire n_4590;
wire n_4602;
wire n_5510;
wire n_5329;
wire n_6251;
wire n_1335;
wire n_3213;
wire n_4394;
wire n_1900;
wire n_3418;
wire n_2614;
wire n_5581;
wire n_1780;
wire n_3865;
wire n_2769;
wire n_4220;
wire n_5812;
wire n_3244;
wire n_3195;
wire n_3997;
wire n_4742;
wire n_2100;
wire n_4948;
wire n_3903;
wire n_3895;
wire n_1194;
wire n_3851;
wire n_4508;
wire n_4934;
wire n_3482;
wire n_2282;
wire n_3654;
wire n_4939;
wire n_4213;
wire n_2430;
wire n_2673;
wire n_2926;
wire n_1534;
wire n_5711;
wire n_3268;
wire n_4703;
wire n_1655;
wire n_3494;
wire n_3615;
wire n_5970;
wire n_3363;
wire n_1186;
wire n_3180;
wire n_5570;
wire n_1743;
wire n_6310;
wire n_1506;
wire n_5061;
wire n_2594;
wire n_1474;
wire n_3150;
wire n_5550;
wire n_4773;
wire n_3853;
wire n_2512;
wire n_4449;
wire n_5219;
wire n_2607;
wire n_4615;
wire n_3911;
wire n_5132;
wire n_4883;
wire n_6249;
wire n_3559;
wire n_5184;
wire n_6440;
wire n_5747;
wire n_4943;
wire n_5821;
wire n_2498;
wire n_4630;
wire n_3812;
wire n_2017;
wire n_1227;
wire n_5326;
wire n_3750;
wire n_5909;
wire n_6050;
wire n_3838;
wire n_5868;
wire n_1954;
wire n_4749;
wire n_1125;
wire n_2687;
wire n_3456;
wire n_3132;
wire n_5618;
wire n_4159;
wire n_4372;
wire n_5528;
wire n_4731;
wire n_4004;
wire n_1134;
wire n_1684;
wire n_4353;
wire n_5593;
wire n_3334;
wire n_3819;
wire n_2023;
wire n_2720;
wire n_3870;
wire n_5740;
wire n_1233;
wire n_5108;
wire n_3653;
wire n_4360;
wire n_6123;
wire n_4897;
wire n_2139;
wire n_3693;
wire n_5477;
wire n_5934;
wire n_5218;
wire n_1138;
wire n_2943;
wire n_5272;
wire n_3135;
wire n_4239;
wire n_3175;
wire n_6273;
wire n_5464;
wire n_6420;
wire n_6474;
wire n_1268;
wire n_3187;
wire n_3830;
wire n_2724;
wire n_5688;
wire n_6141;
wire n_1829;
wire n_1338;
wire n_6234;
wire n_1327;
wire n_5204;
wire n_5400;
wire n_3407;
wire n_3315;
wire n_4470;
wire n_4690;
wire n_3982;
wire n_6311;
wire n_2565;
wire n_4201;
wire n_6288;
wire n_1636;
wire n_1687;
wire n_5303;
wire n_4584;
wire n_3184;
wire n_6290;
wire n_5804;
wire n_4155;
wire n_3890;
wire n_5519;
wire n_5023;
wire n_2032;
wire n_3392;
wire n_4802;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_5971;
wire n_2198;
wire n_1929;
wire n_5095;
wire n_1680;
wire n_1195;
wire n_5902;
wire n_4304;
wire n_4821;
wire n_4975;
wire n_4160;
wire n_2860;
wire n_2448;
wire n_2015;
wire n_4910;
wire n_5064;
wire n_3641;
wire n_5203;
wire n_5065;
wire n_4887;
wire n_5436;
wire n_3996;
wire n_6056;
wire n_2873;
wire n_1576;
wire n_6466;
wire n_3049;
wire n_4015;
wire n_4211;
wire n_4119;
wire n_3620;
wire n_2558;
wire n_2347;
wire n_3884;
wire n_3103;
wire n_3770;
wire n_4591;
wire n_2527;
wire n_5314;
wire n_5044;
wire n_1509;
wire n_1648;
wire n_2944;
wire n_4349;
wire n_1886;
wire n_6228;
wire n_1841;
wire n_5886;
wire n_2685;
wire n_5344;
wire n_1313;
wire n_4223;
wire n_2090;
wire n_5173;
wire n_5585;
wire n_3722;
wire n_5981;
wire n_3802;
wire n_5343;
wire n_5783;
wire n_2215;
wire n_1449;
wire n_1723;
wire n_3129;
wire n_5515;
wire n_4806;
wire n_2116;
wire n_5784;
wire n_5337;
wire n_3592;
wire n_5545;
wire n_1645;
wire n_3186;
wire n_6393;
wire n_6375;
wire n_1943;
wire n_3541;
wire n_1863;
wire n_5209;
wire n_1269;
wire n_2773;
wire n_3097;
wire n_2906;
wire n_5495;
wire n_3910;
wire n_4238;
wire n_1466;
wire n_3667;
wire n_6424;
wire n_3822;
wire n_1276;
wire n_1637;
wire n_2900;
wire n_5799;
wire n_6296;
wire n_3765;
wire n_2216;
wire n_5888;
wire n_4259;
wire n_1620;
wire n_5196;
wire n_5086;
wire n_6025;
wire n_6168;
wire n_3518;
wire n_5885;
wire n_2022;
wire n_3967;
wire n_2373;
wire n_1853;
wire n_2275;
wire n_5398;
wire n_5434;
wire n_5797;
wire n_2899;
wire n_5830;
wire n_5896;
wire n_3351;
wire n_2008;
wire n_5052;
wire n_2859;
wire n_5952;
wire n_6003;
wire n_2564;
wire n_5110;
wire n_5918;
wire n_4799;
wire n_1356;
wire n_2591;
wire n_3965;
wire n_1969;
wire n_5808;
wire n_6119;
wire n_1296;
wire n_4444;
wire n_4676;
wire n_5212;
wire n_1764;
wire n_1250;
wire n_1190;
wire n_5733;
wire n_4598;
wire n_3259;
wire n_5483;
wire n_4533;
wire n_4078;
wire n_1794;
wire n_3779;
wire n_3203;
wire n_3923;
wire n_4392;
wire n_3808;
wire n_4455;
wire n_3093;
wire n_2664;
wire n_1434;
wire n_4129;
wire n_5278;
wire n_2114;
wire n_6204;
wire n_1609;
wire n_5522;
wire n_3530;
wire n_1132;
wire n_5584;
wire n_4548;
wire n_1803;
wire n_5264;
wire n_6321;
wire n_1281;
wire n_4535;
wire n_1447;
wire n_2150;
wire n_6337;
wire n_4999;
wire n_5328;
wire n_2660;
wire n_5447;
wire n_5029;
wire n_5127;
wire n_5006;
wire n_5679;
wire n_4604;
wire n_5123;
wire n_6160;
wire n_3467;
wire n_6156;
wire n_4240;
wire n_2219;
wire n_6116;
wire n_4522;
wire n_1387;
wire n_3371;
wire n_4713;
wire n_1368;
wire n_1154;
wire n_6267;
wire n_2539;
wire n_1701;
wire n_5236;
wire n_5239;
wire n_5307;
wire n_2387;
wire n_3375;
wire n_2397;
wire n_3317;
wire n_3963;
wire n_3461;
wire n_2729;
wire n_1571;
wire n_2529;
wire n_4103;
wire n_4126;
wire n_4710;
wire n_5576;
wire n_3282;
wire n_5144;
wire n_2708;
wire n_5164;
wire n_2748;
wire n_5359;
wire n_5925;
wire n_2224;
wire n_5526;
wire n_5810;
wire n_2233;
wire n_2499;
wire n_6333;
wire n_5172;
wire n_3888;
wire n_4549;
wire n_3309;
wire n_5126;
wire n_1924;
wire n_3024;
wire n_4767;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_5999;
wire n_5147;
wire n_5407;
wire n_1553;
wire n_3542;
wire n_5536;
wire n_6002;
wire n_3374;
wire n_3704;
wire n_2786;
wire n_1905;
wire n_4355;
wire n_2958;
wire n_6140;
wire n_5903;
wire n_2118;
wire n_2259;
wire n_2162;
wire n_4834;
wire n_6336;
wire n_3660;
wire n_2718;
wire n_4712;
wire n_5849;
wire n_1795;
wire n_3634;
wire n_4096;
wire n_2101;
wire n_5378;
wire n_1152;
wire n_3626;
wire n_2599;
wire n_4571;
wire n_5389;
wire n_6166;
wire n_3171;
wire n_6170;
wire n_1733;
wire n_6257;
wire n_3986;
wire n_2853;
wire n_1552;
wire n_4930;
wire n_5345;
wire n_2217;
wire n_3594;
wire n_2866;
wire n_5138;
wire n_3153;
wire n_6202;
wire n_1189;
wire n_4995;
wire n_4039;
wire n_4253;
wire n_4681;
wire n_2623;
wire n_3232;
wire n_5228;
wire n_2178;
wire n_1181;
wire n_3815;
wire n_4375;
wire n_5629;
wire n_5945;
wire n_4205;
wire n_6161;
wire n_3790;
wire n_6147;
wire n_2404;
wire n_5601;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_1203;
wire n_3640;
wire n_2821;
wire n_4768;
wire n_6133;
wire n_6109;
wire n_5985;
wire n_5435;
wire n_5665;
wire n_3299;
wire n_4070;
wire n_4558;
wire n_6436;
wire n_3065;
wire n_2375;
wire n_2572;
wire n_1656;
wire n_2063;
wire n_3082;
wire n_5709;
wire n_4504;
wire n_5176;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_4864;
wire n_3855;
wire n_3357;
wire n_4485;
wire n_1510;
wire n_5003;
wire n_2852;
wire n_2132;
wire n_5567;
wire n_1236;
wire n_3412;
wire n_5765;
wire n_1712;
wire n_6409;
wire n_4537;
wire n_5771;
wire n_5271;
wire n_1184;
wire n_2585;
wire n_2220;
wire n_4005;
wire n_1364;
wire n_3183;
wire n_4323;
wire n_5068;
wire n_4184;
wire n_2468;
wire n_5078;
wire n_3248;
wire n_2606;
wire n_5980;
wire n_4337;
wire n_4826;
wire n_2152;
wire n_5073;
wire n_5420;
wire n_6386;
wire n_5599;
wire n_4952;
wire n_3785;
wire n_3525;
wire n_5508;
wire n_2779;
wire n_1117;
wire n_2547;
wire n_6473;
wire n_1748;
wire n_2935;
wire n_5084;
wire n_2490;
wire n_3127;
wire n_3496;
wire n_3568;
wire n_5789;
wire n_4876;
wire n_5322;
wire n_3841;
wire n_4626;
wire n_1334;
wire n_3879;
wire n_2402;
wire n_1200;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_5590;
wire n_5638;
wire n_4747;
wire n_5152;
wire n_3341;
wire n_4347;
wire n_1852;
wire n_3868;
wire n_4791;
wire n_5497;
wire n_2481;
wire n_4409;
wire n_5361;
wire n_1264;
wire n_2808;
wire n_5010;
wire n_6363;
wire n_3396;
wire n_6007;
wire n_2102;
wire n_3492;
wire n_3558;
wire n_2751;
wire n_1548;
wire n_4824;
wire n_5117;
wire n_2977;
wire n_1682;
wire n_6142;
wire n_3599;
wire n_6244;
wire n_1896;
wire n_1704;
wire n_2234;
wire n_6369;
wire n_5050;
wire n_5608;
wire n_5610;
wire n_4152;
wire n_1352;
wire n_5125;
wire n_2328;
wire n_4587;
wire n_6118;
wire n_6429;
wire n_6158;
wire n_2332;
wire n_1628;
wire n_1773;
wire n_3580;
wire n_2369;
wire n_5474;
wire n_3584;
wire n_4500;
wire n_5845;
wire n_1395;
wire n_4660;
wire n_2823;
wire n_3274;
wire n_2613;
wire n_6049;
wire n_2419;
wire n_5794;
wire n_5299;
wire n_2807;
wire n_4047;
wire n_5905;
wire n_4157;
wire n_3956;
wire n_1431;
wire n_5202;
wire n_5170;
wire n_5724;
wire n_1523;
wire n_1756;
wire n_6108;
wire n_2241;
wire n_2458;
wire n_3401;
wire n_3032;
wire n_5042;
wire n_1750;
wire n_2833;
wire n_3179;
wire n_6382;
wire n_5662;
wire n_1563;
wire n_4051;
wire n_3123;
wire n_1875;
wire n_1615;
wire n_3719;
wire n_5334;
wire n_5595;
wire n_6260;
wire n_5244;
wire n_2635;
wire n_4077;
wire n_3897;
wire n_3475;
wire n_2077;
wire n_2520;
wire n_2193;
wire n_4010;
wire n_4942;
wire n_4255;
wire n_5692;
wire n_2908;
wire n_4561;
wire n_4957;
wire n_2053;
wire n_1580;
wire n_5728;
wire n_2200;
wire n_2304;
wire n_4683;
wire n_6148;
wire n_6404;
wire n_1439;
wire n_2352;
wire n_4839;
wire n_2185;
wire n_2476;
wire n_1266;
wire n_4814;
wire n_2781;
wire n_6217;
wire n_6324;
wire n_2460;
wire n_4694;
wire n_3600;
wire n_4109;
wire n_1870;
wire n_2484;
wire n_2721;
wire n_2308;
wire n_3498;
wire n_4520;
wire n_1428;
wire n_4026;
wire n_2903;
wire n_3659;
wire n_5795;
wire n_4496;
wire n_6048;
wire n_1528;
wire n_3840;
wire n_5889;
wire n_5856;
wire n_3481;
wire n_4719;
wire n_4100;
wire n_3517;
wire n_5722;
wire n_1413;
wire n_2464;
wire n_5498;
wire n_2925;
wire n_2270;
wire n_5034;
wire n_5725;
wire n_1706;
wire n_1592;
wire n_6110;
wire n_1461;
wire n_2695;
wire n_6300;
wire n_5657;
wire n_3656;
wire n_3137;
wire n_3116;
wire n_4426;
wire n_5282;
wire n_5511;
wire n_2414;
wire n_5736;
wire n_5642;
wire n_3316;
wire n_2465;
wire n_3925;
wire n_4089;
wire n_1683;
wire n_4175;
wire n_4458;
wire n_6001;
wire n_3955;
wire n_3158;
wire n_3657;
wire n_5776;
wire n_5826;
wire n_2684;
wire n_2205;
wire n_3284;
wire n_2875;
wire n_1437;
wire n_2747;
wire n_5932;
wire n_4185;
wire n_2064;
wire n_3088;
wire n_1497;
wire n_2002;
wire n_6088;
wire n_4815;
wire n_2545;
wire n_2050;
wire n_3695;
wire n_6239;
wire n_2500;
wire n_1917;
wire n_1444;
wire n_6091;
wire n_4316;
wire n_5453;
wire n_3328;
wire n_2763;
wire n_5136;
wire n_6352;
wire n_2761;
wire n_4020;
wire n_5494;
wire n_6101;
wire n_1920;
wire n_4306;
wire n_6319;
wire n_2997;
wire n_3735;
wire n_2127;
wire n_6188;
wire n_5718;
wire n_5634;
wire n_3228;
wire n_3028;
wire n_5079;
wire n_3706;
wire n_6395;
wire n_1432;
wire n_3322;
wire n_1174;
wire n_6037;
wire n_4512;
wire n_4483;
wire n_3499;
wire n_3552;
wire n_4164;
wire n_1286;
wire n_3784;
wire n_4142;
wire n_6206;
wire n_4621;
wire n_3016;
wire n_1629;
wire n_5706;
wire n_2694;
wire n_6177;
wire n_3609;
wire n_3447;
wire n_3771;
wire n_4678;
wire n_2647;
wire n_1850;
wire n_1670;
wire n_4123;
wire n_2317;
wire n_1384;
wire n_1612;
wire n_5496;
wire n_3113;
wire n_4305;
wire n_2909;
wire n_4007;
wire n_3960;
wire n_1524;
wire n_4707;
wire n_4429;
wire n_1991;
wire n_2566;
wire n_2210;
wire n_5606;
wire n_6322;
wire n_1225;
wire n_2346;
wire n_4695;
wire n_2180;
wire n_3376;
wire n_6313;
wire n_5989;
wire n_2617;
wire n_5870;
wire n_4163;
wire n_2831;
wire n_2865;
wire n_1625;
wire n_4638;
wire n_5530;
wire n_4498;
wire n_2240;
wire n_1797;
wire n_4750;
wire n_3993;
wire n_2120;
wire n_1289;
wire n_1557;
wire n_1567;
wire n_2007;
wire n_2004;
wire n_5424;
wire n_5230;
wire n_2086;
wire n_4832;
wire n_5229;
wire n_3666;
wire n_6374;
wire n_1839;
wire n_5160;
wire n_2330;
wire n_2555;
wire n_1587;
wire n_6356;
wire n_5313;
wire n_2108;
wire n_6462;
wire n_5333;
wire n_5207;
wire n_2535;
wire n_5158;
wire n_2945;
wire n_5154;
wire n_3057;
wire n_4319;
wire n_3760;
wire n_5721;
wire n_1396;
wire n_1923;
wire n_1224;
wire n_5654;
wire n_2196;
wire n_5860;
wire n_1538;
wire n_3773;
wire n_5884;
wire n_2604;
wire n_3462;
wire n_4373;
wire n_2351;
wire n_2437;
wire n_1889;
wire n_1124;
wire n_5839;
wire n_2688;
wire n_4990;
wire n_3302;
wire n_1673;
wire n_5058;
wire n_2085;
wire n_3304;
wire n_1725;
wire n_6231;
wire n_2149;
wire n_2001;
wire n_1800;
wire n_3746;
wire n_3645;
wire n_5823;
wire n_4262;
wire n_4019;
wire n_2735;
wire n_6401;
wire n_2035;
wire n_4436;
wire n_4697;
wire n_1906;
wire n_1647;
wire n_4357;
wire n_4849;
wire n_5101;
wire n_5532;
wire n_4366;
wire n_4139;
wire n_1270;
wire n_5297;
wire n_4340;
wire n_1476;
wire n_2027;
wire n_5611;
wire n_2012;
wire n_3512;
wire n_4720;
wire n_3892;
wire n_1880;
wire n_6225;
wire n_1642;
wire n_5744;
wire n_2447;
wire n_3358;
wire n_5538;
wire n_2894;
wire n_5249;
wire n_5669;
wire n_2587;
wire n_1605;
wire n_6134;
wire n_2099;
wire n_1202;
wire n_5793;
wire n_3410;
wire n_4900;
wire n_6364;
wire n_5715;
wire n_3408;
wire n_3182;
wire n_1879;
wire n_4941;
wire n_1311;
wire n_5966;
wire n_2299;
wire n_2078;
wire n_6284;
wire n_3709;
wire n_3011;
wire n_5383;
wire n_5775;
wire n_2315;
wire n_3623;
wire n_6230;
wire n_5558;
wire n_2157;
wire n_3446;
wire n_5547;
wire n_5572;
wire n_5659;
wire n_5223;
wire n_1770;
wire n_4167;
wire n_6010;
wire n_3058;
wire n_4334;
wire n_6331;
wire n_2211;
wire n_6047;
wire n_5708;
wire n_5817;
wire n_3384;
wire n_4698;
wire n_2225;
wire n_1411;
wire n_5867;
wire n_1501;
wire n_5636;
wire n_5106;
wire n_5800;
wire n_5257;
wire n_4397;
wire n_3611;
wire n_4186;
wire n_2093;
wire n_2675;
wire n_5371;
wire n_4229;
wire n_4294;
wire n_1919;
wire n_4351;
wire n_6226;
wire n_2893;
wire n_6281;
wire n_2009;
wire n_5731;
wire n_4162;
wire n_1416;
wire n_3465;
wire n_1515;
wire n_4127;
wire n_4620;
wire n_1314;
wire n_3059;
wire n_3085;
wire n_2867;
wire n_2229;
wire n_4770;
wire n_3871;
wire n_2388;
wire n_3112;
wire n_5623;
wire n_5921;
wire n_6082;
wire n_3413;
wire n_4580;
wire n_2624;
wire n_1813;
wire n_4581;
wire n_4618;
wire n_5178;
wire n_5853;
wire n_5898;
wire n_5198;
wire n_2898;
wire n_5437;
wire n_2519;
wire n_2231;
wire n_2816;
wire n_2803;
wire n_3402;
wire n_5053;
wire n_1256;
wire n_4670;
wire n_6162;
wire n_5592;
wire n_5484;
wire n_4982;
wire n_5418;
wire n_6079;
wire n_6013;
wire n_5432;
wire n_1769;
wire n_5270;
wire n_1372;
wire n_1847;
wire n_5166;
wire n_5358;
wire n_3805;
wire n_2406;
wire n_4017;
wire n_1586;
wire n_3497;
wire n_5156;
wire n_3382;
wire n_4236;
wire n_4313;
wire n_5548;
wire n_5687;
wire n_3561;
wire n_2543;
wire n_2992;
wire n_1541;
wire n_6008;
wire n_4907;
wire n_4659;
wire n_2128;
wire n_1697;
wire n_1872;
wire n_5822;
wire n_2690;
wire n_3942;
wire n_2020;
wire n_5758;
wire n_1939;
wire n_5366;
wire n_4053;
wire n_5392;
wire n_4279;
wire n_3937;
wire n_6400;
wire n_3303;
wire n_5115;
wire n_5046;
wire n_5139;
wire n_4555;
wire n_5829;
wire n_5686;
wire n_5735;
wire n_3549;
wire n_1481;
wire n_1928;
wire n_4235;
wire n_3972;
wire n_5674;
wire n_2314;
wire n_2126;
wire n_3403;
wire n_1363;
wire n_1691;
wire n_1361;
wire n_5039;
wire n_1693;
wire n_2081;
wire n_5341;
wire n_2993;
wire n_5032;
wire n_3018;
wire n_4820;
wire n_2449;
wire n_2131;
wire n_2526;
wire n_4794;
wire n_1302;
wire n_5041;
wire n_3989;
wire n_5565;
wire n_6350;
wire n_4752;
wire n_4546;
wire n_3918;
wire n_6378;
wire n_3191;
wire n_3051;
wire n_1317;
wire n_3643;
wire n_2615;
wire n_2487;
wire n_3343;
wire n_4415;
wire n_3163;
wire n_6243;
wire n_3786;
wire n_4061;
wire n_4432;
wire n_1912;
wire n_4552;
wire n_3143;
wire n_1876;
wire n_6419;
wire n_4790;
wire n_1811;
wire n_1285;
wire n_5448;
wire n_4263;
wire n_3725;
wire n_5974;
wire n_5852;
wire n_6143;
wire n_1529;
wire n_1824;
wire n_3522;
wire n_4528;
wire n_4888;
wire n_4502;
wire n_5085;
wire n_4335;
wire n_3444;
wire n_4218;
wire n_4705;
wire n_6112;
wire n_6138;
wire n_3009;
wire n_1141;
wire n_4471;
wire n_3297;
wire n_1168;
wire n_5500;
wire n_6045;
wire n_5293;
wire n_6203;
wire n_3000;
wire n_2305;
wire n_1192;
wire n_1290;
wire n_2514;
wire n_4386;
wire n_4547;
wire n_4836;
wire n_5458;
wire n_3545;
wire n_4193;
wire n_5670;
wire n_1336;
wire n_6433;
wire n_6023;
wire n_1358;
wire n_3318;
wire n_5684;
wire n_1397;
wire n_1359;
wire n_3226;
wire n_3702;
wire n_3981;
wire n_4984;
wire n_1532;
wire n_5624;
wire n_3430;
wire n_1685;
wire n_5325;
wire n_2801;
wire n_3225;
wire n_3067;
wire n_6167;
wire n_6189;
wire n_5059;
wire n_1462;
wire n_5825;
wire n_3823;
wire n_4718;
wire n_3185;
wire n_2326;
wire n_5586;
wire n_1398;
wire n_5222;
wire n_1904;
wire n_2966;
wire n_3084;
wire n_4634;
wire n_6335;
wire n_5741;
wire n_1692;
wire n_5875;
wire n_4796;
wire n_6312;
wire n_4560;
wire n_1240;
wire n_3285;
wire n_5045;
wire n_1814;
wire n_4882;
wire n_1808;
wire n_2768;
wire n_1658;
wire n_5038;
wire n_5769;
wire n_3837;
wire n_4841;
wire n_6213;
wire n_3076;
wire n_6264;
wire n_4954;
wire n_4635;
wire n_4521;
wire n_5703;
wire n_3893;
wire n_4272;
wire n_2148;
wire n_2104;
wire n_2653;
wire n_2855;
wire n_6301;
wire n_2618;
wire n_4448;
wire n_3359;
wire n_5501;
wire n_6216;
wire n_2331;
wire n_1600;
wire n_5894;
wire n_4701;
wire n_5248;
wire n_5872;
wire n_4088;
wire n_2136;
wire n_5443;
wire n_6193;
wire n_1913;
wire n_3056;
wire n_4208;
wire n_5363;
wire n_1472;
wire n_1365;
wire n_2443;
wire n_3052;
wire n_4865;
wire n_2066;
wire n_1974;
wire n_1158;
wire n_4589;
wire n_3924;
wire n_1915;
wire n_2534;
wire n_5908;
wire n_4972;
wire n_5597;
wire n_4617;
wire n_3311;
wire n_1160;
wire n_4094;
wire n_4772;
wire n_4857;
wire n_3613;
wire n_1383;
wire n_2057;
wire n_5984;
wire n_6385;
wire n_5533;
wire n_1822;
wire n_6051;
wire n_1804;
wire n_1581;
wire n_5387;
wire n_4776;
wire n_1975;
wire n_3437;
wire n_3744;
wire n_2246;
wire n_2738;
wire n_1851;
wire n_1755;
wire n_5589;
wire n_4702;
wire n_1341;
wire n_4486;
wire n_4946;
wire n_2202;
wire n_5380;
wire n_2262;
wire n_5134;
wire n_1333;
wire n_4506;
wire n_3157;
wire n_4669;
wire n_4226;
wire n_4153;
wire n_6015;
wire n_4329;
wire n_6435;
wire n_4877;
wire n_3442;
wire n_2327;
wire n_4780;
wire n_6411;
wire n_4327;
wire n_5954;
wire n_5412;
wire n_2656;
wire n_6323;
wire n_4168;
wire n_2258;
wire n_4396;
wire n_2039;
wire n_5174;
wire n_4465;
wire n_6174;
wire n_2544;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_3266;
wire n_5468;
wire n_1843;
wire n_2030;
wire n_4576;
wire n_4075;
wire n_5429;
wire n_3593;
wire n_2536;
wire n_1399;
wire n_3685;
wire n_5269;
wire n_4833;
wire n_1903;
wire n_1849;
wire n_3768;
wire n_4224;
wire n_4868;
wire n_5124;
wire n_2676;
wire n_3515;
wire n_3489;
wire n_3181;
wire n_3644;
wire n_5287;
wire n_4387;
wire n_5865;
wire n_2368;
wire n_6437;
wire n_4896;
wire n_1157;
wire n_2065;
wire n_2901;
wire n_5583;
wire n_3818;
wire n_4368;
wire n_1295;
wire n_1983;
wire n_4798;
wire n_1582;
wire n_2201;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_3610;
wire n_5416;
wire n_2569;
wire n_1998;
wire n_1596;
wire n_3077;
wire n_4158;
wire n_4687;
wire n_4756;
wire n_4095;
wire n_2177;
wire n_2123;
wire n_4364;
wire n_3019;
wire n_2235;
wire n_5373;
wire n_4967;
wire n_6067;
wire n_5377;
wire n_2290;
wire n_3272;
wire n_4346;
wire n_2074;
wire n_2897;
wire n_5350;
wire n_6279;
wire n_4668;
wire n_2383;
wire n_5632;
wire n_2640;
wire n_1492;
wire n_6425;
wire n_1478;
wire n_1796;
wire n_3569;
wire n_1614;
wire n_2374;
wire n_4648;
wire n_2598;
wire n_1722;
wire n_5290;
wire n_4179;
wire n_3340;
wire n_2335;
wire n_4785;
wire n_5120;
wire n_2230;
wire n_5535;
wire n_3033;
wire n_2151;
wire n_5382;
wire n_6354;
wire n_4912;
wire n_6320;
wire n_1971;
wire n_5759;
wire n_2479;
wire n_4914;
wire n_2359;
wire n_2360;
wire n_4902;
wire n_4369;
wire n_1392;
wire n_2158;
wire n_6376;
wire n_2571;
wire n_5479;
wire n_6006;
wire n_5598;
wire n_6132;
wire n_2799;
wire n_4708;
wire n_4592;
wire n_1307;
wire n_5578;
wire n_2644;
wire n_4445;
wire n_3211;
wire n_1840;
wire n_2837;
wire n_6089;
wire n_5211;
wire n_1668;
wire n_5861;
wire n_6417;
wire n_1681;
wire n_4031;
wire n_4120;
wire n_3533;
wire n_3896;
wire n_2192;
wire n_4578;
wire n_3323;
wire n_1937;
wire n_3839;
wire n_3509;
wire n_1749;
wire n_2918;
wire n_3353;
wire n_5092;
wire n_1945;
wire n_5430;
wire n_5182;
wire n_2638;
wire n_3939;
wire n_4874;
wire n_1228;
wire n_4840;
wire n_2354;
wire n_5956;
wire n_6027;
wire n_6477;
wire n_4311;
wire n_5766;
wire n_6269;
wire n_1133;
wire n_1926;
wire n_2363;
wire n_2814;
wire n_5094;
wire n_6275;
wire n_3264;
wire n_3204;
wire n_6390;
wire n_2003;
wire n_3727;
wire n_2621;
wire n_2922;
wire n_6306;
wire n_3881;
wire n_1910;
wire n_5446;
wire n_1606;
wire n_5315;
wire n_3711;
wire n_2164;
wire n_1618;
wire n_3748;
wire n_4389;
wire n_3668;
wire n_3197;
wire n_1955;
wire n_4556;
wire n_2413;
wire n_3148;
wire n_4779;
wire n_6122;
wire n_1253;
wire n_1484;
wire n_2686;
wire n_4214;
wire n_4430;
wire n_3151;
wire n_3977;
wire n_3125;
wire n_2812;
wire n_4889;
wire n_4221;
wire n_1638;
wire n_6175;
wire n_5279;
wire n_4650;
wire n_6415;
wire n_2280;
wire n_4428;
wire n_4784;
wire n_2393;
wire n_4766;
wire n_3809;
wire n_1999;
wire n_3810;
wire n_5103;
wire n_5835;
wire n_4968;
wire n_1215;
wire n_3579;
wire n_2777;
wire n_2480;
wire n_5311;
wire n_2283;
wire n_2806;
wire n_6184;
wire n_2813;
wire n_5268;
wire n_4295;
wire n_1716;
wire n_1412;
wire n_6285;
wire n_5773;
wire n_3310;
wire n_4182;
wire n_1401;
wire n_2951;
wire n_5451;
wire n_5452;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_2579;
wire n_2876;
wire n_3301;
wire n_2370;
wire n_5321;
wire n_5215;
wire n_4600;
wire n_2025;
wire n_3451;
wire n_1219;
wire n_4513;
wire n_5635;
wire n_1252;
wire n_2730;
wire n_1927;
wire n_5356;
wire n_4735;
wire n_2767;
wire n_4667;
wire n_5150;
wire n_2826;
wire n_2112;
wire n_6180;
wire n_5613;
wire n_6137;
wire n_2762;
wire n_4774;
wire n_4711;
wire n_3023;
wire n_3224;
wire n_4481;
wire n_3762;
wire n_6410;
wire n_5063;
wire n_4671;
wire n_1326;
wire n_6046;
wire n_4981;
wire n_1799;
wire n_1689;
wire n_1304;
wire n_6465;
wire n_5653;
wire n_2541;
wire n_4879;
wire n_2987;
wire n_5788;
wire n_1702;
wire n_3916;
wire n_3630;
wire n_1558;
wire n_2722;
wire n_5057;
wire n_3618;
wire n_2727;
wire n_5560;
wire n_2719;
wire n_2213;
wire n_5476;
wire n_3521;
wire n_6121;
wire n_2723;
wire n_6077;
wire n_4054;
wire n_1569;
wire n_6000;
wire n_6205;
wire n_4012;
wire n_5582;
wire n_3567;
wire n_4352;
wire n_1988;
wire n_5935;
wire n_6201;
wire n_2401;
wire n_1787;
wire n_3094;
wire n_2166;
wire n_2451;
wire n_4665;
wire n_2631;
wire n_1867;
wire n_5697;
wire n_4252;
wire n_4505;
wire n_4219;
wire n_5119;
wire n_2292;
wire n_6471;
wire n_3560;
wire n_5813;
wire n_1742;
wire n_1818;
wire n_5100;
wire n_3847;
wire n_2203;
wire n_5427;
wire n_4909;
wire n_2693;
wire n_1159;
wire n_2281;
wire n_3202;
wire n_5467;
wire n_2646;
wire n_5346;
wire n_3887;
wire n_3800;
wire n_4435;
wire n_1235;
wire n_6329;
wire n_4755;
wire n_6355;
wire n_3827;
wire n_6145;
wire n_3156;
wire n_4303;
wire n_3457;
wire n_5633;
wire n_1835;
wire n_2697;
wire n_3531;
wire n_2470;
wire n_5726;
wire n_2890;
wire n_4400;
wire n_1519;
wire n_1425;
wire n_4812;
wire n_5415;
wire n_2069;
wire n_2602;
wire n_4090;
wire n_5445;
wire n_6446;
wire n_4996;
wire n_4136;
wire n_5040;
wire n_1156;
wire n_4358;
wire n_2857;
wire n_5031;
wire n_1360;
wire n_5814;
wire n_5374;
wire n_2070;
wire n_3471;
wire n_4098;
wire n_3117;
wire n_3039;
wire n_3900;
wire n_3478;
wire n_3701;
wire n_2766;
wire n_3756;
wire n_3754;
wire n_4156;
wire n_6057;
wire n_5818;
wire n_2416;
wire n_2962;
wire n_3694;
wire n_2052;
wire n_3690;
wire n_6221;
wire n_5876;
wire n_5529;
wire n_3006;
wire n_3348;
wire n_4758;
wire n_2236;
wire n_5317;
wire n_3957;
wire n_2377;
wire n_2577;
wire n_3165;
wire n_4419;
wire n_2795;
wire n_5490;
wire n_3520;
wire n_2632;
wire n_4406;
wire n_5897;
wire n_5331;
wire n_6107;
wire n_4655;
wire n_6080;
wire n_1634;
wire n_5556;
wire n_1452;
wire n_4953;
wire n_6339;
wire n_4570;
wire n_5391;
wire n_5431;
wire n_3966;
wire n_4293;
wire n_6371;
wire n_6014;
wire n_1577;
wire n_1700;
wire n_4542;
wire n_4122;
wire n_5021;
wire n_2819;
wire n_5523;
wire n_5456;
wire n_1140;
wire n_1985;
wire n_4740;
wire n_3007;
wire n_1487;
wire n_6373;
wire n_1237;
wire n_4230;
wire n_2741;
wire n_4333;
wire n_5231;
wire n_5512;
wire n_6406;
wire n_3436;
wire n_6223;
wire n_4460;
wire n_2312;
wire n_2946;
wire n_4040;
wire n_1884;
wire n_1589;
wire n_2717;
wire n_5720;
wire n_4527;
wire n_2877;
wire n_5881;
wire n_1996;
wire n_5857;
wire n_5256;
wire n_3964;
wire n_3110;
wire n_5717;
wire n_1677;
wire n_4384;
wire n_2297;
wire n_3037;
wire n_3188;
wire n_2780;
wire n_1792;
wire n_3250;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_4762;
wire n_5561;
wire n_1877;
wire n_1477;
wire n_3155;
wire n_4938;
wire n_5487;
wire n_4407;
wire n_5961;
wire n_5077;
wire n_5214;
wire n_1249;
wire n_3468;
wire n_2006;
wire n_1990;
wire n_5413;
wire n_3680;
wire n_6227;
wire n_3624;
wire n_6098;
wire n_4989;
wire n_2467;
wire n_5066;
wire n_4292;
wire n_3145;
wire n_5682;
wire n_2662;
wire n_3872;
wire n_5602;
wire n_3801;
wire n_2883;
wire n_1178;
wire n_6163;
wire n_1464;
wire n_1566;
wire n_4092;
wire n_3003;
wire n_4244;
wire n_2277;
wire n_1982;
wire n_2252;
wire n_1695;
wire n_3331;
wire n_2999;
wire n_2910;
wire n_4414;
wire n_2294;
wire n_2295;
wire n_4977;
wire n_4706;
wire n_1602;
wire n_2965;
wire n_6076;
wire n_5347;
wire n_2382;
wire n_2557;
wire n_2505;
wire n_3554;
wire n_6199;
wire n_3730;
wire n_4307;
wire n_4356;
wire n_1935;
wire n_5568;
wire n_3367;
wire n_1146;
wire n_2785;
wire n_5060;
wire n_4929;
wire n_5121;
wire n_1608;
wire n_3776;
wire n_4951;
wire n_5756;
wire n_5162;
wire n_5224;
wire n_2160;
wire n_2699;
wire n_2991;
wire n_6214;
wire n_1436;
wire n_4137;
wire n_1485;
wire n_2239;
wire n_6289;
wire n_3826;
wire n_4365;
wire n_1979;
wire n_3781;
wire n_4215;
wire n_4315;
wire n_2971;
wire n_3072;
wire n_1545;
wire n_3249;
wire n_3797;
wire n_3281;
wire n_3505;
wire n_4427;
wire n_4564;
wire n_2934;
wire n_6430;
wire n_4042;
wire n_5663;
wire n_2525;
wire n_5552;
wire n_4624;
wire n_6043;
wire n_4317;
wire n_3087;
wire n_4925;
wire n_2197;
wire n_1470;
wire n_2098;
wire n_1761;
wire n_4041;
wire n_5672;
wire n_4958;
wire n_5051;
wire n_4297;
wire n_5367;
wire n_5339;
wire n_4709;
wire n_3379;
wire n_4425;
wire n_3390;
wire n_5000;
wire n_1806;
wire n_1539;
wire n_2711;
wire n_3646;
wire n_2209;
wire n_3020;
wire n_3142;
wire n_2612;
wire n_5226;
wire n_2095;
wire n_2486;
wire n_5855;
wire n_5819;
wire n_2521;
wire n_5388;
wire n_1574;
wire n_6186;
wire n_4764;
wire n_4899;
wire n_6283;
wire n_6445;
wire n_4141;
wire n_4614;
wire n_2979;
wire n_4739;
wire n_1300;
wire n_4035;
wire n_4291;
wire n_6372;
wire n_3419;
wire n_4935;
wire n_4880;
wire n_3167;
wire n_5188;
wire n_2986;
wire n_4969;
wire n_2400;
wire n_6467;
wire n_6144;
wire n_5681;
wire n_2507;
wire n_3682;
wire n_3131;
wire n_1495;
wire n_6291;
wire n_1357;
wire n_4566;
wire n_5262;
wire n_2794;
wire n_3672;
wire n_2496;
wire n_4918;
wire n_2974;
wire n_5604;
wire n_2990;
wire n_2923;
wire n_3449;
wire n_1339;
wire n_1544;
wire n_4933;
wire n_4872;
wire n_5910;
wire n_1315;
wire n_4647;
wire n_2340;
wire n_6125;
wire n_2117;
wire n_5990;
wire n_1328;
wire n_4837;
wire n_6218;
wire n_3638;
wire n_2106;
wire n_5880;
wire n_5685;
wire n_6060;
wire n_1263;
wire n_4940;
wire n_4176;
wire n_4454;
wire n_5992;
wire n_5105;
wire n_5807;
wire n_3772;
wire n_2948;
wire n_4322;
wire n_2298;
wire n_2771;
wire n_4336;
wire n_3219;
wire n_5449;
wire n_3867;
wire n_4956;
wire n_2045;
wire n_1535;
wire n_4227;
wire n_2190;
wire n_1972;
wire n_3080;
wire n_2772;
wire n_2778;
wire n_3929;
wire n_1898;
wire n_1254;
wire n_2524;
wire n_3927;
wire n_1941;
wire n_5338;
wire n_5070;
wire n_3564;
wire n_3095;
wire n_1783;
wire n_5842;
wire n_3279;
wire n_1815;
wire n_3344;
wire n_6173;
wire n_4133;
wire n_6093;
wire n_3985;
wire n_6099;
wire n_5939;
wire n_5481;
wire n_5187;
wire n_5762;
wire n_3252;
wire n_1162;
wire n_2578;
wire n_5486;
wire n_5426;
wire n_2745;
wire n_2110;
wire n_6031;
wire n_6064;
wire n_3747;
wire n_1323;
wire n_5846;
wire n_6033;
wire n_3710;
wire n_1429;
wire n_6316;
wire n_3209;
wire n_2026;
wire n_5537;
wire n_3588;
wire n_5220;
wire n_6341;
wire n_2103;
wire n_4497;
wire n_4388;
wire n_3632;
wire n_5200;
wire n_1874;
wire n_4116;
wire n_3377;
wire n_5816;
wire n_1601;
wire n_3414;
wire n_2933;
wire n_3828;
wire n_1367;
wire n_3240;
wire n_2895;
wire n_1694;
wire n_1458;
wire n_2271;
wire n_2356;
wire n_5676;
wire n_5463;
wire n_2261;
wire n_4066;
wire n_2994;
wire n_4980;
wire n_2105;
wire n_2187;
wire n_5780;
wire n_2642;
wire n_5485;
wire n_5737;
wire n_1643;
wire n_1789;
wire n_2415;
wire n_3152;
wire n_3154;
wire n_2344;
wire n_3589;
wire n_2384;
wire n_1376;
wire n_1858;
wire n_3523;
wire n_2815;
wire n_2446;
wire n_3388;
wire n_1172;
wire n_2659;
wire n_3616;
wire n_6039;
wire n_5355;
wire n_4048;
wire n_4084;
wire n_5149;
wire n_1527;
wire n_3174;
wire n_4848;
wire n_5185;
wire n_2849;
wire n_5847;
wire n_5091;
wire n_5936;
wire n_1177;
wire n_3292;
wire n_6442;
wire n_3940;
wire n_6475;
wire n_2502;
wire n_5396;
wire n_4860;
wire n_4438;
wire n_5300;
wire n_3290;
wire n_3585;
wire n_2878;
wire n_1810;
wire n_6342;
wire n_3047;
wire n_2610;
wire n_5917;
wire n_5306;
wire n_3427;
wire n_1188;
wire n_3431;
wire n_2024;
wire n_3783;
wire n_1503;
wire n_1942;
wire n_4326;
wire n_3141;
wire n_2698;
wire n_3930;
wire n_4149;
wire n_5518;
wire n_5531;
wire n_1259;
wire n_4101;
wire n_4792;
wire n_2916;
wire n_3736;
wire n_2611;
wire n_6012;
wire n_4383;
wire n_2709;
wire n_5074;
wire n_2244;
wire n_6387;
wire n_3664;
wire n_1456;
wire n_3907;
wire n_5246;
wire n_2665;
wire n_5544;
wire n_3063;
wire n_4543;
wire n_2881;
wire n_3862;
wire n_2018;
wire n_3134;
wire n_5652;
wire n_5409;
wire n_2581;
wire n_6271;
wire n_5540;
wire n_2237;
wire n_2268;
wire n_2320;
wire n_2255;
wire n_1820;
wire n_3906;
wire n_3474;
wire n_1946;
wire n_3111;
wire n_4212;
wire n_4827;
wire n_1639;
wire n_2154;
wire n_6149;
wire n_3162;
wire n_4599;
wire n_2732;
wire n_3004;
wire n_3333;
wire n_4509;
wire n_3705;
wire n_4783;
wire n_3276;
wire n_2956;
wire n_1415;
wire n_3743;
wire n_4068;
wire n_2153;
wire n_5777;
wire n_2891;
wire n_2457;
wire n_3825;
wire n_4434;
wire n_2737;
wire n_5557;
wire n_1406;
wire n_3591;
wire n_6054;
wire n_2137;
wire n_5442;
wire n_1473;
wire n_3140;
wire n_2125;
wire n_1176;
wire n_3848;
wire n_1897;
wire n_2477;
wire n_4622;
wire n_5549;
wire n_3139;
wire n_4715;
wire n_6250;
wire n_4222;
wire n_5730;
wire n_2206;
wire n_3734;
wire n_3538;
wire n_4716;
wire n_4588;
wire n_2265;
wire n_5054;
wire n_5349;
wire n_1167;
wire n_3231;
wire n_6423;
wire n_3138;
wire n_6303;
wire n_1282;
wire n_2067;
wire n_2517;
wire n_3349;
wire n_4988;
wire n_5128;
wire n_3454;
wire n_6299;
wire n_4143;
wire n_5027;
wire n_4410;
wire n_5026;
wire n_5189;
wire n_1718;
wire n_3229;
wire n_2546;
wire n_4741;
wire n_6383;
wire n_5516;
wire n_1139;
wire n_2345;
wire n_1324;
wire n_4440;
wire n_3649;
wire n_1838;
wire n_3824;
wire n_3439;
wire n_5525;
wire n_1513;
wire n_5836;
wire n_5677;
wire n_6182;
wire n_1788;
wire n_5764;
wire n_2348;
wire n_6171;
wire n_2417;
wire n_2043;
wire n_3601;
wire n_1621;
wire n_2338;
wire n_3571;
wire n_5768;
wire n_6353;
wire n_6472;
wire n_2248;
wire n_3500;
wire n_2850;
wire n_3962;
wire n_6360;
wire n_3846;
wire n_4328;
wire n_5142;
wire n_1433;
wire n_5082;
wire n_1907;
wire n_3994;
wire n_5911;
wire n_5118;
wire n_2135;
wire n_5781;
wire n_5739;
wire n_6075;
wire n_5145;
wire n_4487;
wire n_1165;
wire n_5111;
wire n_4148;
wire n_3066;
wire n_6135;
wire n_2869;
wire n_6422;
wire n_4829;
wire n_2455;
wire n_2874;
wire n_4937;
wire n_4463;
wire n_2284;
wire n_1931;
wire n_6266;
wire n_5748;
wire n_1809;
wire n_3491;
wire n_4844;
wire n_3271;
wire n_5734;
wire n_2667;
wire n_6317;
wire n_6059;
wire n_5247;
wire n_1565;
wire n_2325;
wire n_6041;
wire n_3346;
wire n_5411;
wire n_5422;
wire n_3391;
wire n_1547;
wire n_1542;
wire n_5991;
wire n_1362;
wire n_6343;
wire n_4178;
wire n_4324;
wire n_3288;
wire n_2518;
wire n_6069;
wire n_3045;
wire n_3014;
wire n_5475;
wire n_1951;
wire n_1330;
wire n_5850;
wire n_6307;
wire n_5440;
wire n_1940;
wire n_3767;
wire n_1212;
wire n_1199;
wire n_4852;
wire n_1978;
wire n_1767;
wire n_1443;
wire n_5641;
wire n_1861;
wire n_1564;
wire n_2593;
wire n_1623;
wire n_6413;
wire n_1131;
wire n_3120;
wire n_1554;
wire n_4843;
wire n_6255;
wire n_4761;
wire n_6294;
wire n_2021;
wire n_2713;
wire n_3227;
wire n_2938;
wire n_3342;
wire n_5441;
wire n_2939;
wire n_4036;
wire n_1147;
wire n_5055;
wire n_4380;
wire n_2790;
wire n_2034;
wire n_3102;
wire n_4345;
wire n_1892;
wire n_5761;
wire n_6195;
wire n_2061;
wire n_6038;
wire n_1373;
wire n_3866;
wire n_3803;
wire n_2083;
wire n_2119;
wire n_5976;
wire n_2207;
wire n_4210;
wire n_3485;
wire n_4810;
wire n_3149;
wire n_5871;
wire n_2827;
wire n_5680;
wire n_3278;
wire n_2701;
wire n_2337;
wire n_4045;
wire n_4871;
wire n_2513;
wire n_1369;
wire n_1297;
wire n_1734;
wire n_4461;
wire n_2323;
wire n_6086;
wire n_5915;
wire n_5524;
wire n_5112;
wire n_3042;
wire n_5542;
wire n_5627;
wire n_2561;
wire n_5785;
wire n_2491;
wire n_6438;
wire n_5298;
wire n_1161;
wire n_4363;
wire n_5564;
wire n_5603;
wire n_3551;
wire n_3992;
wire n_4147;
wire n_6451;
wire n_4811;
wire n_5093;
wire n_5710;
wire n_3176;
wire n_2429;
wire n_3326;
wire n_5986;
wire n_3581;
wire n_3423;
wire n_1646;
wire n_4161;
wire n_5137;
wire n_1759;
wire n_2096;
wire n_5912;
wire n_2296;
wire n_6194;
wire n_1911;
wire n_6381;
wire n_2870;
wire n_4869;
wire n_6397;
wire n_4013;
wire n_1211;
wire n_4482;
wire n_3794;
wire n_5283;
wire n_1419;
wire n_4738;
wire n_1193;
wire n_2928;
wire n_3380;
wire n_3557;
wire n_2227;
wire n_2652;
wire n_3596;
wire n_5286;
wire n_2627;
wire n_1827;
wire n_3369;
wire n_5626;
wire n_4086;
wire n_5410;
wire n_4112;
wire n_2501;
wire n_2051;
wire n_1805;
wire n_3737;
wire n_1183;
wire n_3160;
wire n_4744;
wire n_1204;
wire n_1151;
wire n_3286;
wire n_2668;
wire n_1386;
wire n_2931;
wire n_2492;
wire n_5960;
wire n_3636;
wire n_4787;
wire n_4885;
wire n_2927;
wire n_4459;
wire n_1516;
wire n_4551;
wire n_4484;
wire n_5988;
wire n_1499;
wire n_5838;
wire n_2155;
wire n_3938;
wire n_6103;
wire n_6016;
wire n_3114;
wire n_3905;
wire n_1661;
wire n_6261;
wire n_1965;
wire n_5616;
wire n_1757;
wire n_6399;
wire n_4726;
wire n_3617;
wire n_3602;
wire n_4298;
wire n_6181;
wire n_3053;
wire n_5965;
wire n_3894;
wire n_2407;
wire n_2267;
wire n_2302;
wire n_2082;
wire n_2560;
wire n_2453;
wire n_4544;
wire n_4418;
wire n_4595;
wire n_2770;
wire n_2704;
wire n_6246;
wire n_1762;
wire n_4944;
wire n_4468;
wire n_5923;
wire n_6357;
wire n_3421;
wire n_4950;
wire n_3247;
wire n_1454;
wire n_4108;
wire n_4594;
wire n_6359;
wire n_5949;
wire n_1325;
wire n_2754;
wire n_4629;
wire n_4903;
wire n_3041;
wire n_4194;
wire n_3713;
wire n_2692;
wire n_5738;
wire n_3889;
wire n_3325;
wire n_4299;
wire n_1744;
wire n_2324;
wire n_6096;
wire n_4921;
wire n_1819;
wire n_4863;
wire n_2670;
wire n_1745;
wire n_3941;
wire n_3516;
wire n_3933;
wire n_3562;
wire n_1916;
wire n_3873;
wire n_2073;
wire n_4093;
wire n_1947;
wire n_2165;
wire n_2016;
wire n_3793;
wire n_5080;
wire n_5975;
wire n_1791;
wire n_5301;
wire n_6464;
wire n_4817;
wire n_1468;
wire n_4917;
wire n_6017;
wire n_5507;
wire n_1164;
wire n_6340;
wire n_3749;
wire n_5470;
wire n_6315;
wire n_3691;
wire n_4452;
wire n_3501;
wire n_2538;
wire n_1559;
wire n_4446;
wire n_1280;
wire n_2854;
wire n_3258;
wire n_2932;
wire n_6392;
wire n_4280;
wire n_2285;
wire n_5979;
wire n_1934;
wire n_2040;
wire n_3246;
wire n_2186;
wire n_5648;
wire n_1665;
wire n_5335;
wire n_5594;
wire n_3417;
wire n_2725;
wire n_1482;
wire n_4782;
wire n_5393;
wire n_5661;
wire n_4978;
wire n_6292;
wire n_5690;
wire n_2349;
wire n_1902;
wire n_2474;
wire n_6154;
wire n_5963;
wire n_6293;
wire n_1417;
wire n_5455;
wire n_3536;
wire n_1346;
wire n_5873;
wire n_2834;
wire n_6127;
wire n_1123;
wire n_1272;
wire n_2497;
wire n_3040;
wire n_6028;
wire n_6325;
wire n_1410;
wire n_3528;
wire n_3677;
wire n_2657;
wire n_2743;
wire n_5698;
wire n_4662;
wire n_2658;

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_1011),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_477),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_359),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_370),
.Y(n_1119)
);

BUFx10_ASAP7_75t_L g1120 ( 
.A(n_267),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_937),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_31),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_841),
.Y(n_1123)
);

BUFx3_ASAP7_75t_L g1124 ( 
.A(n_815),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_280),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_428),
.Y(n_1126)
);

BUFx10_ASAP7_75t_L g1127 ( 
.A(n_1074),
.Y(n_1127)
);

BUFx2_ASAP7_75t_L g1128 ( 
.A(n_16),
.Y(n_1128)
);

INVx2_ASAP7_75t_SL g1129 ( 
.A(n_839),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_266),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_466),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_96),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_734),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_518),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_624),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_357),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_1054),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_772),
.Y(n_1138)
);

BUFx10_ASAP7_75t_L g1139 ( 
.A(n_819),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_160),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_648),
.Y(n_1141)
);

INVx2_ASAP7_75t_SL g1142 ( 
.A(n_821),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1009),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_210),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_760),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_551),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_523),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_34),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_950),
.Y(n_1149)
);

CKINVDCx20_ASAP7_75t_R g1150 ( 
.A(n_102),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_789),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_272),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_1069),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_624),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_1021),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_385),
.Y(n_1156)
);

BUFx6f_ASAP7_75t_L g1157 ( 
.A(n_507),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_1073),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_1112),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1092),
.Y(n_1160)
);

BUFx10_ASAP7_75t_L g1161 ( 
.A(n_1036),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_205),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_157),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_45),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_895),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_682),
.Y(n_1166)
);

INVx2_ASAP7_75t_SL g1167 ( 
.A(n_51),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_536),
.Y(n_1168)
);

BUFx6f_ASAP7_75t_L g1169 ( 
.A(n_336),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_12),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_906),
.Y(n_1171)
);

INVx1_ASAP7_75t_SL g1172 ( 
.A(n_184),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_443),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_259),
.Y(n_1174)
);

BUFx6f_ASAP7_75t_L g1175 ( 
.A(n_157),
.Y(n_1175)
);

BUFx6f_ASAP7_75t_L g1176 ( 
.A(n_582),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_637),
.Y(n_1177)
);

BUFx8_ASAP7_75t_SL g1178 ( 
.A(n_61),
.Y(n_1178)
);

BUFx3_ASAP7_75t_L g1179 ( 
.A(n_686),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_621),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1114),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_804),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_624),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_236),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_289),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_11),
.Y(n_1186)
);

BUFx6f_ASAP7_75t_L g1187 ( 
.A(n_1067),
.Y(n_1187)
);

CKINVDCx20_ASAP7_75t_R g1188 ( 
.A(n_312),
.Y(n_1188)
);

CKINVDCx20_ASAP7_75t_R g1189 ( 
.A(n_791),
.Y(n_1189)
);

CKINVDCx16_ASAP7_75t_R g1190 ( 
.A(n_385),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_312),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_564),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1022),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_1035),
.Y(n_1194)
);

CKINVDCx20_ASAP7_75t_R g1195 ( 
.A(n_534),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_286),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_1009),
.Y(n_1197)
);

BUFx6f_ASAP7_75t_L g1198 ( 
.A(n_1079),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1070),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_1084),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_699),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_408),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_105),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_813),
.Y(n_1204)
);

INVxp67_ASAP7_75t_L g1205 ( 
.A(n_1032),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_995),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_1077),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_122),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_920),
.Y(n_1209)
);

BUFx10_ASAP7_75t_L g1210 ( 
.A(n_826),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_296),
.Y(n_1211)
);

BUFx10_ASAP7_75t_L g1212 ( 
.A(n_354),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_617),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_697),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_492),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_419),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_216),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_813),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_554),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_295),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_296),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_45),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_794),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1066),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_943),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_662),
.Y(n_1226)
);

INVx2_ASAP7_75t_SL g1227 ( 
.A(n_483),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_413),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_727),
.Y(n_1229)
);

BUFx2_ASAP7_75t_L g1230 ( 
.A(n_243),
.Y(n_1230)
);

BUFx2_ASAP7_75t_L g1231 ( 
.A(n_921),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_1012),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_29),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_1011),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_1070),
.Y(n_1235)
);

CKINVDCx20_ASAP7_75t_R g1236 ( 
.A(n_425),
.Y(n_1236)
);

BUFx10_ASAP7_75t_L g1237 ( 
.A(n_850),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_621),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_318),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_501),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_1022),
.Y(n_1241)
);

CKINVDCx5p33_ASAP7_75t_R g1242 ( 
.A(n_31),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_388),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_828),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_970),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_467),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_546),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_717),
.Y(n_1248)
);

CKINVDCx5p33_ASAP7_75t_R g1249 ( 
.A(n_177),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_940),
.Y(n_1250)
);

CKINVDCx20_ASAP7_75t_R g1251 ( 
.A(n_872),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_1031),
.Y(n_1252)
);

CKINVDCx20_ASAP7_75t_R g1253 ( 
.A(n_705),
.Y(n_1253)
);

BUFx2_ASAP7_75t_L g1254 ( 
.A(n_484),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_377),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_805),
.Y(n_1256)
);

CKINVDCx20_ASAP7_75t_R g1257 ( 
.A(n_44),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_696),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_40),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_943),
.Y(n_1260)
);

CKINVDCx5p33_ASAP7_75t_R g1261 ( 
.A(n_982),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_929),
.Y(n_1262)
);

CKINVDCx5p33_ASAP7_75t_R g1263 ( 
.A(n_400),
.Y(n_1263)
);

BUFx6f_ASAP7_75t_L g1264 ( 
.A(n_89),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_390),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_879),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_588),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_459),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_629),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_768),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_973),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_866),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_737),
.Y(n_1273)
);

INVx1_ASAP7_75t_SL g1274 ( 
.A(n_101),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_528),
.Y(n_1275)
);

CKINVDCx5p33_ASAP7_75t_R g1276 ( 
.A(n_908),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_841),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_859),
.Y(n_1278)
);

CKINVDCx5p33_ASAP7_75t_R g1279 ( 
.A(n_287),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_1112),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_516),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_76),
.Y(n_1282)
);

CKINVDCx5p33_ASAP7_75t_R g1283 ( 
.A(n_608),
.Y(n_1283)
);

CKINVDCx5p33_ASAP7_75t_R g1284 ( 
.A(n_383),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_451),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_222),
.Y(n_1286)
);

INVx1_ASAP7_75t_SL g1287 ( 
.A(n_175),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_872),
.Y(n_1288)
);

CKINVDCx5p33_ASAP7_75t_R g1289 ( 
.A(n_1014),
.Y(n_1289)
);

BUFx6f_ASAP7_75t_L g1290 ( 
.A(n_170),
.Y(n_1290)
);

CKINVDCx20_ASAP7_75t_R g1291 ( 
.A(n_125),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_497),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_308),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_72),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_289),
.Y(n_1295)
);

INVx2_ASAP7_75t_L g1296 ( 
.A(n_976),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_1082),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_1054),
.Y(n_1298)
);

HB1xp67_ASAP7_75t_L g1299 ( 
.A(n_296),
.Y(n_1299)
);

BUFx6f_ASAP7_75t_L g1300 ( 
.A(n_144),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_713),
.Y(n_1301)
);

INVxp67_ASAP7_75t_SL g1302 ( 
.A(n_40),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_578),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_901),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_930),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_56),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1004),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_214),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_959),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_626),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_606),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_785),
.Y(n_1312)
);

CKINVDCx5p33_ASAP7_75t_R g1313 ( 
.A(n_102),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_767),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_378),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1017),
.Y(n_1316)
);

CKINVDCx5p33_ASAP7_75t_R g1317 ( 
.A(n_635),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_1017),
.Y(n_1318)
);

CKINVDCx5p33_ASAP7_75t_R g1319 ( 
.A(n_849),
.Y(n_1319)
);

CKINVDCx5p33_ASAP7_75t_R g1320 ( 
.A(n_351),
.Y(n_1320)
);

BUFx5_ASAP7_75t_L g1321 ( 
.A(n_271),
.Y(n_1321)
);

INVx1_ASAP7_75t_SL g1322 ( 
.A(n_156),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_611),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_771),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_112),
.Y(n_1325)
);

CKINVDCx5p33_ASAP7_75t_R g1326 ( 
.A(n_834),
.Y(n_1326)
);

BUFx10_ASAP7_75t_L g1327 ( 
.A(n_934),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_45),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_274),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_45),
.Y(n_1330)
);

CKINVDCx20_ASAP7_75t_R g1331 ( 
.A(n_942),
.Y(n_1331)
);

CKINVDCx5p33_ASAP7_75t_R g1332 ( 
.A(n_561),
.Y(n_1332)
);

BUFx8_ASAP7_75t_SL g1333 ( 
.A(n_230),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_276),
.Y(n_1334)
);

CKINVDCx5p33_ASAP7_75t_R g1335 ( 
.A(n_817),
.Y(n_1335)
);

CKINVDCx16_ASAP7_75t_R g1336 ( 
.A(n_672),
.Y(n_1336)
);

CKINVDCx5p33_ASAP7_75t_R g1337 ( 
.A(n_286),
.Y(n_1337)
);

BUFx6f_ASAP7_75t_L g1338 ( 
.A(n_463),
.Y(n_1338)
);

CKINVDCx5p33_ASAP7_75t_R g1339 ( 
.A(n_531),
.Y(n_1339)
);

CKINVDCx5p33_ASAP7_75t_R g1340 ( 
.A(n_584),
.Y(n_1340)
);

BUFx3_ASAP7_75t_L g1341 ( 
.A(n_315),
.Y(n_1341)
);

BUFx6f_ASAP7_75t_L g1342 ( 
.A(n_186),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1105),
.Y(n_1343)
);

BUFx3_ASAP7_75t_L g1344 ( 
.A(n_1081),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_523),
.Y(n_1345)
);

CKINVDCx5p33_ASAP7_75t_R g1346 ( 
.A(n_545),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_704),
.Y(n_1347)
);

CKINVDCx5p33_ASAP7_75t_R g1348 ( 
.A(n_607),
.Y(n_1348)
);

BUFx6f_ASAP7_75t_L g1349 ( 
.A(n_1086),
.Y(n_1349)
);

CKINVDCx5p33_ASAP7_75t_R g1350 ( 
.A(n_874),
.Y(n_1350)
);

CKINVDCx5p33_ASAP7_75t_R g1351 ( 
.A(n_846),
.Y(n_1351)
);

CKINVDCx5p33_ASAP7_75t_R g1352 ( 
.A(n_422),
.Y(n_1352)
);

CKINVDCx5p33_ASAP7_75t_R g1353 ( 
.A(n_847),
.Y(n_1353)
);

CKINVDCx16_ASAP7_75t_R g1354 ( 
.A(n_404),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_219),
.Y(n_1355)
);

INVx2_ASAP7_75t_SL g1356 ( 
.A(n_1043),
.Y(n_1356)
);

CKINVDCx5p33_ASAP7_75t_R g1357 ( 
.A(n_713),
.Y(n_1357)
);

CKINVDCx20_ASAP7_75t_R g1358 ( 
.A(n_852),
.Y(n_1358)
);

CKINVDCx16_ASAP7_75t_R g1359 ( 
.A(n_840),
.Y(n_1359)
);

CKINVDCx5p33_ASAP7_75t_R g1360 ( 
.A(n_486),
.Y(n_1360)
);

CKINVDCx5p33_ASAP7_75t_R g1361 ( 
.A(n_1080),
.Y(n_1361)
);

CKINVDCx20_ASAP7_75t_R g1362 ( 
.A(n_629),
.Y(n_1362)
);

BUFx3_ASAP7_75t_L g1363 ( 
.A(n_985),
.Y(n_1363)
);

BUFx6f_ASAP7_75t_L g1364 ( 
.A(n_685),
.Y(n_1364)
);

CKINVDCx5p33_ASAP7_75t_R g1365 ( 
.A(n_631),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1053),
.Y(n_1366)
);

CKINVDCx5p33_ASAP7_75t_R g1367 ( 
.A(n_399),
.Y(n_1367)
);

INVx1_ASAP7_75t_SL g1368 ( 
.A(n_743),
.Y(n_1368)
);

CKINVDCx5p33_ASAP7_75t_R g1369 ( 
.A(n_169),
.Y(n_1369)
);

CKINVDCx5p33_ASAP7_75t_R g1370 ( 
.A(n_997),
.Y(n_1370)
);

CKINVDCx5p33_ASAP7_75t_R g1371 ( 
.A(n_1031),
.Y(n_1371)
);

CKINVDCx5p33_ASAP7_75t_R g1372 ( 
.A(n_239),
.Y(n_1372)
);

CKINVDCx5p33_ASAP7_75t_R g1373 ( 
.A(n_327),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_35),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_917),
.Y(n_1375)
);

BUFx3_ASAP7_75t_L g1376 ( 
.A(n_284),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_219),
.Y(n_1377)
);

INVx1_ASAP7_75t_SL g1378 ( 
.A(n_241),
.Y(n_1378)
);

CKINVDCx20_ASAP7_75t_R g1379 ( 
.A(n_466),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1102),
.Y(n_1380)
);

CKINVDCx5p33_ASAP7_75t_R g1381 ( 
.A(n_270),
.Y(n_1381)
);

CKINVDCx5p33_ASAP7_75t_R g1382 ( 
.A(n_277),
.Y(n_1382)
);

CKINVDCx5p33_ASAP7_75t_R g1383 ( 
.A(n_49),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_25),
.Y(n_1384)
);

CKINVDCx5p33_ASAP7_75t_R g1385 ( 
.A(n_236),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1084),
.Y(n_1386)
);

CKINVDCx5p33_ASAP7_75t_R g1387 ( 
.A(n_1003),
.Y(n_1387)
);

BUFx2_ASAP7_75t_L g1388 ( 
.A(n_4),
.Y(n_1388)
);

CKINVDCx5p33_ASAP7_75t_R g1389 ( 
.A(n_551),
.Y(n_1389)
);

CKINVDCx5p33_ASAP7_75t_R g1390 ( 
.A(n_273),
.Y(n_1390)
);

CKINVDCx5p33_ASAP7_75t_R g1391 ( 
.A(n_461),
.Y(n_1391)
);

CKINVDCx5p33_ASAP7_75t_R g1392 ( 
.A(n_377),
.Y(n_1392)
);

CKINVDCx16_ASAP7_75t_R g1393 ( 
.A(n_462),
.Y(n_1393)
);

INVx1_ASAP7_75t_SL g1394 ( 
.A(n_936),
.Y(n_1394)
);

CKINVDCx14_ASAP7_75t_R g1395 ( 
.A(n_227),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_198),
.Y(n_1396)
);

BUFx6f_ASAP7_75t_L g1397 ( 
.A(n_806),
.Y(n_1397)
);

CKINVDCx5p33_ASAP7_75t_R g1398 ( 
.A(n_287),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_955),
.Y(n_1399)
);

CKINVDCx5p33_ASAP7_75t_R g1400 ( 
.A(n_790),
.Y(n_1400)
);

CKINVDCx5p33_ASAP7_75t_R g1401 ( 
.A(n_642),
.Y(n_1401)
);

CKINVDCx5p33_ASAP7_75t_R g1402 ( 
.A(n_380),
.Y(n_1402)
);

CKINVDCx5p33_ASAP7_75t_R g1403 ( 
.A(n_22),
.Y(n_1403)
);

CKINVDCx20_ASAP7_75t_R g1404 ( 
.A(n_701),
.Y(n_1404)
);

CKINVDCx5p33_ASAP7_75t_R g1405 ( 
.A(n_433),
.Y(n_1405)
);

CKINVDCx5p33_ASAP7_75t_R g1406 ( 
.A(n_1035),
.Y(n_1406)
);

CKINVDCx5p33_ASAP7_75t_R g1407 ( 
.A(n_581),
.Y(n_1407)
);

CKINVDCx5p33_ASAP7_75t_R g1408 ( 
.A(n_186),
.Y(n_1408)
);

CKINVDCx20_ASAP7_75t_R g1409 ( 
.A(n_281),
.Y(n_1409)
);

CKINVDCx5p33_ASAP7_75t_R g1410 ( 
.A(n_669),
.Y(n_1410)
);

CKINVDCx5p33_ASAP7_75t_R g1411 ( 
.A(n_912),
.Y(n_1411)
);

BUFx2_ASAP7_75t_L g1412 ( 
.A(n_54),
.Y(n_1412)
);

CKINVDCx5p33_ASAP7_75t_R g1413 ( 
.A(n_25),
.Y(n_1413)
);

CKINVDCx5p33_ASAP7_75t_R g1414 ( 
.A(n_469),
.Y(n_1414)
);

CKINVDCx5p33_ASAP7_75t_R g1415 ( 
.A(n_283),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_49),
.Y(n_1416)
);

BUFx6f_ASAP7_75t_L g1417 ( 
.A(n_626),
.Y(n_1417)
);

BUFx3_ASAP7_75t_L g1418 ( 
.A(n_846),
.Y(n_1418)
);

BUFx6f_ASAP7_75t_L g1419 ( 
.A(n_398),
.Y(n_1419)
);

CKINVDCx5p33_ASAP7_75t_R g1420 ( 
.A(n_695),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_261),
.Y(n_1421)
);

CKINVDCx5p33_ASAP7_75t_R g1422 ( 
.A(n_125),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_369),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_153),
.Y(n_1424)
);

BUFx3_ASAP7_75t_L g1425 ( 
.A(n_196),
.Y(n_1425)
);

CKINVDCx5p33_ASAP7_75t_R g1426 ( 
.A(n_504),
.Y(n_1426)
);

CKINVDCx5p33_ASAP7_75t_R g1427 ( 
.A(n_462),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1111),
.Y(n_1428)
);

BUFx10_ASAP7_75t_L g1429 ( 
.A(n_483),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_136),
.Y(n_1430)
);

CKINVDCx5p33_ASAP7_75t_R g1431 ( 
.A(n_236),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_982),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1026),
.Y(n_1433)
);

CKINVDCx5p33_ASAP7_75t_R g1434 ( 
.A(n_1011),
.Y(n_1434)
);

CKINVDCx5p33_ASAP7_75t_R g1435 ( 
.A(n_966),
.Y(n_1435)
);

BUFx2_ASAP7_75t_L g1436 ( 
.A(n_770),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_435),
.Y(n_1437)
);

CKINVDCx5p33_ASAP7_75t_R g1438 ( 
.A(n_503),
.Y(n_1438)
);

CKINVDCx5p33_ASAP7_75t_R g1439 ( 
.A(n_369),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_480),
.Y(n_1440)
);

CKINVDCx20_ASAP7_75t_R g1441 ( 
.A(n_240),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_116),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_382),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_563),
.Y(n_1444)
);

CKINVDCx5p33_ASAP7_75t_R g1445 ( 
.A(n_465),
.Y(n_1445)
);

INVx2_ASAP7_75t_L g1446 ( 
.A(n_801),
.Y(n_1446)
);

INVx1_ASAP7_75t_SL g1447 ( 
.A(n_819),
.Y(n_1447)
);

CKINVDCx5p33_ASAP7_75t_R g1448 ( 
.A(n_892),
.Y(n_1448)
);

CKINVDCx5p33_ASAP7_75t_R g1449 ( 
.A(n_622),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_648),
.Y(n_1450)
);

CKINVDCx5p33_ASAP7_75t_R g1451 ( 
.A(n_264),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_363),
.Y(n_1452)
);

CKINVDCx5p33_ASAP7_75t_R g1453 ( 
.A(n_699),
.Y(n_1453)
);

CKINVDCx5p33_ASAP7_75t_R g1454 ( 
.A(n_638),
.Y(n_1454)
);

CKINVDCx5p33_ASAP7_75t_R g1455 ( 
.A(n_244),
.Y(n_1455)
);

CKINVDCx5p33_ASAP7_75t_R g1456 ( 
.A(n_862),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_516),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_631),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_530),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_427),
.Y(n_1460)
);

CKINVDCx5p33_ASAP7_75t_R g1461 ( 
.A(n_415),
.Y(n_1461)
);

CKINVDCx5p33_ASAP7_75t_R g1462 ( 
.A(n_237),
.Y(n_1462)
);

HB1xp67_ASAP7_75t_L g1463 ( 
.A(n_764),
.Y(n_1463)
);

CKINVDCx5p33_ASAP7_75t_R g1464 ( 
.A(n_651),
.Y(n_1464)
);

CKINVDCx5p33_ASAP7_75t_R g1465 ( 
.A(n_172),
.Y(n_1465)
);

CKINVDCx5p33_ASAP7_75t_R g1466 ( 
.A(n_202),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_618),
.Y(n_1467)
);

CKINVDCx5p33_ASAP7_75t_R g1468 ( 
.A(n_405),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_992),
.Y(n_1469)
);

CKINVDCx5p33_ASAP7_75t_R g1470 ( 
.A(n_605),
.Y(n_1470)
);

BUFx5_ASAP7_75t_L g1471 ( 
.A(n_414),
.Y(n_1471)
);

BUFx10_ASAP7_75t_L g1472 ( 
.A(n_712),
.Y(n_1472)
);

CKINVDCx5p33_ASAP7_75t_R g1473 ( 
.A(n_1112),
.Y(n_1473)
);

BUFx10_ASAP7_75t_L g1474 ( 
.A(n_549),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1019),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_498),
.Y(n_1476)
);

INVx1_ASAP7_75t_SL g1477 ( 
.A(n_962),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_30),
.Y(n_1478)
);

CKINVDCx20_ASAP7_75t_R g1479 ( 
.A(n_124),
.Y(n_1479)
);

CKINVDCx5p33_ASAP7_75t_R g1480 ( 
.A(n_565),
.Y(n_1480)
);

CKINVDCx5p33_ASAP7_75t_R g1481 ( 
.A(n_275),
.Y(n_1481)
);

CKINVDCx5p33_ASAP7_75t_R g1482 ( 
.A(n_285),
.Y(n_1482)
);

BUFx2_ASAP7_75t_L g1483 ( 
.A(n_110),
.Y(n_1483)
);

CKINVDCx5p33_ASAP7_75t_R g1484 ( 
.A(n_6),
.Y(n_1484)
);

BUFx10_ASAP7_75t_L g1485 ( 
.A(n_518),
.Y(n_1485)
);

BUFx3_ASAP7_75t_L g1486 ( 
.A(n_1033),
.Y(n_1486)
);

CKINVDCx5p33_ASAP7_75t_R g1487 ( 
.A(n_242),
.Y(n_1487)
);

INVxp67_ASAP7_75t_L g1488 ( 
.A(n_878),
.Y(n_1488)
);

CKINVDCx20_ASAP7_75t_R g1489 ( 
.A(n_695),
.Y(n_1489)
);

CKINVDCx5p33_ASAP7_75t_R g1490 ( 
.A(n_186),
.Y(n_1490)
);

CKINVDCx5p33_ASAP7_75t_R g1491 ( 
.A(n_463),
.Y(n_1491)
);

CKINVDCx5p33_ASAP7_75t_R g1492 ( 
.A(n_424),
.Y(n_1492)
);

CKINVDCx5p33_ASAP7_75t_R g1493 ( 
.A(n_63),
.Y(n_1493)
);

CKINVDCx5p33_ASAP7_75t_R g1494 ( 
.A(n_387),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_428),
.Y(n_1495)
);

CKINVDCx5p33_ASAP7_75t_R g1496 ( 
.A(n_27),
.Y(n_1496)
);

BUFx10_ASAP7_75t_L g1497 ( 
.A(n_80),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_27),
.Y(n_1498)
);

CKINVDCx5p33_ASAP7_75t_R g1499 ( 
.A(n_94),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1074),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_696),
.Y(n_1501)
);

INVx1_ASAP7_75t_SL g1502 ( 
.A(n_412),
.Y(n_1502)
);

CKINVDCx5p33_ASAP7_75t_R g1503 ( 
.A(n_187),
.Y(n_1503)
);

CKINVDCx5p33_ASAP7_75t_R g1504 ( 
.A(n_755),
.Y(n_1504)
);

CKINVDCx5p33_ASAP7_75t_R g1505 ( 
.A(n_997),
.Y(n_1505)
);

INVxp67_ASAP7_75t_L g1506 ( 
.A(n_678),
.Y(n_1506)
);

BUFx6f_ASAP7_75t_L g1507 ( 
.A(n_441),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_124),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_48),
.Y(n_1509)
);

CKINVDCx5p33_ASAP7_75t_R g1510 ( 
.A(n_1037),
.Y(n_1510)
);

CKINVDCx5p33_ASAP7_75t_R g1511 ( 
.A(n_41),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_893),
.Y(n_1512)
);

CKINVDCx5p33_ASAP7_75t_R g1513 ( 
.A(n_44),
.Y(n_1513)
);

CKINVDCx5p33_ASAP7_75t_R g1514 ( 
.A(n_15),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_561),
.Y(n_1515)
);

CKINVDCx5p33_ASAP7_75t_R g1516 ( 
.A(n_378),
.Y(n_1516)
);

INVx1_ASAP7_75t_SL g1517 ( 
.A(n_642),
.Y(n_1517)
);

CKINVDCx5p33_ASAP7_75t_R g1518 ( 
.A(n_358),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_383),
.Y(n_1519)
);

CKINVDCx5p33_ASAP7_75t_R g1520 ( 
.A(n_819),
.Y(n_1520)
);

CKINVDCx20_ASAP7_75t_R g1521 ( 
.A(n_621),
.Y(n_1521)
);

CKINVDCx5p33_ASAP7_75t_R g1522 ( 
.A(n_192),
.Y(n_1522)
);

CKINVDCx5p33_ASAP7_75t_R g1523 ( 
.A(n_574),
.Y(n_1523)
);

BUFx2_ASAP7_75t_L g1524 ( 
.A(n_805),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_279),
.Y(n_1525)
);

CKINVDCx5p33_ASAP7_75t_R g1526 ( 
.A(n_847),
.Y(n_1526)
);

CKINVDCx5p33_ASAP7_75t_R g1527 ( 
.A(n_786),
.Y(n_1527)
);

BUFx2_ASAP7_75t_L g1528 ( 
.A(n_719),
.Y(n_1528)
);

CKINVDCx5p33_ASAP7_75t_R g1529 ( 
.A(n_369),
.Y(n_1529)
);

CKINVDCx5p33_ASAP7_75t_R g1530 ( 
.A(n_83),
.Y(n_1530)
);

CKINVDCx20_ASAP7_75t_R g1531 ( 
.A(n_668),
.Y(n_1531)
);

CKINVDCx5p33_ASAP7_75t_R g1532 ( 
.A(n_423),
.Y(n_1532)
);

CKINVDCx5p33_ASAP7_75t_R g1533 ( 
.A(n_957),
.Y(n_1533)
);

CKINVDCx20_ASAP7_75t_R g1534 ( 
.A(n_659),
.Y(n_1534)
);

CKINVDCx20_ASAP7_75t_R g1535 ( 
.A(n_953),
.Y(n_1535)
);

CKINVDCx5p33_ASAP7_75t_R g1536 ( 
.A(n_165),
.Y(n_1536)
);

CKINVDCx20_ASAP7_75t_R g1537 ( 
.A(n_301),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_50),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_473),
.Y(n_1539)
);

CKINVDCx5p33_ASAP7_75t_R g1540 ( 
.A(n_887),
.Y(n_1540)
);

CKINVDCx5p33_ASAP7_75t_R g1541 ( 
.A(n_422),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_425),
.Y(n_1542)
);

CKINVDCx5p33_ASAP7_75t_R g1543 ( 
.A(n_538),
.Y(n_1543)
);

CKINVDCx5p33_ASAP7_75t_R g1544 ( 
.A(n_506),
.Y(n_1544)
);

CKINVDCx16_ASAP7_75t_R g1545 ( 
.A(n_609),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_822),
.Y(n_1546)
);

HB1xp67_ASAP7_75t_L g1547 ( 
.A(n_999),
.Y(n_1547)
);

CKINVDCx5p33_ASAP7_75t_R g1548 ( 
.A(n_940),
.Y(n_1548)
);

CKINVDCx5p33_ASAP7_75t_R g1549 ( 
.A(n_1064),
.Y(n_1549)
);

CKINVDCx5p33_ASAP7_75t_R g1550 ( 
.A(n_676),
.Y(n_1550)
);

BUFx5_ASAP7_75t_L g1551 ( 
.A(n_93),
.Y(n_1551)
);

CKINVDCx5p33_ASAP7_75t_R g1552 ( 
.A(n_432),
.Y(n_1552)
);

CKINVDCx5p33_ASAP7_75t_R g1553 ( 
.A(n_1075),
.Y(n_1553)
);

CKINVDCx5p33_ASAP7_75t_R g1554 ( 
.A(n_631),
.Y(n_1554)
);

BUFx3_ASAP7_75t_L g1555 ( 
.A(n_552),
.Y(n_1555)
);

BUFx5_ASAP7_75t_L g1556 ( 
.A(n_335),
.Y(n_1556)
);

CKINVDCx14_ASAP7_75t_R g1557 ( 
.A(n_307),
.Y(n_1557)
);

CKINVDCx5p33_ASAP7_75t_R g1558 ( 
.A(n_994),
.Y(n_1558)
);

CKINVDCx5p33_ASAP7_75t_R g1559 ( 
.A(n_596),
.Y(n_1559)
);

CKINVDCx5p33_ASAP7_75t_R g1560 ( 
.A(n_158),
.Y(n_1560)
);

CKINVDCx5p33_ASAP7_75t_R g1561 ( 
.A(n_75),
.Y(n_1561)
);

CKINVDCx5p33_ASAP7_75t_R g1562 ( 
.A(n_551),
.Y(n_1562)
);

INVx1_ASAP7_75t_SL g1563 ( 
.A(n_569),
.Y(n_1563)
);

CKINVDCx5p33_ASAP7_75t_R g1564 ( 
.A(n_1111),
.Y(n_1564)
);

CKINVDCx5p33_ASAP7_75t_R g1565 ( 
.A(n_1032),
.Y(n_1565)
);

CKINVDCx5p33_ASAP7_75t_R g1566 ( 
.A(n_955),
.Y(n_1566)
);

CKINVDCx5p33_ASAP7_75t_R g1567 ( 
.A(n_724),
.Y(n_1567)
);

CKINVDCx5p33_ASAP7_75t_R g1568 ( 
.A(n_780),
.Y(n_1568)
);

BUFx10_ASAP7_75t_L g1569 ( 
.A(n_637),
.Y(n_1569)
);

CKINVDCx5p33_ASAP7_75t_R g1570 ( 
.A(n_1087),
.Y(n_1570)
);

INVx1_ASAP7_75t_SL g1571 ( 
.A(n_80),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_501),
.Y(n_1572)
);

INVx1_ASAP7_75t_SL g1573 ( 
.A(n_1070),
.Y(n_1573)
);

CKINVDCx5p33_ASAP7_75t_R g1574 ( 
.A(n_419),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_274),
.Y(n_1575)
);

CKINVDCx5p33_ASAP7_75t_R g1576 ( 
.A(n_535),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_269),
.Y(n_1577)
);

INVx1_ASAP7_75t_SL g1578 ( 
.A(n_564),
.Y(n_1578)
);

CKINVDCx5p33_ASAP7_75t_R g1579 ( 
.A(n_1072),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_900),
.Y(n_1580)
);

CKINVDCx5p33_ASAP7_75t_R g1581 ( 
.A(n_1071),
.Y(n_1581)
);

CKINVDCx5p33_ASAP7_75t_R g1582 ( 
.A(n_191),
.Y(n_1582)
);

CKINVDCx16_ASAP7_75t_R g1583 ( 
.A(n_217),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_398),
.Y(n_1584)
);

CKINVDCx5p33_ASAP7_75t_R g1585 ( 
.A(n_69),
.Y(n_1585)
);

CKINVDCx5p33_ASAP7_75t_R g1586 ( 
.A(n_941),
.Y(n_1586)
);

CKINVDCx5p33_ASAP7_75t_R g1587 ( 
.A(n_669),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_778),
.Y(n_1588)
);

CKINVDCx5p33_ASAP7_75t_R g1589 ( 
.A(n_1036),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_510),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_781),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_136),
.Y(n_1592)
);

CKINVDCx5p33_ASAP7_75t_R g1593 ( 
.A(n_877),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_611),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1062),
.Y(n_1595)
);

CKINVDCx5p33_ASAP7_75t_R g1596 ( 
.A(n_796),
.Y(n_1596)
);

BUFx10_ASAP7_75t_L g1597 ( 
.A(n_327),
.Y(n_1597)
);

CKINVDCx5p33_ASAP7_75t_R g1598 ( 
.A(n_89),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_822),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_106),
.Y(n_1600)
);

CKINVDCx5p33_ASAP7_75t_R g1601 ( 
.A(n_900),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_504),
.Y(n_1602)
);

CKINVDCx5p33_ASAP7_75t_R g1603 ( 
.A(n_452),
.Y(n_1603)
);

HB1xp67_ASAP7_75t_L g1604 ( 
.A(n_277),
.Y(n_1604)
);

CKINVDCx5p33_ASAP7_75t_R g1605 ( 
.A(n_251),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_985),
.Y(n_1606)
);

CKINVDCx5p33_ASAP7_75t_R g1607 ( 
.A(n_556),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_180),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_499),
.Y(n_1609)
);

CKINVDCx5p33_ASAP7_75t_R g1610 ( 
.A(n_50),
.Y(n_1610)
);

CKINVDCx5p33_ASAP7_75t_R g1611 ( 
.A(n_591),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_636),
.Y(n_1612)
);

CKINVDCx14_ASAP7_75t_R g1613 ( 
.A(n_375),
.Y(n_1613)
);

CKINVDCx16_ASAP7_75t_R g1614 ( 
.A(n_345),
.Y(n_1614)
);

CKINVDCx5p33_ASAP7_75t_R g1615 ( 
.A(n_598),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_185),
.Y(n_1616)
);

CKINVDCx5p33_ASAP7_75t_R g1617 ( 
.A(n_458),
.Y(n_1617)
);

CKINVDCx5p33_ASAP7_75t_R g1618 ( 
.A(n_546),
.Y(n_1618)
);

CKINVDCx20_ASAP7_75t_R g1619 ( 
.A(n_265),
.Y(n_1619)
);

CKINVDCx5p33_ASAP7_75t_R g1620 ( 
.A(n_626),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_59),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1031),
.Y(n_1622)
);

CKINVDCx5p33_ASAP7_75t_R g1623 ( 
.A(n_353),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_258),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_957),
.Y(n_1625)
);

HB1xp67_ASAP7_75t_L g1626 ( 
.A(n_815),
.Y(n_1626)
);

CKINVDCx5p33_ASAP7_75t_R g1627 ( 
.A(n_402),
.Y(n_1627)
);

CKINVDCx5p33_ASAP7_75t_R g1628 ( 
.A(n_250),
.Y(n_1628)
);

CKINVDCx20_ASAP7_75t_R g1629 ( 
.A(n_620),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_289),
.Y(n_1630)
);

INVx1_ASAP7_75t_SL g1631 ( 
.A(n_662),
.Y(n_1631)
);

CKINVDCx5p33_ASAP7_75t_R g1632 ( 
.A(n_352),
.Y(n_1632)
);

CKINVDCx5p33_ASAP7_75t_R g1633 ( 
.A(n_148),
.Y(n_1633)
);

CKINVDCx5p33_ASAP7_75t_R g1634 ( 
.A(n_108),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_183),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_282),
.Y(n_1636)
);

BUFx2_ASAP7_75t_SL g1637 ( 
.A(n_356),
.Y(n_1637)
);

CKINVDCx5p33_ASAP7_75t_R g1638 ( 
.A(n_977),
.Y(n_1638)
);

CKINVDCx5p33_ASAP7_75t_R g1639 ( 
.A(n_866),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_617),
.Y(n_1640)
);

CKINVDCx5p33_ASAP7_75t_R g1641 ( 
.A(n_1078),
.Y(n_1641)
);

CKINVDCx5p33_ASAP7_75t_R g1642 ( 
.A(n_84),
.Y(n_1642)
);

CKINVDCx5p33_ASAP7_75t_R g1643 ( 
.A(n_641),
.Y(n_1643)
);

CKINVDCx5p33_ASAP7_75t_R g1644 ( 
.A(n_268),
.Y(n_1644)
);

CKINVDCx5p33_ASAP7_75t_R g1645 ( 
.A(n_649),
.Y(n_1645)
);

BUFx10_ASAP7_75t_L g1646 ( 
.A(n_800),
.Y(n_1646)
);

CKINVDCx5p33_ASAP7_75t_R g1647 ( 
.A(n_764),
.Y(n_1647)
);

INVxp67_ASAP7_75t_L g1648 ( 
.A(n_69),
.Y(n_1648)
);

CKINVDCx5p33_ASAP7_75t_R g1649 ( 
.A(n_963),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_776),
.Y(n_1650)
);

CKINVDCx5p33_ASAP7_75t_R g1651 ( 
.A(n_129),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_199),
.Y(n_1652)
);

CKINVDCx5p33_ASAP7_75t_R g1653 ( 
.A(n_1010),
.Y(n_1653)
);

CKINVDCx5p33_ASAP7_75t_R g1654 ( 
.A(n_243),
.Y(n_1654)
);

CKINVDCx20_ASAP7_75t_R g1655 ( 
.A(n_70),
.Y(n_1655)
);

INVx3_ASAP7_75t_L g1656 ( 
.A(n_1065),
.Y(n_1656)
);

CKINVDCx5p33_ASAP7_75t_R g1657 ( 
.A(n_787),
.Y(n_1657)
);

INVx1_ASAP7_75t_SL g1658 ( 
.A(n_490),
.Y(n_1658)
);

CKINVDCx16_ASAP7_75t_R g1659 ( 
.A(n_1051),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_375),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_450),
.Y(n_1661)
);

CKINVDCx5p33_ASAP7_75t_R g1662 ( 
.A(n_105),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_57),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_79),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_272),
.Y(n_1665)
);

BUFx2_ASAP7_75t_L g1666 ( 
.A(n_1105),
.Y(n_1666)
);

CKINVDCx5p33_ASAP7_75t_R g1667 ( 
.A(n_1088),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_552),
.Y(n_1668)
);

CKINVDCx5p33_ASAP7_75t_R g1669 ( 
.A(n_332),
.Y(n_1669)
);

INVxp33_ASAP7_75t_SL g1670 ( 
.A(n_273),
.Y(n_1670)
);

CKINVDCx16_ASAP7_75t_R g1671 ( 
.A(n_1002),
.Y(n_1671)
);

CKINVDCx5p33_ASAP7_75t_R g1672 ( 
.A(n_263),
.Y(n_1672)
);

CKINVDCx5p33_ASAP7_75t_R g1673 ( 
.A(n_101),
.Y(n_1673)
);

CKINVDCx5p33_ASAP7_75t_R g1674 ( 
.A(n_813),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_791),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_499),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_825),
.Y(n_1677)
);

CKINVDCx5p33_ASAP7_75t_R g1678 ( 
.A(n_269),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_303),
.Y(n_1679)
);

CKINVDCx5p33_ASAP7_75t_R g1680 ( 
.A(n_902),
.Y(n_1680)
);

CKINVDCx5p33_ASAP7_75t_R g1681 ( 
.A(n_34),
.Y(n_1681)
);

CKINVDCx5p33_ASAP7_75t_R g1682 ( 
.A(n_0),
.Y(n_1682)
);

INVxp67_ASAP7_75t_L g1683 ( 
.A(n_1048),
.Y(n_1683)
);

BUFx3_ASAP7_75t_L g1684 ( 
.A(n_1085),
.Y(n_1684)
);

CKINVDCx5p33_ASAP7_75t_R g1685 ( 
.A(n_176),
.Y(n_1685)
);

BUFx2_ASAP7_75t_L g1686 ( 
.A(n_525),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_949),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_539),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_68),
.Y(n_1689)
);

CKINVDCx5p33_ASAP7_75t_R g1690 ( 
.A(n_1068),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1077),
.Y(n_1691)
);

CKINVDCx20_ASAP7_75t_R g1692 ( 
.A(n_1099),
.Y(n_1692)
);

BUFx3_ASAP7_75t_L g1693 ( 
.A(n_99),
.Y(n_1693)
);

BUFx2_ASAP7_75t_L g1694 ( 
.A(n_1076),
.Y(n_1694)
);

INVx1_ASAP7_75t_SL g1695 ( 
.A(n_752),
.Y(n_1695)
);

CKINVDCx5p33_ASAP7_75t_R g1696 ( 
.A(n_1064),
.Y(n_1696)
);

CKINVDCx5p33_ASAP7_75t_R g1697 ( 
.A(n_221),
.Y(n_1697)
);

CKINVDCx5p33_ASAP7_75t_R g1698 ( 
.A(n_121),
.Y(n_1698)
);

BUFx10_ASAP7_75t_L g1699 ( 
.A(n_262),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1083),
.Y(n_1700)
);

CKINVDCx5p33_ASAP7_75t_R g1701 ( 
.A(n_242),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_324),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_722),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_929),
.Y(n_1704)
);

CKINVDCx5p33_ASAP7_75t_R g1705 ( 
.A(n_303),
.Y(n_1705)
);

CKINVDCx5p33_ASAP7_75t_R g1706 ( 
.A(n_825),
.Y(n_1706)
);

BUFx5_ASAP7_75t_L g1707 ( 
.A(n_1103),
.Y(n_1707)
);

CKINVDCx20_ASAP7_75t_R g1708 ( 
.A(n_9),
.Y(n_1708)
);

CKINVDCx5p33_ASAP7_75t_R g1709 ( 
.A(n_417),
.Y(n_1709)
);

BUFx6f_ASAP7_75t_L g1710 ( 
.A(n_193),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_649),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_802),
.Y(n_1712)
);

CKINVDCx5p33_ASAP7_75t_R g1713 ( 
.A(n_350),
.Y(n_1713)
);

INVxp33_ASAP7_75t_R g1714 ( 
.A(n_340),
.Y(n_1714)
);

CKINVDCx5p33_ASAP7_75t_R g1715 ( 
.A(n_1004),
.Y(n_1715)
);

CKINVDCx5p33_ASAP7_75t_R g1716 ( 
.A(n_863),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_330),
.Y(n_1717)
);

CKINVDCx5p33_ASAP7_75t_R g1718 ( 
.A(n_339),
.Y(n_1718)
);

CKINVDCx5p33_ASAP7_75t_R g1719 ( 
.A(n_90),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1083),
.Y(n_1720)
);

INVx1_ASAP7_75t_SL g1721 ( 
.A(n_528),
.Y(n_1721)
);

CKINVDCx5p33_ASAP7_75t_R g1722 ( 
.A(n_585),
.Y(n_1722)
);

CKINVDCx5p33_ASAP7_75t_R g1723 ( 
.A(n_1003),
.Y(n_1723)
);

CKINVDCx5p33_ASAP7_75t_R g1724 ( 
.A(n_532),
.Y(n_1724)
);

CKINVDCx5p33_ASAP7_75t_R g1725 ( 
.A(n_278),
.Y(n_1725)
);

CKINVDCx5p33_ASAP7_75t_R g1726 ( 
.A(n_270),
.Y(n_1726)
);

CKINVDCx5p33_ASAP7_75t_R g1727 ( 
.A(n_914),
.Y(n_1727)
);

CKINVDCx5p33_ASAP7_75t_R g1728 ( 
.A(n_684),
.Y(n_1728)
);

INVx1_ASAP7_75t_SL g1729 ( 
.A(n_549),
.Y(n_1729)
);

CKINVDCx5p33_ASAP7_75t_R g1730 ( 
.A(n_11),
.Y(n_1730)
);

CKINVDCx5p33_ASAP7_75t_R g1731 ( 
.A(n_1049),
.Y(n_1731)
);

CKINVDCx20_ASAP7_75t_R g1732 ( 
.A(n_602),
.Y(n_1732)
);

CKINVDCx5p33_ASAP7_75t_R g1733 ( 
.A(n_968),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_650),
.Y(n_1734)
);

CKINVDCx5p33_ASAP7_75t_R g1735 ( 
.A(n_120),
.Y(n_1735)
);

CKINVDCx5p33_ASAP7_75t_R g1736 ( 
.A(n_727),
.Y(n_1736)
);

INVxp67_ASAP7_75t_L g1737 ( 
.A(n_430),
.Y(n_1737)
);

INVx1_ASAP7_75t_SL g1738 ( 
.A(n_779),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_215),
.Y(n_1739)
);

CKINVDCx5p33_ASAP7_75t_R g1740 ( 
.A(n_56),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_477),
.Y(n_1741)
);

CKINVDCx20_ASAP7_75t_R g1742 ( 
.A(n_870),
.Y(n_1742)
);

CKINVDCx5p33_ASAP7_75t_R g1743 ( 
.A(n_125),
.Y(n_1743)
);

CKINVDCx5p33_ASAP7_75t_R g1744 ( 
.A(n_218),
.Y(n_1744)
);

CKINVDCx5p33_ASAP7_75t_R g1745 ( 
.A(n_1075),
.Y(n_1745)
);

CKINVDCx5p33_ASAP7_75t_R g1746 ( 
.A(n_899),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_594),
.Y(n_1747)
);

CKINVDCx5p33_ASAP7_75t_R g1748 ( 
.A(n_237),
.Y(n_1748)
);

BUFx2_ASAP7_75t_L g1749 ( 
.A(n_895),
.Y(n_1749)
);

CKINVDCx5p33_ASAP7_75t_R g1750 ( 
.A(n_740),
.Y(n_1750)
);

CKINVDCx20_ASAP7_75t_R g1751 ( 
.A(n_919),
.Y(n_1751)
);

CKINVDCx20_ASAP7_75t_R g1752 ( 
.A(n_405),
.Y(n_1752)
);

CKINVDCx5p33_ASAP7_75t_R g1753 ( 
.A(n_61),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_0),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1120),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1120),
.Y(n_1756)
);

INVxp33_ASAP7_75t_SL g1757 ( 
.A(n_1604),
.Y(n_1757)
);

INVxp33_ASAP7_75t_L g1758 ( 
.A(n_1178),
.Y(n_1758)
);

CKINVDCx5p33_ASAP7_75t_R g1759 ( 
.A(n_1178),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1120),
.Y(n_1760)
);

CKINVDCx20_ASAP7_75t_R g1761 ( 
.A(n_1333),
.Y(n_1761)
);

INVxp67_ASAP7_75t_L g1762 ( 
.A(n_1128),
.Y(n_1762)
);

CKINVDCx5p33_ASAP7_75t_R g1763 ( 
.A(n_1333),
.Y(n_1763)
);

INVxp33_ASAP7_75t_L g1764 ( 
.A(n_1299),
.Y(n_1764)
);

BUFx6f_ASAP7_75t_L g1765 ( 
.A(n_1157),
.Y(n_1765)
);

CKINVDCx20_ASAP7_75t_R g1766 ( 
.A(n_1395),
.Y(n_1766)
);

CKINVDCx20_ASAP7_75t_R g1767 ( 
.A(n_1395),
.Y(n_1767)
);

HB1xp67_ASAP7_75t_L g1768 ( 
.A(n_1230),
.Y(n_1768)
);

OR2x2_ASAP7_75t_L g1769 ( 
.A(n_1583),
.B(n_0),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1321),
.Y(n_1770)
);

INVxp67_ASAP7_75t_SL g1771 ( 
.A(n_1376),
.Y(n_1771)
);

BUFx10_ASAP7_75t_L g1772 ( 
.A(n_1753),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1497),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1497),
.Y(n_1774)
);

NOR2xp33_ASAP7_75t_L g1775 ( 
.A(n_1670),
.B(n_0),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1497),
.Y(n_1776)
);

CKINVDCx16_ASAP7_75t_R g1777 ( 
.A(n_1190),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1699),
.Y(n_1778)
);

INVxp67_ASAP7_75t_L g1779 ( 
.A(n_1388),
.Y(n_1779)
);

INVxp67_ASAP7_75t_SL g1780 ( 
.A(n_1376),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1699),
.Y(n_1781)
);

INVxp67_ASAP7_75t_SL g1782 ( 
.A(n_1425),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1699),
.Y(n_1783)
);

CKINVDCx5p33_ASAP7_75t_R g1784 ( 
.A(n_1557),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1412),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1483),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1152),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1163),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1164),
.Y(n_1789)
);

CKINVDCx14_ASAP7_75t_R g1790 ( 
.A(n_1557),
.Y(n_1790)
);

CKINVDCx5p33_ASAP7_75t_R g1791 ( 
.A(n_1613),
.Y(n_1791)
);

CKINVDCx5p33_ASAP7_75t_R g1792 ( 
.A(n_1613),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1174),
.Y(n_1793)
);

INVxp33_ASAP7_75t_SL g1794 ( 
.A(n_1463),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1203),
.Y(n_1795)
);

CKINVDCx16_ASAP7_75t_R g1796 ( 
.A(n_1336),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1308),
.Y(n_1797)
);

CKINVDCx16_ASAP7_75t_R g1798 ( 
.A(n_1354),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1330),
.Y(n_1799)
);

INVxp67_ASAP7_75t_SL g1800 ( 
.A(n_1425),
.Y(n_1800)
);

CKINVDCx5p33_ASAP7_75t_R g1801 ( 
.A(n_1122),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1355),
.Y(n_1802)
);

INVxp67_ASAP7_75t_SL g1803 ( 
.A(n_1693),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1374),
.Y(n_1804)
);

CKINVDCx20_ASAP7_75t_R g1805 ( 
.A(n_1150),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1384),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1396),
.Y(n_1807)
);

CKINVDCx16_ASAP7_75t_R g1808 ( 
.A(n_1359),
.Y(n_1808)
);

CKINVDCx16_ASAP7_75t_R g1809 ( 
.A(n_1393),
.Y(n_1809)
);

INVx2_ASAP7_75t_L g1810 ( 
.A(n_1321),
.Y(n_1810)
);

INVxp67_ASAP7_75t_SL g1811 ( 
.A(n_1693),
.Y(n_1811)
);

INVx2_ASAP7_75t_L g1812 ( 
.A(n_1321),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1416),
.Y(n_1813)
);

CKINVDCx20_ASAP7_75t_R g1814 ( 
.A(n_1150),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1421),
.Y(n_1815)
);

CKINVDCx20_ASAP7_75t_R g1816 ( 
.A(n_1409),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1424),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1430),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1442),
.Y(n_1819)
);

BUFx6f_ASAP7_75t_L g1820 ( 
.A(n_1157),
.Y(n_1820)
);

CKINVDCx5p33_ASAP7_75t_R g1821 ( 
.A(n_1125),
.Y(n_1821)
);

HB1xp67_ASAP7_75t_L g1822 ( 
.A(n_1547),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1478),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1498),
.Y(n_1824)
);

CKINVDCx5p33_ASAP7_75t_R g1825 ( 
.A(n_1740),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1508),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1509),
.Y(n_1827)
);

HB1xp67_ASAP7_75t_L g1828 ( 
.A(n_1626),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1575),
.Y(n_1829)
);

CKINVDCx16_ASAP7_75t_R g1830 ( 
.A(n_1545),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1577),
.Y(n_1831)
);

INVx2_ASAP7_75t_L g1832 ( 
.A(n_1321),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1600),
.Y(n_1833)
);

INVxp67_ASAP7_75t_L g1834 ( 
.A(n_1231),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1608),
.Y(n_1835)
);

INVxp67_ASAP7_75t_SL g1836 ( 
.A(n_1656),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1621),
.Y(n_1837)
);

CKINVDCx20_ASAP7_75t_R g1838 ( 
.A(n_1409),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1321),
.Y(n_1839)
);

CKINVDCx5p33_ASAP7_75t_R g1840 ( 
.A(n_1130),
.Y(n_1840)
);

CKINVDCx5p33_ASAP7_75t_R g1841 ( 
.A(n_1132),
.Y(n_1841)
);

INVxp67_ASAP7_75t_SL g1842 ( 
.A(n_1656),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1635),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1636),
.Y(n_1844)
);

CKINVDCx16_ASAP7_75t_R g1845 ( 
.A(n_1614),
.Y(n_1845)
);

CKINVDCx20_ASAP7_75t_R g1846 ( 
.A(n_1441),
.Y(n_1846)
);

CKINVDCx16_ASAP7_75t_R g1847 ( 
.A(n_1659),
.Y(n_1847)
);

INVxp67_ASAP7_75t_L g1848 ( 
.A(n_1254),
.Y(n_1848)
);

CKINVDCx20_ASAP7_75t_R g1849 ( 
.A(n_1441),
.Y(n_1849)
);

INVxp67_ASAP7_75t_SL g1850 ( 
.A(n_1656),
.Y(n_1850)
);

CKINVDCx16_ASAP7_75t_R g1851 ( 
.A(n_1671),
.Y(n_1851)
);

NOR2xp33_ASAP7_75t_L g1852 ( 
.A(n_1436),
.B(n_1),
.Y(n_1852)
);

INVxp67_ASAP7_75t_L g1853 ( 
.A(n_1524),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1652),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1663),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1664),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1665),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1689),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1739),
.Y(n_1859)
);

INVxp33_ASAP7_75t_SL g1860 ( 
.A(n_1140),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1754),
.Y(n_1861)
);

CKINVDCx20_ASAP7_75t_R g1862 ( 
.A(n_1479),
.Y(n_1862)
);

INVx2_ASAP7_75t_L g1863 ( 
.A(n_1321),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1167),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1129),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1142),
.Y(n_1866)
);

CKINVDCx5p33_ASAP7_75t_R g1867 ( 
.A(n_1743),
.Y(n_1867)
);

INVxp67_ASAP7_75t_SL g1868 ( 
.A(n_1648),
.Y(n_1868)
);

INVxp67_ASAP7_75t_SL g1869 ( 
.A(n_1196),
.Y(n_1869)
);

CKINVDCx20_ASAP7_75t_R g1870 ( 
.A(n_1479),
.Y(n_1870)
);

BUFx3_ASAP7_75t_L g1871 ( 
.A(n_1321),
.Y(n_1871)
);

INVxp67_ASAP7_75t_SL g1872 ( 
.A(n_1196),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1227),
.Y(n_1873)
);

BUFx3_ASAP7_75t_L g1874 ( 
.A(n_1551),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1356),
.Y(n_1875)
);

CKINVDCx16_ASAP7_75t_R g1876 ( 
.A(n_1127),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1749),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1528),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1666),
.Y(n_1879)
);

INVx2_ASAP7_75t_L g1880 ( 
.A(n_1551),
.Y(n_1880)
);

INVx2_ASAP7_75t_L g1881 ( 
.A(n_1551),
.Y(n_1881)
);

INVx2_ASAP7_75t_L g1882 ( 
.A(n_1871),
.Y(n_1882)
);

AND2x2_ASAP7_75t_L g1883 ( 
.A(n_1762),
.B(n_1686),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_SL g1884 ( 
.A(n_1876),
.B(n_1551),
.Y(n_1884)
);

BUFx6f_ASAP7_75t_L g1885 ( 
.A(n_1765),
.Y(n_1885)
);

INVx2_ASAP7_75t_L g1886 ( 
.A(n_1874),
.Y(n_1886)
);

BUFx6f_ASAP7_75t_L g1887 ( 
.A(n_1765),
.Y(n_1887)
);

AND2x2_ASAP7_75t_L g1888 ( 
.A(n_1762),
.B(n_1694),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1782),
.Y(n_1889)
);

AOI22xp5_ASAP7_75t_L g1890 ( 
.A1(n_1757),
.A2(n_1655),
.B1(n_1619),
.B2(n_1148),
.Y(n_1890)
);

AND2x2_ASAP7_75t_L g1891 ( 
.A(n_1779),
.B(n_1127),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1782),
.Y(n_1892)
);

NOR2xp33_ASAP7_75t_L g1893 ( 
.A(n_1755),
.B(n_1205),
.Y(n_1893)
);

BUFx6f_ASAP7_75t_L g1894 ( 
.A(n_1765),
.Y(n_1894)
);

INVx2_ASAP7_75t_L g1895 ( 
.A(n_1770),
.Y(n_1895)
);

AND2x4_ASAP7_75t_L g1896 ( 
.A(n_1779),
.B(n_1124),
.Y(n_1896)
);

INVx4_ASAP7_75t_L g1897 ( 
.A(n_1772),
.Y(n_1897)
);

AOI22xp5_ASAP7_75t_L g1898 ( 
.A1(n_1794),
.A2(n_1848),
.B1(n_1853),
.B2(n_1834),
.Y(n_1898)
);

INVx2_ASAP7_75t_L g1899 ( 
.A(n_1810),
.Y(n_1899)
);

INVx2_ASAP7_75t_L g1900 ( 
.A(n_1812),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1811),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1811),
.Y(n_1902)
);

AND2x4_ASAP7_75t_L g1903 ( 
.A(n_1834),
.B(n_1124),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1771),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1868),
.B(n_1836),
.Y(n_1905)
);

OAI22x1_ASAP7_75t_L g1906 ( 
.A1(n_1759),
.A2(n_1714),
.B1(n_1162),
.B2(n_1170),
.Y(n_1906)
);

INVx2_ASAP7_75t_L g1907 ( 
.A(n_1832),
.Y(n_1907)
);

INVx2_ASAP7_75t_L g1908 ( 
.A(n_1839),
.Y(n_1908)
);

BUFx6f_ASAP7_75t_L g1909 ( 
.A(n_1820),
.Y(n_1909)
);

BUFx2_ASAP7_75t_L g1910 ( 
.A(n_1801),
.Y(n_1910)
);

AND2x4_ASAP7_75t_L g1911 ( 
.A(n_1848),
.B(n_1179),
.Y(n_1911)
);

CKINVDCx5p33_ASAP7_75t_R g1912 ( 
.A(n_1860),
.Y(n_1912)
);

INVx5_ASAP7_75t_L g1913 ( 
.A(n_1820),
.Y(n_1913)
);

INVx2_ASAP7_75t_L g1914 ( 
.A(n_1863),
.Y(n_1914)
);

HB1xp67_ASAP7_75t_L g1915 ( 
.A(n_1768),
.Y(n_1915)
);

INVx3_ASAP7_75t_L g1916 ( 
.A(n_1772),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1780),
.Y(n_1917)
);

INVx6_ASAP7_75t_L g1918 ( 
.A(n_1777),
.Y(n_1918)
);

AOI22xp5_ASAP7_75t_L g1919 ( 
.A1(n_1853),
.A2(n_1655),
.B1(n_1619),
.B2(n_1184),
.Y(n_1919)
);

BUFx6f_ASAP7_75t_L g1920 ( 
.A(n_1820),
.Y(n_1920)
);

INVxp67_ASAP7_75t_L g1921 ( 
.A(n_1822),
.Y(n_1921)
);

CKINVDCx14_ASAP7_75t_R g1922 ( 
.A(n_1790),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1800),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1803),
.Y(n_1924)
);

INVx2_ASAP7_75t_L g1925 ( 
.A(n_1880),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1842),
.Y(n_1926)
);

INVx2_ASAP7_75t_L g1927 ( 
.A(n_1881),
.Y(n_1927)
);

INVx3_ASAP7_75t_L g1928 ( 
.A(n_1864),
.Y(n_1928)
);

BUFx6f_ASAP7_75t_L g1929 ( 
.A(n_1787),
.Y(n_1929)
);

INVx2_ASAP7_75t_L g1930 ( 
.A(n_1865),
.Y(n_1930)
);

AOI22xp5_ASAP7_75t_L g1931 ( 
.A1(n_1766),
.A2(n_1186),
.B1(n_1208),
.B2(n_1144),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1850),
.Y(n_1932)
);

INVx2_ASAP7_75t_L g1933 ( 
.A(n_1866),
.Y(n_1933)
);

BUFx8_ASAP7_75t_SL g1934 ( 
.A(n_1761),
.Y(n_1934)
);

AOI22xp5_ASAP7_75t_L g1935 ( 
.A1(n_1767),
.A2(n_1222),
.B1(n_1233),
.B2(n_1217),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1756),
.B(n_1242),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1869),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1760),
.B(n_1249),
.Y(n_1938)
);

BUFx12f_ASAP7_75t_L g1939 ( 
.A(n_1763),
.Y(n_1939)
);

XNOR2xp5_ASAP7_75t_L g1940 ( 
.A(n_1805),
.B(n_1358),
.Y(n_1940)
);

OA21x2_ASAP7_75t_L g1941 ( 
.A1(n_1788),
.A2(n_1334),
.B(n_1282),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1872),
.Y(n_1942)
);

AND2x6_ASAP7_75t_L g1943 ( 
.A(n_1773),
.B(n_1179),
.Y(n_1943)
);

INVx2_ASAP7_75t_L g1944 ( 
.A(n_1873),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1875),
.Y(n_1945)
);

BUFx6f_ASAP7_75t_L g1946 ( 
.A(n_1789),
.Y(n_1946)
);

INVx3_ASAP7_75t_L g1947 ( 
.A(n_1774),
.Y(n_1947)
);

INVx3_ASAP7_75t_L g1948 ( 
.A(n_1776),
.Y(n_1948)
);

BUFx8_ASAP7_75t_SL g1949 ( 
.A(n_1814),
.Y(n_1949)
);

INVx3_ASAP7_75t_L g1950 ( 
.A(n_1778),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1793),
.Y(n_1951)
);

INVx5_ASAP7_75t_L g1952 ( 
.A(n_1796),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1795),
.Y(n_1953)
);

AND2x4_ASAP7_75t_L g1954 ( 
.A(n_1877),
.B(n_1341),
.Y(n_1954)
);

AOI22xp5_ASAP7_75t_L g1955 ( 
.A1(n_1764),
.A2(n_1259),
.B1(n_1286),
.B2(n_1279),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1781),
.B(n_1294),
.Y(n_1956)
);

OA21x2_ASAP7_75t_L g1957 ( 
.A1(n_1797),
.A2(n_1334),
.B(n_1282),
.Y(n_1957)
);

NOR2xp33_ASAP7_75t_L g1958 ( 
.A(n_1783),
.B(n_1488),
.Y(n_1958)
);

BUFx3_ASAP7_75t_L g1959 ( 
.A(n_1821),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1799),
.Y(n_1960)
);

AND2x4_ASAP7_75t_L g1961 ( 
.A(n_1878),
.B(n_1341),
.Y(n_1961)
);

OAI22xp5_ASAP7_75t_L g1962 ( 
.A1(n_1798),
.A2(n_1306),
.B1(n_1325),
.B2(n_1313),
.Y(n_1962)
);

AND2x2_ASAP7_75t_L g1963 ( 
.A(n_1828),
.B(n_1127),
.Y(n_1963)
);

AO22x1_ASAP7_75t_L g1964 ( 
.A1(n_1758),
.A2(n_1329),
.B1(n_1337),
.B2(n_1328),
.Y(n_1964)
);

AND2x4_ASAP7_75t_L g1965 ( 
.A(n_1879),
.B(n_1344),
.Y(n_1965)
);

INVx2_ASAP7_75t_L g1966 ( 
.A(n_1802),
.Y(n_1966)
);

AND2x4_ASAP7_75t_L g1967 ( 
.A(n_1785),
.B(n_1344),
.Y(n_1967)
);

OAI22xp5_ASAP7_75t_SL g1968 ( 
.A1(n_1816),
.A2(n_1362),
.B1(n_1379),
.B2(n_1358),
.Y(n_1968)
);

INVx2_ASAP7_75t_L g1969 ( 
.A(n_1804),
.Y(n_1969)
);

AOI22xp5_ASAP7_75t_L g1970 ( 
.A1(n_1825),
.A2(n_1841),
.B1(n_1867),
.B2(n_1840),
.Y(n_1970)
);

BUFx6f_ASAP7_75t_L g1971 ( 
.A(n_1806),
.Y(n_1971)
);

INVx5_ASAP7_75t_L g1972 ( 
.A(n_1808),
.Y(n_1972)
);

OA21x2_ASAP7_75t_L g1973 ( 
.A1(n_1807),
.A2(n_1525),
.B(n_1377),
.Y(n_1973)
);

AND2x4_ASAP7_75t_L g1974 ( 
.A(n_1786),
.B(n_1363),
.Y(n_1974)
);

CKINVDCx6p67_ASAP7_75t_R g1975 ( 
.A(n_1809),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_L g1976 ( 
.A(n_1813),
.B(n_1369),
.Y(n_1976)
);

AND2x4_ASAP7_75t_L g1977 ( 
.A(n_1784),
.B(n_1363),
.Y(n_1977)
);

NOR2xp33_ASAP7_75t_L g1978 ( 
.A(n_1791),
.B(n_1506),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1815),
.Y(n_1979)
);

AND2x4_ASAP7_75t_L g1980 ( 
.A(n_1792),
.B(n_1418),
.Y(n_1980)
);

INVx2_ASAP7_75t_L g1981 ( 
.A(n_1817),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1818),
.Y(n_1982)
);

OA21x2_ASAP7_75t_L g1983 ( 
.A1(n_1819),
.A2(n_1525),
.B(n_1377),
.Y(n_1983)
);

BUFx6f_ASAP7_75t_L g1984 ( 
.A(n_1823),
.Y(n_1984)
);

INVx2_ASAP7_75t_L g1985 ( 
.A(n_1824),
.Y(n_1985)
);

NAND2xp33_ASAP7_75t_L g1986 ( 
.A(n_1826),
.B(n_1551),
.Y(n_1986)
);

INVx2_ASAP7_75t_L g1987 ( 
.A(n_1827),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1829),
.Y(n_1988)
);

INVx2_ASAP7_75t_L g1989 ( 
.A(n_1831),
.Y(n_1989)
);

CKINVDCx16_ASAP7_75t_R g1990 ( 
.A(n_1830),
.Y(n_1990)
);

INVx3_ASAP7_75t_L g1991 ( 
.A(n_1833),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1835),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1837),
.Y(n_1993)
);

INVx2_ASAP7_75t_L g1994 ( 
.A(n_1843),
.Y(n_1994)
);

INVx2_ASAP7_75t_L g1995 ( 
.A(n_1844),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_L g1996 ( 
.A(n_1854),
.B(n_1372),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1855),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1856),
.Y(n_1998)
);

OAI22xp5_ASAP7_75t_L g1999 ( 
.A1(n_1845),
.A2(n_1381),
.B1(n_1383),
.B2(n_1382),
.Y(n_1999)
);

BUFx6f_ASAP7_75t_L g2000 ( 
.A(n_1857),
.Y(n_2000)
);

BUFx6f_ASAP7_75t_L g2001 ( 
.A(n_1858),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1859),
.Y(n_2002)
);

AND2x4_ASAP7_75t_L g2003 ( 
.A(n_1769),
.B(n_1418),
.Y(n_2003)
);

HB1xp67_ASAP7_75t_L g2004 ( 
.A(n_1847),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_L g2005 ( 
.A(n_1861),
.B(n_1852),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1775),
.Y(n_2006)
);

AOI22xp5_ASAP7_75t_L g2007 ( 
.A1(n_1851),
.A2(n_1390),
.B1(n_1398),
.B2(n_1385),
.Y(n_2007)
);

AND2x6_ASAP7_75t_L g2008 ( 
.A(n_1838),
.B(n_1486),
.Y(n_2008)
);

HB1xp67_ASAP7_75t_L g2009 ( 
.A(n_1846),
.Y(n_2009)
);

INVx2_ASAP7_75t_L g2010 ( 
.A(n_1849),
.Y(n_2010)
);

BUFx3_ASAP7_75t_L g2011 ( 
.A(n_1862),
.Y(n_2011)
);

BUFx6f_ASAP7_75t_L g2012 ( 
.A(n_1870),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1782),
.Y(n_2013)
);

BUFx12f_ASAP7_75t_L g2014 ( 
.A(n_1759),
.Y(n_2014)
);

OAI21x1_ASAP7_75t_L g2015 ( 
.A1(n_1787),
.A2(n_1592),
.B(n_1538),
.Y(n_2015)
);

BUFx6f_ASAP7_75t_L g2016 ( 
.A(n_1765),
.Y(n_2016)
);

OAI21x1_ASAP7_75t_L g2017 ( 
.A1(n_1787),
.A2(n_1592),
.B(n_1538),
.Y(n_2017)
);

BUFx6f_ASAP7_75t_L g2018 ( 
.A(n_1765),
.Y(n_2018)
);

AND2x2_ASAP7_75t_L g2019 ( 
.A(n_1762),
.B(n_1139),
.Y(n_2019)
);

INVx2_ASAP7_75t_L g2020 ( 
.A(n_1871),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_L g2021 ( 
.A(n_1762),
.B(n_1403),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1782),
.Y(n_2022)
);

BUFx6f_ASAP7_75t_L g2023 ( 
.A(n_1765),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1782),
.Y(n_2024)
);

INVx2_ASAP7_75t_L g2025 ( 
.A(n_1871),
.Y(n_2025)
);

INVx6_ASAP7_75t_L g2026 ( 
.A(n_1876),
.Y(n_2026)
);

INVx3_ASAP7_75t_L g2027 ( 
.A(n_1772),
.Y(n_2027)
);

INVx2_ASAP7_75t_L g2028 ( 
.A(n_1871),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1782),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1782),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1782),
.Y(n_2031)
);

BUFx6f_ASAP7_75t_L g2032 ( 
.A(n_1765),
.Y(n_2032)
);

AND2x2_ASAP7_75t_L g2033 ( 
.A(n_1762),
.B(n_1139),
.Y(n_2033)
);

INVx2_ASAP7_75t_L g2034 ( 
.A(n_1871),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1782),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_1782),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_1782),
.Y(n_2037)
);

BUFx6f_ASAP7_75t_L g2038 ( 
.A(n_1765),
.Y(n_2038)
);

AND2x4_ASAP7_75t_L g2039 ( 
.A(n_1762),
.B(n_1486),
.Y(n_2039)
);

NAND2xp5_ASAP7_75t_L g2040 ( 
.A(n_1762),
.B(n_1408),
.Y(n_2040)
);

NAND2xp5_ASAP7_75t_L g2041 ( 
.A(n_1762),
.B(n_1413),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1782),
.Y(n_2042)
);

INVx2_ASAP7_75t_L g2043 ( 
.A(n_1871),
.Y(n_2043)
);

CKINVDCx16_ASAP7_75t_R g2044 ( 
.A(n_1876),
.Y(n_2044)
);

OAI22xp5_ASAP7_75t_L g2045 ( 
.A1(n_1762),
.A2(n_1415),
.B1(n_1431),
.B2(n_1422),
.Y(n_2045)
);

HB1xp67_ASAP7_75t_L g2046 ( 
.A(n_1768),
.Y(n_2046)
);

OA21x2_ASAP7_75t_L g2047 ( 
.A1(n_1787),
.A2(n_1624),
.B(n_1616),
.Y(n_2047)
);

NAND2xp33_ASAP7_75t_L g2048 ( 
.A(n_1784),
.B(n_1551),
.Y(n_2048)
);

INVxp67_ASAP7_75t_L g2049 ( 
.A(n_1768),
.Y(n_2049)
);

CKINVDCx8_ASAP7_75t_R g2050 ( 
.A(n_1759),
.Y(n_2050)
);

INVx2_ASAP7_75t_L g2051 ( 
.A(n_1871),
.Y(n_2051)
);

HB1xp67_ASAP7_75t_L g2052 ( 
.A(n_1768),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1782),
.Y(n_2053)
);

INVx6_ASAP7_75t_L g2054 ( 
.A(n_1876),
.Y(n_2054)
);

AND2x2_ASAP7_75t_L g2055 ( 
.A(n_1762),
.B(n_1139),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_1782),
.Y(n_2056)
);

CKINVDCx5p33_ASAP7_75t_R g2057 ( 
.A(n_1860),
.Y(n_2057)
);

NAND2xp5_ASAP7_75t_L g2058 ( 
.A(n_1762),
.B(n_1451),
.Y(n_2058)
);

BUFx6f_ASAP7_75t_L g2059 ( 
.A(n_1765),
.Y(n_2059)
);

BUFx12f_ASAP7_75t_L g2060 ( 
.A(n_1759),
.Y(n_2060)
);

INVx2_ASAP7_75t_L g2061 ( 
.A(n_1871),
.Y(n_2061)
);

AND2x6_ASAP7_75t_L g2062 ( 
.A(n_1755),
.B(n_1555),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_1782),
.Y(n_2063)
);

INVx2_ASAP7_75t_L g2064 ( 
.A(n_1871),
.Y(n_2064)
);

OAI22xp5_ASAP7_75t_L g2065 ( 
.A1(n_1762),
.A2(n_1455),
.B1(n_1465),
.B2(n_1462),
.Y(n_2065)
);

BUFx6f_ASAP7_75t_L g2066 ( 
.A(n_1765),
.Y(n_2066)
);

INVx2_ASAP7_75t_L g2067 ( 
.A(n_1871),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_1782),
.Y(n_2068)
);

OAI22x1_ASAP7_75t_SL g2069 ( 
.A1(n_1805),
.A2(n_1379),
.B1(n_1404),
.B2(n_1362),
.Y(n_2069)
);

BUFx6f_ASAP7_75t_L g2070 ( 
.A(n_1765),
.Y(n_2070)
);

AND2x4_ASAP7_75t_L g2071 ( 
.A(n_1762),
.B(n_1555),
.Y(n_2071)
);

INVx6_ASAP7_75t_L g2072 ( 
.A(n_1876),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_1782),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_1782),
.Y(n_2074)
);

BUFx3_ASAP7_75t_L g2075 ( 
.A(n_1772),
.Y(n_2075)
);

NAND2xp5_ASAP7_75t_L g2076 ( 
.A(n_1762),
.B(n_1466),
.Y(n_2076)
);

INVx2_ASAP7_75t_L g2077 ( 
.A(n_1871),
.Y(n_2077)
);

OAI21x1_ASAP7_75t_L g2078 ( 
.A1(n_1787),
.A2(n_1624),
.B(n_1616),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_L g2079 ( 
.A(n_1762),
.B(n_1481),
.Y(n_2079)
);

INVx2_ASAP7_75t_L g2080 ( 
.A(n_1871),
.Y(n_2080)
);

AND2x2_ASAP7_75t_L g2081 ( 
.A(n_1762),
.B(n_1161),
.Y(n_2081)
);

BUFx6f_ASAP7_75t_L g2082 ( 
.A(n_1765),
.Y(n_2082)
);

BUFx6f_ASAP7_75t_L g2083 ( 
.A(n_1765),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_1782),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_1782),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_1782),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_1782),
.Y(n_2087)
);

INVx2_ASAP7_75t_L g2088 ( 
.A(n_1871),
.Y(n_2088)
);

AND2x2_ASAP7_75t_L g2089 ( 
.A(n_1762),
.B(n_1161),
.Y(n_2089)
);

OA21x2_ASAP7_75t_L g2090 ( 
.A1(n_1787),
.A2(n_1147),
.B(n_1131),
.Y(n_2090)
);

INVx2_ASAP7_75t_L g2091 ( 
.A(n_1871),
.Y(n_2091)
);

INVx2_ASAP7_75t_L g2092 ( 
.A(n_1871),
.Y(n_2092)
);

AND2x2_ASAP7_75t_L g2093 ( 
.A(n_1762),
.B(n_1161),
.Y(n_2093)
);

INVx2_ASAP7_75t_L g2094 ( 
.A(n_1871),
.Y(n_2094)
);

BUFx3_ASAP7_75t_L g2095 ( 
.A(n_1772),
.Y(n_2095)
);

BUFx6f_ASAP7_75t_L g2096 ( 
.A(n_1765),
.Y(n_2096)
);

INVx2_ASAP7_75t_L g2097 ( 
.A(n_1871),
.Y(n_2097)
);

BUFx12f_ASAP7_75t_L g2098 ( 
.A(n_1759),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_1782),
.Y(n_2099)
);

INVx2_ASAP7_75t_L g2100 ( 
.A(n_1871),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_1782),
.Y(n_2101)
);

AND2x2_ASAP7_75t_L g2102 ( 
.A(n_1762),
.B(n_1210),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_1782),
.Y(n_2103)
);

AND2x4_ASAP7_75t_L g2104 ( 
.A(n_1762),
.B(n_1684),
.Y(n_2104)
);

CKINVDCx5p33_ASAP7_75t_R g2105 ( 
.A(n_1949),
.Y(n_2105)
);

NOR2xp33_ASAP7_75t_R g2106 ( 
.A(n_1922),
.B(n_1257),
.Y(n_2106)
);

NOR2xp33_ASAP7_75t_R g2107 ( 
.A(n_1912),
.B(n_1291),
.Y(n_2107)
);

CKINVDCx5p33_ASAP7_75t_R g2108 ( 
.A(n_2057),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_L g2109 ( 
.A(n_1976),
.B(n_1482),
.Y(n_2109)
);

INVx2_ASAP7_75t_L g2110 ( 
.A(n_2015),
.Y(n_2110)
);

INVx2_ASAP7_75t_L g2111 ( 
.A(n_2017),
.Y(n_2111)
);

CKINVDCx5p33_ASAP7_75t_R g2112 ( 
.A(n_1934),
.Y(n_2112)
);

CKINVDCx5p33_ASAP7_75t_R g2113 ( 
.A(n_1975),
.Y(n_2113)
);

CKINVDCx5p33_ASAP7_75t_R g2114 ( 
.A(n_2044),
.Y(n_2114)
);

CKINVDCx5p33_ASAP7_75t_R g2115 ( 
.A(n_1990),
.Y(n_2115)
);

CKINVDCx5p33_ASAP7_75t_R g2116 ( 
.A(n_2026),
.Y(n_2116)
);

CKINVDCx5p33_ASAP7_75t_R g2117 ( 
.A(n_2026),
.Y(n_2117)
);

CKINVDCx5p33_ASAP7_75t_R g2118 ( 
.A(n_2054),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_1930),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_1933),
.Y(n_2120)
);

BUFx3_ASAP7_75t_L g2121 ( 
.A(n_2075),
.Y(n_2121)
);

CKINVDCx5p33_ASAP7_75t_R g2122 ( 
.A(n_2054),
.Y(n_2122)
);

CKINVDCx5p33_ASAP7_75t_R g2123 ( 
.A(n_2072),
.Y(n_2123)
);

AO22x2_ASAP7_75t_L g2124 ( 
.A1(n_1968),
.A2(n_1489),
.B1(n_1521),
.B2(n_1404),
.Y(n_2124)
);

CKINVDCx5p33_ASAP7_75t_R g2125 ( 
.A(n_2072),
.Y(n_2125)
);

BUFx3_ASAP7_75t_L g2126 ( 
.A(n_2095),
.Y(n_2126)
);

CKINVDCx20_ASAP7_75t_R g2127 ( 
.A(n_1910),
.Y(n_2127)
);

CKINVDCx20_ASAP7_75t_R g2128 ( 
.A(n_1910),
.Y(n_2128)
);

INVx2_ASAP7_75t_L g2129 ( 
.A(n_2078),
.Y(n_2129)
);

CKINVDCx20_ASAP7_75t_R g2130 ( 
.A(n_1940),
.Y(n_2130)
);

NOR2xp33_ASAP7_75t_R g2131 ( 
.A(n_2050),
.B(n_1708),
.Y(n_2131)
);

CKINVDCx5p33_ASAP7_75t_R g2132 ( 
.A(n_1939),
.Y(n_2132)
);

CKINVDCx5p33_ASAP7_75t_R g2133 ( 
.A(n_2014),
.Y(n_2133)
);

CKINVDCx5p33_ASAP7_75t_R g2134 ( 
.A(n_2060),
.Y(n_2134)
);

CKINVDCx5p33_ASAP7_75t_R g2135 ( 
.A(n_2098),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_1944),
.Y(n_2136)
);

CKINVDCx5p33_ASAP7_75t_R g2137 ( 
.A(n_1940),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_1928),
.Y(n_2138)
);

INVx2_ASAP7_75t_L g2139 ( 
.A(n_1957),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_1991),
.Y(n_2140)
);

CKINVDCx5p33_ASAP7_75t_R g2141 ( 
.A(n_2011),
.Y(n_2141)
);

CKINVDCx5p33_ASAP7_75t_R g2142 ( 
.A(n_2004),
.Y(n_2142)
);

CKINVDCx5p33_ASAP7_75t_R g2143 ( 
.A(n_1897),
.Y(n_2143)
);

CKINVDCx5p33_ASAP7_75t_R g2144 ( 
.A(n_2069),
.Y(n_2144)
);

AOI22xp5_ASAP7_75t_L g2145 ( 
.A1(n_1891),
.A2(n_1487),
.B1(n_1490),
.B2(n_1484),
.Y(n_2145)
);

CKINVDCx5p33_ASAP7_75t_R g2146 ( 
.A(n_1959),
.Y(n_2146)
);

CKINVDCx5p33_ASAP7_75t_R g2147 ( 
.A(n_1890),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_1937),
.Y(n_2148)
);

HB1xp67_ASAP7_75t_L g2149 ( 
.A(n_1921),
.Y(n_2149)
);

INVx2_ASAP7_75t_L g2150 ( 
.A(n_1973),
.Y(n_2150)
);

CKINVDCx5p33_ASAP7_75t_R g2151 ( 
.A(n_1918),
.Y(n_2151)
);

CKINVDCx5p33_ASAP7_75t_R g2152 ( 
.A(n_1918),
.Y(n_2152)
);

CKINVDCx5p33_ASAP7_75t_R g2153 ( 
.A(n_2009),
.Y(n_2153)
);

BUFx10_ASAP7_75t_L g2154 ( 
.A(n_1978),
.Y(n_2154)
);

CKINVDCx20_ASAP7_75t_R g2155 ( 
.A(n_1915),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_1942),
.Y(n_2156)
);

NOR2xp33_ASAP7_75t_L g2157 ( 
.A(n_1947),
.B(n_1683),
.Y(n_2157)
);

NOR2xp33_ASAP7_75t_R g2158 ( 
.A(n_1916),
.B(n_1489),
.Y(n_2158)
);

CKINVDCx5p33_ASAP7_75t_R g2159 ( 
.A(n_1952),
.Y(n_2159)
);

NOR2xp33_ASAP7_75t_R g2160 ( 
.A(n_2027),
.B(n_1521),
.Y(n_2160)
);

CKINVDCx5p33_ASAP7_75t_R g2161 ( 
.A(n_1952),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_1945),
.Y(n_2162)
);

CKINVDCx5p33_ASAP7_75t_R g2163 ( 
.A(n_1972),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_1941),
.Y(n_2164)
);

CKINVDCx5p33_ASAP7_75t_R g2165 ( 
.A(n_1972),
.Y(n_2165)
);

HB1xp67_ASAP7_75t_L g2166 ( 
.A(n_2046),
.Y(n_2166)
);

INVx1_ASAP7_75t_SL g2167 ( 
.A(n_2052),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_1941),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_1889),
.Y(n_2169)
);

NOR2xp33_ASAP7_75t_R g2170 ( 
.A(n_2008),
.B(n_1531),
.Y(n_2170)
);

CKINVDCx5p33_ASAP7_75t_R g2171 ( 
.A(n_2012),
.Y(n_2171)
);

CKINVDCx5p33_ASAP7_75t_R g2172 ( 
.A(n_2012),
.Y(n_2172)
);

NOR2xp33_ASAP7_75t_R g2173 ( 
.A(n_2008),
.B(n_1531),
.Y(n_2173)
);

INVx1_ASAP7_75t_L g2174 ( 
.A(n_1892),
.Y(n_2174)
);

CKINVDCx5p33_ASAP7_75t_R g2175 ( 
.A(n_1962),
.Y(n_2175)
);

CKINVDCx5p33_ASAP7_75t_R g2176 ( 
.A(n_1999),
.Y(n_2176)
);

NOR2xp33_ASAP7_75t_R g2177 ( 
.A(n_2008),
.B(n_1534),
.Y(n_2177)
);

INVx3_ASAP7_75t_L g2178 ( 
.A(n_1948),
.Y(n_2178)
);

INVx8_ASAP7_75t_L g2179 ( 
.A(n_1943),
.Y(n_2179)
);

CKINVDCx5p33_ASAP7_75t_R g2180 ( 
.A(n_1919),
.Y(n_2180)
);

INVx2_ASAP7_75t_L g2181 ( 
.A(n_1983),
.Y(n_2181)
);

HB1xp67_ASAP7_75t_L g2182 ( 
.A(n_2049),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_1901),
.Y(n_2183)
);

NAND2xp33_ASAP7_75t_R g2184 ( 
.A(n_1891),
.B(n_1493),
.Y(n_2184)
);

NOR2xp33_ASAP7_75t_R g2185 ( 
.A(n_1963),
.B(n_1534),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_1902),
.Y(n_2186)
);

NOR2xp33_ASAP7_75t_L g2187 ( 
.A(n_1950),
.B(n_1737),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_2013),
.Y(n_2188)
);

CKINVDCx5p33_ASAP7_75t_R g2189 ( 
.A(n_2045),
.Y(n_2189)
);

CKINVDCx5p33_ASAP7_75t_R g2190 ( 
.A(n_2065),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_2022),
.Y(n_2191)
);

CKINVDCx5p33_ASAP7_75t_R g2192 ( 
.A(n_1970),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_2024),
.Y(n_2193)
);

CKINVDCx5p33_ASAP7_75t_R g2194 ( 
.A(n_1898),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_2029),
.Y(n_2195)
);

BUFx2_ASAP7_75t_L g2196 ( 
.A(n_1963),
.Y(n_2196)
);

CKINVDCx5p33_ASAP7_75t_R g2197 ( 
.A(n_1955),
.Y(n_2197)
);

NOR2xp33_ASAP7_75t_R g2198 ( 
.A(n_2019),
.B(n_1535),
.Y(n_2198)
);

NAND2xp5_ASAP7_75t_L g2199 ( 
.A(n_1996),
.B(n_1496),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_2030),
.Y(n_2200)
);

CKINVDCx20_ASAP7_75t_R g2201 ( 
.A(n_1931),
.Y(n_2201)
);

CKINVDCx5p33_ASAP7_75t_R g2202 ( 
.A(n_1964),
.Y(n_2202)
);

INVx2_ASAP7_75t_L g2203 ( 
.A(n_2047),
.Y(n_2203)
);

INVx2_ASAP7_75t_L g2204 ( 
.A(n_2090),
.Y(n_2204)
);

BUFx6f_ASAP7_75t_L g2205 ( 
.A(n_1929),
.Y(n_2205)
);

CKINVDCx5p33_ASAP7_75t_R g2206 ( 
.A(n_1935),
.Y(n_2206)
);

CKINVDCx20_ASAP7_75t_R g2207 ( 
.A(n_2007),
.Y(n_2207)
);

NOR2xp33_ASAP7_75t_R g2208 ( 
.A(n_2019),
.B(n_1535),
.Y(n_2208)
);

NOR2xp67_ASAP7_75t_L g2209 ( 
.A(n_1906),
.B(n_1),
.Y(n_2209)
);

CKINVDCx20_ASAP7_75t_R g2210 ( 
.A(n_1883),
.Y(n_2210)
);

CKINVDCx5p33_ASAP7_75t_R g2211 ( 
.A(n_1906),
.Y(n_2211)
);

HB1xp67_ASAP7_75t_L g2212 ( 
.A(n_2033),
.Y(n_2212)
);

CKINVDCx5p33_ASAP7_75t_R g2213 ( 
.A(n_1883),
.Y(n_2213)
);

CKINVDCx5p33_ASAP7_75t_R g2214 ( 
.A(n_1888),
.Y(n_2214)
);

NAND2xp33_ASAP7_75t_R g2215 ( 
.A(n_2033),
.B(n_1499),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_2031),
.Y(n_2216)
);

NAND2xp5_ASAP7_75t_L g2217 ( 
.A(n_2005),
.B(n_1503),
.Y(n_2217)
);

CKINVDCx5p33_ASAP7_75t_R g2218 ( 
.A(n_1888),
.Y(n_2218)
);

CKINVDCx5p33_ASAP7_75t_R g2219 ( 
.A(n_2010),
.Y(n_2219)
);

HB1xp67_ASAP7_75t_L g2220 ( 
.A(n_2055),
.Y(n_2220)
);

HB1xp67_ASAP7_75t_L g2221 ( 
.A(n_2055),
.Y(n_2221)
);

CKINVDCx5p33_ASAP7_75t_R g2222 ( 
.A(n_2081),
.Y(n_2222)
);

INVx2_ASAP7_75t_SL g2223 ( 
.A(n_2081),
.Y(n_2223)
);

NAND2xp33_ASAP7_75t_R g2224 ( 
.A(n_2089),
.B(n_1511),
.Y(n_2224)
);

CKINVDCx20_ASAP7_75t_R g2225 ( 
.A(n_2089),
.Y(n_2225)
);

BUFx3_ASAP7_75t_L g2226 ( 
.A(n_2003),
.Y(n_2226)
);

NOR2xp33_ASAP7_75t_R g2227 ( 
.A(n_2093),
.B(n_1537),
.Y(n_2227)
);

INVx2_ASAP7_75t_L g2228 ( 
.A(n_1929),
.Y(n_2228)
);

CKINVDCx5p33_ASAP7_75t_R g2229 ( 
.A(n_2093),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_2035),
.Y(n_2230)
);

CKINVDCx5p33_ASAP7_75t_R g2231 ( 
.A(n_2102),
.Y(n_2231)
);

CKINVDCx5p33_ASAP7_75t_R g2232 ( 
.A(n_2102),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_2036),
.Y(n_2233)
);

NOR2xp67_ASAP7_75t_L g2234 ( 
.A(n_2021),
.B(n_1),
.Y(n_2234)
);

NOR2xp67_ASAP7_75t_L g2235 ( 
.A(n_2040),
.B(n_1),
.Y(n_2235)
);

CKINVDCx5p33_ASAP7_75t_R g2236 ( 
.A(n_2041),
.Y(n_2236)
);

BUFx6f_ASAP7_75t_L g2237 ( 
.A(n_1946),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_2037),
.Y(n_2238)
);

CKINVDCx20_ASAP7_75t_R g2239 ( 
.A(n_2058),
.Y(n_2239)
);

NAND2xp5_ASAP7_75t_SL g2240 ( 
.A(n_2076),
.B(n_1513),
.Y(n_2240)
);

CKINVDCx5p33_ASAP7_75t_R g2241 ( 
.A(n_2079),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_2042),
.Y(n_2242)
);

CKINVDCx5p33_ASAP7_75t_R g2243 ( 
.A(n_1896),
.Y(n_2243)
);

CKINVDCx5p33_ASAP7_75t_R g2244 ( 
.A(n_2039),
.Y(n_2244)
);

INVx2_ASAP7_75t_L g2245 ( 
.A(n_1946),
.Y(n_2245)
);

BUFx10_ASAP7_75t_L g2246 ( 
.A(n_2071),
.Y(n_2246)
);

OA22x2_ASAP7_75t_L g2247 ( 
.A1(n_2006),
.A2(n_1117),
.B1(n_1118),
.B2(n_1116),
.Y(n_2247)
);

CKINVDCx5p33_ASAP7_75t_R g2248 ( 
.A(n_2104),
.Y(n_2248)
);

INVx1_ASAP7_75t_L g2249 ( 
.A(n_2053),
.Y(n_2249)
);

CKINVDCx20_ASAP7_75t_R g2250 ( 
.A(n_1905),
.Y(n_2250)
);

CKINVDCx5p33_ASAP7_75t_R g2251 ( 
.A(n_1903),
.Y(n_2251)
);

CKINVDCx5p33_ASAP7_75t_R g2252 ( 
.A(n_1911),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_2056),
.Y(n_2253)
);

CKINVDCx5p33_ASAP7_75t_R g2254 ( 
.A(n_1977),
.Y(n_2254)
);

CKINVDCx5p33_ASAP7_75t_R g2255 ( 
.A(n_1980),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_2063),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_2068),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_2073),
.Y(n_2258)
);

NOR2xp67_ASAP7_75t_L g2259 ( 
.A(n_1893),
.B(n_1958),
.Y(n_2259)
);

CKINVDCx5p33_ASAP7_75t_R g2260 ( 
.A(n_2074),
.Y(n_2260)
);

CKINVDCx5p33_ASAP7_75t_R g2261 ( 
.A(n_2084),
.Y(n_2261)
);

NOR2xp33_ASAP7_75t_R g2262 ( 
.A(n_2048),
.B(n_1537),
.Y(n_2262)
);

CKINVDCx5p33_ASAP7_75t_R g2263 ( 
.A(n_2085),
.Y(n_2263)
);

NAND2xp5_ASAP7_75t_L g2264 ( 
.A(n_2086),
.B(n_1514),
.Y(n_2264)
);

INVxp33_ASAP7_75t_L g2265 ( 
.A(n_1967),
.Y(n_2265)
);

NOR2xp33_ASAP7_75t_L g2266 ( 
.A(n_1926),
.B(n_1522),
.Y(n_2266)
);

CKINVDCx20_ASAP7_75t_R g2267 ( 
.A(n_1884),
.Y(n_2267)
);

CKINVDCx5p33_ASAP7_75t_R g2268 ( 
.A(n_2087),
.Y(n_2268)
);

NOR2xp33_ASAP7_75t_R g2269 ( 
.A(n_1943),
.B(n_2062),
.Y(n_2269)
);

INVx1_ASAP7_75t_L g2270 ( 
.A(n_2099),
.Y(n_2270)
);

CKINVDCx5p33_ASAP7_75t_R g2271 ( 
.A(n_2101),
.Y(n_2271)
);

CKINVDCx5p33_ASAP7_75t_R g2272 ( 
.A(n_2103),
.Y(n_2272)
);

CKINVDCx5p33_ASAP7_75t_R g2273 ( 
.A(n_1936),
.Y(n_2273)
);

CKINVDCx5p33_ASAP7_75t_R g2274 ( 
.A(n_1938),
.Y(n_2274)
);

INVx2_ASAP7_75t_L g2275 ( 
.A(n_1971),
.Y(n_2275)
);

INVx1_ASAP7_75t_L g2276 ( 
.A(n_1932),
.Y(n_2276)
);

NOR2xp33_ASAP7_75t_L g2277 ( 
.A(n_1904),
.B(n_1530),
.Y(n_2277)
);

CKINVDCx20_ASAP7_75t_R g2278 ( 
.A(n_1956),
.Y(n_2278)
);

INVx2_ASAP7_75t_L g2279 ( 
.A(n_1971),
.Y(n_2279)
);

CKINVDCx5p33_ASAP7_75t_R g2280 ( 
.A(n_1917),
.Y(n_2280)
);

CKINVDCx5p33_ASAP7_75t_R g2281 ( 
.A(n_1923),
.Y(n_2281)
);

CKINVDCx5p33_ASAP7_75t_R g2282 ( 
.A(n_1924),
.Y(n_2282)
);

CKINVDCx5p33_ASAP7_75t_R g2283 ( 
.A(n_1943),
.Y(n_2283)
);

NOR2xp33_ASAP7_75t_R g2284 ( 
.A(n_2062),
.B(n_1629),
.Y(n_2284)
);

INVx1_ASAP7_75t_L g2285 ( 
.A(n_1984),
.Y(n_2285)
);

CKINVDCx20_ASAP7_75t_R g2286 ( 
.A(n_1984),
.Y(n_2286)
);

CKINVDCx5p33_ASAP7_75t_R g2287 ( 
.A(n_2062),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_2000),
.Y(n_2288)
);

CKINVDCx5p33_ASAP7_75t_R g2289 ( 
.A(n_1974),
.Y(n_2289)
);

BUFx2_ASAP7_75t_L g2290 ( 
.A(n_1954),
.Y(n_2290)
);

INVx2_ASAP7_75t_L g2291 ( 
.A(n_2000),
.Y(n_2291)
);

CKINVDCx5p33_ASAP7_75t_R g2292 ( 
.A(n_1961),
.Y(n_2292)
);

INVx2_ASAP7_75t_L g2293 ( 
.A(n_2001),
.Y(n_2293)
);

CKINVDCx5p33_ASAP7_75t_R g2294 ( 
.A(n_1965),
.Y(n_2294)
);

BUFx6f_ASAP7_75t_L g2295 ( 
.A(n_2001),
.Y(n_2295)
);

CKINVDCx20_ASAP7_75t_R g2296 ( 
.A(n_1951),
.Y(n_2296)
);

CKINVDCx5p33_ASAP7_75t_R g2297 ( 
.A(n_1966),
.Y(n_2297)
);

NAND2xp5_ASAP7_75t_L g2298 ( 
.A(n_1953),
.B(n_1536),
.Y(n_2298)
);

CKINVDCx5p33_ASAP7_75t_R g2299 ( 
.A(n_1969),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_1981),
.Y(n_2300)
);

INVx3_ASAP7_75t_L g2301 ( 
.A(n_1985),
.Y(n_2301)
);

HB1xp67_ASAP7_75t_L g2302 ( 
.A(n_1987),
.Y(n_2302)
);

CKINVDCx5p33_ASAP7_75t_R g2303 ( 
.A(n_1989),
.Y(n_2303)
);

INVx2_ASAP7_75t_L g2304 ( 
.A(n_1994),
.Y(n_2304)
);

CKINVDCx5p33_ASAP7_75t_R g2305 ( 
.A(n_1995),
.Y(n_2305)
);

INVxp67_ASAP7_75t_L g2306 ( 
.A(n_1960),
.Y(n_2306)
);

CKINVDCx5p33_ASAP7_75t_R g2307 ( 
.A(n_1979),
.Y(n_2307)
);

CKINVDCx5p33_ASAP7_75t_R g2308 ( 
.A(n_1982),
.Y(n_2308)
);

INVx1_ASAP7_75t_L g2309 ( 
.A(n_1988),
.Y(n_2309)
);

INVx1_ASAP7_75t_L g2310 ( 
.A(n_1992),
.Y(n_2310)
);

CKINVDCx5p33_ASAP7_75t_R g2311 ( 
.A(n_1993),
.Y(n_2311)
);

NAND2xp5_ASAP7_75t_L g2312 ( 
.A(n_1997),
.B(n_1560),
.Y(n_2312)
);

CKINVDCx5p33_ASAP7_75t_R g2313 ( 
.A(n_1998),
.Y(n_2313)
);

CKINVDCx5p33_ASAP7_75t_R g2314 ( 
.A(n_2002),
.Y(n_2314)
);

CKINVDCx5p33_ASAP7_75t_R g2315 ( 
.A(n_1895),
.Y(n_2315)
);

CKINVDCx5p33_ASAP7_75t_R g2316 ( 
.A(n_1899),
.Y(n_2316)
);

NAND2xp33_ASAP7_75t_R g2317 ( 
.A(n_1900),
.B(n_1561),
.Y(n_2317)
);

NAND2xp33_ASAP7_75t_L g2318 ( 
.A(n_1882),
.B(n_1551),
.Y(n_2318)
);

INVxp67_ASAP7_75t_L g2319 ( 
.A(n_1986),
.Y(n_2319)
);

HB1xp67_ASAP7_75t_L g2320 ( 
.A(n_1907),
.Y(n_2320)
);

BUFx2_ASAP7_75t_L g2321 ( 
.A(n_1908),
.Y(n_2321)
);

CKINVDCx5p33_ASAP7_75t_R g2322 ( 
.A(n_1914),
.Y(n_2322)
);

CKINVDCx5p33_ASAP7_75t_R g2323 ( 
.A(n_1925),
.Y(n_2323)
);

CKINVDCx5p33_ASAP7_75t_R g2324 ( 
.A(n_1927),
.Y(n_2324)
);

CKINVDCx5p33_ASAP7_75t_R g2325 ( 
.A(n_1886),
.Y(n_2325)
);

BUFx2_ASAP7_75t_L g2326 ( 
.A(n_2020),
.Y(n_2326)
);

INVx2_ASAP7_75t_L g2327 ( 
.A(n_2025),
.Y(n_2327)
);

CKINVDCx5p33_ASAP7_75t_R g2328 ( 
.A(n_2028),
.Y(n_2328)
);

CKINVDCx20_ASAP7_75t_R g2329 ( 
.A(n_1913),
.Y(n_2329)
);

CKINVDCx5p33_ASAP7_75t_R g2330 ( 
.A(n_2034),
.Y(n_2330)
);

CKINVDCx5p33_ASAP7_75t_R g2331 ( 
.A(n_2043),
.Y(n_2331)
);

INVx1_ASAP7_75t_L g2332 ( 
.A(n_2051),
.Y(n_2332)
);

CKINVDCx5p33_ASAP7_75t_R g2333 ( 
.A(n_2061),
.Y(n_2333)
);

OAI21x1_ASAP7_75t_L g2334 ( 
.A1(n_2064),
.A2(n_1147),
.B(n_1131),
.Y(n_2334)
);

BUFx6f_ASAP7_75t_SL g2335 ( 
.A(n_1885),
.Y(n_2335)
);

CKINVDCx5p33_ASAP7_75t_R g2336 ( 
.A(n_2067),
.Y(n_2336)
);

BUFx6f_ASAP7_75t_L g2337 ( 
.A(n_1885),
.Y(n_2337)
);

INVx2_ASAP7_75t_L g2338 ( 
.A(n_2077),
.Y(n_2338)
);

BUFx6f_ASAP7_75t_L g2339 ( 
.A(n_1887),
.Y(n_2339)
);

CKINVDCx5p33_ASAP7_75t_R g2340 ( 
.A(n_2080),
.Y(n_2340)
);

NOR2xp33_ASAP7_75t_R g2341 ( 
.A(n_2088),
.B(n_1629),
.Y(n_2341)
);

CKINVDCx5p33_ASAP7_75t_R g2342 ( 
.A(n_2091),
.Y(n_2342)
);

CKINVDCx5p33_ASAP7_75t_R g2343 ( 
.A(n_2092),
.Y(n_2343)
);

INVx3_ASAP7_75t_L g2344 ( 
.A(n_2094),
.Y(n_2344)
);

NOR2xp33_ASAP7_75t_R g2345 ( 
.A(n_2097),
.B(n_1752),
.Y(n_2345)
);

CKINVDCx5p33_ASAP7_75t_R g2346 ( 
.A(n_2100),
.Y(n_2346)
);

INVx2_ASAP7_75t_L g2347 ( 
.A(n_1913),
.Y(n_2347)
);

CKINVDCx5p33_ASAP7_75t_R g2348 ( 
.A(n_1887),
.Y(n_2348)
);

INVx1_ASAP7_75t_L g2349 ( 
.A(n_1894),
.Y(n_2349)
);

INVx2_ASAP7_75t_L g2350 ( 
.A(n_1894),
.Y(n_2350)
);

CKINVDCx5p33_ASAP7_75t_R g2351 ( 
.A(n_1909),
.Y(n_2351)
);

NAND2xp33_ASAP7_75t_R g2352 ( 
.A(n_1909),
.B(n_1582),
.Y(n_2352)
);

CKINVDCx5p33_ASAP7_75t_R g2353 ( 
.A(n_1920),
.Y(n_2353)
);

INVx1_ASAP7_75t_L g2354 ( 
.A(n_1920),
.Y(n_2354)
);

NAND2xp5_ASAP7_75t_L g2355 ( 
.A(n_2016),
.B(n_1585),
.Y(n_2355)
);

INVx1_ASAP7_75t_L g2356 ( 
.A(n_2016),
.Y(n_2356)
);

HB1xp67_ASAP7_75t_L g2357 ( 
.A(n_2018),
.Y(n_2357)
);

INVx2_ASAP7_75t_L g2358 ( 
.A(n_2018),
.Y(n_2358)
);

CKINVDCx5p33_ASAP7_75t_R g2359 ( 
.A(n_2023),
.Y(n_2359)
);

BUFx6f_ASAP7_75t_L g2360 ( 
.A(n_2023),
.Y(n_2360)
);

NAND2xp33_ASAP7_75t_R g2361 ( 
.A(n_2032),
.B(n_1598),
.Y(n_2361)
);

CKINVDCx5p33_ASAP7_75t_R g2362 ( 
.A(n_2032),
.Y(n_2362)
);

BUFx6f_ASAP7_75t_L g2363 ( 
.A(n_2038),
.Y(n_2363)
);

CKINVDCx5p33_ASAP7_75t_R g2364 ( 
.A(n_2038),
.Y(n_2364)
);

CKINVDCx20_ASAP7_75t_R g2365 ( 
.A(n_2059),
.Y(n_2365)
);

CKINVDCx20_ASAP7_75t_R g2366 ( 
.A(n_2059),
.Y(n_2366)
);

CKINVDCx5p33_ASAP7_75t_R g2367 ( 
.A(n_2066),
.Y(n_2367)
);

CKINVDCx5p33_ASAP7_75t_R g2368 ( 
.A(n_2066),
.Y(n_2368)
);

CKINVDCx5p33_ASAP7_75t_R g2369 ( 
.A(n_2070),
.Y(n_2369)
);

NOR2xp33_ASAP7_75t_R g2370 ( 
.A(n_2070),
.B(n_1752),
.Y(n_2370)
);

CKINVDCx5p33_ASAP7_75t_R g2371 ( 
.A(n_2082),
.Y(n_2371)
);

BUFx3_ASAP7_75t_L g2372 ( 
.A(n_2082),
.Y(n_2372)
);

INVx1_ASAP7_75t_L g2373 ( 
.A(n_2083),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_2083),
.Y(n_2374)
);

NOR2xp33_ASAP7_75t_L g2375 ( 
.A(n_2096),
.B(n_1605),
.Y(n_2375)
);

CKINVDCx5p33_ASAP7_75t_R g2376 ( 
.A(n_2096),
.Y(n_2376)
);

CKINVDCx5p33_ASAP7_75t_R g2377 ( 
.A(n_1949),
.Y(n_2377)
);

INVx1_ASAP7_75t_L g2378 ( 
.A(n_1930),
.Y(n_2378)
);

INVx1_ASAP7_75t_L g2379 ( 
.A(n_1930),
.Y(n_2379)
);

INVx2_ASAP7_75t_L g2380 ( 
.A(n_2015),
.Y(n_2380)
);

INVx3_ASAP7_75t_L g2381 ( 
.A(n_1941),
.Y(n_2381)
);

CKINVDCx20_ASAP7_75t_R g2382 ( 
.A(n_1949),
.Y(n_2382)
);

CKINVDCx5p33_ASAP7_75t_R g2383 ( 
.A(n_1949),
.Y(n_2383)
);

NAND2xp5_ASAP7_75t_L g2384 ( 
.A(n_1976),
.B(n_1610),
.Y(n_2384)
);

HB1xp67_ASAP7_75t_L g2385 ( 
.A(n_1921),
.Y(n_2385)
);

INVx2_ASAP7_75t_L g2386 ( 
.A(n_2015),
.Y(n_2386)
);

INVx1_ASAP7_75t_L g2387 ( 
.A(n_1930),
.Y(n_2387)
);

NAND2xp33_ASAP7_75t_R g2388 ( 
.A(n_1912),
.B(n_1628),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_1930),
.Y(n_2389)
);

CKINVDCx5p33_ASAP7_75t_R g2390 ( 
.A(n_1949),
.Y(n_2390)
);

INVx3_ASAP7_75t_L g2391 ( 
.A(n_1941),
.Y(n_2391)
);

INVx1_ASAP7_75t_L g2392 ( 
.A(n_1930),
.Y(n_2392)
);

INVx1_ASAP7_75t_L g2393 ( 
.A(n_1930),
.Y(n_2393)
);

CKINVDCx20_ASAP7_75t_R g2394 ( 
.A(n_1949),
.Y(n_2394)
);

INVx1_ASAP7_75t_L g2395 ( 
.A(n_1930),
.Y(n_2395)
);

INVx1_ASAP7_75t_L g2396 ( 
.A(n_1930),
.Y(n_2396)
);

INVx2_ASAP7_75t_L g2397 ( 
.A(n_2015),
.Y(n_2397)
);

CKINVDCx5p33_ASAP7_75t_R g2398 ( 
.A(n_1949),
.Y(n_2398)
);

HB1xp67_ASAP7_75t_L g2399 ( 
.A(n_1921),
.Y(n_2399)
);

INVx3_ASAP7_75t_L g2400 ( 
.A(n_1941),
.Y(n_2400)
);

NOR2xp33_ASAP7_75t_R g2401 ( 
.A(n_1922),
.B(n_1188),
.Y(n_2401)
);

INVx3_ASAP7_75t_L g2402 ( 
.A(n_1941),
.Y(n_2402)
);

INVx1_ASAP7_75t_L g2403 ( 
.A(n_1930),
.Y(n_2403)
);

BUFx3_ASAP7_75t_L g2404 ( 
.A(n_2075),
.Y(n_2404)
);

CKINVDCx5p33_ASAP7_75t_R g2405 ( 
.A(n_1949),
.Y(n_2405)
);

INVx1_ASAP7_75t_L g2406 ( 
.A(n_1930),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_1930),
.Y(n_2407)
);

CKINVDCx5p33_ASAP7_75t_R g2408 ( 
.A(n_1949),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_1930),
.Y(n_2409)
);

INVx1_ASAP7_75t_L g2410 ( 
.A(n_1930),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_2148),
.Y(n_2411)
);

INVx4_ASAP7_75t_L g2412 ( 
.A(n_2143),
.Y(n_2412)
);

BUFx6f_ASAP7_75t_L g2413 ( 
.A(n_2121),
.Y(n_2413)
);

AND2x4_ASAP7_75t_L g2414 ( 
.A(n_2223),
.B(n_1302),
.Y(n_2414)
);

INVx1_ASAP7_75t_L g2415 ( 
.A(n_2156),
.Y(n_2415)
);

NOR2xp33_ASAP7_75t_L g2416 ( 
.A(n_2236),
.B(n_1189),
.Y(n_2416)
);

INVxp67_ASAP7_75t_L g2417 ( 
.A(n_2149),
.Y(n_2417)
);

AND2x6_ASAP7_75t_L g2418 ( 
.A(n_2164),
.B(n_2168),
.Y(n_2418)
);

AND2x2_ASAP7_75t_L g2419 ( 
.A(n_2167),
.B(n_1195),
.Y(n_2419)
);

INVx2_ASAP7_75t_L g2420 ( 
.A(n_2334),
.Y(n_2420)
);

NAND2x1p5_ASAP7_75t_L g2421 ( 
.A(n_2126),
.B(n_1368),
.Y(n_2421)
);

INVx2_ASAP7_75t_SL g2422 ( 
.A(n_2370),
.Y(n_2422)
);

AND2x4_ASAP7_75t_L g2423 ( 
.A(n_2178),
.B(n_1119),
.Y(n_2423)
);

HB1xp67_ASAP7_75t_L g2424 ( 
.A(n_2166),
.Y(n_2424)
);

OR2x6_ASAP7_75t_L g2425 ( 
.A(n_2124),
.B(n_1637),
.Y(n_2425)
);

BUFx6f_ASAP7_75t_L g2426 ( 
.A(n_2404),
.Y(n_2426)
);

INVx3_ASAP7_75t_L g2427 ( 
.A(n_2246),
.Y(n_2427)
);

CKINVDCx5p33_ASAP7_75t_R g2428 ( 
.A(n_2131),
.Y(n_2428)
);

NAND2xp5_ASAP7_75t_SL g2429 ( 
.A(n_2269),
.B(n_1633),
.Y(n_2429)
);

AND2x2_ASAP7_75t_L g2430 ( 
.A(n_2385),
.B(n_1236),
.Y(n_2430)
);

INVx5_ASAP7_75t_L g2431 ( 
.A(n_2179),
.Y(n_2431)
);

INVx1_ASAP7_75t_L g2432 ( 
.A(n_2276),
.Y(n_2432)
);

AND2x6_ASAP7_75t_L g2433 ( 
.A(n_2169),
.B(n_1684),
.Y(n_2433)
);

AND2x2_ASAP7_75t_L g2434 ( 
.A(n_2399),
.B(n_1251),
.Y(n_2434)
);

NOR2xp33_ASAP7_75t_L g2435 ( 
.A(n_2241),
.B(n_1253),
.Y(n_2435)
);

NAND2xp5_ASAP7_75t_SL g2436 ( 
.A(n_2273),
.B(n_1634),
.Y(n_2436)
);

INVx1_ASAP7_75t_L g2437 ( 
.A(n_2302),
.Y(n_2437)
);

INVx2_ASAP7_75t_L g2438 ( 
.A(n_2381),
.Y(n_2438)
);

INVx1_ASAP7_75t_L g2439 ( 
.A(n_2174),
.Y(n_2439)
);

INVx1_ASAP7_75t_L g2440 ( 
.A(n_2183),
.Y(n_2440)
);

INVx2_ASAP7_75t_L g2441 ( 
.A(n_2381),
.Y(n_2441)
);

INVx1_ASAP7_75t_L g2442 ( 
.A(n_2186),
.Y(n_2442)
);

NOR2xp33_ASAP7_75t_L g2443 ( 
.A(n_2182),
.B(n_2274),
.Y(n_2443)
);

INVx4_ASAP7_75t_SL g2444 ( 
.A(n_2335),
.Y(n_2444)
);

AND2x2_ASAP7_75t_L g2445 ( 
.A(n_2196),
.B(n_1331),
.Y(n_2445)
);

BUFx10_ASAP7_75t_L g2446 ( 
.A(n_2113),
.Y(n_2446)
);

INVx1_ASAP7_75t_L g2447 ( 
.A(n_2188),
.Y(n_2447)
);

INVx1_ASAP7_75t_L g2448 ( 
.A(n_2191),
.Y(n_2448)
);

NAND2xp5_ASAP7_75t_L g2449 ( 
.A(n_2217),
.B(n_1642),
.Y(n_2449)
);

INVx4_ASAP7_75t_SL g2450 ( 
.A(n_2335),
.Y(n_2450)
);

NOR2xp33_ASAP7_75t_L g2451 ( 
.A(n_2212),
.B(n_1692),
.Y(n_2451)
);

NOR2xp33_ASAP7_75t_L g2452 ( 
.A(n_2220),
.B(n_2221),
.Y(n_2452)
);

NAND2xp5_ASAP7_75t_L g2453 ( 
.A(n_2306),
.B(n_1644),
.Y(n_2453)
);

INVxp33_ASAP7_75t_L g2454 ( 
.A(n_2107),
.Y(n_2454)
);

INVx4_ASAP7_75t_L g2455 ( 
.A(n_2116),
.Y(n_2455)
);

INVx1_ASAP7_75t_L g2456 ( 
.A(n_2193),
.Y(n_2456)
);

INVxp33_ASAP7_75t_L g2457 ( 
.A(n_2341),
.Y(n_2457)
);

INVx1_ASAP7_75t_L g2458 ( 
.A(n_2195),
.Y(n_2458)
);

BUFx6f_ASAP7_75t_L g2459 ( 
.A(n_2205),
.Y(n_2459)
);

INVx2_ASAP7_75t_L g2460 ( 
.A(n_2391),
.Y(n_2460)
);

AND2x4_ASAP7_75t_L g2461 ( 
.A(n_2178),
.B(n_1135),
.Y(n_2461)
);

OR2x2_ASAP7_75t_L g2462 ( 
.A(n_2213),
.B(n_1394),
.Y(n_2462)
);

BUFx3_ASAP7_75t_L g2463 ( 
.A(n_2365),
.Y(n_2463)
);

INVx1_ASAP7_75t_L g2464 ( 
.A(n_2200),
.Y(n_2464)
);

BUFx6f_ASAP7_75t_L g2465 ( 
.A(n_2205),
.Y(n_2465)
);

AOI22xp33_ASAP7_75t_L g2466 ( 
.A1(n_2247),
.A2(n_1654),
.B1(n_1662),
.B2(n_1651),
.Y(n_2466)
);

BUFx3_ASAP7_75t_L g2467 ( 
.A(n_2366),
.Y(n_2467)
);

INVx2_ASAP7_75t_SL g2468 ( 
.A(n_2246),
.Y(n_2468)
);

INVx1_ASAP7_75t_L g2469 ( 
.A(n_2216),
.Y(n_2469)
);

INVx1_ASAP7_75t_L g2470 ( 
.A(n_2230),
.Y(n_2470)
);

INVx2_ASAP7_75t_L g2471 ( 
.A(n_2391),
.Y(n_2471)
);

AOI22xp33_ASAP7_75t_L g2472 ( 
.A1(n_2266),
.A2(n_1673),
.B1(n_1678),
.B2(n_1672),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_2233),
.Y(n_2473)
);

NOR2xp33_ASAP7_75t_L g2474 ( 
.A(n_2222),
.B(n_1732),
.Y(n_2474)
);

INVx2_ASAP7_75t_L g2475 ( 
.A(n_2400),
.Y(n_2475)
);

INVx1_ASAP7_75t_L g2476 ( 
.A(n_2238),
.Y(n_2476)
);

INVx1_ASAP7_75t_L g2477 ( 
.A(n_2242),
.Y(n_2477)
);

INVxp33_ASAP7_75t_L g2478 ( 
.A(n_2345),
.Y(n_2478)
);

NOR2xp33_ASAP7_75t_L g2479 ( 
.A(n_2229),
.B(n_1742),
.Y(n_2479)
);

AND2x2_ASAP7_75t_L g2480 ( 
.A(n_2214),
.B(n_1751),
.Y(n_2480)
);

INVx5_ASAP7_75t_L g2481 ( 
.A(n_2179),
.Y(n_2481)
);

INVx1_ASAP7_75t_L g2482 ( 
.A(n_2249),
.Y(n_2482)
);

INVx1_ASAP7_75t_L g2483 ( 
.A(n_2253),
.Y(n_2483)
);

INVx1_ASAP7_75t_L g2484 ( 
.A(n_2256),
.Y(n_2484)
);

AND2x2_ASAP7_75t_L g2485 ( 
.A(n_2218),
.B(n_1210),
.Y(n_2485)
);

HB1xp67_ASAP7_75t_L g2486 ( 
.A(n_2155),
.Y(n_2486)
);

INVx1_ASAP7_75t_L g2487 ( 
.A(n_2257),
.Y(n_2487)
);

XOR2xp5_ASAP7_75t_L g2488 ( 
.A(n_2130),
.B(n_1681),
.Y(n_2488)
);

INVx4_ASAP7_75t_L g2489 ( 
.A(n_2117),
.Y(n_2489)
);

INVx1_ASAP7_75t_SL g2490 ( 
.A(n_2127),
.Y(n_2490)
);

NAND2xp5_ASAP7_75t_L g2491 ( 
.A(n_2145),
.B(n_1682),
.Y(n_2491)
);

INVx4_ASAP7_75t_L g2492 ( 
.A(n_2118),
.Y(n_2492)
);

INVx1_ASAP7_75t_L g2493 ( 
.A(n_2258),
.Y(n_2493)
);

CKINVDCx5p33_ASAP7_75t_R g2494 ( 
.A(n_2106),
.Y(n_2494)
);

CKINVDCx5p33_ASAP7_75t_R g2495 ( 
.A(n_2105),
.Y(n_2495)
);

INVx1_ASAP7_75t_L g2496 ( 
.A(n_2270),
.Y(n_2496)
);

INVx3_ASAP7_75t_L g2497 ( 
.A(n_2122),
.Y(n_2497)
);

INVx1_ASAP7_75t_L g2498 ( 
.A(n_2309),
.Y(n_2498)
);

NAND2xp5_ASAP7_75t_L g2499 ( 
.A(n_2109),
.B(n_1685),
.Y(n_2499)
);

INVx1_ASAP7_75t_L g2500 ( 
.A(n_2310),
.Y(n_2500)
);

INVx4_ASAP7_75t_SL g2501 ( 
.A(n_2226),
.Y(n_2501)
);

BUFx3_ASAP7_75t_L g2502 ( 
.A(n_2329),
.Y(n_2502)
);

INVx1_ASAP7_75t_L g2503 ( 
.A(n_2162),
.Y(n_2503)
);

INVx1_ASAP7_75t_L g2504 ( 
.A(n_2320),
.Y(n_2504)
);

INVxp67_ASAP7_75t_SL g2505 ( 
.A(n_2286),
.Y(n_2505)
);

INVx1_ASAP7_75t_L g2506 ( 
.A(n_2119),
.Y(n_2506)
);

XNOR2xp5_ASAP7_75t_L g2507 ( 
.A(n_2124),
.B(n_1697),
.Y(n_2507)
);

INVx2_ASAP7_75t_L g2508 ( 
.A(n_2400),
.Y(n_2508)
);

INVx1_ASAP7_75t_L g2509 ( 
.A(n_2120),
.Y(n_2509)
);

BUFx2_ASAP7_75t_L g2510 ( 
.A(n_2185),
.Y(n_2510)
);

AND2x4_ASAP7_75t_L g2511 ( 
.A(n_2240),
.B(n_1143),
.Y(n_2511)
);

INVx2_ASAP7_75t_SL g2512 ( 
.A(n_2284),
.Y(n_2512)
);

INVx4_ASAP7_75t_L g2513 ( 
.A(n_2123),
.Y(n_2513)
);

NAND2xp5_ASAP7_75t_SL g2514 ( 
.A(n_2307),
.B(n_1698),
.Y(n_2514)
);

INVx2_ASAP7_75t_L g2515 ( 
.A(n_2402),
.Y(n_2515)
);

BUFx2_ASAP7_75t_L g2516 ( 
.A(n_2198),
.Y(n_2516)
);

BUFx6f_ASAP7_75t_L g2517 ( 
.A(n_2205),
.Y(n_2517)
);

INVx1_ASAP7_75t_L g2518 ( 
.A(n_2136),
.Y(n_2518)
);

INVx5_ASAP7_75t_L g2519 ( 
.A(n_2179),
.Y(n_2519)
);

CKINVDCx11_ASAP7_75t_R g2520 ( 
.A(n_2382),
.Y(n_2520)
);

INVx2_ASAP7_75t_L g2521 ( 
.A(n_2402),
.Y(n_2521)
);

AO22x2_ASAP7_75t_L g2522 ( 
.A1(n_2204),
.A2(n_1477),
.B1(n_1502),
.B2(n_1447),
.Y(n_2522)
);

INVx1_ASAP7_75t_L g2523 ( 
.A(n_2378),
.Y(n_2523)
);

INVx1_ASAP7_75t_SL g2524 ( 
.A(n_2128),
.Y(n_2524)
);

AOI22xp33_ASAP7_75t_L g2525 ( 
.A1(n_2277),
.A2(n_1719),
.B1(n_1725),
.B2(n_1701),
.Y(n_2525)
);

BUFx6f_ASAP7_75t_L g2526 ( 
.A(n_2237),
.Y(n_2526)
);

BUFx3_ASAP7_75t_L g2527 ( 
.A(n_2394),
.Y(n_2527)
);

INVx2_ASAP7_75t_SL g2528 ( 
.A(n_2142),
.Y(n_2528)
);

INVx1_ASAP7_75t_SL g2529 ( 
.A(n_2208),
.Y(n_2529)
);

NAND2xp5_ASAP7_75t_SL g2530 ( 
.A(n_2308),
.B(n_1726),
.Y(n_2530)
);

INVx1_ASAP7_75t_L g2531 ( 
.A(n_2379),
.Y(n_2531)
);

AND2x2_ASAP7_75t_L g2532 ( 
.A(n_2250),
.B(n_1210),
.Y(n_2532)
);

BUFx2_ASAP7_75t_L g2533 ( 
.A(n_2227),
.Y(n_2533)
);

AOI22xp33_ASAP7_75t_L g2534 ( 
.A1(n_2260),
.A2(n_1735),
.B1(n_1744),
.B2(n_1730),
.Y(n_2534)
);

INVx3_ASAP7_75t_L g2535 ( 
.A(n_2125),
.Y(n_2535)
);

INVx1_ASAP7_75t_L g2536 ( 
.A(n_2387),
.Y(n_2536)
);

BUFx6f_ASAP7_75t_L g2537 ( 
.A(n_2237),
.Y(n_2537)
);

INVx2_ASAP7_75t_L g2538 ( 
.A(n_2139),
.Y(n_2538)
);

INVx3_ASAP7_75t_L g2539 ( 
.A(n_2301),
.Y(n_2539)
);

INVx1_ASAP7_75t_L g2540 ( 
.A(n_2389),
.Y(n_2540)
);

AND2x2_ASAP7_75t_L g2541 ( 
.A(n_2231),
.B(n_1212),
.Y(n_2541)
);

NAND2xp5_ASAP7_75t_L g2542 ( 
.A(n_2199),
.B(n_1748),
.Y(n_2542)
);

NAND2xp5_ASAP7_75t_SL g2543 ( 
.A(n_2311),
.B(n_1172),
.Y(n_2543)
);

INVx2_ASAP7_75t_L g2544 ( 
.A(n_2150),
.Y(n_2544)
);

INVx1_ASAP7_75t_L g2545 ( 
.A(n_2392),
.Y(n_2545)
);

INVx1_ASAP7_75t_L g2546 ( 
.A(n_2393),
.Y(n_2546)
);

INVx2_ASAP7_75t_L g2547 ( 
.A(n_2181),
.Y(n_2547)
);

NAND2xp5_ASAP7_75t_L g2548 ( 
.A(n_2384),
.B(n_1121),
.Y(n_2548)
);

NOR2xp33_ASAP7_75t_L g2549 ( 
.A(n_2232),
.B(n_1123),
.Y(n_2549)
);

OAI22xp33_ASAP7_75t_L g2550 ( 
.A1(n_2210),
.A2(n_1133),
.B1(n_1134),
.B2(n_1126),
.Y(n_2550)
);

AND2x2_ASAP7_75t_L g2551 ( 
.A(n_2297),
.B(n_1212),
.Y(n_2551)
);

INVx4_ASAP7_75t_L g2552 ( 
.A(n_2151),
.Y(n_2552)
);

INVx1_ASAP7_75t_L g2553 ( 
.A(n_2395),
.Y(n_2553)
);

OR2x2_ASAP7_75t_L g2554 ( 
.A(n_2180),
.B(n_1517),
.Y(n_2554)
);

INVx1_ASAP7_75t_L g2555 ( 
.A(n_2396),
.Y(n_2555)
);

OR2x2_ASAP7_75t_L g2556 ( 
.A(n_2147),
.B(n_1563),
.Y(n_2556)
);

BUFx6f_ASAP7_75t_L g2557 ( 
.A(n_2237),
.Y(n_2557)
);

AND2x2_ASAP7_75t_L g2558 ( 
.A(n_2299),
.B(n_1212),
.Y(n_2558)
);

INVx1_ASAP7_75t_L g2559 ( 
.A(n_2403),
.Y(n_2559)
);

AOI22xp33_ASAP7_75t_L g2560 ( 
.A1(n_2261),
.A2(n_1237),
.B1(n_1429),
.B2(n_1327),
.Y(n_2560)
);

INVx1_ASAP7_75t_L g2561 ( 
.A(n_2406),
.Y(n_2561)
);

CKINVDCx6p67_ASAP7_75t_R g2562 ( 
.A(n_2296),
.Y(n_2562)
);

CKINVDCx5p33_ASAP7_75t_R g2563 ( 
.A(n_2377),
.Y(n_2563)
);

INVx2_ASAP7_75t_L g2564 ( 
.A(n_2203),
.Y(n_2564)
);

NAND2xp33_ASAP7_75t_L g2565 ( 
.A(n_2283),
.B(n_1471),
.Y(n_2565)
);

INVx1_ASAP7_75t_L g2566 ( 
.A(n_2407),
.Y(n_2566)
);

INVx2_ASAP7_75t_L g2567 ( 
.A(n_2301),
.Y(n_2567)
);

NAND2xp5_ASAP7_75t_SL g2568 ( 
.A(n_2313),
.B(n_1274),
.Y(n_2568)
);

BUFx6f_ASAP7_75t_SL g2569 ( 
.A(n_2112),
.Y(n_2569)
);

NAND2xp5_ASAP7_75t_SL g2570 ( 
.A(n_2314),
.B(n_2303),
.Y(n_2570)
);

NAND2xp5_ASAP7_75t_SL g2571 ( 
.A(n_2305),
.B(n_1287),
.Y(n_2571)
);

BUFx6f_ASAP7_75t_L g2572 ( 
.A(n_2295),
.Y(n_2572)
);

NOR2xp33_ASAP7_75t_L g2573 ( 
.A(n_2278),
.B(n_1136),
.Y(n_2573)
);

NOR2xp33_ASAP7_75t_L g2574 ( 
.A(n_2265),
.B(n_1137),
.Y(n_2574)
);

AOI22xp33_ASAP7_75t_L g2575 ( 
.A1(n_2263),
.A2(n_2268),
.B1(n_2272),
.B2(n_2271),
.Y(n_2575)
);

BUFx2_ASAP7_75t_L g2576 ( 
.A(n_2158),
.Y(n_2576)
);

BUFx6f_ASAP7_75t_L g2577 ( 
.A(n_2295),
.Y(n_2577)
);

INVx3_ASAP7_75t_L g2578 ( 
.A(n_2159),
.Y(n_2578)
);

INVx3_ASAP7_75t_L g2579 ( 
.A(n_2161),
.Y(n_2579)
);

OR2x6_ASAP7_75t_L g2580 ( 
.A(n_2209),
.B(n_1273),
.Y(n_2580)
);

BUFx3_ASAP7_75t_L g2581 ( 
.A(n_2152),
.Y(n_2581)
);

INVx1_ASAP7_75t_L g2582 ( 
.A(n_2409),
.Y(n_2582)
);

INVx3_ASAP7_75t_L g2583 ( 
.A(n_2163),
.Y(n_2583)
);

NAND2xp5_ASAP7_75t_L g2584 ( 
.A(n_2298),
.B(n_1138),
.Y(n_2584)
);

INVx1_ASAP7_75t_L g2585 ( 
.A(n_2410),
.Y(n_2585)
);

INVx2_ASAP7_75t_L g2586 ( 
.A(n_2295),
.Y(n_2586)
);

INVx1_ASAP7_75t_L g2587 ( 
.A(n_2321),
.Y(n_2587)
);

OAI21xp33_ASAP7_75t_SL g2588 ( 
.A1(n_2312),
.A2(n_1378),
.B(n_1322),
.Y(n_2588)
);

INVx1_ASAP7_75t_L g2589 ( 
.A(n_2300),
.Y(n_2589)
);

INVx1_ASAP7_75t_L g2590 ( 
.A(n_2304),
.Y(n_2590)
);

NAND2xp5_ASAP7_75t_L g2591 ( 
.A(n_2259),
.B(n_1141),
.Y(n_2591)
);

HB1xp67_ASAP7_75t_L g2592 ( 
.A(n_2317),
.Y(n_2592)
);

NAND2xp5_ASAP7_75t_L g2593 ( 
.A(n_2264),
.B(n_1145),
.Y(n_2593)
);

INVx2_ASAP7_75t_L g2594 ( 
.A(n_2110),
.Y(n_2594)
);

BUFx4f_ASAP7_75t_L g2595 ( 
.A(n_2290),
.Y(n_2595)
);

INVx3_ASAP7_75t_L g2596 ( 
.A(n_2165),
.Y(n_2596)
);

INVx3_ASAP7_75t_L g2597 ( 
.A(n_2146),
.Y(n_2597)
);

AOI22xp33_ASAP7_75t_L g2598 ( 
.A1(n_2280),
.A2(n_1237),
.B1(n_1429),
.B2(n_1327),
.Y(n_2598)
);

BUFx6f_ASAP7_75t_L g2599 ( 
.A(n_2348),
.Y(n_2599)
);

INVx3_ASAP7_75t_L g2600 ( 
.A(n_2132),
.Y(n_2600)
);

INVx1_ASAP7_75t_L g2601 ( 
.A(n_2326),
.Y(n_2601)
);

OAI22xp5_ASAP7_75t_L g2602 ( 
.A1(n_2281),
.A2(n_1571),
.B1(n_1151),
.B2(n_1153),
.Y(n_2602)
);

NOR2xp33_ASAP7_75t_L g2603 ( 
.A(n_2239),
.B(n_1146),
.Y(n_2603)
);

INVx3_ASAP7_75t_L g2604 ( 
.A(n_2133),
.Y(n_2604)
);

BUFx3_ASAP7_75t_L g2605 ( 
.A(n_2134),
.Y(n_2605)
);

NAND2xp5_ASAP7_75t_L g2606 ( 
.A(n_2157),
.B(n_2187),
.Y(n_2606)
);

INVxp33_ASAP7_75t_L g2607 ( 
.A(n_2160),
.Y(n_2607)
);

INVx1_ASAP7_75t_L g2608 ( 
.A(n_2140),
.Y(n_2608)
);

INVx2_ASAP7_75t_L g2609 ( 
.A(n_2111),
.Y(n_2609)
);

AND2x4_ASAP7_75t_L g2610 ( 
.A(n_2138),
.B(n_1149),
.Y(n_2610)
);

INVx2_ASAP7_75t_L g2611 ( 
.A(n_2129),
.Y(n_2611)
);

INVx2_ASAP7_75t_L g2612 ( 
.A(n_2380),
.Y(n_2612)
);

AOI22xp33_ASAP7_75t_L g2613 ( 
.A1(n_2282),
.A2(n_1237),
.B1(n_1429),
.B2(n_1327),
.Y(n_2613)
);

NAND2xp5_ASAP7_75t_L g2614 ( 
.A(n_2315),
.B(n_1155),
.Y(n_2614)
);

AND2x2_ASAP7_75t_SL g2615 ( 
.A(n_2170),
.B(n_1273),
.Y(n_2615)
);

INVx2_ASAP7_75t_L g2616 ( 
.A(n_2386),
.Y(n_2616)
);

INVx2_ASAP7_75t_L g2617 ( 
.A(n_2397),
.Y(n_2617)
);

NAND2xp5_ASAP7_75t_SL g2618 ( 
.A(n_2287),
.B(n_1156),
.Y(n_2618)
);

AND2x2_ASAP7_75t_L g2619 ( 
.A(n_2225),
.B(n_1472),
.Y(n_2619)
);

INVx1_ASAP7_75t_SL g2620 ( 
.A(n_2401),
.Y(n_2620)
);

NOR2xp33_ASAP7_75t_L g2621 ( 
.A(n_2243),
.B(n_1158),
.Y(n_2621)
);

INVx2_ASAP7_75t_L g2622 ( 
.A(n_2327),
.Y(n_2622)
);

AOI22xp33_ASAP7_75t_L g2623 ( 
.A1(n_2234),
.A2(n_1474),
.B1(n_1485),
.B2(n_1472),
.Y(n_2623)
);

INVx1_ASAP7_75t_L g2624 ( 
.A(n_2332),
.Y(n_2624)
);

INVx2_ASAP7_75t_L g2625 ( 
.A(n_2338),
.Y(n_2625)
);

INVx1_ASAP7_75t_SL g2626 ( 
.A(n_2316),
.Y(n_2626)
);

AND2x2_ASAP7_75t_L g2627 ( 
.A(n_2189),
.B(n_1472),
.Y(n_2627)
);

INVx2_ASAP7_75t_L g2628 ( 
.A(n_2344),
.Y(n_2628)
);

BUFx6f_ASAP7_75t_L g2629 ( 
.A(n_2351),
.Y(n_2629)
);

NAND2xp5_ASAP7_75t_SL g2630 ( 
.A(n_2202),
.B(n_1159),
.Y(n_2630)
);

AND2x4_ASAP7_75t_L g2631 ( 
.A(n_2235),
.B(n_1154),
.Y(n_2631)
);

NOR2xp33_ASAP7_75t_L g2632 ( 
.A(n_2244),
.B(n_1165),
.Y(n_2632)
);

NAND2xp5_ASAP7_75t_SL g2633 ( 
.A(n_2322),
.B(n_1166),
.Y(n_2633)
);

AND2x6_ASAP7_75t_L g2634 ( 
.A(n_2344),
.B(n_1157),
.Y(n_2634)
);

NAND2xp5_ASAP7_75t_L g2635 ( 
.A(n_2323),
.B(n_1168),
.Y(n_2635)
);

NAND2xp5_ASAP7_75t_L g2636 ( 
.A(n_2324),
.B(n_1171),
.Y(n_2636)
);

NAND2xp5_ASAP7_75t_L g2637 ( 
.A(n_2325),
.B(n_1173),
.Y(n_2637)
);

NOR2xp33_ASAP7_75t_L g2638 ( 
.A(n_2248),
.B(n_1180),
.Y(n_2638)
);

INVx4_ASAP7_75t_L g2639 ( 
.A(n_2135),
.Y(n_2639)
);

BUFx3_ASAP7_75t_L g2640 ( 
.A(n_2171),
.Y(n_2640)
);

INVx1_ASAP7_75t_L g2641 ( 
.A(n_2355),
.Y(n_2641)
);

HB1xp67_ASAP7_75t_L g2642 ( 
.A(n_2352),
.Y(n_2642)
);

OR2x6_ASAP7_75t_L g2643 ( 
.A(n_2173),
.B(n_1296),
.Y(n_2643)
);

INVx3_ASAP7_75t_L g2644 ( 
.A(n_2115),
.Y(n_2644)
);

INVx1_ASAP7_75t_L g2645 ( 
.A(n_2328),
.Y(n_2645)
);

BUFx3_ASAP7_75t_L g2646 ( 
.A(n_2172),
.Y(n_2646)
);

INVx2_ASAP7_75t_L g2647 ( 
.A(n_2228),
.Y(n_2647)
);

BUFx10_ASAP7_75t_L g2648 ( 
.A(n_2383),
.Y(n_2648)
);

NAND2xp5_ASAP7_75t_L g2649 ( 
.A(n_2330),
.B(n_1182),
.Y(n_2649)
);

INVx1_ASAP7_75t_L g2650 ( 
.A(n_2331),
.Y(n_2650)
);

OR2x6_ASAP7_75t_L g2651 ( 
.A(n_2177),
.B(n_1296),
.Y(n_2651)
);

INVx1_ASAP7_75t_L g2652 ( 
.A(n_2333),
.Y(n_2652)
);

NAND2xp5_ASAP7_75t_L g2653 ( 
.A(n_2336),
.B(n_2340),
.Y(n_2653)
);

INVx1_ASAP7_75t_L g2654 ( 
.A(n_2342),
.Y(n_2654)
);

INVx1_ASAP7_75t_L g2655 ( 
.A(n_2343),
.Y(n_2655)
);

BUFx3_ASAP7_75t_L g2656 ( 
.A(n_2390),
.Y(n_2656)
);

AND2x4_ASAP7_75t_L g2657 ( 
.A(n_2346),
.B(n_1160),
.Y(n_2657)
);

INVx1_ASAP7_75t_L g2658 ( 
.A(n_2285),
.Y(n_2658)
);

INVx3_ASAP7_75t_L g2659 ( 
.A(n_2114),
.Y(n_2659)
);

NOR2xp33_ASAP7_75t_L g2660 ( 
.A(n_2251),
.B(n_2252),
.Y(n_2660)
);

NAND2xp5_ASAP7_75t_L g2661 ( 
.A(n_2154),
.B(n_1183),
.Y(n_2661)
);

INVx2_ASAP7_75t_L g2662 ( 
.A(n_2245),
.Y(n_2662)
);

AND2x2_ASAP7_75t_L g2663 ( 
.A(n_2190),
.B(n_2154),
.Y(n_2663)
);

INVx4_ASAP7_75t_SL g2664 ( 
.A(n_2361),
.Y(n_2664)
);

NOR2xp33_ASAP7_75t_L g2665 ( 
.A(n_2289),
.B(n_2292),
.Y(n_2665)
);

AND2x6_ASAP7_75t_L g2666 ( 
.A(n_2288),
.B(n_1157),
.Y(n_2666)
);

BUFx3_ASAP7_75t_L g2667 ( 
.A(n_2398),
.Y(n_2667)
);

AND2x6_ASAP7_75t_L g2668 ( 
.A(n_2275),
.B(n_1169),
.Y(n_2668)
);

INVx4_ASAP7_75t_L g2669 ( 
.A(n_2108),
.Y(n_2669)
);

NAND2x1p5_ASAP7_75t_L g2670 ( 
.A(n_2347),
.B(n_1573),
.Y(n_2670)
);

INVx4_ASAP7_75t_L g2671 ( 
.A(n_2405),
.Y(n_2671)
);

INVx1_ASAP7_75t_L g2672 ( 
.A(n_2375),
.Y(n_2672)
);

INVxp67_ASAP7_75t_SL g2673 ( 
.A(n_2388),
.Y(n_2673)
);

BUFx10_ASAP7_75t_L g2674 ( 
.A(n_2408),
.Y(n_2674)
);

NAND2xp5_ASAP7_75t_SL g2675 ( 
.A(n_2262),
.B(n_1185),
.Y(n_2675)
);

INVxp67_ASAP7_75t_L g2676 ( 
.A(n_2184),
.Y(n_2676)
);

NAND3x1_ASAP7_75t_L g2677 ( 
.A(n_2144),
.B(n_1181),
.C(n_1177),
.Y(n_2677)
);

INVx2_ASAP7_75t_L g2678 ( 
.A(n_2279),
.Y(n_2678)
);

NAND2xp5_ASAP7_75t_L g2679 ( 
.A(n_2175),
.B(n_1191),
.Y(n_2679)
);

INVx1_ASAP7_75t_L g2680 ( 
.A(n_2291),
.Y(n_2680)
);

AND2x2_ASAP7_75t_L g2681 ( 
.A(n_2176),
.B(n_2197),
.Y(n_2681)
);

NAND2xp5_ASAP7_75t_SL g2682 ( 
.A(n_2319),
.B(n_1192),
.Y(n_2682)
);

HB1xp67_ASAP7_75t_L g2683 ( 
.A(n_2215),
.Y(n_2683)
);

INVx2_ASAP7_75t_L g2684 ( 
.A(n_2293),
.Y(n_2684)
);

INVx1_ASAP7_75t_SL g2685 ( 
.A(n_2153),
.Y(n_2685)
);

INVx1_ASAP7_75t_L g2686 ( 
.A(n_2357),
.Y(n_2686)
);

BUFx6f_ASAP7_75t_L g2687 ( 
.A(n_2353),
.Y(n_2687)
);

INVx1_ASAP7_75t_SL g2688 ( 
.A(n_2141),
.Y(n_2688)
);

NAND2xp5_ASAP7_75t_L g2689 ( 
.A(n_2206),
.B(n_1194),
.Y(n_2689)
);

INVx1_ASAP7_75t_L g2690 ( 
.A(n_2318),
.Y(n_2690)
);

BUFx2_ASAP7_75t_L g2691 ( 
.A(n_2294),
.Y(n_2691)
);

NAND2xp5_ASAP7_75t_SL g2692 ( 
.A(n_2219),
.B(n_1197),
.Y(n_2692)
);

BUFx6f_ASAP7_75t_L g2693 ( 
.A(n_2359),
.Y(n_2693)
);

AND2x2_ASAP7_75t_SL g2694 ( 
.A(n_2201),
.B(n_1307),
.Y(n_2694)
);

NOR2xp33_ASAP7_75t_L g2695 ( 
.A(n_2194),
.B(n_1200),
.Y(n_2695)
);

INVx1_ASAP7_75t_L g2696 ( 
.A(n_2376),
.Y(n_2696)
);

CKINVDCx5p33_ASAP7_75t_R g2697 ( 
.A(n_2224),
.Y(n_2697)
);

AND2x4_ASAP7_75t_L g2698 ( 
.A(n_2267),
.B(n_1193),
.Y(n_2698)
);

INVx1_ASAP7_75t_L g2699 ( 
.A(n_2362),
.Y(n_2699)
);

AND2x4_ASAP7_75t_L g2700 ( 
.A(n_2254),
.B(n_1199),
.Y(n_2700)
);

INVx2_ASAP7_75t_L g2701 ( 
.A(n_2372),
.Y(n_2701)
);

INVxp67_ASAP7_75t_L g2702 ( 
.A(n_2255),
.Y(n_2702)
);

INVx1_ASAP7_75t_L g2703 ( 
.A(n_2364),
.Y(n_2703)
);

INVx1_ASAP7_75t_L g2704 ( 
.A(n_2367),
.Y(n_2704)
);

CKINVDCx20_ASAP7_75t_R g2705 ( 
.A(n_2207),
.Y(n_2705)
);

INVx1_ASAP7_75t_L g2706 ( 
.A(n_2368),
.Y(n_2706)
);

AND2x6_ASAP7_75t_L g2707 ( 
.A(n_2337),
.B(n_1169),
.Y(n_2707)
);

NAND2xp5_ASAP7_75t_L g2708 ( 
.A(n_2192),
.B(n_1201),
.Y(n_2708)
);

INVx2_ASAP7_75t_L g2709 ( 
.A(n_2337),
.Y(n_2709)
);

NAND2xp5_ASAP7_75t_L g2710 ( 
.A(n_2369),
.B(n_1204),
.Y(n_2710)
);

INVx4_ASAP7_75t_SL g2711 ( 
.A(n_2211),
.Y(n_2711)
);

INVx6_ASAP7_75t_L g2712 ( 
.A(n_2337),
.Y(n_2712)
);

CKINVDCx5p33_ASAP7_75t_R g2713 ( 
.A(n_2137),
.Y(n_2713)
);

INVx1_ASAP7_75t_L g2714 ( 
.A(n_2371),
.Y(n_2714)
);

NAND2xp5_ASAP7_75t_L g2715 ( 
.A(n_2339),
.B(n_1206),
.Y(n_2715)
);

INVx1_ASAP7_75t_L g2716 ( 
.A(n_2349),
.Y(n_2716)
);

BUFx4f_ASAP7_75t_L g2717 ( 
.A(n_2354),
.Y(n_2717)
);

BUFx10_ASAP7_75t_L g2718 ( 
.A(n_2356),
.Y(n_2718)
);

NOR2xp33_ASAP7_75t_L g2719 ( 
.A(n_2373),
.B(n_1207),
.Y(n_2719)
);

INVx2_ASAP7_75t_L g2720 ( 
.A(n_2339),
.Y(n_2720)
);

NAND2xp5_ASAP7_75t_SL g2721 ( 
.A(n_2339),
.B(n_1209),
.Y(n_2721)
);

BUFx3_ASAP7_75t_L g2722 ( 
.A(n_2374),
.Y(n_2722)
);

INVx1_ASAP7_75t_L g2723 ( 
.A(n_2350),
.Y(n_2723)
);

INVx1_ASAP7_75t_L g2724 ( 
.A(n_2358),
.Y(n_2724)
);

AO21x1_ASAP7_75t_L g2725 ( 
.A1(n_2360),
.A2(n_1213),
.B(n_1202),
.Y(n_2725)
);

NAND2xp5_ASAP7_75t_L g2726 ( 
.A(n_2360),
.B(n_1211),
.Y(n_2726)
);

INVx2_ASAP7_75t_SL g2727 ( 
.A(n_2360),
.Y(n_2727)
);

OR2x2_ASAP7_75t_SL g2728 ( 
.A(n_2363),
.B(n_1214),
.Y(n_2728)
);

NAND2x1p5_ASAP7_75t_L g2729 ( 
.A(n_2363),
.B(n_1578),
.Y(n_2729)
);

NAND2xp5_ASAP7_75t_L g2730 ( 
.A(n_2363),
.B(n_1216),
.Y(n_2730)
);

INVx2_ASAP7_75t_L g2731 ( 
.A(n_2334),
.Y(n_2731)
);

NAND2xp33_ASAP7_75t_L g2732 ( 
.A(n_2269),
.B(n_1471),
.Y(n_2732)
);

AOI22xp5_ASAP7_75t_L g2733 ( 
.A1(n_2250),
.A2(n_1218),
.B1(n_1220),
.B2(n_1219),
.Y(n_2733)
);

INVx1_ASAP7_75t_L g2734 ( 
.A(n_2148),
.Y(n_2734)
);

AND2x2_ASAP7_75t_L g2735 ( 
.A(n_2167),
.B(n_1474),
.Y(n_2735)
);

NAND2xp5_ASAP7_75t_SL g2736 ( 
.A(n_2269),
.B(n_1221),
.Y(n_2736)
);

INVx3_ASAP7_75t_L g2737 ( 
.A(n_2121),
.Y(n_2737)
);

INVx1_ASAP7_75t_L g2738 ( 
.A(n_2148),
.Y(n_2738)
);

INVx4_ASAP7_75t_L g2739 ( 
.A(n_2143),
.Y(n_2739)
);

INVx1_ASAP7_75t_L g2740 ( 
.A(n_2148),
.Y(n_2740)
);

NAND2xp5_ASAP7_75t_SL g2741 ( 
.A(n_2269),
.B(n_1223),
.Y(n_2741)
);

INVx3_ASAP7_75t_L g2742 ( 
.A(n_2121),
.Y(n_2742)
);

NAND2xp5_ASAP7_75t_L g2743 ( 
.A(n_2217),
.B(n_1225),
.Y(n_2743)
);

INVx1_ASAP7_75t_L g2744 ( 
.A(n_2148),
.Y(n_2744)
);

INVx1_ASAP7_75t_L g2745 ( 
.A(n_2148),
.Y(n_2745)
);

AND2x2_ASAP7_75t_L g2746 ( 
.A(n_2167),
.B(n_1474),
.Y(n_2746)
);

INVx1_ASAP7_75t_L g2747 ( 
.A(n_2148),
.Y(n_2747)
);

NOR2x1_ASAP7_75t_L g2748 ( 
.A(n_2121),
.B(n_1215),
.Y(n_2748)
);

BUFx2_ASAP7_75t_L g2749 ( 
.A(n_2155),
.Y(n_2749)
);

INVx2_ASAP7_75t_L g2750 ( 
.A(n_2334),
.Y(n_2750)
);

INVx1_ASAP7_75t_L g2751 ( 
.A(n_2148),
.Y(n_2751)
);

OAI221xp5_ASAP7_75t_L g2752 ( 
.A1(n_2145),
.A2(n_1695),
.B1(n_1721),
.B2(n_1658),
.C(n_1631),
.Y(n_2752)
);

NAND2xp5_ASAP7_75t_L g2753 ( 
.A(n_2217),
.B(n_1226),
.Y(n_2753)
);

NOR2xp33_ASAP7_75t_L g2754 ( 
.A(n_2236),
.B(n_1228),
.Y(n_2754)
);

INVx2_ASAP7_75t_L g2755 ( 
.A(n_2334),
.Y(n_2755)
);

OR2x2_ASAP7_75t_L g2756 ( 
.A(n_2167),
.B(n_1729),
.Y(n_2756)
);

NAND2xp5_ASAP7_75t_L g2757 ( 
.A(n_2217),
.B(n_1229),
.Y(n_2757)
);

INVx3_ASAP7_75t_L g2758 ( 
.A(n_2121),
.Y(n_2758)
);

BUFx10_ASAP7_75t_L g2759 ( 
.A(n_2143),
.Y(n_2759)
);

BUFx3_ASAP7_75t_L g2760 ( 
.A(n_2365),
.Y(n_2760)
);

CKINVDCx5p33_ASAP7_75t_R g2761 ( 
.A(n_2131),
.Y(n_2761)
);

NOR2xp33_ASAP7_75t_SL g2762 ( 
.A(n_2167),
.B(n_1485),
.Y(n_2762)
);

INVx3_ASAP7_75t_L g2763 ( 
.A(n_2121),
.Y(n_2763)
);

CKINVDCx5p33_ASAP7_75t_R g2764 ( 
.A(n_2131),
.Y(n_2764)
);

BUFx6f_ASAP7_75t_L g2765 ( 
.A(n_2121),
.Y(n_2765)
);

INVx2_ASAP7_75t_L g2766 ( 
.A(n_2334),
.Y(n_2766)
);

NAND2xp5_ASAP7_75t_L g2767 ( 
.A(n_2217),
.B(n_1232),
.Y(n_2767)
);

AND2x2_ASAP7_75t_L g2768 ( 
.A(n_2167),
.B(n_1485),
.Y(n_2768)
);

NAND2xp5_ASAP7_75t_L g2769 ( 
.A(n_2217),
.B(n_1234),
.Y(n_2769)
);

NOR2xp33_ASAP7_75t_L g2770 ( 
.A(n_2236),
.B(n_1235),
.Y(n_2770)
);

NAND2xp5_ASAP7_75t_SL g2771 ( 
.A(n_2269),
.B(n_1240),
.Y(n_2771)
);

NOR2xp33_ASAP7_75t_L g2772 ( 
.A(n_2236),
.B(n_1241),
.Y(n_2772)
);

AOI22xp33_ASAP7_75t_L g2773 ( 
.A1(n_2212),
.A2(n_1597),
.B1(n_1646),
.B2(n_1569),
.Y(n_2773)
);

INVx2_ASAP7_75t_L g2774 ( 
.A(n_2334),
.Y(n_2774)
);

INVx1_ASAP7_75t_L g2775 ( 
.A(n_2148),
.Y(n_2775)
);

CKINVDCx8_ASAP7_75t_R g2776 ( 
.A(n_2112),
.Y(n_2776)
);

AND2x2_ASAP7_75t_L g2777 ( 
.A(n_2167),
.B(n_1569),
.Y(n_2777)
);

INVx1_ASAP7_75t_SL g2778 ( 
.A(n_2167),
.Y(n_2778)
);

NAND2xp5_ASAP7_75t_L g2779 ( 
.A(n_2217),
.B(n_1244),
.Y(n_2779)
);

BUFx6f_ASAP7_75t_L g2780 ( 
.A(n_2121),
.Y(n_2780)
);

BUFx3_ASAP7_75t_L g2781 ( 
.A(n_2365),
.Y(n_2781)
);

INVx5_ASAP7_75t_L g2782 ( 
.A(n_2179),
.Y(n_2782)
);

NAND2xp5_ASAP7_75t_L g2783 ( 
.A(n_2217),
.B(n_1245),
.Y(n_2783)
);

AND2x2_ASAP7_75t_SL g2784 ( 
.A(n_2166),
.B(n_1307),
.Y(n_2784)
);

AOI22xp5_ASAP7_75t_L g2785 ( 
.A1(n_2250),
.A2(n_1248),
.B1(n_1252),
.B2(n_1247),
.Y(n_2785)
);

NOR2xp33_ASAP7_75t_L g2786 ( 
.A(n_2236),
.B(n_1255),
.Y(n_2786)
);

NOR2xp33_ASAP7_75t_L g2787 ( 
.A(n_2236),
.B(n_1256),
.Y(n_2787)
);

AND2x6_ASAP7_75t_L g2788 ( 
.A(n_2164),
.B(n_1169),
.Y(n_2788)
);

AND2x4_ASAP7_75t_L g2789 ( 
.A(n_2223),
.B(n_1224),
.Y(n_2789)
);

INVx4_ASAP7_75t_SL g2790 ( 
.A(n_2121),
.Y(n_2790)
);

INVx2_ASAP7_75t_L g2791 ( 
.A(n_2334),
.Y(n_2791)
);

INVx2_ASAP7_75t_L g2792 ( 
.A(n_2334),
.Y(n_2792)
);

BUFx6f_ASAP7_75t_L g2793 ( 
.A(n_2121),
.Y(n_2793)
);

BUFx10_ASAP7_75t_L g2794 ( 
.A(n_2143),
.Y(n_2794)
);

AND2x6_ASAP7_75t_L g2795 ( 
.A(n_2164),
.B(n_1169),
.Y(n_2795)
);

INVx1_ASAP7_75t_L g2796 ( 
.A(n_2148),
.Y(n_2796)
);

NAND2xp5_ASAP7_75t_L g2797 ( 
.A(n_2217),
.B(n_1258),
.Y(n_2797)
);

BUFx3_ASAP7_75t_L g2798 ( 
.A(n_2365),
.Y(n_2798)
);

INVx3_ASAP7_75t_L g2799 ( 
.A(n_2121),
.Y(n_2799)
);

INVx2_ASAP7_75t_L g2800 ( 
.A(n_2538),
.Y(n_2800)
);

NAND2xp5_ASAP7_75t_L g2801 ( 
.A(n_2778),
.B(n_2411),
.Y(n_2801)
);

NAND2xp5_ASAP7_75t_L g2802 ( 
.A(n_2415),
.B(n_1261),
.Y(n_2802)
);

NAND2xp33_ASAP7_75t_L g2803 ( 
.A(n_2418),
.B(n_1262),
.Y(n_2803)
);

NAND2xp5_ASAP7_75t_L g2804 ( 
.A(n_2432),
.B(n_1263),
.Y(n_2804)
);

NAND2xp5_ASAP7_75t_L g2805 ( 
.A(n_2498),
.B(n_1267),
.Y(n_2805)
);

INVx1_ASAP7_75t_L g2806 ( 
.A(n_2437),
.Y(n_2806)
);

NAND2xp5_ASAP7_75t_L g2807 ( 
.A(n_2500),
.B(n_1268),
.Y(n_2807)
);

INVx1_ASAP7_75t_L g2808 ( 
.A(n_2734),
.Y(n_2808)
);

INVx2_ASAP7_75t_L g2809 ( 
.A(n_2544),
.Y(n_2809)
);

NAND2xp5_ASAP7_75t_SL g2810 ( 
.A(n_2762),
.B(n_1269),
.Y(n_2810)
);

NAND2xp5_ASAP7_75t_SL g2811 ( 
.A(n_2575),
.B(n_1276),
.Y(n_2811)
);

INVx1_ASAP7_75t_SL g2812 ( 
.A(n_2424),
.Y(n_2812)
);

INVx2_ASAP7_75t_L g2813 ( 
.A(n_2547),
.Y(n_2813)
);

INVx1_ASAP7_75t_L g2814 ( 
.A(n_2738),
.Y(n_2814)
);

INVx3_ASAP7_75t_L g2815 ( 
.A(n_2431),
.Y(n_2815)
);

NOR2xp33_ASAP7_75t_L g2816 ( 
.A(n_2689),
.B(n_1277),
.Y(n_2816)
);

INVx2_ASAP7_75t_L g2817 ( 
.A(n_2564),
.Y(n_2817)
);

INVx2_ASAP7_75t_SL g2818 ( 
.A(n_2759),
.Y(n_2818)
);

INVx3_ASAP7_75t_L g2819 ( 
.A(n_2431),
.Y(n_2819)
);

NAND2xp5_ASAP7_75t_L g2820 ( 
.A(n_2503),
.B(n_1278),
.Y(n_2820)
);

OAI22xp33_ASAP7_75t_L g2821 ( 
.A1(n_2562),
.A2(n_1283),
.B1(n_1284),
.B2(n_1280),
.Y(n_2821)
);

INVx2_ASAP7_75t_L g2822 ( 
.A(n_2740),
.Y(n_2822)
);

INVx2_ASAP7_75t_L g2823 ( 
.A(n_2744),
.Y(n_2823)
);

INVx1_ASAP7_75t_L g2824 ( 
.A(n_2745),
.Y(n_2824)
);

AOI21xp5_ASAP7_75t_L g2825 ( 
.A1(n_2594),
.A2(n_1239),
.B(n_1238),
.Y(n_2825)
);

INVx2_ASAP7_75t_L g2826 ( 
.A(n_2747),
.Y(n_2826)
);

NOR2xp33_ASAP7_75t_L g2827 ( 
.A(n_2443),
.B(n_1289),
.Y(n_2827)
);

INVx1_ASAP7_75t_L g2828 ( 
.A(n_2751),
.Y(n_2828)
);

NAND2xp5_ASAP7_75t_SL g2829 ( 
.A(n_2784),
.B(n_1293),
.Y(n_2829)
);

NOR2xp33_ASAP7_75t_L g2830 ( 
.A(n_2708),
.B(n_2474),
.Y(n_2830)
);

NOR2xp33_ASAP7_75t_L g2831 ( 
.A(n_2479),
.B(n_2417),
.Y(n_2831)
);

INVx3_ASAP7_75t_L g2832 ( 
.A(n_2431),
.Y(n_2832)
);

INVx1_ASAP7_75t_L g2833 ( 
.A(n_2775),
.Y(n_2833)
);

HB1xp67_ASAP7_75t_L g2834 ( 
.A(n_2419),
.Y(n_2834)
);

NAND2xp5_ASAP7_75t_L g2835 ( 
.A(n_2439),
.B(n_1297),
.Y(n_2835)
);

INVx1_ASAP7_75t_L g2836 ( 
.A(n_2796),
.Y(n_2836)
);

INVxp67_ASAP7_75t_L g2837 ( 
.A(n_2756),
.Y(n_2837)
);

NAND2xp5_ASAP7_75t_L g2838 ( 
.A(n_2440),
.B(n_1298),
.Y(n_2838)
);

OAI22xp5_ASAP7_75t_L g2839 ( 
.A1(n_2522),
.A2(n_2728),
.B1(n_2447),
.B2(n_2448),
.Y(n_2839)
);

NAND2xp5_ASAP7_75t_L g2840 ( 
.A(n_2442),
.B(n_1301),
.Y(n_2840)
);

NAND2xp5_ASAP7_75t_L g2841 ( 
.A(n_2456),
.B(n_1303),
.Y(n_2841)
);

INVx1_ASAP7_75t_L g2842 ( 
.A(n_2458),
.Y(n_2842)
);

OR2x6_ASAP7_75t_L g2843 ( 
.A(n_2643),
.B(n_1309),
.Y(n_2843)
);

NAND2xp5_ASAP7_75t_SL g2844 ( 
.A(n_2626),
.B(n_1304),
.Y(n_2844)
);

NAND2xp5_ASAP7_75t_L g2845 ( 
.A(n_2464),
.B(n_1312),
.Y(n_2845)
);

INVxp67_ASAP7_75t_L g2846 ( 
.A(n_2749),
.Y(n_2846)
);

A2O1A1Ixp33_ASAP7_75t_L g2847 ( 
.A1(n_2588),
.A2(n_1399),
.B(n_1423),
.C(n_1309),
.Y(n_2847)
);

AND2x2_ASAP7_75t_L g2848 ( 
.A(n_2694),
.B(n_1569),
.Y(n_2848)
);

NOR2xp33_ASAP7_75t_L g2849 ( 
.A(n_2416),
.B(n_1314),
.Y(n_2849)
);

NAND2xp5_ASAP7_75t_SL g2850 ( 
.A(n_2615),
.B(n_1317),
.Y(n_2850)
);

INVx3_ASAP7_75t_L g2851 ( 
.A(n_2481),
.Y(n_2851)
);

NAND2xp5_ASAP7_75t_L g2852 ( 
.A(n_2469),
.B(n_1318),
.Y(n_2852)
);

NAND2xp5_ASAP7_75t_L g2853 ( 
.A(n_2470),
.B(n_1319),
.Y(n_2853)
);

NAND2xp33_ASAP7_75t_L g2854 ( 
.A(n_2418),
.B(n_1320),
.Y(n_2854)
);

INVx2_ASAP7_75t_SL g2855 ( 
.A(n_2759),
.Y(n_2855)
);

AOI22xp33_ASAP7_75t_L g2856 ( 
.A1(n_2425),
.A2(n_1646),
.B1(n_1597),
.B2(n_1326),
.Y(n_2856)
);

NOR3xp33_ASAP7_75t_L g2857 ( 
.A(n_2752),
.B(n_1738),
.C(n_1246),
.Y(n_2857)
);

NAND2xp5_ASAP7_75t_L g2858 ( 
.A(n_2473),
.B(n_1323),
.Y(n_2858)
);

AND2x2_ASAP7_75t_SL g2859 ( 
.A(n_2510),
.B(n_1399),
.Y(n_2859)
);

HB1xp67_ASAP7_75t_L g2860 ( 
.A(n_2749),
.Y(n_2860)
);

NAND2xp5_ASAP7_75t_L g2861 ( 
.A(n_2476),
.B(n_1332),
.Y(n_2861)
);

AND2x2_ASAP7_75t_SL g2862 ( 
.A(n_2510),
.B(n_1423),
.Y(n_2862)
);

NAND2xp5_ASAP7_75t_SL g2863 ( 
.A(n_2735),
.B(n_2746),
.Y(n_2863)
);

NAND2xp33_ASAP7_75t_L g2864 ( 
.A(n_2418),
.B(n_1335),
.Y(n_2864)
);

NAND2xp5_ASAP7_75t_SL g2865 ( 
.A(n_2768),
.B(n_1339),
.Y(n_2865)
);

NAND2xp5_ASAP7_75t_L g2866 ( 
.A(n_2477),
.B(n_1340),
.Y(n_2866)
);

NAND2xp5_ASAP7_75t_SL g2867 ( 
.A(n_2777),
.B(n_1345),
.Y(n_2867)
);

OAI22xp5_ASAP7_75t_L g2868 ( 
.A1(n_2522),
.A2(n_1446),
.B1(n_1475),
.B2(n_1428),
.Y(n_2868)
);

NAND2xp33_ASAP7_75t_L g2869 ( 
.A(n_2459),
.B(n_1346),
.Y(n_2869)
);

OAI22xp5_ASAP7_75t_L g2870 ( 
.A1(n_2482),
.A2(n_1446),
.B1(n_1475),
.B2(n_1428),
.Y(n_2870)
);

NAND2xp5_ASAP7_75t_L g2871 ( 
.A(n_2483),
.B(n_2484),
.Y(n_2871)
);

NAND2xp5_ASAP7_75t_SL g2872 ( 
.A(n_2550),
.B(n_1347),
.Y(n_2872)
);

NAND2xp5_ASAP7_75t_SL g2873 ( 
.A(n_2421),
.B(n_1348),
.Y(n_2873)
);

NOR2xp33_ASAP7_75t_L g2874 ( 
.A(n_2435),
.B(n_1350),
.Y(n_2874)
);

NAND2xp5_ASAP7_75t_SL g2875 ( 
.A(n_2602),
.B(n_1351),
.Y(n_2875)
);

INVx1_ASAP7_75t_L g2876 ( 
.A(n_2487),
.Y(n_2876)
);

NAND2xp5_ASAP7_75t_SL g2877 ( 
.A(n_2685),
.B(n_1352),
.Y(n_2877)
);

NOR2xp33_ASAP7_75t_L g2878 ( 
.A(n_2451),
.B(n_1353),
.Y(n_2878)
);

INVx2_ASAP7_75t_L g2879 ( 
.A(n_2493),
.Y(n_2879)
);

NOR2xp33_ASAP7_75t_L g2880 ( 
.A(n_2556),
.B(n_1357),
.Y(n_2880)
);

OAI21xp33_ASAP7_75t_L g2881 ( 
.A1(n_2606),
.A2(n_1361),
.B(n_1360),
.Y(n_2881)
);

NAND2xp5_ASAP7_75t_L g2882 ( 
.A(n_2496),
.B(n_1365),
.Y(n_2882)
);

NOR2xp67_ASAP7_75t_L g2883 ( 
.A(n_2412),
.B(n_294),
.Y(n_2883)
);

INVx1_ASAP7_75t_L g2884 ( 
.A(n_2504),
.Y(n_2884)
);

NAND2xp5_ASAP7_75t_L g2885 ( 
.A(n_2449),
.B(n_1367),
.Y(n_2885)
);

BUFx3_ASAP7_75t_L g2886 ( 
.A(n_2463),
.Y(n_2886)
);

NAND2xp5_ASAP7_75t_L g2887 ( 
.A(n_2641),
.B(n_1370),
.Y(n_2887)
);

CKINVDCx5p33_ASAP7_75t_R g2888 ( 
.A(n_2520),
.Y(n_2888)
);

INVxp67_ASAP7_75t_L g2889 ( 
.A(n_2486),
.Y(n_2889)
);

INVx2_ASAP7_75t_L g2890 ( 
.A(n_2609),
.Y(n_2890)
);

INVx2_ASAP7_75t_L g2891 ( 
.A(n_2611),
.Y(n_2891)
);

CKINVDCx5p33_ASAP7_75t_R g2892 ( 
.A(n_2569),
.Y(n_2892)
);

AOI22xp33_ASAP7_75t_L g2893 ( 
.A1(n_2425),
.A2(n_2695),
.B1(n_2698),
.B2(n_2434),
.Y(n_2893)
);

NAND2xp5_ASAP7_75t_L g2894 ( 
.A(n_2452),
.B(n_1371),
.Y(n_2894)
);

INVx1_ASAP7_75t_L g2895 ( 
.A(n_2506),
.Y(n_2895)
);

NAND2xp5_ASAP7_75t_L g2896 ( 
.A(n_2453),
.B(n_1373),
.Y(n_2896)
);

NAND2xp5_ASAP7_75t_L g2897 ( 
.A(n_2414),
.B(n_2789),
.Y(n_2897)
);

NAND2xp5_ASAP7_75t_SL g2898 ( 
.A(n_2516),
.B(n_1387),
.Y(n_2898)
);

NOR2xp33_ASAP7_75t_L g2899 ( 
.A(n_2554),
.B(n_1389),
.Y(n_2899)
);

O2A1O1Ixp33_ASAP7_75t_L g2900 ( 
.A1(n_2499),
.A2(n_1250),
.B(n_1260),
.C(n_1243),
.Y(n_2900)
);

INVx2_ASAP7_75t_SL g2901 ( 
.A(n_2794),
.Y(n_2901)
);

NAND2x1_ASAP7_75t_L g2902 ( 
.A(n_2707),
.B(n_1176),
.Y(n_2902)
);

AND3x1_ASAP7_75t_L g2903 ( 
.A(n_2681),
.B(n_2604),
.C(n_2600),
.Y(n_2903)
);

INVx1_ASAP7_75t_L g2904 ( 
.A(n_2509),
.Y(n_2904)
);

AOI22xp33_ASAP7_75t_L g2905 ( 
.A1(n_2698),
.A2(n_1646),
.B1(n_1597),
.B2(n_1392),
.Y(n_2905)
);

NAND2xp33_ASAP7_75t_L g2906 ( 
.A(n_2459),
.B(n_1405),
.Y(n_2906)
);

AND2x2_ASAP7_75t_L g2907 ( 
.A(n_2532),
.B(n_1391),
.Y(n_2907)
);

NAND2xp5_ASAP7_75t_L g2908 ( 
.A(n_2414),
.B(n_1400),
.Y(n_2908)
);

AOI22xp33_ASAP7_75t_L g2909 ( 
.A1(n_2430),
.A2(n_1402),
.B1(n_1406),
.B2(n_1401),
.Y(n_2909)
);

NOR2xp33_ASAP7_75t_L g2910 ( 
.A(n_2529),
.B(n_1407),
.Y(n_2910)
);

NAND2xp5_ASAP7_75t_L g2911 ( 
.A(n_2789),
.B(n_1410),
.Y(n_2911)
);

NOR2xp33_ASAP7_75t_R g2912 ( 
.A(n_2495),
.B(n_2563),
.Y(n_2912)
);

AND2x2_ASAP7_75t_L g2913 ( 
.A(n_2445),
.B(n_2551),
.Y(n_2913)
);

OAI22xp5_ASAP7_75t_L g2914 ( 
.A1(n_2518),
.A2(n_1519),
.B1(n_1650),
.B2(n_1476),
.Y(n_2914)
);

AOI22xp33_ASAP7_75t_L g2915 ( 
.A1(n_2549),
.A2(n_1414),
.B1(n_1420),
.B2(n_1411),
.Y(n_2915)
);

BUFx3_ASAP7_75t_L g2916 ( 
.A(n_2467),
.Y(n_2916)
);

NOR2xp33_ASAP7_75t_SL g2917 ( 
.A(n_2669),
.B(n_1426),
.Y(n_2917)
);

NOR2xp67_ASAP7_75t_L g2918 ( 
.A(n_2739),
.B(n_294),
.Y(n_2918)
);

INVx2_ASAP7_75t_L g2919 ( 
.A(n_2612),
.Y(n_2919)
);

NAND2xp33_ASAP7_75t_L g2920 ( 
.A(n_2465),
.B(n_1456),
.Y(n_2920)
);

INVx3_ASAP7_75t_L g2921 ( 
.A(n_2481),
.Y(n_2921)
);

NOR2xp33_ASAP7_75t_L g2922 ( 
.A(n_2462),
.B(n_1427),
.Y(n_2922)
);

NOR2xp33_ASAP7_75t_L g2923 ( 
.A(n_2619),
.B(n_1434),
.Y(n_2923)
);

NOR2xp33_ASAP7_75t_L g2924 ( 
.A(n_2627),
.B(n_1435),
.Y(n_2924)
);

AND2x2_ASAP7_75t_L g2925 ( 
.A(n_2558),
.B(n_1438),
.Y(n_2925)
);

NOR2xp33_ASAP7_75t_L g2926 ( 
.A(n_2570),
.B(n_1439),
.Y(n_2926)
);

BUFx6f_ASAP7_75t_L g2927 ( 
.A(n_2465),
.Y(n_2927)
);

NAND2xp5_ASAP7_75t_L g2928 ( 
.A(n_2542),
.B(n_1445),
.Y(n_2928)
);

BUFx6f_ASAP7_75t_SL g2929 ( 
.A(n_2527),
.Y(n_2929)
);

INVx2_ASAP7_75t_L g2930 ( 
.A(n_2616),
.Y(n_2930)
);

INVx2_ASAP7_75t_SL g2931 ( 
.A(n_2794),
.Y(n_2931)
);

AND2x2_ASAP7_75t_L g2932 ( 
.A(n_2754),
.B(n_1448),
.Y(n_2932)
);

NAND2xp5_ASAP7_75t_L g2933 ( 
.A(n_2472),
.B(n_1449),
.Y(n_2933)
);

INVx2_ASAP7_75t_L g2934 ( 
.A(n_2617),
.Y(n_2934)
);

NAND2xp5_ASAP7_75t_L g2935 ( 
.A(n_2525),
.B(n_1453),
.Y(n_2935)
);

AND2x6_ASAP7_75t_L g2936 ( 
.A(n_2517),
.B(n_1176),
.Y(n_2936)
);

AOI22xp33_ASAP7_75t_L g2937 ( 
.A1(n_2507),
.A2(n_1461),
.B1(n_1464),
.B2(n_1454),
.Y(n_2937)
);

AOI221xp5_ASAP7_75t_L g2938 ( 
.A1(n_2466),
.A2(n_1473),
.B1(n_1480),
.B2(n_1470),
.C(n_1468),
.Y(n_2938)
);

AOI22xp5_ASAP7_75t_L g2939 ( 
.A1(n_2573),
.A2(n_1492),
.B1(n_1494),
.B2(n_1491),
.Y(n_2939)
);

INVx2_ASAP7_75t_L g2940 ( 
.A(n_2523),
.Y(n_2940)
);

BUFx5_ASAP7_75t_L g2941 ( 
.A(n_2707),
.Y(n_2941)
);

NAND2xp33_ASAP7_75t_L g2942 ( 
.A(n_2517),
.B(n_1518),
.Y(n_2942)
);

NAND2xp5_ASAP7_75t_L g2943 ( 
.A(n_2534),
.B(n_1504),
.Y(n_2943)
);

AND2x2_ASAP7_75t_SL g2944 ( 
.A(n_2516),
.B(n_1476),
.Y(n_2944)
);

INVx1_ASAP7_75t_L g2945 ( 
.A(n_2531),
.Y(n_2945)
);

NAND2xp5_ASAP7_75t_SL g2946 ( 
.A(n_2533),
.B(n_1505),
.Y(n_2946)
);

INVx3_ASAP7_75t_L g2947 ( 
.A(n_2481),
.Y(n_2947)
);

AOI22xp5_ASAP7_75t_L g2948 ( 
.A1(n_2603),
.A2(n_1516),
.B1(n_1520),
.B2(n_1510),
.Y(n_2948)
);

NAND2xp5_ASAP7_75t_L g2949 ( 
.A(n_2631),
.B(n_1523),
.Y(n_2949)
);

NOR2xp33_ASAP7_75t_L g2950 ( 
.A(n_2533),
.B(n_1526),
.Y(n_2950)
);

NAND2xp5_ASAP7_75t_L g2951 ( 
.A(n_2631),
.B(n_1527),
.Y(n_2951)
);

INVx1_ASAP7_75t_L g2952 ( 
.A(n_2536),
.Y(n_2952)
);

HB1xp67_ASAP7_75t_L g2953 ( 
.A(n_2760),
.Y(n_2953)
);

NAND2xp5_ASAP7_75t_L g2954 ( 
.A(n_2743),
.B(n_1529),
.Y(n_2954)
);

NAND2xp5_ASAP7_75t_L g2955 ( 
.A(n_2753),
.B(n_1532),
.Y(n_2955)
);

INVx1_ASAP7_75t_L g2956 ( 
.A(n_2540),
.Y(n_2956)
);

NAND2xp5_ASAP7_75t_SL g2957 ( 
.A(n_2653),
.B(n_1533),
.Y(n_2957)
);

INVx2_ASAP7_75t_L g2958 ( 
.A(n_2545),
.Y(n_2958)
);

NAND2xp5_ASAP7_75t_SL g2959 ( 
.A(n_2670),
.B(n_1540),
.Y(n_2959)
);

BUFx3_ASAP7_75t_L g2960 ( 
.A(n_2781),
.Y(n_2960)
);

INVx1_ASAP7_75t_L g2961 ( 
.A(n_2546),
.Y(n_2961)
);

AND2x4_ASAP7_75t_L g2962 ( 
.A(n_2519),
.B(n_1265),
.Y(n_2962)
);

OAI22xp33_ASAP7_75t_L g2963 ( 
.A1(n_2733),
.A2(n_1543),
.B1(n_1544),
.B2(n_1541),
.Y(n_2963)
);

NAND2xp5_ASAP7_75t_L g2964 ( 
.A(n_2757),
.B(n_2767),
.Y(n_2964)
);

NAND2xp5_ASAP7_75t_SL g2965 ( 
.A(n_2528),
.B(n_2770),
.Y(n_2965)
);

INVx2_ASAP7_75t_L g2966 ( 
.A(n_2553),
.Y(n_2966)
);

NAND2xp5_ASAP7_75t_L g2967 ( 
.A(n_2769),
.B(n_1548),
.Y(n_2967)
);

INVx2_ASAP7_75t_L g2968 ( 
.A(n_2555),
.Y(n_2968)
);

INVx1_ASAP7_75t_L g2969 ( 
.A(n_2559),
.Y(n_2969)
);

NAND2xp5_ASAP7_75t_L g2970 ( 
.A(n_2779),
.B(n_2783),
.Y(n_2970)
);

NOR2xp33_ASAP7_75t_L g2971 ( 
.A(n_2436),
.B(n_1549),
.Y(n_2971)
);

NOR2xp33_ASAP7_75t_L g2972 ( 
.A(n_2772),
.B(n_2786),
.Y(n_2972)
);

AND2x6_ASAP7_75t_SL g2973 ( 
.A(n_2643),
.B(n_1266),
.Y(n_2973)
);

NOR2xp33_ASAP7_75t_L g2974 ( 
.A(n_2787),
.B(n_1550),
.Y(n_2974)
);

INVx1_ASAP7_75t_L g2975 ( 
.A(n_2561),
.Y(n_2975)
);

INVx3_ASAP7_75t_L g2976 ( 
.A(n_2519),
.Y(n_2976)
);

NAND2xp5_ASAP7_75t_SL g2977 ( 
.A(n_2576),
.B(n_1552),
.Y(n_2977)
);

NOR2xp33_ASAP7_75t_L g2978 ( 
.A(n_2679),
.B(n_1553),
.Y(n_2978)
);

INVx2_ASAP7_75t_L g2979 ( 
.A(n_2566),
.Y(n_2979)
);

NAND2xp5_ASAP7_75t_L g2980 ( 
.A(n_2582),
.B(n_1554),
.Y(n_2980)
);

INVx1_ASAP7_75t_L g2981 ( 
.A(n_2585),
.Y(n_2981)
);

CKINVDCx20_ASAP7_75t_R g2982 ( 
.A(n_2776),
.Y(n_2982)
);

AOI22xp5_ASAP7_75t_L g2983 ( 
.A1(n_2785),
.A2(n_1559),
.B1(n_1562),
.B2(n_1558),
.Y(n_2983)
);

AOI22xp5_ASAP7_75t_L g2984 ( 
.A1(n_2480),
.A2(n_1565),
.B1(n_1566),
.B2(n_1564),
.Y(n_2984)
);

NAND2xp5_ASAP7_75t_L g2985 ( 
.A(n_2589),
.B(n_1567),
.Y(n_2985)
);

BUFx6f_ASAP7_75t_L g2986 ( 
.A(n_2526),
.Y(n_2986)
);

NOR2xp33_ASAP7_75t_L g2987 ( 
.A(n_2490),
.B(n_1568),
.Y(n_2987)
);

NAND2xp5_ASAP7_75t_SL g2988 ( 
.A(n_2576),
.B(n_1570),
.Y(n_2988)
);

A2O1A1Ixp33_ASAP7_75t_L g2989 ( 
.A1(n_2797),
.A2(n_1650),
.B(n_1675),
.C(n_1519),
.Y(n_2989)
);

NAND2xp5_ASAP7_75t_L g2990 ( 
.A(n_2511),
.B(n_1574),
.Y(n_2990)
);

NAND2xp5_ASAP7_75t_L g2991 ( 
.A(n_2511),
.B(n_1576),
.Y(n_2991)
);

NAND2xp5_ASAP7_75t_L g2992 ( 
.A(n_2593),
.B(n_1579),
.Y(n_2992)
);

OR2x2_ASAP7_75t_L g2993 ( 
.A(n_2524),
.B(n_1581),
.Y(n_2993)
);

NAND2xp5_ASAP7_75t_L g2994 ( 
.A(n_2548),
.B(n_1587),
.Y(n_2994)
);

NAND2xp5_ASAP7_75t_L g2995 ( 
.A(n_2584),
.B(n_1589),
.Y(n_2995)
);

INVx1_ASAP7_75t_L g2996 ( 
.A(n_2423),
.Y(n_2996)
);

AND2x2_ASAP7_75t_SL g2997 ( 
.A(n_2642),
.B(n_1675),
.Y(n_2997)
);

INVx2_ASAP7_75t_L g2998 ( 
.A(n_2608),
.Y(n_2998)
);

BUFx6f_ASAP7_75t_L g2999 ( 
.A(n_2526),
.Y(n_2999)
);

NAND2xp5_ASAP7_75t_L g3000 ( 
.A(n_2610),
.B(n_1593),
.Y(n_3000)
);

NOR2xp33_ASAP7_75t_L g3001 ( 
.A(n_2676),
.B(n_1586),
.Y(n_3001)
);

NAND2xp5_ASAP7_75t_L g3002 ( 
.A(n_2610),
.B(n_1596),
.Y(n_3002)
);

NAND2xp5_ASAP7_75t_SL g3003 ( 
.A(n_2729),
.B(n_1601),
.Y(n_3003)
);

NAND2xp5_ASAP7_75t_L g3004 ( 
.A(n_2491),
.B(n_2672),
.Y(n_3004)
);

NAND2xp5_ASAP7_75t_L g3005 ( 
.A(n_2624),
.B(n_1603),
.Y(n_3005)
);

NAND2xp5_ASAP7_75t_L g3006 ( 
.A(n_2433),
.B(n_1611),
.Y(n_3006)
);

O2A1O1Ixp5_ASAP7_75t_L g3007 ( 
.A1(n_2725),
.A2(n_1734),
.B(n_1271),
.C(n_1272),
.Y(n_3007)
);

AOI22xp33_ASAP7_75t_L g3008 ( 
.A1(n_2507),
.A2(n_1615),
.B1(n_1617),
.B2(n_1607),
.Y(n_3008)
);

NOR2xp33_ASAP7_75t_L g3009 ( 
.A(n_2457),
.B(n_1618),
.Y(n_3009)
);

INVxp67_ASAP7_75t_SL g3010 ( 
.A(n_2798),
.Y(n_3010)
);

AND2x4_ASAP7_75t_L g3011 ( 
.A(n_2519),
.B(n_1270),
.Y(n_3011)
);

INVx1_ASAP7_75t_L g3012 ( 
.A(n_2423),
.Y(n_3012)
);

NAND2xp5_ASAP7_75t_L g3013 ( 
.A(n_2433),
.B(n_1620),
.Y(n_3013)
);

NAND2xp5_ASAP7_75t_SL g3014 ( 
.A(n_2782),
.B(n_1623),
.Y(n_3014)
);

BUFx12f_ASAP7_75t_L g3015 ( 
.A(n_2648),
.Y(n_3015)
);

NAND2xp5_ASAP7_75t_L g3016 ( 
.A(n_2433),
.B(n_1627),
.Y(n_3016)
);

NAND2xp5_ASAP7_75t_L g3017 ( 
.A(n_2461),
.B(n_1632),
.Y(n_3017)
);

NAND2xp5_ASAP7_75t_L g3018 ( 
.A(n_2461),
.B(n_1638),
.Y(n_3018)
);

INVx2_ASAP7_75t_L g3019 ( 
.A(n_2438),
.Y(n_3019)
);

AOI22xp33_ASAP7_75t_L g3020 ( 
.A1(n_2700),
.A2(n_1641),
.B1(n_1643),
.B2(n_1639),
.Y(n_3020)
);

INVx2_ASAP7_75t_L g3021 ( 
.A(n_2441),
.Y(n_3021)
);

OAI22xp33_ASAP7_75t_L g3022 ( 
.A1(n_2651),
.A2(n_1647),
.B1(n_1649),
.B2(n_1645),
.Y(n_3022)
);

NAND2xp5_ASAP7_75t_L g3023 ( 
.A(n_2657),
.B(n_1653),
.Y(n_3023)
);

OAI22xp5_ASAP7_75t_L g3024 ( 
.A1(n_2651),
.A2(n_1734),
.B1(n_1176),
.B2(n_1198),
.Y(n_3024)
);

AOI22xp33_ASAP7_75t_L g3025 ( 
.A1(n_2700),
.A2(n_1667),
.B1(n_1669),
.B2(n_1657),
.Y(n_3025)
);

AOI22xp33_ASAP7_75t_L g3026 ( 
.A1(n_2601),
.A2(n_1680),
.B1(n_1690),
.B2(n_1674),
.Y(n_3026)
);

NAND2xp5_ASAP7_75t_SL g3027 ( 
.A(n_2782),
.B(n_1696),
.Y(n_3027)
);

NAND2xp5_ASAP7_75t_L g3028 ( 
.A(n_2657),
.B(n_1705),
.Y(n_3028)
);

OAI21xp5_ASAP7_75t_L g3029 ( 
.A1(n_2460),
.A2(n_2475),
.B(n_2471),
.Y(n_3029)
);

INVx1_ASAP7_75t_L g3030 ( 
.A(n_2587),
.Y(n_3030)
);

INVx1_ASAP7_75t_L g3031 ( 
.A(n_2590),
.Y(n_3031)
);

NOR2xp33_ASAP7_75t_L g3032 ( 
.A(n_2478),
.B(n_1706),
.Y(n_3032)
);

INVx2_ASAP7_75t_L g3033 ( 
.A(n_2508),
.Y(n_3033)
);

AOI221xp5_ASAP7_75t_L g3034 ( 
.A1(n_2574),
.A2(n_2485),
.B1(n_2568),
.B2(n_2543),
.C(n_2571),
.Y(n_3034)
);

INVx2_ASAP7_75t_L g3035 ( 
.A(n_2515),
.Y(n_3035)
);

INVx2_ASAP7_75t_SL g3036 ( 
.A(n_2599),
.Y(n_3036)
);

INVx2_ASAP7_75t_SL g3037 ( 
.A(n_2599),
.Y(n_3037)
);

NOR2xp33_ASAP7_75t_SL g3038 ( 
.A(n_2639),
.B(n_1709),
.Y(n_3038)
);

NOR3x1_ASAP7_75t_L g3039 ( 
.A(n_2673),
.B(n_1741),
.C(n_1720),
.Y(n_3039)
);

NAND2xp5_ASAP7_75t_SL g3040 ( 
.A(n_2782),
.B(n_2592),
.Y(n_3040)
);

BUFx3_ASAP7_75t_L g3041 ( 
.A(n_2629),
.Y(n_3041)
);

INVx1_ASAP7_75t_L g3042 ( 
.A(n_2622),
.Y(n_3042)
);

OA22x2_ASAP7_75t_L g3043 ( 
.A1(n_2683),
.A2(n_1722),
.B1(n_1723),
.B2(n_1718),
.Y(n_3043)
);

A2O1A1Ixp33_ASAP7_75t_L g3044 ( 
.A1(n_2591),
.A2(n_1281),
.B(n_1285),
.C(n_1275),
.Y(n_3044)
);

NAND2xp5_ASAP7_75t_L g3045 ( 
.A(n_2541),
.B(n_1713),
.Y(n_3045)
);

AOI22xp33_ASAP7_75t_L g3046 ( 
.A1(n_2645),
.A2(n_1716),
.B1(n_1724),
.B2(n_1715),
.Y(n_3046)
);

INVx2_ASAP7_75t_L g3047 ( 
.A(n_2521),
.Y(n_3047)
);

CKINVDCx5p33_ASAP7_75t_R g3048 ( 
.A(n_2648),
.Y(n_3048)
);

NAND2xp5_ASAP7_75t_L g3049 ( 
.A(n_2773),
.B(n_1727),
.Y(n_3049)
);

NAND2xp5_ASAP7_75t_L g3050 ( 
.A(n_2614),
.B(n_1728),
.Y(n_3050)
);

INVx1_ASAP7_75t_L g3051 ( 
.A(n_2625),
.Y(n_3051)
);

AOI22xp5_ASAP7_75t_L g3052 ( 
.A1(n_2621),
.A2(n_1733),
.B1(n_1736),
.B2(n_1731),
.Y(n_3052)
);

AOI22xp33_ASAP7_75t_L g3053 ( 
.A1(n_2650),
.A2(n_1746),
.B1(n_1750),
.B2(n_1745),
.Y(n_3053)
);

OR2x2_ASAP7_75t_L g3054 ( 
.A(n_2488),
.B(n_1288),
.Y(n_3054)
);

INVx2_ASAP7_75t_L g3055 ( 
.A(n_2567),
.Y(n_3055)
);

NAND2xp5_ASAP7_75t_L g3056 ( 
.A(n_2635),
.B(n_1292),
.Y(n_3056)
);

AOI22xp33_ASAP7_75t_L g3057 ( 
.A1(n_2652),
.A2(n_1556),
.B1(n_1707),
.B2(n_1471),
.Y(n_3057)
);

NAND2xp5_ASAP7_75t_L g3058 ( 
.A(n_2636),
.B(n_1295),
.Y(n_3058)
);

NOR2xp33_ASAP7_75t_L g3059 ( 
.A(n_2514),
.B(n_1305),
.Y(n_3059)
);

NAND2xp5_ASAP7_75t_L g3060 ( 
.A(n_2623),
.B(n_1310),
.Y(n_3060)
);

INVx1_ASAP7_75t_L g3061 ( 
.A(n_2686),
.Y(n_3061)
);

NAND2xp5_ASAP7_75t_SL g3062 ( 
.A(n_2661),
.B(n_1175),
.Y(n_3062)
);

NAND2xp33_ASAP7_75t_L g3063 ( 
.A(n_2537),
.B(n_1471),
.Y(n_3063)
);

NAND2xp5_ASAP7_75t_L g3064 ( 
.A(n_2637),
.B(n_1311),
.Y(n_3064)
);

NAND2xp5_ASAP7_75t_L g3065 ( 
.A(n_2649),
.B(n_1315),
.Y(n_3065)
);

NAND2xp5_ASAP7_75t_SL g3066 ( 
.A(n_2595),
.B(n_2598),
.Y(n_3066)
);

NAND2xp5_ASAP7_75t_L g3067 ( 
.A(n_2560),
.B(n_2613),
.Y(n_3067)
);

NAND2xp5_ASAP7_75t_SL g3068 ( 
.A(n_2629),
.B(n_2687),
.Y(n_3068)
);

AOI22xp33_ASAP7_75t_L g3069 ( 
.A1(n_2654),
.A2(n_1556),
.B1(n_1707),
.B2(n_1471),
.Y(n_3069)
);

NAND2xp5_ASAP7_75t_L g3070 ( 
.A(n_2655),
.B(n_1316),
.Y(n_3070)
);

INVxp67_ASAP7_75t_L g3071 ( 
.A(n_2691),
.Y(n_3071)
);

NOR2xp33_ASAP7_75t_L g3072 ( 
.A(n_2530),
.B(n_1324),
.Y(n_3072)
);

INVx1_ASAP7_75t_L g3073 ( 
.A(n_2715),
.Y(n_3073)
);

NAND2xp5_ASAP7_75t_SL g3074 ( 
.A(n_2687),
.B(n_1175),
.Y(n_3074)
);

OR2x6_ASAP7_75t_L g3075 ( 
.A(n_2455),
.B(n_1343),
.Y(n_3075)
);

OAI22xp5_ASAP7_75t_L g3076 ( 
.A1(n_2690),
.A2(n_1176),
.B1(n_1198),
.B2(n_1187),
.Y(n_3076)
);

OAI21xp5_ASAP7_75t_L g3077 ( 
.A1(n_2420),
.A2(n_1375),
.B(n_1366),
.Y(n_3077)
);

AOI22x1_ASAP7_75t_L g3078 ( 
.A1(n_2731),
.A2(n_1187),
.B1(n_1338),
.B2(n_1198),
.Y(n_3078)
);

INVx1_ASAP7_75t_L g3079 ( 
.A(n_2726),
.Y(n_3079)
);

INVx2_ASAP7_75t_L g3080 ( 
.A(n_2658),
.Y(n_3080)
);

INVx1_ASAP7_75t_L g3081 ( 
.A(n_2730),
.Y(n_3081)
);

INVx2_ASAP7_75t_SL g3082 ( 
.A(n_2693),
.Y(n_3082)
);

NAND2xp5_ASAP7_75t_L g3083 ( 
.A(n_2682),
.B(n_1380),
.Y(n_3083)
);

INVx2_ASAP7_75t_L g3084 ( 
.A(n_2750),
.Y(n_3084)
);

AOI22xp5_ASAP7_75t_L g3085 ( 
.A1(n_2632),
.A2(n_1432),
.B1(n_1433),
.B2(n_1386),
.Y(n_3085)
);

INVx1_ASAP7_75t_L g3086 ( 
.A(n_2748),
.Y(n_3086)
);

NOR2xp33_ASAP7_75t_L g3087 ( 
.A(n_2607),
.B(n_1437),
.Y(n_3087)
);

NAND2xp33_ASAP7_75t_L g3088 ( 
.A(n_2537),
.B(n_1471),
.Y(n_3088)
);

INVx1_ASAP7_75t_L g3089 ( 
.A(n_2628),
.Y(n_3089)
);

NAND2xp5_ASAP7_75t_L g3090 ( 
.A(n_2638),
.B(n_1440),
.Y(n_3090)
);

NAND2xp5_ASAP7_75t_L g3091 ( 
.A(n_2675),
.B(n_1443),
.Y(n_3091)
);

INVx2_ASAP7_75t_L g3092 ( 
.A(n_2755),
.Y(n_3092)
);

AOI22xp5_ASAP7_75t_L g3093 ( 
.A1(n_2428),
.A2(n_1450),
.B1(n_1452),
.B2(n_1444),
.Y(n_3093)
);

INVx2_ASAP7_75t_L g3094 ( 
.A(n_2766),
.Y(n_3094)
);

NOR2xp33_ASAP7_75t_SL g3095 ( 
.A(n_2761),
.B(n_2764),
.Y(n_3095)
);

INVx1_ASAP7_75t_L g3096 ( 
.A(n_2539),
.Y(n_3096)
);

OAI22xp5_ASAP7_75t_L g3097 ( 
.A1(n_2774),
.A2(n_1187),
.B1(n_1338),
.B2(n_1198),
.Y(n_3097)
);

NAND2xp5_ASAP7_75t_SL g3098 ( 
.A(n_2693),
.B(n_1175),
.Y(n_3098)
);

INVx2_ASAP7_75t_L g3099 ( 
.A(n_2791),
.Y(n_3099)
);

INVx1_ASAP7_75t_L g3100 ( 
.A(n_2721),
.Y(n_3100)
);

NAND2xp5_ASAP7_75t_L g3101 ( 
.A(n_2663),
.B(n_1457),
.Y(n_3101)
);

BUFx8_ASAP7_75t_L g3102 ( 
.A(n_2605),
.Y(n_3102)
);

INVx2_ASAP7_75t_L g3103 ( 
.A(n_2792),
.Y(n_3103)
);

INVx2_ASAP7_75t_L g3104 ( 
.A(n_2557),
.Y(n_3104)
);

NAND2xp5_ASAP7_75t_L g3105 ( 
.A(n_2633),
.B(n_1458),
.Y(n_3105)
);

NAND2xp5_ASAP7_75t_L g3106 ( 
.A(n_2692),
.B(n_1459),
.Y(n_3106)
);

NAND2xp5_ASAP7_75t_L g3107 ( 
.A(n_2710),
.B(n_1460),
.Y(n_3107)
);

NAND2xp5_ASAP7_75t_L g3108 ( 
.A(n_2719),
.B(n_1467),
.Y(n_3108)
);

NOR3xp33_ASAP7_75t_L g3109 ( 
.A(n_2620),
.B(n_1687),
.C(n_1679),
.Y(n_3109)
);

BUFx3_ASAP7_75t_L g3110 ( 
.A(n_2413),
.Y(n_3110)
);

INVx2_ASAP7_75t_L g3111 ( 
.A(n_2557),
.Y(n_3111)
);

INVx1_ASAP7_75t_L g3112 ( 
.A(n_2716),
.Y(n_3112)
);

NAND2xp5_ASAP7_75t_L g3113 ( 
.A(n_2630),
.B(n_1469),
.Y(n_3113)
);

AOI22xp5_ASAP7_75t_L g3114 ( 
.A1(n_2660),
.A2(n_1495),
.B1(n_1501),
.B2(n_1500),
.Y(n_3114)
);

INVx2_ASAP7_75t_L g3115 ( 
.A(n_2572),
.Y(n_3115)
);

NOR2xp67_ASAP7_75t_L g3116 ( 
.A(n_2671),
.B(n_294),
.Y(n_3116)
);

OAI22xp33_ASAP7_75t_L g3117 ( 
.A1(n_2454),
.A2(n_1515),
.B1(n_1539),
.B2(n_1512),
.Y(n_3117)
);

INVx1_ASAP7_75t_L g3118 ( 
.A(n_2580),
.Y(n_3118)
);

INVx2_ASAP7_75t_L g3119 ( 
.A(n_2572),
.Y(n_3119)
);

INVxp67_ASAP7_75t_L g3120 ( 
.A(n_2691),
.Y(n_3120)
);

NAND2xp5_ASAP7_75t_L g3121 ( 
.A(n_2597),
.B(n_1542),
.Y(n_3121)
);

AOI22xp33_ASAP7_75t_SL g3122 ( 
.A1(n_2697),
.A2(n_1556),
.B1(n_1707),
.B2(n_1471),
.Y(n_3122)
);

BUFx6f_ASAP7_75t_L g3123 ( 
.A(n_2577),
.Y(n_3123)
);

INVx8_ASAP7_75t_L g3124 ( 
.A(n_2413),
.Y(n_3124)
);

INVx1_ASAP7_75t_L g3125 ( 
.A(n_2580),
.Y(n_3125)
);

NOR2xp33_ASAP7_75t_L g3126 ( 
.A(n_2702),
.B(n_1546),
.Y(n_3126)
);

NAND2xp5_ASAP7_75t_SL g3127 ( 
.A(n_2688),
.B(n_1175),
.Y(n_3127)
);

NAND2xp5_ASAP7_75t_L g3128 ( 
.A(n_2512),
.B(n_1572),
.Y(n_3128)
);

NAND2xp5_ASAP7_75t_L g3129 ( 
.A(n_2618),
.B(n_1580),
.Y(n_3129)
);

OR2x2_ASAP7_75t_L g3130 ( 
.A(n_2488),
.B(n_1584),
.Y(n_3130)
);

NAND2xp5_ASAP7_75t_SL g3131 ( 
.A(n_2577),
.B(n_1264),
.Y(n_3131)
);

AOI22xp33_ASAP7_75t_L g3132 ( 
.A1(n_2468),
.A2(n_1707),
.B1(n_1556),
.B2(n_1590),
.Y(n_3132)
);

NAND2xp5_ASAP7_75t_L g3133 ( 
.A(n_2426),
.B(n_2780),
.Y(n_3133)
);

NAND2xp5_ASAP7_75t_L g3134 ( 
.A(n_2426),
.B(n_1588),
.Y(n_3134)
);

NAND2xp5_ASAP7_75t_SL g3135 ( 
.A(n_2765),
.B(n_1264),
.Y(n_3135)
);

NAND2xp5_ASAP7_75t_L g3136 ( 
.A(n_2765),
.B(n_1591),
.Y(n_3136)
);

BUFx3_ASAP7_75t_L g3137 ( 
.A(n_2780),
.Y(n_3137)
);

NAND2xp5_ASAP7_75t_SL g3138 ( 
.A(n_2793),
.B(n_1264),
.Y(n_3138)
);

NAND2xp5_ASAP7_75t_L g3139 ( 
.A(n_2793),
.B(n_1594),
.Y(n_3139)
);

INVx1_ASAP7_75t_L g3140 ( 
.A(n_2701),
.Y(n_3140)
);

INVxp67_ASAP7_75t_L g3141 ( 
.A(n_2505),
.Y(n_3141)
);

INVx2_ASAP7_75t_L g3142 ( 
.A(n_2586),
.Y(n_3142)
);

NAND2xp5_ASAP7_75t_L g3143 ( 
.A(n_2422),
.B(n_1595),
.Y(n_3143)
);

AOI22xp33_ASAP7_75t_L g3144 ( 
.A1(n_2696),
.A2(n_1707),
.B1(n_1556),
.B2(n_1602),
.Y(n_3144)
);

NAND2xp5_ASAP7_75t_L g3145 ( 
.A(n_2737),
.B(n_1599),
.Y(n_3145)
);

INVx1_ASAP7_75t_L g3146 ( 
.A(n_2680),
.Y(n_3146)
);

NAND2xp5_ASAP7_75t_SL g3147 ( 
.A(n_2664),
.B(n_1264),
.Y(n_3147)
);

NOR2x1_ASAP7_75t_L g3148 ( 
.A(n_2656),
.B(n_1606),
.Y(n_3148)
);

NAND2xp5_ASAP7_75t_L g3149 ( 
.A(n_2742),
.B(n_1609),
.Y(n_3149)
);

HB1xp67_ASAP7_75t_L g3150 ( 
.A(n_2640),
.Y(n_3150)
);

NAND2xp5_ASAP7_75t_L g3151 ( 
.A(n_2758),
.B(n_1612),
.Y(n_3151)
);

BUFx6f_ASAP7_75t_L g3152 ( 
.A(n_2707),
.Y(n_3152)
);

INVx2_ASAP7_75t_SL g3153 ( 
.A(n_2581),
.Y(n_3153)
);

INVx1_ASAP7_75t_L g3154 ( 
.A(n_2718),
.Y(n_3154)
);

NAND2xp5_ASAP7_75t_SL g3155 ( 
.A(n_2664),
.B(n_1290),
.Y(n_3155)
);

AOI22xp5_ASAP7_75t_L g3156 ( 
.A1(n_2665),
.A2(n_1622),
.B1(n_1630),
.B2(n_1625),
.Y(n_3156)
);

INVx1_ASAP7_75t_L g3157 ( 
.A(n_2699),
.Y(n_3157)
);

NOR2xp33_ASAP7_75t_L g3158 ( 
.A(n_2644),
.B(n_1640),
.Y(n_3158)
);

O2A1O1Ixp33_ASAP7_75t_L g3159 ( 
.A1(n_2429),
.A2(n_1660),
.B(n_1668),
.C(n_1661),
.Y(n_3159)
);

AOI22xp5_ASAP7_75t_L g3160 ( 
.A1(n_2494),
.A2(n_1676),
.B1(n_1688),
.B2(n_1677),
.Y(n_3160)
);

NAND2xp5_ASAP7_75t_L g3161 ( 
.A(n_2763),
.B(n_1691),
.Y(n_3161)
);

INVx3_ASAP7_75t_L g3162 ( 
.A(n_2712),
.Y(n_3162)
);

NAND2xp5_ASAP7_75t_SL g3163 ( 
.A(n_2717),
.B(n_1290),
.Y(n_3163)
);

BUFx6f_ASAP7_75t_L g3164 ( 
.A(n_2712),
.Y(n_3164)
);

NOR2xp33_ASAP7_75t_L g3165 ( 
.A(n_2659),
.B(n_2497),
.Y(n_3165)
);

NAND2xp5_ASAP7_75t_SL g3166 ( 
.A(n_2489),
.B(n_2492),
.Y(n_3166)
);

INVx2_ASAP7_75t_SL g3167 ( 
.A(n_2646),
.Y(n_3167)
);

BUFx6f_ASAP7_75t_L g3168 ( 
.A(n_2788),
.Y(n_3168)
);

NAND3xp33_ASAP7_75t_L g3169 ( 
.A(n_2565),
.B(n_1338),
.C(n_1187),
.Y(n_3169)
);

INVx1_ASAP7_75t_L g3170 ( 
.A(n_2703),
.Y(n_3170)
);

OR2x2_ASAP7_75t_SL g3171 ( 
.A(n_2444),
.B(n_1700),
.Y(n_3171)
);

OAI21xp5_ASAP7_75t_L g3172 ( 
.A1(n_2647),
.A2(n_2678),
.B(n_2662),
.Y(n_3172)
);

INVx2_ASAP7_75t_L g3173 ( 
.A(n_2684),
.Y(n_3173)
);

NAND2xp5_ASAP7_75t_L g3174 ( 
.A(n_2799),
.B(n_1702),
.Y(n_3174)
);

NAND2xp5_ASAP7_75t_SL g3175 ( 
.A(n_2513),
.B(n_1290),
.Y(n_3175)
);

INVx2_ASAP7_75t_L g3176 ( 
.A(n_2727),
.Y(n_3176)
);

NAND2xp5_ASAP7_75t_SL g3177 ( 
.A(n_2552),
.B(n_1290),
.Y(n_3177)
);

INVxp33_ASAP7_75t_L g3178 ( 
.A(n_2502),
.Y(n_3178)
);

INVx2_ASAP7_75t_L g3179 ( 
.A(n_2634),
.Y(n_3179)
);

NAND2xp5_ASAP7_75t_L g3180 ( 
.A(n_2704),
.B(n_1703),
.Y(n_3180)
);

AOI22xp5_ASAP7_75t_L g3181 ( 
.A1(n_2535),
.A2(n_1704),
.B1(n_1712),
.B2(n_1711),
.Y(n_3181)
);

NAND2xp5_ASAP7_75t_L g3182 ( 
.A(n_2706),
.B(n_1717),
.Y(n_3182)
);

NAND2xp5_ASAP7_75t_SL g3183 ( 
.A(n_2427),
.B(n_1300),
.Y(n_3183)
);

NAND2xp5_ASAP7_75t_L g3184 ( 
.A(n_2714),
.B(n_1747),
.Y(n_3184)
);

INVx2_ASAP7_75t_SL g3185 ( 
.A(n_2444),
.Y(n_3185)
);

NOR2xp67_ASAP7_75t_L g3186 ( 
.A(n_2667),
.B(n_295),
.Y(n_3186)
);

NAND2xp33_ASAP7_75t_L g3187 ( 
.A(n_2795),
.B(n_1556),
.Y(n_3187)
);

INVx2_ASAP7_75t_L g3188 ( 
.A(n_2634),
.Y(n_3188)
);

AND2x2_ASAP7_75t_L g3189 ( 
.A(n_2450),
.B(n_1556),
.Y(n_3189)
);

NAND2xp5_ASAP7_75t_SL g3190 ( 
.A(n_2790),
.B(n_1300),
.Y(n_3190)
);

AOI22xp33_ASAP7_75t_L g3191 ( 
.A1(n_2578),
.A2(n_1707),
.B1(n_1338),
.B2(n_1364),
.Y(n_3191)
);

INVx1_ASAP7_75t_L g3192 ( 
.A(n_2723),
.Y(n_3192)
);

HB1xp67_ASAP7_75t_L g3193 ( 
.A(n_2450),
.Y(n_3193)
);

NOR3xp33_ASAP7_75t_L g3194 ( 
.A(n_2736),
.B(n_1707),
.C(n_290),
.Y(n_3194)
);

NAND2xp5_ASAP7_75t_L g3195 ( 
.A(n_2790),
.B(n_2),
.Y(n_3195)
);

NOR2xp33_ASAP7_75t_L g3196 ( 
.A(n_2713),
.B(n_288),
.Y(n_3196)
);

NAND2xp5_ASAP7_75t_L g3197 ( 
.A(n_2741),
.B(n_2),
.Y(n_3197)
);

INVx2_ASAP7_75t_L g3198 ( 
.A(n_2634),
.Y(n_3198)
);

INVx1_ASAP7_75t_L g3199 ( 
.A(n_2724),
.Y(n_3199)
);

NAND2xp5_ASAP7_75t_L g3200 ( 
.A(n_2771),
.B(n_2),
.Y(n_3200)
);

NOR2xp67_ASAP7_75t_SL g3201 ( 
.A(n_2579),
.B(n_1300),
.Y(n_3201)
);

NAND2xp5_ASAP7_75t_L g3202 ( 
.A(n_2501),
.B(n_2),
.Y(n_3202)
);

NOR2xp33_ASAP7_75t_L g3203 ( 
.A(n_2583),
.B(n_288),
.Y(n_3203)
);

AOI21xp5_ASAP7_75t_L g3204 ( 
.A1(n_2709),
.A2(n_1342),
.B(n_1300),
.Y(n_3204)
);

AND2x2_ASAP7_75t_L g3205 ( 
.A(n_2501),
.B(n_288),
.Y(n_3205)
);

NAND2xp5_ASAP7_75t_L g3206 ( 
.A(n_2596),
.B(n_3),
.Y(n_3206)
);

NAND3xp33_ASAP7_75t_L g3207 ( 
.A(n_2732),
.B(n_1364),
.C(n_1349),
.Y(n_3207)
);

NOR2xp33_ASAP7_75t_L g3208 ( 
.A(n_2705),
.B(n_290),
.Y(n_3208)
);

BUFx3_ASAP7_75t_L g3209 ( 
.A(n_2674),
.Y(n_3209)
);

INVx2_ASAP7_75t_SL g3210 ( 
.A(n_2674),
.Y(n_3210)
);

INVx1_ASAP7_75t_L g3211 ( 
.A(n_2722),
.Y(n_3211)
);

INVx2_ASAP7_75t_L g3212 ( 
.A(n_2720),
.Y(n_3212)
);

NAND2xp5_ASAP7_75t_SL g3213 ( 
.A(n_2446),
.B(n_1342),
.Y(n_3213)
);

AND2x2_ASAP7_75t_L g3214 ( 
.A(n_2711),
.B(n_290),
.Y(n_3214)
);

NOR3xp33_ASAP7_75t_L g3215 ( 
.A(n_2677),
.B(n_2711),
.C(n_2446),
.Y(n_3215)
);

INVx2_ASAP7_75t_L g3216 ( 
.A(n_2788),
.Y(n_3216)
);

INVx2_ASAP7_75t_L g3217 ( 
.A(n_2788),
.Y(n_3217)
);

NOR2xp33_ASAP7_75t_L g3218 ( 
.A(n_2795),
.B(n_291),
.Y(n_3218)
);

INVx2_ASAP7_75t_L g3219 ( 
.A(n_2795),
.Y(n_3219)
);

NAND2xp5_ASAP7_75t_L g3220 ( 
.A(n_2666),
.B(n_3),
.Y(n_3220)
);

NAND2xp5_ASAP7_75t_SL g3221 ( 
.A(n_2666),
.B(n_1342),
.Y(n_3221)
);

NAND2xp5_ASAP7_75t_L g3222 ( 
.A(n_2666),
.B(n_3),
.Y(n_3222)
);

AOI22xp33_ASAP7_75t_L g3223 ( 
.A1(n_2668),
.A2(n_1349),
.B1(n_1397),
.B2(n_1364),
.Y(n_3223)
);

INVx2_ASAP7_75t_L g3224 ( 
.A(n_2668),
.Y(n_3224)
);

INVx1_ASAP7_75t_L g3225 ( 
.A(n_2668),
.Y(n_3225)
);

INVx2_ASAP7_75t_SL g3226 ( 
.A(n_2759),
.Y(n_3226)
);

NOR2xp33_ASAP7_75t_L g3227 ( 
.A(n_2778),
.B(n_291),
.Y(n_3227)
);

OR2x2_ASAP7_75t_L g3228 ( 
.A(n_2778),
.B(n_291),
.Y(n_3228)
);

AOI22xp5_ASAP7_75t_L g3229 ( 
.A1(n_2778),
.A2(n_1710),
.B1(n_1342),
.B2(n_1364),
.Y(n_3229)
);

INVx2_ASAP7_75t_L g3230 ( 
.A(n_2538),
.Y(n_3230)
);

NAND2xp5_ASAP7_75t_L g3231 ( 
.A(n_2778),
.B(n_3),
.Y(n_3231)
);

INVx1_ASAP7_75t_L g3232 ( 
.A(n_2437),
.Y(n_3232)
);

NAND2xp33_ASAP7_75t_L g3233 ( 
.A(n_2418),
.B(n_1710),
.Y(n_3233)
);

AOI22xp33_ASAP7_75t_L g3234 ( 
.A1(n_2694),
.A2(n_1397),
.B1(n_1417),
.B2(n_1349),
.Y(n_3234)
);

INVx2_ASAP7_75t_L g3235 ( 
.A(n_2538),
.Y(n_3235)
);

A2O1A1Ixp33_ASAP7_75t_SL g3236 ( 
.A1(n_2754),
.A2(n_1397),
.B(n_1417),
.C(n_1349),
.Y(n_3236)
);

NOR2xp33_ASAP7_75t_L g3237 ( 
.A(n_2778),
.B(n_292),
.Y(n_3237)
);

NAND2xp5_ASAP7_75t_L g3238 ( 
.A(n_2778),
.B(n_4),
.Y(n_3238)
);

NOR3xp33_ASAP7_75t_L g3239 ( 
.A(n_2443),
.B(n_293),
.C(n_292),
.Y(n_3239)
);

NAND2xp5_ASAP7_75t_L g3240 ( 
.A(n_2778),
.B(n_4),
.Y(n_3240)
);

INVx1_ASAP7_75t_L g3241 ( 
.A(n_2437),
.Y(n_3241)
);

NAND2xp5_ASAP7_75t_L g3242 ( 
.A(n_2778),
.B(n_4),
.Y(n_3242)
);

NOR2xp33_ASAP7_75t_L g3243 ( 
.A(n_2778),
.B(n_292),
.Y(n_3243)
);

INVx2_ASAP7_75t_L g3244 ( 
.A(n_2538),
.Y(n_3244)
);

INVx1_ASAP7_75t_L g3245 ( 
.A(n_2437),
.Y(n_3245)
);

AND2x2_ASAP7_75t_L g3246 ( 
.A(n_2778),
.B(n_1105),
.Y(n_3246)
);

INVx2_ASAP7_75t_L g3247 ( 
.A(n_2538),
.Y(n_3247)
);

NAND2xp5_ASAP7_75t_SL g3248 ( 
.A(n_2778),
.B(n_1710),
.Y(n_3248)
);

INVx2_ASAP7_75t_L g3249 ( 
.A(n_2538),
.Y(n_3249)
);

INVx2_ASAP7_75t_SL g3250 ( 
.A(n_2759),
.Y(n_3250)
);

INVx2_ASAP7_75t_L g3251 ( 
.A(n_2538),
.Y(n_3251)
);

OAI22xp5_ASAP7_75t_L g3252 ( 
.A1(n_2522),
.A2(n_1417),
.B1(n_1419),
.B2(n_1397),
.Y(n_3252)
);

INVx3_ASAP7_75t_L g3253 ( 
.A(n_2431),
.Y(n_3253)
);

NAND2xp5_ASAP7_75t_L g3254 ( 
.A(n_2498),
.B(n_1710),
.Y(n_3254)
);

INVx1_ASAP7_75t_L g3255 ( 
.A(n_2437),
.Y(n_3255)
);

NAND2xp5_ASAP7_75t_L g3256 ( 
.A(n_2498),
.B(n_1417),
.Y(n_3256)
);

INVx1_ASAP7_75t_L g3257 ( 
.A(n_2437),
.Y(n_3257)
);

INVx1_ASAP7_75t_L g3258 ( 
.A(n_2437),
.Y(n_3258)
);

INVx2_ASAP7_75t_L g3259 ( 
.A(n_2538),
.Y(n_3259)
);

CKINVDCx11_ASAP7_75t_R g3260 ( 
.A(n_2520),
.Y(n_3260)
);

INVxp67_ASAP7_75t_L g3261 ( 
.A(n_2778),
.Y(n_3261)
);

AOI21x1_ASAP7_75t_L g3262 ( 
.A1(n_2420),
.A2(n_1507),
.B(n_1419),
.Y(n_3262)
);

AND2x2_ASAP7_75t_L g3263 ( 
.A(n_2778),
.B(n_1106),
.Y(n_3263)
);

INVx2_ASAP7_75t_L g3264 ( 
.A(n_2538),
.Y(n_3264)
);

NOR2xp67_ASAP7_75t_L g3265 ( 
.A(n_2412),
.B(n_293),
.Y(n_3265)
);

CKINVDCx5p33_ASAP7_75t_R g3266 ( 
.A(n_2520),
.Y(n_3266)
);

NAND2xp5_ASAP7_75t_L g3267 ( 
.A(n_2498),
.B(n_1419),
.Y(n_3267)
);

NAND2xp5_ASAP7_75t_L g3268 ( 
.A(n_2498),
.B(n_1419),
.Y(n_3268)
);

INVx3_ASAP7_75t_L g3269 ( 
.A(n_2431),
.Y(n_3269)
);

INVx1_ASAP7_75t_L g3270 ( 
.A(n_2437),
.Y(n_3270)
);

BUFx3_ASAP7_75t_L g3271 ( 
.A(n_2463),
.Y(n_3271)
);

NAND2xp5_ASAP7_75t_L g3272 ( 
.A(n_2498),
.B(n_1507),
.Y(n_3272)
);

INVx2_ASAP7_75t_L g3273 ( 
.A(n_2538),
.Y(n_3273)
);

INVx1_ASAP7_75t_L g3274 ( 
.A(n_2437),
.Y(n_3274)
);

INVx1_ASAP7_75t_L g3275 ( 
.A(n_2437),
.Y(n_3275)
);

INVxp33_ASAP7_75t_SL g3276 ( 
.A(n_2762),
.Y(n_3276)
);

O2A1O1Ixp5_ASAP7_75t_L g3277 ( 
.A1(n_2725),
.A2(n_1507),
.B(n_295),
.C(n_297),
.Y(n_3277)
);

NAND2xp5_ASAP7_75t_L g3278 ( 
.A(n_2498),
.B(n_1507),
.Y(n_3278)
);

INVx8_ASAP7_75t_L g3279 ( 
.A(n_2433),
.Y(n_3279)
);

INVx2_ASAP7_75t_L g3280 ( 
.A(n_2538),
.Y(n_3280)
);

NAND2xp5_ASAP7_75t_L g3281 ( 
.A(n_2498),
.B(n_5),
.Y(n_3281)
);

NOR3xp33_ASAP7_75t_L g3282 ( 
.A(n_2443),
.B(n_298),
.C(n_297),
.Y(n_3282)
);

NAND2xp5_ASAP7_75t_L g3283 ( 
.A(n_2498),
.B(n_5),
.Y(n_3283)
);

NAND2xp5_ASAP7_75t_L g3284 ( 
.A(n_2498),
.B(n_5),
.Y(n_3284)
);

AOI22xp33_ASAP7_75t_L g3285 ( 
.A1(n_2694),
.A2(n_7),
.B1(n_5),
.B2(n_6),
.Y(n_3285)
);

AOI22xp5_ASAP7_75t_L g3286 ( 
.A1(n_2778),
.A2(n_297),
.B1(n_298),
.B2(n_293),
.Y(n_3286)
);

INVx2_ASAP7_75t_L g3287 ( 
.A(n_2538),
.Y(n_3287)
);

AOI22xp5_ASAP7_75t_L g3288 ( 
.A1(n_2778),
.A2(n_299),
.B1(n_300),
.B2(n_298),
.Y(n_3288)
);

NAND2xp5_ASAP7_75t_L g3289 ( 
.A(n_2498),
.B(n_6),
.Y(n_3289)
);

NAND2xp5_ASAP7_75t_L g3290 ( 
.A(n_2498),
.B(n_6),
.Y(n_3290)
);

NOR2xp33_ASAP7_75t_L g3291 ( 
.A(n_2778),
.B(n_299),
.Y(n_3291)
);

INVxp67_ASAP7_75t_SL g3292 ( 
.A(n_2778),
.Y(n_3292)
);

NAND2xp5_ASAP7_75t_L g3293 ( 
.A(n_2498),
.B(n_7),
.Y(n_3293)
);

INVx1_ASAP7_75t_L g3294 ( 
.A(n_2437),
.Y(n_3294)
);

NAND2xp5_ASAP7_75t_L g3295 ( 
.A(n_2498),
.B(n_7),
.Y(n_3295)
);

NOR2xp33_ASAP7_75t_L g3296 ( 
.A(n_2778),
.B(n_299),
.Y(n_3296)
);

NAND2xp5_ASAP7_75t_L g3297 ( 
.A(n_2498),
.B(n_7),
.Y(n_3297)
);

NAND2xp5_ASAP7_75t_L g3298 ( 
.A(n_2498),
.B(n_8),
.Y(n_3298)
);

NAND2xp33_ASAP7_75t_L g3299 ( 
.A(n_2418),
.B(n_8),
.Y(n_3299)
);

INVx2_ASAP7_75t_L g3300 ( 
.A(n_2538),
.Y(n_3300)
);

NAND2xp5_ASAP7_75t_SL g3301 ( 
.A(n_2778),
.B(n_300),
.Y(n_3301)
);

NOR2x1p5_ASAP7_75t_SL g3302 ( 
.A(n_2420),
.B(n_8),
.Y(n_3302)
);

INVx2_ASAP7_75t_L g3303 ( 
.A(n_2538),
.Y(n_3303)
);

NAND2xp5_ASAP7_75t_SL g3304 ( 
.A(n_2778),
.B(n_300),
.Y(n_3304)
);

AOI22xp33_ASAP7_75t_L g3305 ( 
.A1(n_2694),
.A2(n_10),
.B1(n_8),
.B2(n_9),
.Y(n_3305)
);

INVx2_ASAP7_75t_SL g3306 ( 
.A(n_2759),
.Y(n_3306)
);

AND2x2_ASAP7_75t_L g3307 ( 
.A(n_2778),
.B(n_1099),
.Y(n_3307)
);

NOR2xp33_ASAP7_75t_L g3308 ( 
.A(n_2778),
.B(n_301),
.Y(n_3308)
);

NOR2xp33_ASAP7_75t_L g3309 ( 
.A(n_2778),
.B(n_301),
.Y(n_3309)
);

NAND2x1_ASAP7_75t_L g3310 ( 
.A(n_2707),
.B(n_9),
.Y(n_3310)
);

OAI22xp5_ASAP7_75t_L g3311 ( 
.A1(n_2522),
.A2(n_303),
.B1(n_304),
.B2(n_302),
.Y(n_3311)
);

NAND2xp5_ASAP7_75t_L g3312 ( 
.A(n_2498),
.B(n_9),
.Y(n_3312)
);

INVx1_ASAP7_75t_L g3313 ( 
.A(n_2437),
.Y(n_3313)
);

AND2x2_ASAP7_75t_L g3314 ( 
.A(n_2778),
.B(n_1102),
.Y(n_3314)
);

NOR2xp33_ASAP7_75t_L g3315 ( 
.A(n_2778),
.B(n_302),
.Y(n_3315)
);

O2A1O1Ixp33_ASAP7_75t_L g3316 ( 
.A1(n_2588),
.A2(n_304),
.B(n_305),
.C(n_302),
.Y(n_3316)
);

INVxp33_ASAP7_75t_L g3317 ( 
.A(n_2419),
.Y(n_3317)
);

AOI22xp33_ASAP7_75t_L g3318 ( 
.A1(n_2694),
.A2(n_12),
.B1(n_10),
.B2(n_11),
.Y(n_3318)
);

INVx2_ASAP7_75t_L g3319 ( 
.A(n_2538),
.Y(n_3319)
);

INVx1_ASAP7_75t_L g3320 ( 
.A(n_2437),
.Y(n_3320)
);

NAND2xp5_ASAP7_75t_L g3321 ( 
.A(n_2498),
.B(n_10),
.Y(n_3321)
);

NOR2xp33_ASAP7_75t_L g3322 ( 
.A(n_2778),
.B(n_304),
.Y(n_3322)
);

O2A1O1Ixp33_ASAP7_75t_L g3323 ( 
.A1(n_2588),
.A2(n_306),
.B(n_307),
.C(n_305),
.Y(n_3323)
);

INVx1_ASAP7_75t_L g3324 ( 
.A(n_2437),
.Y(n_3324)
);

AOI22xp33_ASAP7_75t_L g3325 ( 
.A1(n_2694),
.A2(n_12),
.B1(n_10),
.B2(n_11),
.Y(n_3325)
);

AND2x2_ASAP7_75t_L g3326 ( 
.A(n_2778),
.B(n_1107),
.Y(n_3326)
);

NAND2xp33_ASAP7_75t_L g3327 ( 
.A(n_2418),
.B(n_12),
.Y(n_3327)
);

NAND2xp5_ASAP7_75t_L g3328 ( 
.A(n_2498),
.B(n_13),
.Y(n_3328)
);

NAND2xp5_ASAP7_75t_L g3329 ( 
.A(n_2498),
.B(n_13),
.Y(n_3329)
);

AOI22xp5_ASAP7_75t_L g3330 ( 
.A1(n_2778),
.A2(n_306),
.B1(n_307),
.B2(n_305),
.Y(n_3330)
);

INVx8_ASAP7_75t_L g3331 ( 
.A(n_2433),
.Y(n_3331)
);

INVx2_ASAP7_75t_L g3332 ( 
.A(n_2538),
.Y(n_3332)
);

NAND2xp5_ASAP7_75t_L g3333 ( 
.A(n_2498),
.B(n_13),
.Y(n_3333)
);

INVx2_ASAP7_75t_L g3334 ( 
.A(n_2538),
.Y(n_3334)
);

NAND2xp5_ASAP7_75t_L g3335 ( 
.A(n_2498),
.B(n_13),
.Y(n_3335)
);

NAND2xp5_ASAP7_75t_L g3336 ( 
.A(n_2498),
.B(n_14),
.Y(n_3336)
);

INVx1_ASAP7_75t_L g3337 ( 
.A(n_2437),
.Y(n_3337)
);

NOR2xp33_ASAP7_75t_L g3338 ( 
.A(n_2778),
.B(n_306),
.Y(n_3338)
);

INVx1_ASAP7_75t_L g3339 ( 
.A(n_2437),
.Y(n_3339)
);

NOR2xp33_ASAP7_75t_L g3340 ( 
.A(n_2778),
.B(n_308),
.Y(n_3340)
);

NAND2xp5_ASAP7_75t_SL g3341 ( 
.A(n_2778),
.B(n_308),
.Y(n_3341)
);

NAND2xp5_ASAP7_75t_L g3342 ( 
.A(n_2498),
.B(n_14),
.Y(n_3342)
);

NOR2xp33_ASAP7_75t_L g3343 ( 
.A(n_2778),
.B(n_309),
.Y(n_3343)
);

AOI22xp5_ASAP7_75t_L g3344 ( 
.A1(n_2778),
.A2(n_310),
.B1(n_311),
.B2(n_309),
.Y(n_3344)
);

AND2x6_ASAP7_75t_L g3345 ( 
.A(n_2538),
.B(n_309),
.Y(n_3345)
);

NAND2xp5_ASAP7_75t_SL g3346 ( 
.A(n_2778),
.B(n_310),
.Y(n_3346)
);

NAND2xp5_ASAP7_75t_L g3347 ( 
.A(n_2498),
.B(n_14),
.Y(n_3347)
);

NOR2xp33_ASAP7_75t_L g3348 ( 
.A(n_2778),
.B(n_310),
.Y(n_3348)
);

NAND2xp5_ASAP7_75t_L g3349 ( 
.A(n_2498),
.B(n_14),
.Y(n_3349)
);

AND2x2_ASAP7_75t_L g3350 ( 
.A(n_2778),
.B(n_1099),
.Y(n_3350)
);

NAND2xp5_ASAP7_75t_L g3351 ( 
.A(n_2498),
.B(n_15),
.Y(n_3351)
);

NAND2xp5_ASAP7_75t_L g3352 ( 
.A(n_2498),
.B(n_15),
.Y(n_3352)
);

NOR2xp33_ASAP7_75t_L g3353 ( 
.A(n_2778),
.B(n_311),
.Y(n_3353)
);

INVx2_ASAP7_75t_L g3354 ( 
.A(n_2538),
.Y(n_3354)
);

INVx1_ASAP7_75t_L g3355 ( 
.A(n_2437),
.Y(n_3355)
);

NOR2x1p5_ASAP7_75t_L g3356 ( 
.A(n_2562),
.B(n_311),
.Y(n_3356)
);

NAND2xp5_ASAP7_75t_SL g3357 ( 
.A(n_2778),
.B(n_312),
.Y(n_3357)
);

INVx1_ASAP7_75t_SL g3358 ( 
.A(n_2778),
.Y(n_3358)
);

NAND2xp5_ASAP7_75t_SL g3359 ( 
.A(n_2778),
.B(n_313),
.Y(n_3359)
);

BUFx6f_ASAP7_75t_L g3360 ( 
.A(n_2459),
.Y(n_3360)
);

OAI22xp5_ASAP7_75t_L g3361 ( 
.A1(n_2522),
.A2(n_314),
.B1(n_315),
.B2(n_313),
.Y(n_3361)
);

INVx2_ASAP7_75t_L g3362 ( 
.A(n_2538),
.Y(n_3362)
);

NAND2xp5_ASAP7_75t_SL g3363 ( 
.A(n_2778),
.B(n_313),
.Y(n_3363)
);

INVx1_ASAP7_75t_L g3364 ( 
.A(n_2437),
.Y(n_3364)
);

INVx1_ASAP7_75t_L g3365 ( 
.A(n_2437),
.Y(n_3365)
);

NAND2xp5_ASAP7_75t_L g3366 ( 
.A(n_2498),
.B(n_15),
.Y(n_3366)
);

INVx1_ASAP7_75t_L g3367 ( 
.A(n_2437),
.Y(n_3367)
);

O2A1O1Ixp33_ASAP7_75t_L g3368 ( 
.A1(n_2588),
.A2(n_315),
.B(n_316),
.C(n_314),
.Y(n_3368)
);

NAND2xp5_ASAP7_75t_L g3369 ( 
.A(n_2498),
.B(n_16),
.Y(n_3369)
);

NOR2xp33_ASAP7_75t_L g3370 ( 
.A(n_2778),
.B(n_314),
.Y(n_3370)
);

AOI22xp5_ASAP7_75t_L g3371 ( 
.A1(n_2778),
.A2(n_317),
.B1(n_318),
.B2(n_316),
.Y(n_3371)
);

NOR2xp33_ASAP7_75t_L g3372 ( 
.A(n_2778),
.B(n_316),
.Y(n_3372)
);

INVx2_ASAP7_75t_L g3373 ( 
.A(n_2538),
.Y(n_3373)
);

NAND2xp5_ASAP7_75t_SL g3374 ( 
.A(n_2778),
.B(n_317),
.Y(n_3374)
);

INVxp67_ASAP7_75t_L g3375 ( 
.A(n_2778),
.Y(n_3375)
);

BUFx6f_ASAP7_75t_L g3376 ( 
.A(n_2459),
.Y(n_3376)
);

BUFx3_ASAP7_75t_L g3377 ( 
.A(n_2463),
.Y(n_3377)
);

NAND2xp5_ASAP7_75t_L g3378 ( 
.A(n_2498),
.B(n_16),
.Y(n_3378)
);

NAND2xp5_ASAP7_75t_L g3379 ( 
.A(n_2498),
.B(n_16),
.Y(n_3379)
);

NAND2xp5_ASAP7_75t_L g3380 ( 
.A(n_2498),
.B(n_17),
.Y(n_3380)
);

BUFx3_ASAP7_75t_L g3381 ( 
.A(n_2463),
.Y(n_3381)
);

BUFx12f_ASAP7_75t_L g3382 ( 
.A(n_2520),
.Y(n_3382)
);

AOI22xp33_ASAP7_75t_L g3383 ( 
.A1(n_2694),
.A2(n_19),
.B1(n_17),
.B2(n_18),
.Y(n_3383)
);

NAND2xp5_ASAP7_75t_SL g3384 ( 
.A(n_2778),
.B(n_317),
.Y(n_3384)
);

OR2x2_ASAP7_75t_L g3385 ( 
.A(n_2778),
.B(n_318),
.Y(n_3385)
);

INVx1_ASAP7_75t_L g3386 ( 
.A(n_2437),
.Y(n_3386)
);

NAND2xp5_ASAP7_75t_SL g3387 ( 
.A(n_2778),
.B(n_319),
.Y(n_3387)
);

NAND2xp5_ASAP7_75t_SL g3388 ( 
.A(n_2778),
.B(n_319),
.Y(n_3388)
);

NOR2xp33_ASAP7_75t_L g3389 ( 
.A(n_2778),
.B(n_319),
.Y(n_3389)
);

AOI22xp33_ASAP7_75t_L g3390 ( 
.A1(n_2694),
.A2(n_19),
.B1(n_17),
.B2(n_18),
.Y(n_3390)
);

NAND2xp5_ASAP7_75t_L g3391 ( 
.A(n_2498),
.B(n_17),
.Y(n_3391)
);

NAND2xp5_ASAP7_75t_L g3392 ( 
.A(n_2498),
.B(n_18),
.Y(n_3392)
);

NAND2xp5_ASAP7_75t_L g3393 ( 
.A(n_2498),
.B(n_18),
.Y(n_3393)
);

NOR2xp33_ASAP7_75t_L g3394 ( 
.A(n_2778),
.B(n_320),
.Y(n_3394)
);

INVxp33_ASAP7_75t_L g3395 ( 
.A(n_2419),
.Y(n_3395)
);

INVx1_ASAP7_75t_L g3396 ( 
.A(n_2437),
.Y(n_3396)
);

INVx2_ASAP7_75t_L g3397 ( 
.A(n_2538),
.Y(n_3397)
);

INVxp67_ASAP7_75t_L g3398 ( 
.A(n_2778),
.Y(n_3398)
);

INVx1_ASAP7_75t_L g3399 ( 
.A(n_2437),
.Y(n_3399)
);

INVx2_ASAP7_75t_SL g3400 ( 
.A(n_2759),
.Y(n_3400)
);

NAND2xp5_ASAP7_75t_SL g3401 ( 
.A(n_2778),
.B(n_320),
.Y(n_3401)
);

NAND2xp5_ASAP7_75t_L g3402 ( 
.A(n_2498),
.B(n_19),
.Y(n_3402)
);

NAND2xp5_ASAP7_75t_L g3403 ( 
.A(n_2498),
.B(n_19),
.Y(n_3403)
);

NAND2xp33_ASAP7_75t_L g3404 ( 
.A(n_2418),
.B(n_20),
.Y(n_3404)
);

NAND2xp5_ASAP7_75t_L g3405 ( 
.A(n_2498),
.B(n_20),
.Y(n_3405)
);

NOR2xp33_ASAP7_75t_L g3406 ( 
.A(n_2778),
.B(n_320),
.Y(n_3406)
);

OR2x2_ASAP7_75t_L g3407 ( 
.A(n_2778),
.B(n_321),
.Y(n_3407)
);

INVx1_ASAP7_75t_L g3408 ( 
.A(n_2437),
.Y(n_3408)
);

INVx2_ASAP7_75t_SL g3409 ( 
.A(n_2759),
.Y(n_3409)
);

INVx1_ASAP7_75t_L g3410 ( 
.A(n_2437),
.Y(n_3410)
);

NAND2xp5_ASAP7_75t_SL g3411 ( 
.A(n_2778),
.B(n_321),
.Y(n_3411)
);

AND2x2_ASAP7_75t_L g3412 ( 
.A(n_2778),
.B(n_1098),
.Y(n_3412)
);

INVx2_ASAP7_75t_SL g3413 ( 
.A(n_2759),
.Y(n_3413)
);

BUFx6f_ASAP7_75t_L g3414 ( 
.A(n_2459),
.Y(n_3414)
);

BUFx3_ASAP7_75t_L g3415 ( 
.A(n_2463),
.Y(n_3415)
);

BUFx6f_ASAP7_75t_SL g3416 ( 
.A(n_2527),
.Y(n_3416)
);

INVx3_ASAP7_75t_L g3417 ( 
.A(n_2431),
.Y(n_3417)
);

INVx1_ASAP7_75t_L g3418 ( 
.A(n_2437),
.Y(n_3418)
);

NOR2xp33_ASAP7_75t_L g3419 ( 
.A(n_2778),
.B(n_321),
.Y(n_3419)
);

AOI22xp33_ASAP7_75t_L g3420 ( 
.A1(n_2694),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.Y(n_3420)
);

NAND2xp5_ASAP7_75t_L g3421 ( 
.A(n_2498),
.B(n_20),
.Y(n_3421)
);

NAND2xp5_ASAP7_75t_SL g3422 ( 
.A(n_2778),
.B(n_323),
.Y(n_3422)
);

NOR3xp33_ASAP7_75t_L g3423 ( 
.A(n_2443),
.B(n_324),
.C(n_323),
.Y(n_3423)
);

NAND2xp5_ASAP7_75t_L g3424 ( 
.A(n_2498),
.B(n_21),
.Y(n_3424)
);

NAND2xp5_ASAP7_75t_L g3425 ( 
.A(n_2498),
.B(n_21),
.Y(n_3425)
);

O2A1O1Ixp33_ASAP7_75t_L g3426 ( 
.A1(n_2588),
.A2(n_323),
.B(n_324),
.C(n_322),
.Y(n_3426)
);

AOI22xp33_ASAP7_75t_L g3427 ( 
.A1(n_2694),
.A2(n_23),
.B1(n_21),
.B2(n_22),
.Y(n_3427)
);

NAND2xp5_ASAP7_75t_SL g3428 ( 
.A(n_2778),
.B(n_322),
.Y(n_3428)
);

NAND2xp5_ASAP7_75t_L g3429 ( 
.A(n_2498),
.B(n_22),
.Y(n_3429)
);

INVx2_ASAP7_75t_L g3430 ( 
.A(n_2538),
.Y(n_3430)
);

NAND2xp5_ASAP7_75t_L g3431 ( 
.A(n_2498),
.B(n_23),
.Y(n_3431)
);

NAND3xp33_ASAP7_75t_L g3432 ( 
.A(n_2575),
.B(n_325),
.C(n_322),
.Y(n_3432)
);

INVx2_ASAP7_75t_SL g3433 ( 
.A(n_2759),
.Y(n_3433)
);

A2O1A1Ixp33_ASAP7_75t_L g3434 ( 
.A1(n_2588),
.A2(n_326),
.B(n_327),
.C(n_325),
.Y(n_3434)
);

NAND2xp5_ASAP7_75t_L g3435 ( 
.A(n_2498),
.B(n_23),
.Y(n_3435)
);

AND2x4_ASAP7_75t_L g3436 ( 
.A(n_2778),
.B(n_325),
.Y(n_3436)
);

INVx1_ASAP7_75t_L g3437 ( 
.A(n_2437),
.Y(n_3437)
);

NAND2xp5_ASAP7_75t_L g3438 ( 
.A(n_2498),
.B(n_23),
.Y(n_3438)
);

INVx2_ASAP7_75t_L g3439 ( 
.A(n_2538),
.Y(n_3439)
);

INVx1_ASAP7_75t_SL g3440 ( 
.A(n_2778),
.Y(n_3440)
);

NAND2xp5_ASAP7_75t_L g3441 ( 
.A(n_2498),
.B(n_24),
.Y(n_3441)
);

INVx1_ASAP7_75t_L g3442 ( 
.A(n_2437),
.Y(n_3442)
);

OR2x2_ASAP7_75t_L g3443 ( 
.A(n_2778),
.B(n_326),
.Y(n_3443)
);

INVx1_ASAP7_75t_L g3444 ( 
.A(n_2437),
.Y(n_3444)
);

INVx1_ASAP7_75t_L g3445 ( 
.A(n_2437),
.Y(n_3445)
);

OAI22xp33_ASAP7_75t_L g3446 ( 
.A1(n_2762),
.A2(n_328),
.B1(n_329),
.B2(n_326),
.Y(n_3446)
);

NAND2xp5_ASAP7_75t_L g3447 ( 
.A(n_2498),
.B(n_24),
.Y(n_3447)
);

NAND2xp5_ASAP7_75t_L g3448 ( 
.A(n_2498),
.B(n_24),
.Y(n_3448)
);

NAND2xp5_ASAP7_75t_SL g3449 ( 
.A(n_2778),
.B(n_328),
.Y(n_3449)
);

INVx3_ASAP7_75t_L g3450 ( 
.A(n_2431),
.Y(n_3450)
);

AOI22xp5_ASAP7_75t_L g3451 ( 
.A1(n_2778),
.A2(n_329),
.B1(n_330),
.B2(n_328),
.Y(n_3451)
);

INVx2_ASAP7_75t_L g3452 ( 
.A(n_2538),
.Y(n_3452)
);

NAND2xp5_ASAP7_75t_SL g3453 ( 
.A(n_2778),
.B(n_329),
.Y(n_3453)
);

NAND2xp5_ASAP7_75t_SL g3454 ( 
.A(n_2778),
.B(n_330),
.Y(n_3454)
);

O2A1O1Ixp33_ASAP7_75t_L g3455 ( 
.A1(n_2588),
.A2(n_332),
.B(n_333),
.C(n_331),
.Y(n_3455)
);

INVxp67_ASAP7_75t_SL g3456 ( 
.A(n_2778),
.Y(n_3456)
);

A2O1A1Ixp33_ASAP7_75t_L g3457 ( 
.A1(n_2964),
.A2(n_26),
.B(n_24),
.C(n_25),
.Y(n_3457)
);

NOR2xp33_ASAP7_75t_L g3458 ( 
.A(n_3317),
.B(n_331),
.Y(n_3458)
);

O2A1O1Ixp33_ASAP7_75t_SL g3459 ( 
.A1(n_3252),
.A2(n_2868),
.B(n_3248),
.C(n_3127),
.Y(n_3459)
);

NAND2xp5_ASAP7_75t_L g3460 ( 
.A(n_2830),
.B(n_331),
.Y(n_3460)
);

NAND2xp5_ASAP7_75t_L g3461 ( 
.A(n_2897),
.B(n_332),
.Y(n_3461)
);

NAND2xp5_ASAP7_75t_L g3462 ( 
.A(n_2970),
.B(n_333),
.Y(n_3462)
);

CKINVDCx10_ASAP7_75t_R g3463 ( 
.A(n_2929),
.Y(n_3463)
);

NAND2xp5_ASAP7_75t_L g3464 ( 
.A(n_2801),
.B(n_333),
.Y(n_3464)
);

BUFx6f_ASAP7_75t_L g3465 ( 
.A(n_2927),
.Y(n_3465)
);

NAND2xp5_ASAP7_75t_L g3466 ( 
.A(n_2837),
.B(n_2834),
.Y(n_3466)
);

NAND2xp5_ASAP7_75t_SL g3467 ( 
.A(n_2859),
.B(n_2862),
.Y(n_3467)
);

AOI21xp5_ASAP7_75t_L g3468 ( 
.A1(n_3233),
.A2(n_335),
.B(n_334),
.Y(n_3468)
);

AOI21xp5_ASAP7_75t_L g3469 ( 
.A1(n_3097),
.A2(n_335),
.B(n_334),
.Y(n_3469)
);

A2O1A1Ixp33_ASAP7_75t_L g3470 ( 
.A1(n_2900),
.A2(n_27),
.B(n_25),
.C(n_26),
.Y(n_3470)
);

AOI21xp5_ASAP7_75t_L g3471 ( 
.A1(n_3097),
.A2(n_336),
.B(n_334),
.Y(n_3471)
);

NAND2xp5_ASAP7_75t_L g3472 ( 
.A(n_3004),
.B(n_336),
.Y(n_3472)
);

OAI321xp33_ASAP7_75t_L g3473 ( 
.A1(n_3252),
.A2(n_28),
.A3(n_30),
.B1(n_26),
.B2(n_27),
.C(n_29),
.Y(n_3473)
);

INVx2_ASAP7_75t_L g3474 ( 
.A(n_2822),
.Y(n_3474)
);

INVx1_ASAP7_75t_L g3475 ( 
.A(n_2806),
.Y(n_3475)
);

AOI21xp5_ASAP7_75t_L g3476 ( 
.A1(n_3004),
.A2(n_338),
.B(n_337),
.Y(n_3476)
);

A2O1A1Ixp33_ASAP7_75t_L g3477 ( 
.A1(n_3299),
.A2(n_29),
.B(n_26),
.C(n_28),
.Y(n_3477)
);

AOI21xp5_ASAP7_75t_L g3478 ( 
.A1(n_3029),
.A2(n_338),
.B(n_337),
.Y(n_3478)
);

AOI21xp5_ASAP7_75t_L g3479 ( 
.A1(n_3084),
.A2(n_338),
.B(n_337),
.Y(n_3479)
);

INVx2_ASAP7_75t_L g3480 ( 
.A(n_2823),
.Y(n_3480)
);

HB1xp67_ASAP7_75t_L g3481 ( 
.A(n_3358),
.Y(n_3481)
);

AOI22xp5_ASAP7_75t_L g3482 ( 
.A1(n_2831),
.A2(n_2972),
.B1(n_2827),
.B2(n_2899),
.Y(n_3482)
);

AND2x4_ASAP7_75t_L g3483 ( 
.A(n_2903),
.B(n_339),
.Y(n_3483)
);

NAND2xp5_ASAP7_75t_L g3484 ( 
.A(n_2871),
.B(n_339),
.Y(n_3484)
);

INVx1_ASAP7_75t_L g3485 ( 
.A(n_2884),
.Y(n_3485)
);

AOI21xp5_ASAP7_75t_L g3486 ( 
.A1(n_3092),
.A2(n_341),
.B(n_340),
.Y(n_3486)
);

OAI21xp33_ASAP7_75t_L g3487 ( 
.A1(n_3038),
.A2(n_28),
.B(n_29),
.Y(n_3487)
);

NAND2xp5_ASAP7_75t_SL g3488 ( 
.A(n_2944),
.B(n_340),
.Y(n_3488)
);

AOI21x1_ASAP7_75t_L g3489 ( 
.A1(n_3262),
.A2(n_342),
.B(n_341),
.Y(n_3489)
);

AOI21xp5_ASAP7_75t_L g3490 ( 
.A1(n_3094),
.A2(n_342),
.B(n_341),
.Y(n_3490)
);

NAND2xp5_ASAP7_75t_SL g3491 ( 
.A(n_2917),
.B(n_342),
.Y(n_3491)
);

BUFx6f_ASAP7_75t_L g3492 ( 
.A(n_2927),
.Y(n_3492)
);

AOI21xp5_ASAP7_75t_L g3493 ( 
.A1(n_3099),
.A2(n_344),
.B(n_343),
.Y(n_3493)
);

AOI22xp33_ASAP7_75t_L g3494 ( 
.A1(n_2857),
.A2(n_344),
.B1(n_345),
.B2(n_343),
.Y(n_3494)
);

NAND2xp33_ASAP7_75t_L g3495 ( 
.A(n_3279),
.B(n_3331),
.Y(n_3495)
);

BUFx8_ASAP7_75t_SL g3496 ( 
.A(n_3382),
.Y(n_3496)
);

NAND2xp5_ASAP7_75t_SL g3497 ( 
.A(n_3440),
.B(n_343),
.Y(n_3497)
);

NAND2xp5_ASAP7_75t_L g3498 ( 
.A(n_2871),
.B(n_344),
.Y(n_3498)
);

AND2x4_ASAP7_75t_L g3499 ( 
.A(n_2826),
.B(n_345),
.Y(n_3499)
);

OAI21xp5_ASAP7_75t_L g3500 ( 
.A1(n_2887),
.A2(n_2885),
.B(n_2992),
.Y(n_3500)
);

OAI21xp33_ASAP7_75t_L g3501 ( 
.A1(n_2868),
.A2(n_28),
.B(n_30),
.Y(n_3501)
);

AOI21xp5_ASAP7_75t_L g3502 ( 
.A1(n_3103),
.A2(n_3404),
.B(n_3327),
.Y(n_3502)
);

BUFx6f_ASAP7_75t_L g3503 ( 
.A(n_2927),
.Y(n_3503)
);

INVx1_ASAP7_75t_L g3504 ( 
.A(n_3232),
.Y(n_3504)
);

OAI22xp5_ASAP7_75t_L g3505 ( 
.A1(n_2843),
.A2(n_347),
.B1(n_348),
.B2(n_346),
.Y(n_3505)
);

NAND2xp5_ASAP7_75t_L g3506 ( 
.A(n_3241),
.B(n_346),
.Y(n_3506)
);

INVx2_ASAP7_75t_L g3507 ( 
.A(n_2879),
.Y(n_3507)
);

OR2x2_ASAP7_75t_L g3508 ( 
.A(n_3054),
.B(n_3130),
.Y(n_3508)
);

NAND2xp5_ASAP7_75t_L g3509 ( 
.A(n_3245),
.B(n_346),
.Y(n_3509)
);

NAND2xp5_ASAP7_75t_L g3510 ( 
.A(n_3255),
.B(n_347),
.Y(n_3510)
);

AND2x2_ASAP7_75t_L g3511 ( 
.A(n_2913),
.B(n_347),
.Y(n_3511)
);

NAND2xp5_ASAP7_75t_L g3512 ( 
.A(n_3257),
.B(n_348),
.Y(n_3512)
);

OAI21xp33_ASAP7_75t_L g3513 ( 
.A1(n_2880),
.A2(n_30),
.B(n_31),
.Y(n_3513)
);

AOI21xp5_ASAP7_75t_L g3514 ( 
.A1(n_3062),
.A2(n_349),
.B(n_348),
.Y(n_3514)
);

INVx2_ASAP7_75t_L g3515 ( 
.A(n_2940),
.Y(n_3515)
);

AND2x2_ASAP7_75t_L g3516 ( 
.A(n_2848),
.B(n_349),
.Y(n_3516)
);

NAND2xp5_ASAP7_75t_SL g3517 ( 
.A(n_3022),
.B(n_349),
.Y(n_3517)
);

NAND2xp5_ASAP7_75t_L g3518 ( 
.A(n_3258),
.B(n_350),
.Y(n_3518)
);

AOI21xp5_ASAP7_75t_L g3519 ( 
.A1(n_3254),
.A2(n_351),
.B(n_350),
.Y(n_3519)
);

NAND2xp5_ASAP7_75t_L g3520 ( 
.A(n_3270),
.B(n_351),
.Y(n_3520)
);

BUFx6f_ASAP7_75t_L g3521 ( 
.A(n_2986),
.Y(n_3521)
);

A2O1A1Ixp33_ASAP7_75t_L g3522 ( 
.A1(n_3316),
.A2(n_33),
.B(n_31),
.C(n_32),
.Y(n_3522)
);

NAND2xp5_ASAP7_75t_L g3523 ( 
.A(n_3274),
.B(n_352),
.Y(n_3523)
);

AOI21xp5_ASAP7_75t_L g3524 ( 
.A1(n_3254),
.A2(n_353),
.B(n_352),
.Y(n_3524)
);

OAI22xp5_ASAP7_75t_L g3525 ( 
.A1(n_2843),
.A2(n_354),
.B1(n_355),
.B2(n_353),
.Y(n_3525)
);

INVx2_ASAP7_75t_L g3526 ( 
.A(n_2958),
.Y(n_3526)
);

BUFx6f_ASAP7_75t_L g3527 ( 
.A(n_2986),
.Y(n_3527)
);

A2O1A1Ixp33_ASAP7_75t_L g3528 ( 
.A1(n_3323),
.A2(n_34),
.B(n_32),
.C(n_33),
.Y(n_3528)
);

AOI21xp5_ASAP7_75t_L g3529 ( 
.A1(n_3256),
.A2(n_355),
.B(n_354),
.Y(n_3529)
);

INVx4_ASAP7_75t_L g3530 ( 
.A(n_3279),
.Y(n_3530)
);

AOI21xp5_ASAP7_75t_L g3531 ( 
.A1(n_3256),
.A2(n_356),
.B(n_355),
.Y(n_3531)
);

AND2x2_ASAP7_75t_L g3532 ( 
.A(n_3292),
.B(n_356),
.Y(n_3532)
);

NAND2xp5_ASAP7_75t_SL g3533 ( 
.A(n_3276),
.B(n_357),
.Y(n_3533)
);

AOI21xp5_ASAP7_75t_L g3534 ( 
.A1(n_3267),
.A2(n_358),
.B(n_357),
.Y(n_3534)
);

BUFx2_ASAP7_75t_L g3535 ( 
.A(n_3261),
.Y(n_3535)
);

NAND2xp5_ASAP7_75t_L g3536 ( 
.A(n_3275),
.B(n_358),
.Y(n_3536)
);

INVxp67_ASAP7_75t_L g3537 ( 
.A(n_3456),
.Y(n_3537)
);

OAI21xp5_ASAP7_75t_L g3538 ( 
.A1(n_2887),
.A2(n_32),
.B(n_33),
.Y(n_3538)
);

NAND2xp5_ASAP7_75t_SL g3539 ( 
.A(n_2997),
.B(n_359),
.Y(n_3539)
);

OAI22xp5_ASAP7_75t_L g3540 ( 
.A1(n_2843),
.A2(n_360),
.B1(n_361),
.B2(n_359),
.Y(n_3540)
);

OAI22xp5_ASAP7_75t_L g3541 ( 
.A1(n_2839),
.A2(n_361),
.B1(n_362),
.B2(n_360),
.Y(n_3541)
);

INVx2_ASAP7_75t_L g3542 ( 
.A(n_2966),
.Y(n_3542)
);

OR2x2_ASAP7_75t_L g3543 ( 
.A(n_2812),
.B(n_3375),
.Y(n_3543)
);

INVx1_ASAP7_75t_L g3544 ( 
.A(n_3294),
.Y(n_3544)
);

AOI21xp5_ASAP7_75t_L g3545 ( 
.A1(n_3267),
.A2(n_3272),
.B(n_3268),
.Y(n_3545)
);

NOR2xp33_ASAP7_75t_L g3546 ( 
.A(n_3395),
.B(n_360),
.Y(n_3546)
);

NOR2xp33_ASAP7_75t_L g3547 ( 
.A(n_3067),
.B(n_361),
.Y(n_3547)
);

AND2x2_ASAP7_75t_L g3548 ( 
.A(n_2922),
.B(n_362),
.Y(n_3548)
);

NAND2xp5_ASAP7_75t_L g3549 ( 
.A(n_3313),
.B(n_362),
.Y(n_3549)
);

INVx2_ASAP7_75t_L g3550 ( 
.A(n_2968),
.Y(n_3550)
);

INVxp67_ASAP7_75t_L g3551 ( 
.A(n_3075),
.Y(n_3551)
);

NAND2xp5_ASAP7_75t_L g3552 ( 
.A(n_3320),
.B(n_363),
.Y(n_3552)
);

AOI21xp5_ASAP7_75t_L g3553 ( 
.A1(n_3268),
.A2(n_364),
.B(n_363),
.Y(n_3553)
);

NAND2xp5_ASAP7_75t_L g3554 ( 
.A(n_3324),
.B(n_364),
.Y(n_3554)
);

INVx1_ASAP7_75t_SL g3555 ( 
.A(n_3075),
.Y(n_3555)
);

NAND2xp5_ASAP7_75t_L g3556 ( 
.A(n_3337),
.B(n_364),
.Y(n_3556)
);

NOR2xp33_ASAP7_75t_L g3557 ( 
.A(n_2846),
.B(n_365),
.Y(n_3557)
);

INVxp67_ASAP7_75t_L g3558 ( 
.A(n_3075),
.Y(n_3558)
);

AO21x1_ASAP7_75t_L g3559 ( 
.A1(n_3311),
.A2(n_366),
.B(n_365),
.Y(n_3559)
);

AO21x1_ASAP7_75t_L g3560 ( 
.A1(n_3311),
.A2(n_366),
.B(n_365),
.Y(n_3560)
);

AND2x2_ASAP7_75t_SL g3561 ( 
.A(n_2803),
.B(n_366),
.Y(n_3561)
);

OAI21xp5_ASAP7_75t_L g3562 ( 
.A1(n_2885),
.A2(n_32),
.B(n_33),
.Y(n_3562)
);

O2A1O1Ixp33_ASAP7_75t_L g3563 ( 
.A1(n_3434),
.A2(n_368),
.B(n_370),
.C(n_367),
.Y(n_3563)
);

INVx2_ASAP7_75t_L g3564 ( 
.A(n_2979),
.Y(n_3564)
);

OAI22xp5_ASAP7_75t_L g3565 ( 
.A1(n_2839),
.A2(n_368),
.B1(n_370),
.B2(n_367),
.Y(n_3565)
);

NAND2xp5_ASAP7_75t_L g3566 ( 
.A(n_3339),
.B(n_367),
.Y(n_3566)
);

INVx2_ASAP7_75t_SL g3567 ( 
.A(n_3124),
.Y(n_3567)
);

INVx2_ASAP7_75t_L g3568 ( 
.A(n_2800),
.Y(n_3568)
);

NOR2xp33_ASAP7_75t_SL g3569 ( 
.A(n_2982),
.B(n_368),
.Y(n_3569)
);

INVx1_ASAP7_75t_L g3570 ( 
.A(n_3355),
.Y(n_3570)
);

O2A1O1Ixp33_ASAP7_75t_L g3571 ( 
.A1(n_2847),
.A2(n_372),
.B(n_373),
.C(n_371),
.Y(n_3571)
);

NAND2xp5_ASAP7_75t_L g3572 ( 
.A(n_3364),
.B(n_371),
.Y(n_3572)
);

OAI21xp5_ASAP7_75t_L g3573 ( 
.A1(n_2992),
.A2(n_34),
.B(n_35),
.Y(n_3573)
);

NOR2xp33_ASAP7_75t_SL g3574 ( 
.A(n_2888),
.B(n_371),
.Y(n_3574)
);

INVx4_ASAP7_75t_L g3575 ( 
.A(n_3279),
.Y(n_3575)
);

INVx1_ASAP7_75t_L g3576 ( 
.A(n_3365),
.Y(n_3576)
);

AOI22xp5_ASAP7_75t_L g3577 ( 
.A1(n_2878),
.A2(n_373),
.B1(n_374),
.B2(n_372),
.Y(n_3577)
);

HB1xp67_ASAP7_75t_L g3578 ( 
.A(n_3398),
.Y(n_3578)
);

NAND2xp5_ASAP7_75t_L g3579 ( 
.A(n_3367),
.B(n_372),
.Y(n_3579)
);

NAND2xp5_ASAP7_75t_L g3580 ( 
.A(n_3386),
.B(n_373),
.Y(n_3580)
);

BUFx6f_ASAP7_75t_L g3581 ( 
.A(n_2986),
.Y(n_3581)
);

INVx1_ASAP7_75t_L g3582 ( 
.A(n_3396),
.Y(n_3582)
);

NAND2xp5_ASAP7_75t_SL g3583 ( 
.A(n_2821),
.B(n_374),
.Y(n_3583)
);

AOI21x1_ASAP7_75t_L g3584 ( 
.A1(n_3272),
.A2(n_375),
.B(n_374),
.Y(n_3584)
);

AOI21xp5_ASAP7_75t_L g3585 ( 
.A1(n_3278),
.A2(n_377),
.B(n_376),
.Y(n_3585)
);

INVx2_ASAP7_75t_L g3586 ( 
.A(n_2809),
.Y(n_3586)
);

AOI22xp5_ASAP7_75t_L g3587 ( 
.A1(n_2849),
.A2(n_378),
.B1(n_379),
.B2(n_376),
.Y(n_3587)
);

NOR2xp67_ASAP7_75t_L g3588 ( 
.A(n_3015),
.B(n_376),
.Y(n_3588)
);

NAND2xp5_ASAP7_75t_L g3589 ( 
.A(n_3399),
.B(n_379),
.Y(n_3589)
);

AND2x2_ASAP7_75t_L g3590 ( 
.A(n_2925),
.B(n_379),
.Y(n_3590)
);

OAI21xp5_ASAP7_75t_L g3591 ( 
.A1(n_2995),
.A2(n_35),
.B(n_36),
.Y(n_3591)
);

INVx2_ASAP7_75t_SL g3592 ( 
.A(n_3124),
.Y(n_3592)
);

AOI21xp5_ASAP7_75t_L g3593 ( 
.A1(n_3278),
.A2(n_381),
.B(n_380),
.Y(n_3593)
);

AOI21xp5_ASAP7_75t_L g3594 ( 
.A1(n_3078),
.A2(n_381),
.B(n_380),
.Y(n_3594)
);

NAND2xp5_ASAP7_75t_L g3595 ( 
.A(n_3408),
.B(n_381),
.Y(n_3595)
);

NAND2xp5_ASAP7_75t_L g3596 ( 
.A(n_3410),
.B(n_382),
.Y(n_3596)
);

BUFx2_ASAP7_75t_L g3597 ( 
.A(n_3102),
.Y(n_3597)
);

O2A1O1Ixp33_ASAP7_75t_L g3598 ( 
.A1(n_3455),
.A2(n_383),
.B(n_384),
.C(n_382),
.Y(n_3598)
);

AOI21xp5_ASAP7_75t_L g3599 ( 
.A1(n_3187),
.A2(n_3077),
.B(n_2807),
.Y(n_3599)
);

AND2x4_ASAP7_75t_L g3600 ( 
.A(n_3073),
.B(n_384),
.Y(n_3600)
);

INVx1_ASAP7_75t_L g3601 ( 
.A(n_3418),
.Y(n_3601)
);

NAND2xp5_ASAP7_75t_L g3602 ( 
.A(n_3437),
.B(n_384),
.Y(n_3602)
);

NAND2xp5_ASAP7_75t_L g3603 ( 
.A(n_3442),
.B(n_3444),
.Y(n_3603)
);

BUFx2_ASAP7_75t_L g3604 ( 
.A(n_3102),
.Y(n_3604)
);

AO21x1_ASAP7_75t_L g3605 ( 
.A1(n_3361),
.A2(n_386),
.B(n_385),
.Y(n_3605)
);

INVx1_ASAP7_75t_L g3606 ( 
.A(n_3445),
.Y(n_3606)
);

INVx1_ASAP7_75t_L g3607 ( 
.A(n_3030),
.Y(n_3607)
);

INVx4_ASAP7_75t_L g3608 ( 
.A(n_3331),
.Y(n_3608)
);

INVx3_ASAP7_75t_L g3609 ( 
.A(n_2815),
.Y(n_3609)
);

HB1xp67_ASAP7_75t_L g3610 ( 
.A(n_3071),
.Y(n_3610)
);

AO21x1_ASAP7_75t_L g3611 ( 
.A1(n_3361),
.A2(n_387),
.B(n_386),
.Y(n_3611)
);

INVx2_ASAP7_75t_L g3612 ( 
.A(n_2813),
.Y(n_3612)
);

BUFx4f_ASAP7_75t_L g3613 ( 
.A(n_3331),
.Y(n_3613)
);

NAND3xp33_ASAP7_75t_SL g3614 ( 
.A(n_3266),
.B(n_35),
.C(n_36),
.Y(n_3614)
);

A2O1A1Ixp33_ASAP7_75t_L g3615 ( 
.A1(n_3368),
.A2(n_3426),
.B(n_3302),
.C(n_3007),
.Y(n_3615)
);

INVx1_ASAP7_75t_L g3616 ( 
.A(n_3061),
.Y(n_3616)
);

BUFx3_ASAP7_75t_L g3617 ( 
.A(n_3041),
.Y(n_3617)
);

NAND2xp5_ASAP7_75t_L g3618 ( 
.A(n_2808),
.B(n_386),
.Y(n_3618)
);

INVx2_ASAP7_75t_L g3619 ( 
.A(n_2817),
.Y(n_3619)
);

BUFx6f_ASAP7_75t_L g3620 ( 
.A(n_2999),
.Y(n_3620)
);

AOI21xp5_ASAP7_75t_L g3621 ( 
.A1(n_2805),
.A2(n_388),
.B(n_387),
.Y(n_3621)
);

NAND2xp5_ASAP7_75t_L g3622 ( 
.A(n_2814),
.B(n_388),
.Y(n_3622)
);

NAND2xp5_ASAP7_75t_L g3623 ( 
.A(n_2824),
.B(n_389),
.Y(n_3623)
);

NAND2xp5_ASAP7_75t_SL g3624 ( 
.A(n_3024),
.B(n_389),
.Y(n_3624)
);

AOI21x1_ASAP7_75t_L g3625 ( 
.A1(n_3216),
.A2(n_390),
.B(n_389),
.Y(n_3625)
);

A2O1A1Ixp33_ASAP7_75t_L g3626 ( 
.A1(n_2825),
.A2(n_38),
.B(n_36),
.C(n_37),
.Y(n_3626)
);

NOR2xp33_ASAP7_75t_L g3627 ( 
.A(n_2907),
.B(n_390),
.Y(n_3627)
);

HB1xp67_ASAP7_75t_L g3628 ( 
.A(n_3120),
.Y(n_3628)
);

BUFx6f_ASAP7_75t_L g3629 ( 
.A(n_2999),
.Y(n_3629)
);

NAND2xp5_ASAP7_75t_SL g3630 ( 
.A(n_3024),
.B(n_391),
.Y(n_3630)
);

OR2x2_ASAP7_75t_L g3631 ( 
.A(n_2990),
.B(n_391),
.Y(n_3631)
);

NAND2xp5_ASAP7_75t_L g3632 ( 
.A(n_2828),
.B(n_391),
.Y(n_3632)
);

NAND2xp5_ASAP7_75t_L g3633 ( 
.A(n_2833),
.B(n_392),
.Y(n_3633)
);

NOR2xp67_ASAP7_75t_L g3634 ( 
.A(n_2818),
.B(n_392),
.Y(n_3634)
);

INVx2_ASAP7_75t_L g3635 ( 
.A(n_3230),
.Y(n_3635)
);

INVxp67_ASAP7_75t_L g3636 ( 
.A(n_3148),
.Y(n_3636)
);

AOI21x1_ASAP7_75t_L g3637 ( 
.A1(n_3217),
.A2(n_393),
.B(n_392),
.Y(n_3637)
);

AOI21xp5_ASAP7_75t_L g3638 ( 
.A1(n_2805),
.A2(n_394),
.B(n_393),
.Y(n_3638)
);

BUFx6f_ASAP7_75t_L g3639 ( 
.A(n_2999),
.Y(n_3639)
);

AOI21xp5_ASAP7_75t_L g3640 ( 
.A1(n_2807),
.A2(n_394),
.B(n_393),
.Y(n_3640)
);

NAND2xp5_ASAP7_75t_L g3641 ( 
.A(n_2836),
.B(n_394),
.Y(n_3641)
);

AOI21xp5_ASAP7_75t_L g3642 ( 
.A1(n_2820),
.A2(n_396),
.B(n_395),
.Y(n_3642)
);

OAI21xp33_ASAP7_75t_L g3643 ( 
.A1(n_3087),
.A2(n_36),
.B(n_37),
.Y(n_3643)
);

NAND2xp5_ASAP7_75t_SL g3644 ( 
.A(n_3168),
.B(n_395),
.Y(n_3644)
);

O2A1O1Ixp33_ASAP7_75t_SL g3645 ( 
.A1(n_3310),
.A2(n_396),
.B(n_397),
.C(n_395),
.Y(n_3645)
);

O2A1O1Ixp33_ASAP7_75t_L g3646 ( 
.A1(n_3044),
.A2(n_397),
.B(n_398),
.C(n_396),
.Y(n_3646)
);

NAND2xp5_ASAP7_75t_SL g3647 ( 
.A(n_3168),
.B(n_397),
.Y(n_3647)
);

OAI21xp5_ASAP7_75t_L g3648 ( 
.A1(n_2995),
.A2(n_37),
.B(n_38),
.Y(n_3648)
);

O2A1O1Ixp33_ASAP7_75t_L g3649 ( 
.A1(n_2863),
.A2(n_400),
.B(n_401),
.C(n_399),
.Y(n_3649)
);

AOI21xp5_ASAP7_75t_L g3650 ( 
.A1(n_2820),
.A2(n_400),
.B(n_399),
.Y(n_3650)
);

AOI21xp5_ASAP7_75t_L g3651 ( 
.A1(n_2835),
.A2(n_2840),
.B(n_2838),
.Y(n_3651)
);

OAI22xp5_ASAP7_75t_L g3652 ( 
.A1(n_2893),
.A2(n_402),
.B1(n_403),
.B2(n_401),
.Y(n_3652)
);

AO21x1_ASAP7_75t_L g3653 ( 
.A1(n_3218),
.A2(n_402),
.B(n_401),
.Y(n_3653)
);

AOI21xp5_ASAP7_75t_L g3654 ( 
.A1(n_2835),
.A2(n_404),
.B(n_403),
.Y(n_3654)
);

NOR2xp33_ASAP7_75t_L g3655 ( 
.A(n_2829),
.B(n_403),
.Y(n_3655)
);

INVx2_ASAP7_75t_L g3656 ( 
.A(n_3235),
.Y(n_3656)
);

O2A1O1Ixp33_ASAP7_75t_L g3657 ( 
.A1(n_2989),
.A2(n_405),
.B(n_406),
.C(n_404),
.Y(n_3657)
);

AOI21xp5_ASAP7_75t_L g3658 ( 
.A1(n_2838),
.A2(n_407),
.B(n_406),
.Y(n_3658)
);

NAND2xp5_ASAP7_75t_SL g3659 ( 
.A(n_3168),
.B(n_406),
.Y(n_3659)
);

AND2x2_ASAP7_75t_SL g3660 ( 
.A(n_2854),
.B(n_407),
.Y(n_3660)
);

NAND2xp5_ASAP7_75t_L g3661 ( 
.A(n_2842),
.B(n_407),
.Y(n_3661)
);

CKINVDCx5p33_ASAP7_75t_R g3662 ( 
.A(n_3260),
.Y(n_3662)
);

NOR2xp33_ASAP7_75t_L g3663 ( 
.A(n_2923),
.B(n_408),
.Y(n_3663)
);

INVxp67_ASAP7_75t_L g3664 ( 
.A(n_3228),
.Y(n_3664)
);

AOI21xp5_ASAP7_75t_L g3665 ( 
.A1(n_2840),
.A2(n_409),
.B(n_408),
.Y(n_3665)
);

OAI22xp5_ASAP7_75t_L g3666 ( 
.A1(n_3285),
.A2(n_410),
.B1(n_411),
.B2(n_409),
.Y(n_3666)
);

INVx11_ASAP7_75t_L g3667 ( 
.A(n_3345),
.Y(n_3667)
);

AO21x1_ASAP7_75t_L g3668 ( 
.A1(n_2864),
.A2(n_410),
.B(n_409),
.Y(n_3668)
);

AOI21xp5_ASAP7_75t_L g3669 ( 
.A1(n_2841),
.A2(n_411),
.B(n_410),
.Y(n_3669)
);

INVx3_ASAP7_75t_L g3670 ( 
.A(n_2815),
.Y(n_3670)
);

NOR2xp33_ASAP7_75t_SL g3671 ( 
.A(n_3048),
.B(n_411),
.Y(n_3671)
);

NAND2xp5_ASAP7_75t_L g3672 ( 
.A(n_2876),
.B(n_412),
.Y(n_3672)
);

HB1xp67_ASAP7_75t_L g3673 ( 
.A(n_3150),
.Y(n_3673)
);

AND2x2_ASAP7_75t_L g3674 ( 
.A(n_2932),
.B(n_412),
.Y(n_3674)
);

NAND2xp5_ASAP7_75t_SL g3675 ( 
.A(n_3152),
.B(n_2883),
.Y(n_3675)
);

NAND2xp5_ASAP7_75t_L g3676 ( 
.A(n_2895),
.B(n_413),
.Y(n_3676)
);

NOR2xp33_ASAP7_75t_L g3677 ( 
.A(n_2889),
.B(n_413),
.Y(n_3677)
);

AOI21xp5_ASAP7_75t_L g3678 ( 
.A1(n_2841),
.A2(n_415),
.B(n_414),
.Y(n_3678)
);

NAND2xp5_ASAP7_75t_L g3679 ( 
.A(n_2904),
.B(n_414),
.Y(n_3679)
);

A2O1A1Ixp33_ASAP7_75t_L g3680 ( 
.A1(n_3159),
.A2(n_39),
.B(n_37),
.C(n_38),
.Y(n_3680)
);

INVx1_ASAP7_75t_L g3681 ( 
.A(n_2945),
.Y(n_3681)
);

OAI321xp33_ASAP7_75t_L g3682 ( 
.A1(n_3446),
.A2(n_40),
.A3(n_42),
.B1(n_38),
.B2(n_39),
.C(n_41),
.Y(n_3682)
);

AOI21xp5_ASAP7_75t_L g3683 ( 
.A1(n_2845),
.A2(n_416),
.B(n_415),
.Y(n_3683)
);

NAND2xp5_ASAP7_75t_L g3684 ( 
.A(n_2952),
.B(n_416),
.Y(n_3684)
);

NOR2xp33_ASAP7_75t_L g3685 ( 
.A(n_3066),
.B(n_416),
.Y(n_3685)
);

AOI21xp5_ASAP7_75t_L g3686 ( 
.A1(n_2845),
.A2(n_418),
.B(n_417),
.Y(n_3686)
);

OAI21xp5_ASAP7_75t_L g3687 ( 
.A1(n_2994),
.A2(n_39),
.B(n_40),
.Y(n_3687)
);

AOI21xp5_ASAP7_75t_L g3688 ( 
.A1(n_2852),
.A2(n_418),
.B(n_417),
.Y(n_3688)
);

INVx1_ASAP7_75t_L g3689 ( 
.A(n_2956),
.Y(n_3689)
);

BUFx2_ASAP7_75t_L g3690 ( 
.A(n_2973),
.Y(n_3690)
);

AOI21xp5_ASAP7_75t_L g3691 ( 
.A1(n_2852),
.A2(n_419),
.B(n_418),
.Y(n_3691)
);

NOR2xp33_ASAP7_75t_L g3692 ( 
.A(n_2874),
.B(n_2924),
.Y(n_3692)
);

NAND2xp5_ASAP7_75t_L g3693 ( 
.A(n_2961),
.B(n_420),
.Y(n_3693)
);

NAND2xp5_ASAP7_75t_L g3694 ( 
.A(n_2969),
.B(n_420),
.Y(n_3694)
);

NAND2xp5_ASAP7_75t_L g3695 ( 
.A(n_2975),
.B(n_420),
.Y(n_3695)
);

NOR2xp33_ASAP7_75t_L g3696 ( 
.A(n_2860),
.B(n_421),
.Y(n_3696)
);

INVx2_ASAP7_75t_L g3697 ( 
.A(n_3244),
.Y(n_3697)
);

INVx1_ASAP7_75t_L g3698 ( 
.A(n_2981),
.Y(n_3698)
);

OAI21x1_ASAP7_75t_SL g3699 ( 
.A1(n_3281),
.A2(n_422),
.B(n_421),
.Y(n_3699)
);

HB1xp67_ASAP7_75t_L g3700 ( 
.A(n_3436),
.Y(n_3700)
);

NOR2xp67_ASAP7_75t_L g3701 ( 
.A(n_2855),
.B(n_421),
.Y(n_3701)
);

NAND2xp5_ASAP7_75t_L g3702 ( 
.A(n_2990),
.B(n_423),
.Y(n_3702)
);

AOI21xp5_ASAP7_75t_L g3703 ( 
.A1(n_2853),
.A2(n_424),
.B(n_423),
.Y(n_3703)
);

INVx2_ASAP7_75t_SL g3704 ( 
.A(n_3124),
.Y(n_3704)
);

AOI21xp5_ASAP7_75t_L g3705 ( 
.A1(n_2853),
.A2(n_425),
.B(n_424),
.Y(n_3705)
);

NAND2x1_ASAP7_75t_L g3706 ( 
.A(n_2936),
.B(n_426),
.Y(n_3706)
);

INVx1_ASAP7_75t_L g3707 ( 
.A(n_3031),
.Y(n_3707)
);

NAND2x1p5_ASAP7_75t_L g3708 ( 
.A(n_3209),
.B(n_426),
.Y(n_3708)
);

O2A1O1Ixp33_ASAP7_75t_L g3709 ( 
.A1(n_3301),
.A2(n_427),
.B(n_428),
.C(n_426),
.Y(n_3709)
);

OAI22xp5_ASAP7_75t_L g3710 ( 
.A1(n_3305),
.A2(n_429),
.B1(n_430),
.B2(n_427),
.Y(n_3710)
);

OAI21xp33_ASAP7_75t_L g3711 ( 
.A1(n_3090),
.A2(n_39),
.B(n_41),
.Y(n_3711)
);

AOI21xp5_ASAP7_75t_L g3712 ( 
.A1(n_2858),
.A2(n_430),
.B(n_429),
.Y(n_3712)
);

NAND2xp5_ASAP7_75t_L g3713 ( 
.A(n_2991),
.B(n_429),
.Y(n_3713)
);

NAND2xp5_ASAP7_75t_L g3714 ( 
.A(n_2991),
.B(n_431),
.Y(n_3714)
);

AOI22xp33_ASAP7_75t_L g3715 ( 
.A1(n_3109),
.A2(n_432),
.B1(n_433),
.B2(n_431),
.Y(n_3715)
);

NAND2xp5_ASAP7_75t_L g3716 ( 
.A(n_2858),
.B(n_431),
.Y(n_3716)
);

INVx1_ASAP7_75t_L g3717 ( 
.A(n_2998),
.Y(n_3717)
);

AOI21xp5_ASAP7_75t_L g3718 ( 
.A1(n_2861),
.A2(n_433),
.B(n_432),
.Y(n_3718)
);

INVx1_ASAP7_75t_L g3719 ( 
.A(n_3281),
.Y(n_3719)
);

INVxp33_ASAP7_75t_SL g3720 ( 
.A(n_2912),
.Y(n_3720)
);

INVx2_ASAP7_75t_L g3721 ( 
.A(n_3247),
.Y(n_3721)
);

NAND2x1p5_ASAP7_75t_L g3722 ( 
.A(n_2901),
.B(n_2931),
.Y(n_3722)
);

AOI21xp5_ASAP7_75t_L g3723 ( 
.A1(n_2861),
.A2(n_435),
.B(n_434),
.Y(n_3723)
);

AOI22x1_ASAP7_75t_L g3724 ( 
.A1(n_3219),
.A2(n_435),
.B1(n_436),
.B2(n_434),
.Y(n_3724)
);

AOI22xp5_ASAP7_75t_L g3725 ( 
.A1(n_2974),
.A2(n_436),
.B1(n_437),
.B2(n_434),
.Y(n_3725)
);

A2O1A1Ixp33_ASAP7_75t_L g3726 ( 
.A1(n_3432),
.A2(n_43),
.B(n_41),
.C(n_42),
.Y(n_3726)
);

OAI21xp5_ASAP7_75t_L g3727 ( 
.A1(n_2994),
.A2(n_42),
.B(n_43),
.Y(n_3727)
);

NOR2x1p5_ASAP7_75t_SL g3728 ( 
.A(n_2941),
.B(n_436),
.Y(n_3728)
);

NAND2xp5_ASAP7_75t_SL g3729 ( 
.A(n_3152),
.B(n_437),
.Y(n_3729)
);

AOI21xp5_ASAP7_75t_L g3730 ( 
.A1(n_2866),
.A2(n_438),
.B(n_437),
.Y(n_3730)
);

NAND2xp5_ASAP7_75t_L g3731 ( 
.A(n_2866),
.B(n_2882),
.Y(n_3731)
);

AOI22xp33_ASAP7_75t_L g3732 ( 
.A1(n_3239),
.A2(n_439),
.B1(n_440),
.B2(n_438),
.Y(n_3732)
);

BUFx2_ASAP7_75t_L g3733 ( 
.A(n_3345),
.Y(n_3733)
);

NAND2xp5_ASAP7_75t_L g3734 ( 
.A(n_2882),
.B(n_438),
.Y(n_3734)
);

AOI21xp5_ASAP7_75t_L g3735 ( 
.A1(n_2980),
.A2(n_440),
.B(n_439),
.Y(n_3735)
);

AOI21xp5_ASAP7_75t_L g3736 ( 
.A1(n_2980),
.A2(n_440),
.B(n_439),
.Y(n_3736)
);

AOI21xp5_ASAP7_75t_L g3737 ( 
.A1(n_2985),
.A2(n_442),
.B(n_441),
.Y(n_3737)
);

NAND2xp5_ASAP7_75t_SL g3738 ( 
.A(n_3152),
.B(n_441),
.Y(n_3738)
);

BUFx6f_ASAP7_75t_L g3739 ( 
.A(n_3123),
.Y(n_3739)
);

NAND2xp5_ASAP7_75t_L g3740 ( 
.A(n_3034),
.B(n_442),
.Y(n_3740)
);

BUFx2_ASAP7_75t_L g3741 ( 
.A(n_3345),
.Y(n_3741)
);

OAI21xp5_ASAP7_75t_L g3742 ( 
.A1(n_2985),
.A2(n_42),
.B(n_43),
.Y(n_3742)
);

INVx1_ASAP7_75t_L g3743 ( 
.A(n_3283),
.Y(n_3743)
);

AOI22xp5_ASAP7_75t_L g3744 ( 
.A1(n_2816),
.A2(n_443),
.B1(n_444),
.B2(n_442),
.Y(n_3744)
);

INVx2_ASAP7_75t_L g3745 ( 
.A(n_3249),
.Y(n_3745)
);

AOI21xp5_ASAP7_75t_L g3746 ( 
.A1(n_3005),
.A2(n_444),
.B(n_443),
.Y(n_3746)
);

AO21x1_ASAP7_75t_L g3747 ( 
.A1(n_3076),
.A2(n_445),
.B(n_444),
.Y(n_3747)
);

AOI22xp5_ASAP7_75t_L g3748 ( 
.A1(n_2978),
.A2(n_446),
.B1(n_447),
.B2(n_445),
.Y(n_3748)
);

AOI21xp5_ASAP7_75t_L g3749 ( 
.A1(n_3005),
.A2(n_446),
.B(n_445),
.Y(n_3749)
);

AOI21xp5_ASAP7_75t_L g3750 ( 
.A1(n_3108),
.A2(n_447),
.B(n_446),
.Y(n_3750)
);

AOI21x1_ASAP7_75t_L g3751 ( 
.A1(n_3147),
.A2(n_448),
.B(n_447),
.Y(n_3751)
);

AOI21xp5_ASAP7_75t_L g3752 ( 
.A1(n_3172),
.A2(n_449),
.B(n_448),
.Y(n_3752)
);

NOR2xp33_ASAP7_75t_L g3753 ( 
.A(n_2850),
.B(n_448),
.Y(n_3753)
);

INVx1_ASAP7_75t_L g3754 ( 
.A(n_3283),
.Y(n_3754)
);

OAI22xp5_ASAP7_75t_L g3755 ( 
.A1(n_3318),
.A2(n_450),
.B1(n_451),
.B2(n_449),
.Y(n_3755)
);

AOI21xp5_ASAP7_75t_L g3756 ( 
.A1(n_2890),
.A2(n_450),
.B(n_449),
.Y(n_3756)
);

INVx1_ASAP7_75t_L g3757 ( 
.A(n_3284),
.Y(n_3757)
);

OAI21xp5_ASAP7_75t_L g3758 ( 
.A1(n_2928),
.A2(n_43),
.B(n_44),
.Y(n_3758)
);

AOI21xp5_ASAP7_75t_L g3759 ( 
.A1(n_2891),
.A2(n_452),
.B(n_451),
.Y(n_3759)
);

AOI21xp5_ASAP7_75t_L g3760 ( 
.A1(n_2919),
.A2(n_453),
.B(n_452),
.Y(n_3760)
);

INVx2_ASAP7_75t_L g3761 ( 
.A(n_3251),
.Y(n_3761)
);

AOI21xp5_ASAP7_75t_L g3762 ( 
.A1(n_2930),
.A2(n_454),
.B(n_453),
.Y(n_3762)
);

AND2x4_ASAP7_75t_L g3763 ( 
.A(n_3079),
.B(n_453),
.Y(n_3763)
);

NAND2xp5_ASAP7_75t_L g3764 ( 
.A(n_3101),
.B(n_454),
.Y(n_3764)
);

AOI21xp5_ASAP7_75t_L g3765 ( 
.A1(n_2934),
.A2(n_455),
.B(n_454),
.Y(n_3765)
);

BUFx6f_ASAP7_75t_L g3766 ( 
.A(n_3123),
.Y(n_3766)
);

INVx6_ASAP7_75t_L g3767 ( 
.A(n_2886),
.Y(n_3767)
);

AOI21xp5_ASAP7_75t_L g3768 ( 
.A1(n_3204),
.A2(n_456),
.B(n_455),
.Y(n_3768)
);

AOI21xp5_ASAP7_75t_L g3769 ( 
.A1(n_3056),
.A2(n_3064),
.B(n_3058),
.Y(n_3769)
);

NAND2xp5_ASAP7_75t_SL g3770 ( 
.A(n_2918),
.B(n_455),
.Y(n_3770)
);

O2A1O1Ixp33_ASAP7_75t_L g3771 ( 
.A1(n_3304),
.A2(n_457),
.B(n_458),
.C(n_456),
.Y(n_3771)
);

AO21x1_ASAP7_75t_L g3772 ( 
.A1(n_3076),
.A2(n_457),
.B(n_456),
.Y(n_3772)
);

AND2x2_ASAP7_75t_L g3773 ( 
.A(n_3436),
.B(n_457),
.Y(n_3773)
);

NAND2x1p5_ASAP7_75t_L g3774 ( 
.A(n_3226),
.B(n_458),
.Y(n_3774)
);

AOI21xp5_ASAP7_75t_L g3775 ( 
.A1(n_3065),
.A2(n_460),
.B(n_459),
.Y(n_3775)
);

OAI22xp5_ASAP7_75t_L g3776 ( 
.A1(n_3325),
.A2(n_460),
.B1(n_461),
.B2(n_459),
.Y(n_3776)
);

AOI22xp5_ASAP7_75t_L g3777 ( 
.A1(n_2963),
.A2(n_461),
.B1(n_462),
.B2(n_460),
.Y(n_3777)
);

NAND2xp5_ASAP7_75t_L g3778 ( 
.A(n_3081),
.B(n_463),
.Y(n_3778)
);

AO21x1_ASAP7_75t_L g3779 ( 
.A1(n_2870),
.A2(n_465),
.B(n_464),
.Y(n_3779)
);

INVx2_ASAP7_75t_L g3780 ( 
.A(n_3259),
.Y(n_3780)
);

NOR2xp33_ASAP7_75t_L g3781 ( 
.A(n_3141),
.B(n_464),
.Y(n_3781)
);

AOI21xp5_ASAP7_75t_L g3782 ( 
.A1(n_3236),
.A2(n_465),
.B(n_464),
.Y(n_3782)
);

NAND2xp5_ASAP7_75t_SL g3783 ( 
.A(n_3265),
.B(n_466),
.Y(n_3783)
);

INVx2_ASAP7_75t_L g3784 ( 
.A(n_3264),
.Y(n_3784)
);

OAI21xp5_ASAP7_75t_L g3785 ( 
.A1(n_2954),
.A2(n_44),
.B(n_46),
.Y(n_3785)
);

NOR3xp33_ASAP7_75t_SL g3786 ( 
.A(n_2892),
.B(n_468),
.C(n_467),
.Y(n_3786)
);

AOI22xp33_ASAP7_75t_L g3787 ( 
.A1(n_3282),
.A2(n_3423),
.B1(n_2937),
.B2(n_3008),
.Y(n_3787)
);

HB1xp67_ASAP7_75t_L g3788 ( 
.A(n_3036),
.Y(n_3788)
);

NAND2xp5_ASAP7_75t_L g3789 ( 
.A(n_3085),
.B(n_467),
.Y(n_3789)
);

NAND2xp33_ASAP7_75t_L g3790 ( 
.A(n_2941),
.B(n_468),
.Y(n_3790)
);

NAND2xp5_ASAP7_75t_L g3791 ( 
.A(n_3157),
.B(n_468),
.Y(n_3791)
);

BUFx6f_ASAP7_75t_L g3792 ( 
.A(n_3123),
.Y(n_3792)
);

AOI21xp5_ASAP7_75t_L g3793 ( 
.A1(n_3273),
.A2(n_470),
.B(n_469),
.Y(n_3793)
);

NAND2xp5_ASAP7_75t_L g3794 ( 
.A(n_3170),
.B(n_469),
.Y(n_3794)
);

O2A1O1Ixp33_ASAP7_75t_L g3795 ( 
.A1(n_3341),
.A2(n_471),
.B(n_472),
.C(n_470),
.Y(n_3795)
);

OAI21xp5_ASAP7_75t_L g3796 ( 
.A1(n_2955),
.A2(n_2967),
.B(n_2896),
.Y(n_3796)
);

NAND2xp5_ASAP7_75t_L g3797 ( 
.A(n_3107),
.B(n_470),
.Y(n_3797)
);

INVx2_ASAP7_75t_L g3798 ( 
.A(n_3280),
.Y(n_3798)
);

NAND2xp5_ASAP7_75t_L g3799 ( 
.A(n_2996),
.B(n_471),
.Y(n_3799)
);

AOI22xp5_ASAP7_75t_L g3800 ( 
.A1(n_2987),
.A2(n_2939),
.B1(n_2948),
.B2(n_3052),
.Y(n_3800)
);

AOI21xp5_ASAP7_75t_L g3801 ( 
.A1(n_3287),
.A2(n_472),
.B(n_471),
.Y(n_3801)
);

NAND2xp5_ASAP7_75t_L g3802 ( 
.A(n_3012),
.B(n_472),
.Y(n_3802)
);

CKINVDCx10_ASAP7_75t_R g3803 ( 
.A(n_2929),
.Y(n_3803)
);

BUFx2_ASAP7_75t_L g3804 ( 
.A(n_3345),
.Y(n_3804)
);

INVx1_ASAP7_75t_L g3805 ( 
.A(n_3284),
.Y(n_3805)
);

AND2x2_ASAP7_75t_L g3806 ( 
.A(n_3246),
.B(n_473),
.Y(n_3806)
);

NAND3xp33_ASAP7_75t_L g3807 ( 
.A(n_2856),
.B(n_3277),
.C(n_3122),
.Y(n_3807)
);

BUFx6f_ASAP7_75t_L g3808 ( 
.A(n_3360),
.Y(n_3808)
);

NAND2xp5_ASAP7_75t_L g3809 ( 
.A(n_3000),
.B(n_473),
.Y(n_3809)
);

INVx1_ASAP7_75t_L g3810 ( 
.A(n_3289),
.Y(n_3810)
);

NAND2xp5_ASAP7_75t_SL g3811 ( 
.A(n_2962),
.B(n_474),
.Y(n_3811)
);

INVx2_ASAP7_75t_L g3812 ( 
.A(n_3300),
.Y(n_3812)
);

O2A1O1Ixp5_ASAP7_75t_L g3813 ( 
.A1(n_3155),
.A2(n_475),
.B(n_476),
.C(n_474),
.Y(n_3813)
);

INVx1_ASAP7_75t_L g3814 ( 
.A(n_3289),
.Y(n_3814)
);

INVx3_ASAP7_75t_L g3815 ( 
.A(n_2819),
.Y(n_3815)
);

INVx4_ASAP7_75t_L g3816 ( 
.A(n_2936),
.Y(n_3816)
);

AOI21xp5_ASAP7_75t_L g3817 ( 
.A1(n_3303),
.A2(n_475),
.B(n_474),
.Y(n_3817)
);

A2O1A1Ixp33_ASAP7_75t_L g3818 ( 
.A1(n_2881),
.A2(n_48),
.B(n_46),
.C(n_47),
.Y(n_3818)
);

NAND2xp5_ASAP7_75t_L g3819 ( 
.A(n_3000),
.B(n_475),
.Y(n_3819)
);

OAI21xp5_ASAP7_75t_L g3820 ( 
.A1(n_3050),
.A2(n_46),
.B(n_47),
.Y(n_3820)
);

A2O1A1Ixp33_ASAP7_75t_L g3821 ( 
.A1(n_3194),
.A2(n_48),
.B(n_46),
.C(n_47),
.Y(n_3821)
);

NOR3xp33_ASAP7_75t_L g3822 ( 
.A(n_2965),
.B(n_477),
.C(n_476),
.Y(n_3822)
);

INVx1_ASAP7_75t_L g3823 ( 
.A(n_3290),
.Y(n_3823)
);

OAI22xp5_ASAP7_75t_L g3824 ( 
.A1(n_3383),
.A2(n_478),
.B1(n_479),
.B2(n_476),
.Y(n_3824)
);

OAI21xp5_ASAP7_75t_L g3825 ( 
.A1(n_3290),
.A2(n_47),
.B(n_48),
.Y(n_3825)
);

NOR2xp33_ASAP7_75t_L g3826 ( 
.A(n_2865),
.B(n_478),
.Y(n_3826)
);

NOR2xp33_ASAP7_75t_L g3827 ( 
.A(n_2867),
.B(n_478),
.Y(n_3827)
);

AOI21xp5_ASAP7_75t_L g3828 ( 
.A1(n_3319),
.A2(n_480),
.B(n_479),
.Y(n_3828)
);

NOR3xp33_ASAP7_75t_L g3829 ( 
.A(n_2873),
.B(n_480),
.C(n_479),
.Y(n_3829)
);

NAND2xp5_ASAP7_75t_SL g3830 ( 
.A(n_2962),
.B(n_481),
.Y(n_3830)
);

OR2x6_ASAP7_75t_L g3831 ( 
.A(n_3356),
.B(n_481),
.Y(n_3831)
);

NAND2xp5_ASAP7_75t_L g3832 ( 
.A(n_3002),
.B(n_481),
.Y(n_3832)
);

AOI21xp5_ASAP7_75t_L g3833 ( 
.A1(n_3332),
.A2(n_483),
.B(n_482),
.Y(n_3833)
);

AND2x4_ASAP7_75t_L g3834 ( 
.A(n_3250),
.B(n_482),
.Y(n_3834)
);

OAI21xp5_ASAP7_75t_L g3835 ( 
.A1(n_3293),
.A2(n_49),
.B(n_50),
.Y(n_3835)
);

NAND2xp5_ASAP7_75t_L g3836 ( 
.A(n_3002),
.B(n_482),
.Y(n_3836)
);

AOI21xp33_ASAP7_75t_L g3837 ( 
.A1(n_2950),
.A2(n_485),
.B(n_484),
.Y(n_3837)
);

AOI21xp5_ASAP7_75t_L g3838 ( 
.A1(n_3334),
.A2(n_485),
.B(n_484),
.Y(n_3838)
);

CKINVDCx10_ASAP7_75t_R g3839 ( 
.A(n_3416),
.Y(n_3839)
);

NAND2xp5_ASAP7_75t_SL g3840 ( 
.A(n_3011),
.B(n_485),
.Y(n_3840)
);

NAND2xp5_ASAP7_75t_L g3841 ( 
.A(n_3070),
.B(n_3059),
.Y(n_3841)
);

AOI21xp5_ASAP7_75t_L g3842 ( 
.A1(n_3354),
.A2(n_3452),
.B(n_3439),
.Y(n_3842)
);

NAND2xp5_ASAP7_75t_L g3843 ( 
.A(n_3072),
.B(n_486),
.Y(n_3843)
);

AOI21xp5_ASAP7_75t_L g3844 ( 
.A1(n_3362),
.A2(n_487),
.B(n_486),
.Y(n_3844)
);

INVx2_ASAP7_75t_L g3845 ( 
.A(n_3373),
.Y(n_3845)
);

AOI21xp5_ASAP7_75t_L g3846 ( 
.A1(n_3397),
.A2(n_3430),
.B(n_3021),
.Y(n_3846)
);

NOR2xp33_ASAP7_75t_R g3847 ( 
.A(n_3416),
.B(n_50),
.Y(n_3847)
);

OR2x6_ASAP7_75t_L g3848 ( 
.A(n_3306),
.B(n_487),
.Y(n_3848)
);

NAND2xp5_ASAP7_75t_SL g3849 ( 
.A(n_3011),
.B(n_487),
.Y(n_3849)
);

OAI21xp5_ASAP7_75t_L g3850 ( 
.A1(n_3293),
.A2(n_49),
.B(n_51),
.Y(n_3850)
);

INVx2_ASAP7_75t_SL g3851 ( 
.A(n_3400),
.Y(n_3851)
);

AOI21xp5_ASAP7_75t_L g3852 ( 
.A1(n_3019),
.A2(n_489),
.B(n_488),
.Y(n_3852)
);

AOI21xp5_ASAP7_75t_L g3853 ( 
.A1(n_3033),
.A2(n_489),
.B(n_488),
.Y(n_3853)
);

AOI21xp5_ASAP7_75t_L g3854 ( 
.A1(n_3035),
.A2(n_489),
.B(n_488),
.Y(n_3854)
);

AO21x2_ASAP7_75t_L g3855 ( 
.A1(n_3295),
.A2(n_491),
.B(n_490),
.Y(n_3855)
);

INVx1_ASAP7_75t_L g3856 ( 
.A(n_3295),
.Y(n_3856)
);

A2O1A1Ixp33_ASAP7_75t_L g3857 ( 
.A1(n_3203),
.A2(n_53),
.B(n_51),
.C(n_52),
.Y(n_3857)
);

AOI22xp33_ASAP7_75t_L g3858 ( 
.A1(n_3043),
.A2(n_491),
.B1(n_492),
.B2(n_490),
.Y(n_3858)
);

O2A1O1Ixp33_ASAP7_75t_L g3859 ( 
.A1(n_3346),
.A2(n_492),
.B(n_493),
.C(n_491),
.Y(n_3859)
);

O2A1O1Ixp5_ASAP7_75t_L g3860 ( 
.A1(n_3040),
.A2(n_494),
.B(n_495),
.C(n_493),
.Y(n_3860)
);

HB1xp67_ASAP7_75t_L g3861 ( 
.A(n_3037),
.Y(n_3861)
);

INVx2_ASAP7_75t_L g3862 ( 
.A(n_3080),
.Y(n_3862)
);

AOI22xp33_ASAP7_75t_L g3863 ( 
.A1(n_3043),
.A2(n_494),
.B1(n_495),
.B2(n_493),
.Y(n_3863)
);

NAND2xp5_ASAP7_75t_L g3864 ( 
.A(n_3114),
.B(n_494),
.Y(n_3864)
);

OAI21xp5_ASAP7_75t_L g3865 ( 
.A1(n_3297),
.A2(n_51),
.B(n_52),
.Y(n_3865)
);

OAI21xp5_ASAP7_75t_L g3866 ( 
.A1(n_3297),
.A2(n_52),
.B(n_53),
.Y(n_3866)
);

NAND2xp5_ASAP7_75t_L g3867 ( 
.A(n_3156),
.B(n_495),
.Y(n_3867)
);

NAND2xp5_ASAP7_75t_L g3868 ( 
.A(n_3060),
.B(n_496),
.Y(n_3868)
);

AOI21xp5_ASAP7_75t_L g3869 ( 
.A1(n_3047),
.A2(n_497),
.B(n_496),
.Y(n_3869)
);

NAND2xp5_ASAP7_75t_L g3870 ( 
.A(n_2908),
.B(n_496),
.Y(n_3870)
);

INVx2_ASAP7_75t_L g3871 ( 
.A(n_3112),
.Y(n_3871)
);

NAND2xp5_ASAP7_75t_L g3872 ( 
.A(n_2911),
.B(n_497),
.Y(n_3872)
);

BUFx6f_ASAP7_75t_L g3873 ( 
.A(n_3360),
.Y(n_3873)
);

NAND2xp5_ASAP7_75t_L g3874 ( 
.A(n_2894),
.B(n_498),
.Y(n_3874)
);

OAI21xp5_ASAP7_75t_L g3875 ( 
.A1(n_3298),
.A2(n_52),
.B(n_53),
.Y(n_3875)
);

BUFx3_ASAP7_75t_L g3876 ( 
.A(n_2916),
.Y(n_3876)
);

HB1xp67_ASAP7_75t_L g3877 ( 
.A(n_3082),
.Y(n_3877)
);

INVx3_ASAP7_75t_L g3878 ( 
.A(n_2819),
.Y(n_3878)
);

AOI21xp5_ASAP7_75t_L g3879 ( 
.A1(n_3142),
.A2(n_499),
.B(n_498),
.Y(n_3879)
);

BUFx6f_ASAP7_75t_L g3880 ( 
.A(n_3360),
.Y(n_3880)
);

NAND2xp5_ASAP7_75t_SL g3881 ( 
.A(n_2941),
.B(n_500),
.Y(n_3881)
);

INVx3_ASAP7_75t_L g3882 ( 
.A(n_2832),
.Y(n_3882)
);

AOI21xp5_ASAP7_75t_L g3883 ( 
.A1(n_3212),
.A2(n_501),
.B(n_500),
.Y(n_3883)
);

INVx1_ASAP7_75t_L g3884 ( 
.A(n_3298),
.Y(n_3884)
);

INVx1_ASAP7_75t_L g3885 ( 
.A(n_3312),
.Y(n_3885)
);

AND2x2_ASAP7_75t_L g3886 ( 
.A(n_3263),
.B(n_500),
.Y(n_3886)
);

INVx2_ASAP7_75t_L g3887 ( 
.A(n_3042),
.Y(n_3887)
);

AOI22xp5_ASAP7_75t_L g3888 ( 
.A1(n_2984),
.A2(n_503),
.B1(n_504),
.B2(n_502),
.Y(n_3888)
);

NOR2xp33_ASAP7_75t_L g3889 ( 
.A(n_2959),
.B(n_3118),
.Y(n_3889)
);

NOR2xp33_ASAP7_75t_SL g3890 ( 
.A(n_3095),
.B(n_502),
.Y(n_3890)
);

OAI321xp33_ASAP7_75t_L g3891 ( 
.A1(n_3390),
.A2(n_55),
.A3(n_57),
.B1(n_53),
.B2(n_54),
.C(n_56),
.Y(n_3891)
);

NAND2xp5_ASAP7_75t_L g3892 ( 
.A(n_3126),
.B(n_502),
.Y(n_3892)
);

AOI21xp5_ASAP7_75t_L g3893 ( 
.A1(n_3051),
.A2(n_505),
.B(n_503),
.Y(n_3893)
);

AOI21xp5_ASAP7_75t_L g3894 ( 
.A1(n_3312),
.A2(n_506),
.B(n_505),
.Y(n_3894)
);

BUFx6f_ASAP7_75t_L g3895 ( 
.A(n_3376),
.Y(n_3895)
);

NAND2xp5_ASAP7_75t_L g3896 ( 
.A(n_3180),
.B(n_505),
.Y(n_3896)
);

BUFx3_ASAP7_75t_L g3897 ( 
.A(n_2960),
.Y(n_3897)
);

AOI21xp5_ASAP7_75t_L g3898 ( 
.A1(n_3321),
.A2(n_507),
.B(n_506),
.Y(n_3898)
);

NAND2xp5_ASAP7_75t_L g3899 ( 
.A(n_3182),
.B(n_507),
.Y(n_3899)
);

O2A1O1Ixp33_ASAP7_75t_L g3900 ( 
.A1(n_3357),
.A2(n_509),
.B(n_510),
.C(n_508),
.Y(n_3900)
);

OAI22xp5_ASAP7_75t_L g3901 ( 
.A1(n_3420),
.A2(n_509),
.B1(n_510),
.B2(n_508),
.Y(n_3901)
);

AOI22x1_ASAP7_75t_L g3902 ( 
.A1(n_3179),
.A2(n_509),
.B1(n_511),
.B2(n_508),
.Y(n_3902)
);

INVx8_ASAP7_75t_L g3903 ( 
.A(n_3345),
.Y(n_3903)
);

BUFx3_ASAP7_75t_L g3904 ( 
.A(n_3271),
.Y(n_3904)
);

NOR2xp67_ASAP7_75t_L g3905 ( 
.A(n_3409),
.B(n_511),
.Y(n_3905)
);

INVx2_ASAP7_75t_L g3906 ( 
.A(n_3146),
.Y(n_3906)
);

INVx3_ASAP7_75t_L g3907 ( 
.A(n_2832),
.Y(n_3907)
);

BUFx2_ASAP7_75t_SL g3908 ( 
.A(n_3413),
.Y(n_3908)
);

CKINVDCx5p33_ASAP7_75t_R g3909 ( 
.A(n_3377),
.Y(n_3909)
);

NAND2xp5_ASAP7_75t_L g3910 ( 
.A(n_3184),
.B(n_511),
.Y(n_3910)
);

NAND2xp5_ASAP7_75t_SL g3911 ( 
.A(n_2941),
.B(n_512),
.Y(n_3911)
);

INVx4_ASAP7_75t_L g3912 ( 
.A(n_2936),
.Y(n_3912)
);

AND2x2_ASAP7_75t_L g3913 ( 
.A(n_3307),
.B(n_512),
.Y(n_3913)
);

NOR2xp33_ASAP7_75t_L g3914 ( 
.A(n_3125),
.B(n_512),
.Y(n_3914)
);

AO21x1_ASAP7_75t_L g3915 ( 
.A1(n_2870),
.A2(n_514),
.B(n_513),
.Y(n_3915)
);

A2O1A1Ixp33_ASAP7_75t_L g3916 ( 
.A1(n_3321),
.A2(n_56),
.B(n_54),
.C(n_55),
.Y(n_3916)
);

A2O1A1Ixp33_ASAP7_75t_L g3917 ( 
.A1(n_3328),
.A2(n_57),
.B(n_54),
.C(n_55),
.Y(n_3917)
);

NAND2xp5_ASAP7_75t_L g3918 ( 
.A(n_3181),
.B(n_513),
.Y(n_3918)
);

INVx3_ASAP7_75t_L g3919 ( 
.A(n_2851),
.Y(n_3919)
);

AOI21xp5_ASAP7_75t_L g3920 ( 
.A1(n_3328),
.A2(n_514),
.B(n_513),
.Y(n_3920)
);

AOI21xp5_ASAP7_75t_L g3921 ( 
.A1(n_3329),
.A2(n_515),
.B(n_514),
.Y(n_3921)
);

INVx2_ASAP7_75t_L g3922 ( 
.A(n_3192),
.Y(n_3922)
);

AOI21xp5_ASAP7_75t_L g3923 ( 
.A1(n_3329),
.A2(n_516),
.B(n_515),
.Y(n_3923)
);

AOI21xp5_ASAP7_75t_L g3924 ( 
.A1(n_3333),
.A2(n_517),
.B(n_515),
.Y(n_3924)
);

AOI22xp5_ASAP7_75t_L g3925 ( 
.A1(n_3020),
.A2(n_518),
.B1(n_519),
.B2(n_517),
.Y(n_3925)
);

BUFx3_ASAP7_75t_L g3926 ( 
.A(n_3381),
.Y(n_3926)
);

AOI21xp5_ASAP7_75t_L g3927 ( 
.A1(n_3333),
.A2(n_519),
.B(n_517),
.Y(n_3927)
);

NAND2xp5_ASAP7_75t_L g3928 ( 
.A(n_2949),
.B(n_519),
.Y(n_3928)
);

AOI21xp5_ASAP7_75t_L g3929 ( 
.A1(n_3335),
.A2(n_521),
.B(n_520),
.Y(n_3929)
);

AOI21xp5_ASAP7_75t_L g3930 ( 
.A1(n_3335),
.A2(n_521),
.B(n_520),
.Y(n_3930)
);

BUFx6f_ASAP7_75t_L g3931 ( 
.A(n_3376),
.Y(n_3931)
);

AOI21xp5_ASAP7_75t_L g3932 ( 
.A1(n_3336),
.A2(n_521),
.B(n_520),
.Y(n_3932)
);

INVx3_ASAP7_75t_L g3933 ( 
.A(n_2851),
.Y(n_3933)
);

OAI21xp5_ASAP7_75t_L g3934 ( 
.A1(n_3336),
.A2(n_55),
.B(n_57),
.Y(n_3934)
);

OAI321xp33_ASAP7_75t_L g3935 ( 
.A1(n_3427),
.A2(n_60),
.A3(n_62),
.B1(n_58),
.B2(n_59),
.C(n_61),
.Y(n_3935)
);

NAND2xp5_ASAP7_75t_L g3936 ( 
.A(n_2951),
.B(n_2909),
.Y(n_3936)
);

NAND2xp5_ASAP7_75t_SL g3937 ( 
.A(n_2941),
.B(n_522),
.Y(n_3937)
);

AND2x2_ASAP7_75t_L g3938 ( 
.A(n_3314),
.B(n_522),
.Y(n_3938)
);

A2O1A1Ixp33_ASAP7_75t_L g3939 ( 
.A1(n_3342),
.A2(n_60),
.B(n_58),
.C(n_59),
.Y(n_3939)
);

AOI21xp5_ASAP7_75t_L g3940 ( 
.A1(n_3342),
.A2(n_523),
.B(n_522),
.Y(n_3940)
);

INVx1_ASAP7_75t_L g3941 ( 
.A(n_3347),
.Y(n_3941)
);

AOI21xp5_ASAP7_75t_L g3942 ( 
.A1(n_3347),
.A2(n_525),
.B(n_524),
.Y(n_3942)
);

AOI21xp5_ASAP7_75t_L g3943 ( 
.A1(n_3349),
.A2(n_525),
.B(n_524),
.Y(n_3943)
);

NOR3xp33_ASAP7_75t_L g3944 ( 
.A(n_3117),
.B(n_526),
.C(n_524),
.Y(n_3944)
);

OAI22xp5_ASAP7_75t_L g3945 ( 
.A1(n_3234),
.A2(n_527),
.B1(n_528),
.B2(n_526),
.Y(n_3945)
);

AND2x2_ASAP7_75t_L g3946 ( 
.A(n_3326),
.B(n_526),
.Y(n_3946)
);

NOR2xp33_ASAP7_75t_L g3947 ( 
.A(n_3045),
.B(n_527),
.Y(n_3947)
);

AOI21xp5_ASAP7_75t_L g3948 ( 
.A1(n_3349),
.A2(n_529),
.B(n_527),
.Y(n_3948)
);

O2A1O1Ixp33_ASAP7_75t_L g3949 ( 
.A1(n_3359),
.A2(n_530),
.B(n_531),
.C(n_529),
.Y(n_3949)
);

INVx2_ASAP7_75t_L g3950 ( 
.A(n_3199),
.Y(n_3950)
);

INVx3_ASAP7_75t_L g3951 ( 
.A(n_2921),
.Y(n_3951)
);

O2A1O1Ixp5_ASAP7_75t_L g3952 ( 
.A1(n_3213),
.A2(n_530),
.B(n_531),
.C(n_529),
.Y(n_3952)
);

A2O1A1Ixp33_ASAP7_75t_L g3953 ( 
.A1(n_3351),
.A2(n_60),
.B(n_58),
.C(n_59),
.Y(n_3953)
);

OAI21xp5_ASAP7_75t_L g3954 ( 
.A1(n_3351),
.A2(n_58),
.B(n_60),
.Y(n_3954)
);

OA21x2_ASAP7_75t_L g3955 ( 
.A1(n_3352),
.A2(n_533),
.B(n_532),
.Y(n_3955)
);

AOI21xp5_ASAP7_75t_L g3956 ( 
.A1(n_3352),
.A2(n_533),
.B(n_532),
.Y(n_3956)
);

NOR2xp33_ASAP7_75t_L g3957 ( 
.A(n_2993),
.B(n_533),
.Y(n_3957)
);

INVx2_ASAP7_75t_L g3958 ( 
.A(n_3173),
.Y(n_3958)
);

A2O1A1Ixp33_ASAP7_75t_L g3959 ( 
.A1(n_3366),
.A2(n_3369),
.B(n_3379),
.C(n_3378),
.Y(n_3959)
);

O2A1O1Ixp33_ASAP7_75t_L g3960 ( 
.A1(n_3363),
.A2(n_535),
.B(n_536),
.C(n_534),
.Y(n_3960)
);

NAND2xp5_ASAP7_75t_L g3961 ( 
.A(n_3158),
.B(n_534),
.Y(n_3961)
);

AOI21xp5_ASAP7_75t_L g3962 ( 
.A1(n_3366),
.A2(n_536),
.B(n_535),
.Y(n_3962)
);

NOR3xp33_ASAP7_75t_L g3963 ( 
.A(n_2810),
.B(n_538),
.C(n_537),
.Y(n_3963)
);

INVx3_ASAP7_75t_L g3964 ( 
.A(n_2921),
.Y(n_3964)
);

HB1xp67_ASAP7_75t_L g3965 ( 
.A(n_3153),
.Y(n_3965)
);

O2A1O1Ixp5_ASAP7_75t_L g3966 ( 
.A1(n_3074),
.A2(n_538),
.B(n_539),
.C(n_537),
.Y(n_3966)
);

NOR3xp33_ASAP7_75t_L g3967 ( 
.A(n_3374),
.B(n_539),
.C(n_537),
.Y(n_3967)
);

NAND2xp5_ASAP7_75t_SL g3968 ( 
.A(n_2941),
.B(n_540),
.Y(n_3968)
);

INVx2_ASAP7_75t_L g3969 ( 
.A(n_3055),
.Y(n_3969)
);

BUFx6f_ASAP7_75t_L g3970 ( 
.A(n_3376),
.Y(n_3970)
);

OAI21xp5_ASAP7_75t_L g3971 ( 
.A1(n_3369),
.A2(n_61),
.B(n_62),
.Y(n_3971)
);

AOI21x1_ASAP7_75t_L g3972 ( 
.A1(n_3201),
.A2(n_541),
.B(n_540),
.Y(n_3972)
);

A2O1A1Ixp33_ASAP7_75t_L g3973 ( 
.A1(n_3378),
.A2(n_64),
.B(n_62),
.C(n_63),
.Y(n_3973)
);

AOI21xp5_ASAP7_75t_L g3974 ( 
.A1(n_3379),
.A2(n_541),
.B(n_540),
.Y(n_3974)
);

BUFx4f_ASAP7_75t_L g3975 ( 
.A(n_2936),
.Y(n_3975)
);

AOI21xp5_ASAP7_75t_L g3976 ( 
.A1(n_3380),
.A2(n_3392),
.B(n_3391),
.Y(n_3976)
);

NAND2xp5_ASAP7_75t_L g3977 ( 
.A(n_3380),
.B(n_541),
.Y(n_3977)
);

NAND2xp5_ASAP7_75t_L g3978 ( 
.A(n_3391),
.B(n_542),
.Y(n_3978)
);

OAI21xp33_ASAP7_75t_L g3979 ( 
.A1(n_2905),
.A2(n_3093),
.B(n_3160),
.Y(n_3979)
);

HB1xp67_ASAP7_75t_L g3980 ( 
.A(n_3167),
.Y(n_3980)
);

NAND2xp5_ASAP7_75t_L g3981 ( 
.A(n_3392),
.B(n_542),
.Y(n_3981)
);

NOR2x1p5_ASAP7_75t_L g3982 ( 
.A(n_3415),
.B(n_542),
.Y(n_3982)
);

AOI21xp5_ASAP7_75t_L g3983 ( 
.A1(n_3393),
.A2(n_3403),
.B(n_3402),
.Y(n_3983)
);

INVx2_ASAP7_75t_L g3984 ( 
.A(n_3089),
.Y(n_3984)
);

NAND2xp5_ASAP7_75t_L g3985 ( 
.A(n_3393),
.B(n_543),
.Y(n_3985)
);

NAND2xp5_ASAP7_75t_L g3986 ( 
.A(n_3402),
.B(n_543),
.Y(n_3986)
);

OAI21xp5_ASAP7_75t_L g3987 ( 
.A1(n_3403),
.A2(n_62),
.B(n_63),
.Y(n_3987)
);

OAI321xp33_ASAP7_75t_L g3988 ( 
.A1(n_3286),
.A2(n_65),
.A3(n_67),
.B1(n_63),
.B2(n_64),
.C(n_66),
.Y(n_3988)
);

NAND2xp5_ASAP7_75t_SL g3989 ( 
.A(n_3006),
.B(n_543),
.Y(n_3989)
);

OAI21xp5_ASAP7_75t_L g3990 ( 
.A1(n_3405),
.A2(n_64),
.B(n_65),
.Y(n_3990)
);

NOR2xp33_ASAP7_75t_R g3991 ( 
.A(n_3433),
.B(n_65),
.Y(n_3991)
);

O2A1O1Ixp33_ASAP7_75t_L g3992 ( 
.A1(n_3384),
.A2(n_545),
.B(n_546),
.C(n_544),
.Y(n_3992)
);

NAND2xp5_ASAP7_75t_L g3993 ( 
.A(n_3405),
.B(n_544),
.Y(n_3993)
);

NAND2xp5_ASAP7_75t_L g3994 ( 
.A(n_3421),
.B(n_544),
.Y(n_3994)
);

OAI21xp5_ASAP7_75t_L g3995 ( 
.A1(n_3421),
.A2(n_64),
.B(n_65),
.Y(n_3995)
);

INVx1_ASAP7_75t_L g3996 ( 
.A(n_3424),
.Y(n_3996)
);

AOI21xp5_ASAP7_75t_L g3997 ( 
.A1(n_3424),
.A2(n_547),
.B(n_545),
.Y(n_3997)
);

NAND2xp5_ASAP7_75t_L g3998 ( 
.A(n_3425),
.B(n_547),
.Y(n_3998)
);

AOI21xp5_ASAP7_75t_L g3999 ( 
.A1(n_3425),
.A2(n_548),
.B(n_547),
.Y(n_3999)
);

AND2x2_ASAP7_75t_L g4000 ( 
.A(n_3350),
.B(n_3412),
.Y(n_4000)
);

NOR2x1_ASAP7_75t_L g4001 ( 
.A(n_2947),
.B(n_548),
.Y(n_4001)
);

NAND2xp5_ASAP7_75t_L g4002 ( 
.A(n_3429),
.B(n_548),
.Y(n_4002)
);

NAND2xp5_ASAP7_75t_L g4003 ( 
.A(n_3429),
.B(n_549),
.Y(n_4003)
);

INVx2_ASAP7_75t_L g4004 ( 
.A(n_3431),
.Y(n_4004)
);

INVx1_ASAP7_75t_L g4005 ( 
.A(n_3431),
.Y(n_4005)
);

NOR2xp33_ASAP7_75t_L g4006 ( 
.A(n_2811),
.B(n_550),
.Y(n_4006)
);

INVx1_ASAP7_75t_L g4007 ( 
.A(n_3435),
.Y(n_4007)
);

INVx4_ASAP7_75t_L g4008 ( 
.A(n_2936),
.Y(n_4008)
);

OAI22xp5_ASAP7_75t_L g4009 ( 
.A1(n_2914),
.A2(n_552),
.B1(n_553),
.B2(n_550),
.Y(n_4009)
);

NAND2xp5_ASAP7_75t_L g4010 ( 
.A(n_3435),
.B(n_550),
.Y(n_4010)
);

NOR2xp33_ASAP7_75t_L g4011 ( 
.A(n_3023),
.B(n_553),
.Y(n_4011)
);

INVx2_ASAP7_75t_L g4012 ( 
.A(n_3438),
.Y(n_4012)
);

NAND2xp5_ASAP7_75t_L g4013 ( 
.A(n_3438),
.B(n_553),
.Y(n_4013)
);

AOI21xp5_ASAP7_75t_L g4014 ( 
.A1(n_3441),
.A2(n_555),
.B(n_554),
.Y(n_4014)
);

BUFx6f_ASAP7_75t_L g4015 ( 
.A(n_3414),
.Y(n_4015)
);

AOI21xp5_ASAP7_75t_L g4016 ( 
.A1(n_3441),
.A2(n_555),
.B(n_554),
.Y(n_4016)
);

AOI21xp5_ASAP7_75t_L g4017 ( 
.A1(n_3447),
.A2(n_556),
.B(n_555),
.Y(n_4017)
);

NAND2xp5_ASAP7_75t_SL g4018 ( 
.A(n_3006),
.B(n_556),
.Y(n_4018)
);

AOI21xp5_ASAP7_75t_L g4019 ( 
.A1(n_3447),
.A2(n_3448),
.B(n_3088),
.Y(n_4019)
);

AOI222xp33_ASAP7_75t_L g4020 ( 
.A1(n_3208),
.A2(n_560),
.B1(n_558),
.B2(n_561),
.C1(n_559),
.C2(n_557),
.Y(n_4020)
);

AOI21xp5_ASAP7_75t_L g4021 ( 
.A1(n_3448),
.A2(n_558),
.B(n_557),
.Y(n_4021)
);

AOI21xp5_ASAP7_75t_L g4022 ( 
.A1(n_3063),
.A2(n_558),
.B(n_557),
.Y(n_4022)
);

INVx2_ASAP7_75t_L g4023 ( 
.A(n_3414),
.Y(n_4023)
);

O2A1O1Ixp33_ASAP7_75t_L g4024 ( 
.A1(n_3387),
.A2(n_560),
.B(n_562),
.C(n_559),
.Y(n_4024)
);

AO21x1_ASAP7_75t_L g4025 ( 
.A1(n_2914),
.A2(n_560),
.B(n_559),
.Y(n_4025)
);

OAI22xp5_ASAP7_75t_L g4026 ( 
.A1(n_3028),
.A2(n_563),
.B1(n_564),
.B2(n_562),
.Y(n_4026)
);

AOI21xp5_ASAP7_75t_L g4027 ( 
.A1(n_3131),
.A2(n_563),
.B(n_562),
.Y(n_4027)
);

OAI21xp5_ASAP7_75t_L g4028 ( 
.A1(n_3769),
.A2(n_3128),
.B(n_3143),
.Y(n_4028)
);

NAND2xp5_ASAP7_75t_L g4029 ( 
.A(n_3979),
.B(n_3025),
.Y(n_4029)
);

INVxp67_ASAP7_75t_L g4030 ( 
.A(n_3535),
.Y(n_4030)
);

OAI22xp5_ASAP7_75t_L g4031 ( 
.A1(n_3667),
.A2(n_3171),
.B1(n_3186),
.B2(n_3288),
.Y(n_4031)
);

NOR2xp33_ASAP7_75t_SL g4032 ( 
.A(n_3720),
.B(n_3215),
.Y(n_4032)
);

NOR2xp33_ASAP7_75t_L g4033 ( 
.A(n_3482),
.B(n_3178),
.Y(n_4033)
);

A2O1A1Ixp33_ASAP7_75t_L g4034 ( 
.A1(n_3598),
.A2(n_3116),
.B(n_3237),
.C(n_3227),
.Y(n_4034)
);

OAI22xp5_ASAP7_75t_L g4035 ( 
.A1(n_3561),
.A2(n_3344),
.B1(n_3371),
.B2(n_3330),
.Y(n_4035)
);

NOR2xp33_ASAP7_75t_L g4036 ( 
.A(n_3508),
.B(n_2953),
.Y(n_4036)
);

CKINVDCx8_ASAP7_75t_R g4037 ( 
.A(n_3463),
.Y(n_4037)
);

O2A1O1Ixp33_ASAP7_75t_L g4038 ( 
.A1(n_3500),
.A2(n_3401),
.B(n_3411),
.C(n_3388),
.Y(n_4038)
);

INVx1_ASAP7_75t_L g4039 ( 
.A(n_3603),
.Y(n_4039)
);

BUFx6f_ASAP7_75t_L g4040 ( 
.A(n_3975),
.Y(n_4040)
);

INVx2_ASAP7_75t_L g4041 ( 
.A(n_3474),
.Y(n_4041)
);

INVx1_ASAP7_75t_SL g4042 ( 
.A(n_3908),
.Y(n_4042)
);

AOI22xp33_ASAP7_75t_L g4043 ( 
.A1(n_3660),
.A2(n_3453),
.B1(n_3454),
.B2(n_3449),
.Y(n_4043)
);

NOR2xp33_ASAP7_75t_R g4044 ( 
.A(n_3662),
.B(n_3210),
.Y(n_4044)
);

OR2x6_ASAP7_75t_SL g4045 ( 
.A(n_3909),
.B(n_3385),
.Y(n_4045)
);

BUFx4_ASAP7_75t_SL g4046 ( 
.A(n_3831),
.Y(n_4046)
);

NAND2xp5_ASAP7_75t_SL g4047 ( 
.A(n_3975),
.B(n_3414),
.Y(n_4047)
);

NAND2xp5_ASAP7_75t_L g4048 ( 
.A(n_3719),
.B(n_2938),
.Y(n_4048)
);

NAND2xp5_ASAP7_75t_SL g4049 ( 
.A(n_3555),
.B(n_3013),
.Y(n_4049)
);

AND2x2_ASAP7_75t_L g4050 ( 
.A(n_3511),
.B(n_3039),
.Y(n_4050)
);

NAND2xp5_ASAP7_75t_SL g4051 ( 
.A(n_3733),
.B(n_3013),
.Y(n_4051)
);

NAND3xp33_ASAP7_75t_L g4052 ( 
.A(n_3786),
.B(n_3863),
.C(n_3858),
.Y(n_4052)
);

NAND2xp5_ASAP7_75t_SL g4053 ( 
.A(n_3741),
.B(n_3016),
.Y(n_4053)
);

OAI22xp5_ASAP7_75t_L g4054 ( 
.A1(n_3903),
.A2(n_3451),
.B1(n_3443),
.B2(n_3407),
.Y(n_4054)
);

OAI21x1_ASAP7_75t_L g4055 ( 
.A1(n_3545),
.A2(n_3198),
.B(n_3188),
.Y(n_4055)
);

NAND2xp5_ASAP7_75t_SL g4056 ( 
.A(n_3804),
.B(n_3016),
.Y(n_4056)
);

OA21x2_ASAP7_75t_L g4057 ( 
.A1(n_3959),
.A2(n_3169),
.B(n_3229),
.Y(n_4057)
);

O2A1O1Ixp5_ASAP7_75t_L g4058 ( 
.A1(n_3467),
.A2(n_3190),
.B(n_3098),
.C(n_3422),
.Y(n_4058)
);

O2A1O1Ixp33_ASAP7_75t_L g4059 ( 
.A1(n_3841),
.A2(n_3428),
.B(n_2872),
.C(n_2875),
.Y(n_4059)
);

A2O1A1Ixp33_ASAP7_75t_L g4060 ( 
.A1(n_3468),
.A2(n_3291),
.B(n_3308),
.C(n_3296),
.Y(n_4060)
);

BUFx2_ASAP7_75t_L g4061 ( 
.A(n_3903),
.Y(n_4061)
);

OAI22xp5_ASAP7_75t_L g4062 ( 
.A1(n_3551),
.A2(n_3348),
.B1(n_3353),
.B2(n_3343),
.Y(n_4062)
);

AOI21xp5_ASAP7_75t_L g4063 ( 
.A1(n_3790),
.A2(n_3183),
.B(n_3207),
.Y(n_4063)
);

AOI221xp5_ASAP7_75t_L g4064 ( 
.A1(n_3627),
.A2(n_3651),
.B1(n_3796),
.B2(n_3731),
.C(n_4011),
.Y(n_4064)
);

NAND2xp5_ASAP7_75t_L g4065 ( 
.A(n_3743),
.B(n_3017),
.Y(n_4065)
);

NAND2xp5_ASAP7_75t_L g4066 ( 
.A(n_3754),
.B(n_3018),
.Y(n_4066)
);

OR2x6_ASAP7_75t_L g4067 ( 
.A(n_3831),
.B(n_3185),
.Y(n_4067)
);

NAND2xp5_ASAP7_75t_SL g4068 ( 
.A(n_3816),
.B(n_3243),
.Y(n_4068)
);

CKINVDCx16_ASAP7_75t_R g4069 ( 
.A(n_3991),
.Y(n_4069)
);

A2O1A1Ixp33_ASAP7_75t_L g4070 ( 
.A1(n_3513),
.A2(n_3315),
.B(n_3322),
.C(n_3309),
.Y(n_4070)
);

INVx1_ASAP7_75t_L g4071 ( 
.A(n_3475),
.Y(n_4071)
);

AND2x6_ASAP7_75t_L g4072 ( 
.A(n_3499),
.B(n_2947),
.Y(n_4072)
);

INVx1_ASAP7_75t_SL g4073 ( 
.A(n_3543),
.Y(n_4073)
);

AOI21xp5_ASAP7_75t_L g4074 ( 
.A1(n_3502),
.A2(n_3983),
.B(n_3976),
.Y(n_4074)
);

AOI22xp33_ASAP7_75t_L g4075 ( 
.A1(n_3692),
.A2(n_3340),
.B1(n_3370),
.B2(n_3338),
.Y(n_4075)
);

OAI22xp5_ASAP7_75t_L g4076 ( 
.A1(n_3558),
.A2(n_3389),
.B1(n_3394),
.B2(n_3372),
.Y(n_4076)
);

BUFx6f_ASAP7_75t_L g4077 ( 
.A(n_3465),
.Y(n_4077)
);

AND2x2_ASAP7_75t_L g4078 ( 
.A(n_3590),
.B(n_3406),
.Y(n_4078)
);

BUFx8_ASAP7_75t_L g4079 ( 
.A(n_3597),
.Y(n_4079)
);

HB1xp67_ASAP7_75t_L g4080 ( 
.A(n_3481),
.Y(n_4080)
);

INVxp67_ASAP7_75t_L g4081 ( 
.A(n_3578),
.Y(n_4081)
);

OAI22xp5_ASAP7_75t_L g4082 ( 
.A1(n_3600),
.A2(n_3419),
.B1(n_3238),
.B2(n_3240),
.Y(n_4082)
);

BUFx3_ASAP7_75t_L g4083 ( 
.A(n_3617),
.Y(n_4083)
);

INVx3_ASAP7_75t_L g4084 ( 
.A(n_3816),
.Y(n_4084)
);

NAND2xp5_ASAP7_75t_SL g4085 ( 
.A(n_3912),
.B(n_2976),
.Y(n_4085)
);

NAND2xp5_ASAP7_75t_SL g4086 ( 
.A(n_3912),
.B(n_2976),
.Y(n_4086)
);

CKINVDCx5p33_ASAP7_75t_R g4087 ( 
.A(n_3496),
.Y(n_4087)
);

OR2x2_ASAP7_75t_L g4088 ( 
.A(n_3480),
.B(n_3231),
.Y(n_4088)
);

INVx2_ASAP7_75t_L g4089 ( 
.A(n_3507),
.Y(n_4089)
);

INVx1_ASAP7_75t_L g4090 ( 
.A(n_3485),
.Y(n_4090)
);

HB1xp67_ASAP7_75t_L g4091 ( 
.A(n_3610),
.Y(n_4091)
);

INVx2_ASAP7_75t_SL g4092 ( 
.A(n_3604),
.Y(n_4092)
);

AOI22xp5_ASAP7_75t_L g4093 ( 
.A1(n_3800),
.A2(n_3196),
.B1(n_2910),
.B2(n_3032),
.Y(n_4093)
);

OAI22xp5_ASAP7_75t_L g4094 ( 
.A1(n_3600),
.A2(n_3242),
.B1(n_3206),
.B2(n_2915),
.Y(n_4094)
);

BUFx2_ASAP7_75t_L g4095 ( 
.A(n_3876),
.Y(n_4095)
);

NAND2xp5_ASAP7_75t_SL g4096 ( 
.A(n_4008),
.B(n_3253),
.Y(n_4096)
);

BUFx12f_ASAP7_75t_L g4097 ( 
.A(n_3767),
.Y(n_4097)
);

NOR2xp33_ASAP7_75t_L g4098 ( 
.A(n_3690),
.B(n_3010),
.Y(n_4098)
);

AOI21xp5_ASAP7_75t_L g4099 ( 
.A1(n_3599),
.A2(n_3111),
.B(n_3104),
.Y(n_4099)
);

AOI21xp5_ASAP7_75t_L g4100 ( 
.A1(n_3459),
.A2(n_3119),
.B(n_3115),
.Y(n_4100)
);

O2A1O1Ixp33_ASAP7_75t_L g4101 ( 
.A1(n_3488),
.A2(n_3049),
.B(n_2933),
.C(n_2935),
.Y(n_4101)
);

NAND2xp33_ASAP7_75t_SL g4102 ( 
.A(n_4008),
.B(n_3193),
.Y(n_4102)
);

INVx1_ASAP7_75t_L g4103 ( 
.A(n_3504),
.Y(n_4103)
);

NOR2xp33_ASAP7_75t_L g4104 ( 
.A(n_3936),
.B(n_2877),
.Y(n_4104)
);

INVx3_ASAP7_75t_SL g4105 ( 
.A(n_3767),
.Y(n_4105)
);

NAND2xp5_ASAP7_75t_L g4106 ( 
.A(n_3757),
.B(n_2802),
.Y(n_4106)
);

AND2x2_ASAP7_75t_L g4107 ( 
.A(n_3773),
.B(n_3205),
.Y(n_4107)
);

A2O1A1Ixp33_ASAP7_75t_L g4108 ( 
.A1(n_3563),
.A2(n_3571),
.B(n_3487),
.C(n_3501),
.Y(n_4108)
);

INVx1_ASAP7_75t_L g4109 ( 
.A(n_3544),
.Y(n_4109)
);

NAND2xp5_ASAP7_75t_L g4110 ( 
.A(n_3805),
.B(n_2804),
.Y(n_4110)
);

OAI21x1_ASAP7_75t_L g4111 ( 
.A1(n_3489),
.A2(n_3225),
.B(n_3138),
.Y(n_4111)
);

NAND2xp5_ASAP7_75t_L g4112 ( 
.A(n_3810),
.B(n_3121),
.Y(n_4112)
);

NAND2xp5_ASAP7_75t_L g4113 ( 
.A(n_3814),
.B(n_2983),
.Y(n_4113)
);

BUFx2_ASAP7_75t_L g4114 ( 
.A(n_3897),
.Y(n_4114)
);

OAI22xp5_ASAP7_75t_L g4115 ( 
.A1(n_3763),
.A2(n_3026),
.B1(n_3053),
.B2(n_3046),
.Y(n_4115)
);

AOI21xp5_ASAP7_75t_L g4116 ( 
.A1(n_4019),
.A2(n_3177),
.B(n_3175),
.Y(n_4116)
);

INVx1_ASAP7_75t_L g4117 ( 
.A(n_3570),
.Y(n_4117)
);

AOI21xp5_ASAP7_75t_L g4118 ( 
.A1(n_3594),
.A2(n_3615),
.B(n_4004),
.Y(n_4118)
);

OAI22xp5_ASAP7_75t_L g4119 ( 
.A1(n_3763),
.A2(n_3848),
.B1(n_3477),
.B2(n_3787),
.Y(n_4119)
);

NAND2xp5_ASAP7_75t_L g4120 ( 
.A(n_3823),
.B(n_3165),
.Y(n_4120)
);

INVx2_ASAP7_75t_L g4121 ( 
.A(n_3515),
.Y(n_4121)
);

NOR2xp33_ASAP7_75t_L g4122 ( 
.A(n_3636),
.B(n_2844),
.Y(n_4122)
);

NAND2xp5_ASAP7_75t_SL g4123 ( 
.A(n_3483),
.B(n_3253),
.Y(n_4123)
);

INVx1_ASAP7_75t_L g4124 ( 
.A(n_3576),
.Y(n_4124)
);

AOI21xp5_ASAP7_75t_L g4125 ( 
.A1(n_4012),
.A2(n_3135),
.B(n_3163),
.Y(n_4125)
);

AOI21xp5_ASAP7_75t_L g4126 ( 
.A1(n_3856),
.A2(n_3003),
.B(n_2906),
.Y(n_4126)
);

NAND2xp5_ASAP7_75t_SL g4127 ( 
.A(n_3483),
.B(n_3634),
.Y(n_4127)
);

CKINVDCx11_ASAP7_75t_R g4128 ( 
.A(n_3904),
.Y(n_4128)
);

BUFx12f_ASAP7_75t_L g4129 ( 
.A(n_3982),
.Y(n_4129)
);

NOR2xp33_ASAP7_75t_L g4130 ( 
.A(n_3539),
.B(n_2926),
.Y(n_4130)
);

NOR2xp33_ASAP7_75t_L g4131 ( 
.A(n_3663),
.B(n_2971),
.Y(n_4131)
);

INVx2_ASAP7_75t_L g4132 ( 
.A(n_3526),
.Y(n_4132)
);

NAND2xp5_ASAP7_75t_L g4133 ( 
.A(n_3884),
.B(n_3091),
.Y(n_4133)
);

INVx1_ASAP7_75t_L g4134 ( 
.A(n_3582),
.Y(n_4134)
);

A2O1A1Ixp33_ASAP7_75t_L g4135 ( 
.A1(n_3657),
.A2(n_3197),
.B(n_3200),
.C(n_3100),
.Y(n_4135)
);

AOI21xp5_ASAP7_75t_L g4136 ( 
.A1(n_3885),
.A2(n_2920),
.B(n_2869),
.Y(n_4136)
);

O2A1O1Ixp33_ASAP7_75t_L g4137 ( 
.A1(n_3470),
.A2(n_2943),
.B(n_2957),
.C(n_3202),
.Y(n_4137)
);

INVx2_ASAP7_75t_SL g4138 ( 
.A(n_3803),
.Y(n_4138)
);

A2O1A1Ixp33_ASAP7_75t_L g4139 ( 
.A1(n_3538),
.A2(n_3189),
.B(n_3086),
.C(n_3195),
.Y(n_4139)
);

NOR2xp33_ASAP7_75t_L g4140 ( 
.A(n_3516),
.B(n_2898),
.Y(n_4140)
);

NOR3xp33_ASAP7_75t_SL g4141 ( 
.A(n_3614),
.B(n_3166),
.C(n_3009),
.Y(n_4141)
);

INVx2_ASAP7_75t_L g4142 ( 
.A(n_3542),
.Y(n_4142)
);

NOR2xp33_ASAP7_75t_L g4143 ( 
.A(n_3466),
.B(n_2946),
.Y(n_4143)
);

INVx3_ASAP7_75t_L g4144 ( 
.A(n_3530),
.Y(n_4144)
);

OAI22xp5_ASAP7_75t_L g4145 ( 
.A1(n_3848),
.A2(n_3149),
.B1(n_3151),
.B2(n_3145),
.Y(n_4145)
);

AND2x2_ASAP7_75t_L g4146 ( 
.A(n_3674),
.B(n_3214),
.Y(n_4146)
);

A2O1A1Ixp33_ASAP7_75t_L g4147 ( 
.A1(n_3562),
.A2(n_3417),
.B(n_3450),
.C(n_3269),
.Y(n_4147)
);

BUFx12f_ASAP7_75t_L g4148 ( 
.A(n_3708),
.Y(n_4148)
);

INVx1_ASAP7_75t_L g4149 ( 
.A(n_3601),
.Y(n_4149)
);

A2O1A1Ixp33_ASAP7_75t_L g4150 ( 
.A1(n_3573),
.A2(n_3417),
.B(n_3450),
.C(n_3269),
.Y(n_4150)
);

AOI21xp5_ASAP7_75t_L g4151 ( 
.A1(n_3941),
.A2(n_2942),
.B(n_3221),
.Y(n_4151)
);

NAND2xp5_ASAP7_75t_L g4152 ( 
.A(n_3996),
.B(n_3105),
.Y(n_4152)
);

INVx1_ASAP7_75t_L g4153 ( 
.A(n_3606),
.Y(n_4153)
);

INVx1_ASAP7_75t_L g4154 ( 
.A(n_3616),
.Y(n_4154)
);

AND2x2_ASAP7_75t_L g4155 ( 
.A(n_4000),
.B(n_3110),
.Y(n_4155)
);

AND2x4_ASAP7_75t_L g4156 ( 
.A(n_3530),
.B(n_3211),
.Y(n_4156)
);

INVx5_ASAP7_75t_L g4157 ( 
.A(n_3465),
.Y(n_4157)
);

NAND2xp5_ASAP7_75t_SL g4158 ( 
.A(n_3701),
.B(n_3164),
.Y(n_4158)
);

O2A1O1Ixp33_ASAP7_75t_SL g4159 ( 
.A1(n_3706),
.A2(n_2902),
.B(n_3222),
.C(n_3220),
.Y(n_4159)
);

AOI21xp5_ASAP7_75t_L g4160 ( 
.A1(n_4005),
.A2(n_3224),
.B(n_3027),
.Y(n_4160)
);

AOI21xp5_ASAP7_75t_L g4161 ( 
.A1(n_4007),
.A2(n_3014),
.B(n_3176),
.Y(n_4161)
);

AOI22xp5_ASAP7_75t_L g4162 ( 
.A1(n_3944),
.A2(n_3001),
.B1(n_2988),
.B2(n_2977),
.Y(n_4162)
);

INVx1_ASAP7_75t_SL g4163 ( 
.A(n_3926),
.Y(n_4163)
);

INVx2_ASAP7_75t_L g4164 ( 
.A(n_3550),
.Y(n_4164)
);

OAI22xp5_ASAP7_75t_L g4165 ( 
.A1(n_3537),
.A2(n_3174),
.B1(n_3161),
.B2(n_3136),
.Y(n_4165)
);

INVx1_ASAP7_75t_L g4166 ( 
.A(n_3607),
.Y(n_4166)
);

OAI22xp5_ASAP7_75t_L g4167 ( 
.A1(n_3777),
.A2(n_3139),
.B1(n_3134),
.B2(n_3144),
.Y(n_4167)
);

INVxp67_ASAP7_75t_L g4168 ( 
.A(n_3569),
.Y(n_4168)
);

OAI22xp5_ASAP7_75t_SL g4169 ( 
.A1(n_3774),
.A2(n_3154),
.B1(n_3137),
.B2(n_3133),
.Y(n_4169)
);

NOR2xp67_ASAP7_75t_SL g4170 ( 
.A(n_3575),
.B(n_3068),
.Y(n_4170)
);

NAND3xp33_ASAP7_75t_L g4171 ( 
.A(n_3829),
.B(n_3191),
.C(n_3069),
.Y(n_4171)
);

AOI21xp5_ASAP7_75t_L g4172 ( 
.A1(n_3842),
.A2(n_3057),
.B(n_3083),
.Y(n_4172)
);

AOI21xp5_ASAP7_75t_L g4173 ( 
.A1(n_3846),
.A2(n_3140),
.B(n_3106),
.Y(n_4173)
);

AOI21xp5_ASAP7_75t_L g4174 ( 
.A1(n_3881),
.A2(n_3096),
.B(n_3129),
.Y(n_4174)
);

INVx5_ASAP7_75t_L g4175 ( 
.A(n_3465),
.Y(n_4175)
);

AOI21xp5_ASAP7_75t_L g4176 ( 
.A1(n_3911),
.A2(n_3132),
.B(n_3113),
.Y(n_4176)
);

INVx2_ASAP7_75t_L g4177 ( 
.A(n_3564),
.Y(n_4177)
);

OR2x6_ASAP7_75t_L g4178 ( 
.A(n_3575),
.B(n_3164),
.Y(n_4178)
);

INVx2_ASAP7_75t_SL g4179 ( 
.A(n_3839),
.Y(n_4179)
);

AOI22xp33_ASAP7_75t_L g4180 ( 
.A1(n_3822),
.A2(n_3162),
.B1(n_3164),
.B2(n_3223),
.Y(n_4180)
);

INVx2_ASAP7_75t_L g4181 ( 
.A(n_3862),
.Y(n_4181)
);

INVx1_ASAP7_75t_L g4182 ( 
.A(n_3681),
.Y(n_4182)
);

INVx1_ASAP7_75t_L g4183 ( 
.A(n_3689),
.Y(n_4183)
);

INVx2_ASAP7_75t_SL g4184 ( 
.A(n_3722),
.Y(n_4184)
);

AND2x4_ASAP7_75t_L g4185 ( 
.A(n_3608),
.B(n_3162),
.Y(n_4185)
);

BUFx6f_ASAP7_75t_L g4186 ( 
.A(n_3492),
.Y(n_4186)
);

INVx1_ASAP7_75t_L g4187 ( 
.A(n_3698),
.Y(n_4187)
);

OAI22xp5_ASAP7_75t_L g4188 ( 
.A1(n_3732),
.A2(n_3577),
.B1(n_3725),
.B2(n_3499),
.Y(n_4188)
);

O2A1O1Ixp33_ASAP7_75t_L g4189 ( 
.A1(n_3583),
.A2(n_566),
.B(n_567),
.C(n_565),
.Y(n_4189)
);

NAND2xp5_ASAP7_75t_L g4190 ( 
.A(n_3547),
.B(n_565),
.Y(n_4190)
);

NAND2xp5_ASAP7_75t_L g4191 ( 
.A(n_3947),
.B(n_566),
.Y(n_4191)
);

INVx1_ASAP7_75t_L g4192 ( 
.A(n_3707),
.Y(n_4192)
);

OR2x2_ASAP7_75t_L g4193 ( 
.A(n_3717),
.B(n_566),
.Y(n_4193)
);

OAI22xp5_ASAP7_75t_L g4194 ( 
.A1(n_3587),
.A2(n_568),
.B1(n_569),
.B2(n_567),
.Y(n_4194)
);

OAI22xp5_ASAP7_75t_L g4195 ( 
.A1(n_3961),
.A2(n_568),
.B1(n_569),
.B2(n_567),
.Y(n_4195)
);

NOR2xp33_ASAP7_75t_L g4196 ( 
.A(n_3957),
.B(n_568),
.Y(n_4196)
);

INVxp67_ASAP7_75t_L g4197 ( 
.A(n_3673),
.Y(n_4197)
);

NAND2x1p5_ASAP7_75t_L g4198 ( 
.A(n_3613),
.B(n_574),
.Y(n_4198)
);

BUFx4f_ASAP7_75t_L g4199 ( 
.A(n_3834),
.Y(n_4199)
);

NOR2xp33_ASAP7_75t_L g4200 ( 
.A(n_3664),
.B(n_570),
.Y(n_4200)
);

AND2x2_ASAP7_75t_L g4201 ( 
.A(n_3806),
.B(n_1103),
.Y(n_4201)
);

OAI22xp5_ASAP7_75t_L g4202 ( 
.A1(n_3484),
.A2(n_571),
.B1(n_572),
.B2(n_570),
.Y(n_4202)
);

O2A1O1Ixp33_ASAP7_75t_SL g4203 ( 
.A1(n_3624),
.A2(n_1104),
.B(n_1106),
.C(n_1103),
.Y(n_4203)
);

OAI21x1_ASAP7_75t_L g4204 ( 
.A1(n_3584),
.A2(n_571),
.B(n_570),
.Y(n_4204)
);

INVx2_ASAP7_75t_L g4205 ( 
.A(n_3871),
.Y(n_4205)
);

BUFx6f_ASAP7_75t_L g4206 ( 
.A(n_3492),
.Y(n_4206)
);

BUFx3_ASAP7_75t_L g4207 ( 
.A(n_3567),
.Y(n_4207)
);

NOR2xp33_ASAP7_75t_R g4208 ( 
.A(n_3613),
.B(n_571),
.Y(n_4208)
);

INVx1_ASAP7_75t_SL g4209 ( 
.A(n_3965),
.Y(n_4209)
);

NAND2xp5_ASAP7_75t_L g4210 ( 
.A(n_3462),
.B(n_572),
.Y(n_4210)
);

INVx1_ASAP7_75t_L g4211 ( 
.A(n_3906),
.Y(n_4211)
);

AND2x2_ASAP7_75t_L g4212 ( 
.A(n_3886),
.B(n_1107),
.Y(n_4212)
);

NAND2xp5_ASAP7_75t_L g4213 ( 
.A(n_3740),
.B(n_572),
.Y(n_4213)
);

AND2x4_ASAP7_75t_L g4214 ( 
.A(n_3608),
.B(n_573),
.Y(n_4214)
);

NOR2xp33_ASAP7_75t_L g4215 ( 
.A(n_3631),
.B(n_573),
.Y(n_4215)
);

OAI22xp5_ASAP7_75t_L g4216 ( 
.A1(n_3498),
.A2(n_574),
.B1(n_575),
.B2(n_573),
.Y(n_4216)
);

OAI22xp5_ASAP7_75t_SL g4217 ( 
.A1(n_3834),
.A2(n_576),
.B1(n_577),
.B2(n_575),
.Y(n_4217)
);

OR2x6_ASAP7_75t_L g4218 ( 
.A(n_3905),
.B(n_575),
.Y(n_4218)
);

NOR3xp33_ASAP7_75t_L g4219 ( 
.A(n_3533),
.B(n_577),
.C(n_576),
.Y(n_4219)
);

INVx2_ASAP7_75t_L g4220 ( 
.A(n_3887),
.Y(n_4220)
);

INVx2_ASAP7_75t_L g4221 ( 
.A(n_3922),
.Y(n_4221)
);

NAND2xp5_ASAP7_75t_L g4222 ( 
.A(n_3472),
.B(n_576),
.Y(n_4222)
);

AOI21xp5_ASAP7_75t_L g4223 ( 
.A1(n_3937),
.A2(n_3968),
.B(n_3977),
.Y(n_4223)
);

NAND2xp33_ASAP7_75t_SL g4224 ( 
.A(n_3847),
.B(n_3541),
.Y(n_4224)
);

AOI22xp5_ASAP7_75t_L g4225 ( 
.A1(n_3685),
.A2(n_578),
.B1(n_579),
.B2(n_577),
.Y(n_4225)
);

A2O1A1Ixp33_ASAP7_75t_L g4226 ( 
.A1(n_3591),
.A2(n_579),
.B(n_580),
.C(n_578),
.Y(n_4226)
);

INVx1_ASAP7_75t_SL g4227 ( 
.A(n_3980),
.Y(n_4227)
);

INVx1_ASAP7_75t_L g4228 ( 
.A(n_3950),
.Y(n_4228)
);

OAI22xp5_ASAP7_75t_L g4229 ( 
.A1(n_3744),
.A2(n_580),
.B1(n_581),
.B2(n_579),
.Y(n_4229)
);

INVxp67_ASAP7_75t_SL g4230 ( 
.A(n_3700),
.Y(n_4230)
);

OR2x2_ASAP7_75t_L g4231 ( 
.A(n_3984),
.B(n_580),
.Y(n_4231)
);

O2A1O1Ixp33_ASAP7_75t_L g4232 ( 
.A1(n_3522),
.A2(n_582),
.B(n_583),
.C(n_581),
.Y(n_4232)
);

NOR2xp33_ASAP7_75t_L g4233 ( 
.A(n_3460),
.B(n_582),
.Y(n_4233)
);

BUFx2_ASAP7_75t_L g4234 ( 
.A(n_3592),
.Y(n_4234)
);

AND2x2_ASAP7_75t_L g4235 ( 
.A(n_3913),
.B(n_1100),
.Y(n_4235)
);

INVx4_ASAP7_75t_L g4236 ( 
.A(n_3492),
.Y(n_4236)
);

NAND2xp5_ASAP7_75t_SL g4237 ( 
.A(n_3890),
.B(n_583),
.Y(n_4237)
);

OAI22xp5_ASAP7_75t_SL g4238 ( 
.A1(n_3715),
.A2(n_3851),
.B1(n_3494),
.B2(n_3677),
.Y(n_4238)
);

AOI21xp5_ASAP7_75t_L g4239 ( 
.A1(n_3978),
.A2(n_584),
.B(n_583),
.Y(n_4239)
);

O2A1O1Ixp33_ASAP7_75t_L g4240 ( 
.A1(n_3528),
.A2(n_585),
.B(n_586),
.C(n_584),
.Y(n_4240)
);

BUFx2_ASAP7_75t_L g4241 ( 
.A(n_3704),
.Y(n_4241)
);

NAND2xp5_ASAP7_75t_L g4242 ( 
.A(n_3789),
.B(n_585),
.Y(n_4242)
);

NOR2xp33_ASAP7_75t_L g4243 ( 
.A(n_3628),
.B(n_586),
.Y(n_4243)
);

NAND2xp5_ASAP7_75t_SL g4244 ( 
.A(n_3473),
.B(n_586),
.Y(n_4244)
);

O2A1O1Ixp33_ASAP7_75t_L g4245 ( 
.A1(n_3497),
.A2(n_588),
.B(n_589),
.C(n_587),
.Y(n_4245)
);

CKINVDCx14_ASAP7_75t_R g4246 ( 
.A(n_3788),
.Y(n_4246)
);

NAND2xp5_ASAP7_75t_L g4247 ( 
.A(n_3864),
.B(n_587),
.Y(n_4247)
);

AOI22xp5_ASAP7_75t_L g4248 ( 
.A1(n_3517),
.A2(n_588),
.B1(n_589),
.B2(n_587),
.Y(n_4248)
);

AND2x2_ASAP7_75t_L g4249 ( 
.A(n_3938),
.B(n_1108),
.Y(n_4249)
);

INVx3_ASAP7_75t_L g4250 ( 
.A(n_3503),
.Y(n_4250)
);

A2O1A1Ixp33_ASAP7_75t_SL g4251 ( 
.A1(n_4006),
.A2(n_68),
.B(n_66),
.C(n_67),
.Y(n_4251)
);

A2O1A1Ixp33_ASAP7_75t_L g4252 ( 
.A1(n_3648),
.A2(n_3687),
.B(n_3727),
.C(n_3825),
.Y(n_4252)
);

HB1xp67_ASAP7_75t_L g4253 ( 
.A(n_3861),
.Y(n_4253)
);

A2O1A1Ixp33_ASAP7_75t_L g4254 ( 
.A1(n_3835),
.A2(n_590),
.B(n_591),
.C(n_589),
.Y(n_4254)
);

AOI21xp5_ASAP7_75t_L g4255 ( 
.A1(n_3981),
.A2(n_591),
.B(n_590),
.Y(n_4255)
);

NAND2xp5_ASAP7_75t_SL g4256 ( 
.A(n_3668),
.B(n_590),
.Y(n_4256)
);

NOR2xp33_ASAP7_75t_R g4257 ( 
.A(n_3671),
.B(n_592),
.Y(n_4257)
);

AOI21xp5_ASAP7_75t_L g4258 ( 
.A1(n_3985),
.A2(n_593),
.B(n_592),
.Y(n_4258)
);

BUFx2_ASAP7_75t_L g4259 ( 
.A(n_3877),
.Y(n_4259)
);

OAI22xp5_ASAP7_75t_L g4260 ( 
.A1(n_3748),
.A2(n_593),
.B1(n_594),
.B2(n_592),
.Y(n_4260)
);

O2A1O1Ixp33_ASAP7_75t_L g4261 ( 
.A1(n_3892),
.A2(n_594),
.B(n_595),
.C(n_593),
.Y(n_4261)
);

AOI22xp33_ASAP7_75t_L g4262 ( 
.A1(n_3967),
.A2(n_596),
.B1(n_597),
.B2(n_595),
.Y(n_4262)
);

AO21x2_ASAP7_75t_L g4263 ( 
.A1(n_3699),
.A2(n_596),
.B(n_595),
.Y(n_4263)
);

NAND2xp5_ASAP7_75t_L g4264 ( 
.A(n_3867),
.B(n_597),
.Y(n_4264)
);

NOR2xp33_ASAP7_75t_L g4265 ( 
.A(n_3548),
.B(n_3889),
.Y(n_4265)
);

OAI21xp5_ASAP7_75t_L g4266 ( 
.A1(n_3807),
.A2(n_598),
.B(n_597),
.Y(n_4266)
);

INVx2_ASAP7_75t_L g4267 ( 
.A(n_3568),
.Y(n_4267)
);

NAND2xp5_ASAP7_75t_L g4268 ( 
.A(n_3797),
.B(n_598),
.Y(n_4268)
);

NAND2xp5_ASAP7_75t_L g4269 ( 
.A(n_3764),
.B(n_599),
.Y(n_4269)
);

O2A1O1Ixp33_ASAP7_75t_L g4270 ( 
.A1(n_3821),
.A2(n_600),
.B(n_601),
.C(n_599),
.Y(n_4270)
);

NAND2xp5_ASAP7_75t_L g4271 ( 
.A(n_3702),
.B(n_599),
.Y(n_4271)
);

O2A1O1Ixp33_ASAP7_75t_L g4272 ( 
.A1(n_3857),
.A2(n_601),
.B(n_602),
.C(n_600),
.Y(n_4272)
);

INVx2_ASAP7_75t_SL g4273 ( 
.A(n_3609),
.Y(n_4273)
);

O2A1O1Ixp33_ASAP7_75t_L g4274 ( 
.A1(n_3680),
.A2(n_601),
.B(n_602),
.C(n_600),
.Y(n_4274)
);

INVx3_ASAP7_75t_L g4275 ( 
.A(n_3503),
.Y(n_4275)
);

NAND2xp5_ASAP7_75t_SL g4276 ( 
.A(n_3503),
.B(n_603),
.Y(n_4276)
);

BUFx6f_ASAP7_75t_L g4277 ( 
.A(n_3521),
.Y(n_4277)
);

INVx3_ASAP7_75t_L g4278 ( 
.A(n_3521),
.Y(n_4278)
);

OAI22x1_ASAP7_75t_L g4279 ( 
.A1(n_4001),
.A2(n_604),
.B1(n_605),
.B2(n_603),
.Y(n_4279)
);

BUFx3_ASAP7_75t_L g4280 ( 
.A(n_3609),
.Y(n_4280)
);

AOI21x1_ASAP7_75t_L g4281 ( 
.A1(n_3675),
.A2(n_604),
.B(n_603),
.Y(n_4281)
);

AND2x2_ASAP7_75t_L g4282 ( 
.A(n_3946),
.B(n_1107),
.Y(n_4282)
);

O2A1O1Ixp33_ASAP7_75t_L g4283 ( 
.A1(n_3843),
.A2(n_605),
.B(n_606),
.C(n_604),
.Y(n_4283)
);

AOI22xp33_ASAP7_75t_L g4284 ( 
.A1(n_3963),
.A2(n_607),
.B1(n_608),
.B2(n_606),
.Y(n_4284)
);

OAI22xp5_ASAP7_75t_L g4285 ( 
.A1(n_3888),
.A2(n_608),
.B1(n_609),
.B2(n_607),
.Y(n_4285)
);

NOR2xp33_ASAP7_75t_L g4286 ( 
.A(n_3696),
.B(n_3713),
.Y(n_4286)
);

NAND2xp5_ASAP7_75t_L g4287 ( 
.A(n_3714),
.B(n_609),
.Y(n_4287)
);

AOI21xp5_ASAP7_75t_L g4288 ( 
.A1(n_3986),
.A2(n_611),
.B(n_610),
.Y(n_4288)
);

AOI21xp5_ASAP7_75t_L g4289 ( 
.A1(n_3993),
.A2(n_612),
.B(n_610),
.Y(n_4289)
);

BUFx2_ASAP7_75t_L g4290 ( 
.A(n_3670),
.Y(n_4290)
);

AND2x4_ASAP7_75t_L g4291 ( 
.A(n_3670),
.B(n_610),
.Y(n_4291)
);

INVx2_ASAP7_75t_L g4292 ( 
.A(n_3586),
.Y(n_4292)
);

O2A1O1Ixp5_ASAP7_75t_L g4293 ( 
.A1(n_3770),
.A2(n_613),
.B(n_614),
.C(n_612),
.Y(n_4293)
);

O2A1O1Ixp33_ASAP7_75t_L g4294 ( 
.A1(n_3457),
.A2(n_613),
.B(n_614),
.C(n_612),
.Y(n_4294)
);

CKINVDCx20_ASAP7_75t_R g4295 ( 
.A(n_3532),
.Y(n_4295)
);

BUFx6f_ASAP7_75t_L g4296 ( 
.A(n_3521),
.Y(n_4296)
);

INVx1_ASAP7_75t_L g4297 ( 
.A(n_3506),
.Y(n_4297)
);

NOR2xp33_ASAP7_75t_L g4298 ( 
.A(n_3458),
.B(n_613),
.Y(n_4298)
);

BUFx2_ASAP7_75t_L g4299 ( 
.A(n_3815),
.Y(n_4299)
);

CKINVDCx5p33_ASAP7_75t_R g4300 ( 
.A(n_3505),
.Y(n_4300)
);

INVx2_ASAP7_75t_SL g4301 ( 
.A(n_3815),
.Y(n_4301)
);

AND2x4_ASAP7_75t_L g4302 ( 
.A(n_3878),
.B(n_614),
.Y(n_4302)
);

CKINVDCx16_ASAP7_75t_R g4303 ( 
.A(n_3574),
.Y(n_4303)
);

BUFx8_ASAP7_75t_L g4304 ( 
.A(n_3969),
.Y(n_4304)
);

INVx2_ASAP7_75t_SL g4305 ( 
.A(n_3878),
.Y(n_4305)
);

INVx1_ASAP7_75t_L g4306 ( 
.A(n_3509),
.Y(n_4306)
);

OAI22xp5_ASAP7_75t_L g4307 ( 
.A1(n_3742),
.A2(n_616),
.B1(n_617),
.B2(n_615),
.Y(n_4307)
);

AOI21xp5_ASAP7_75t_L g4308 ( 
.A1(n_3994),
.A2(n_616),
.B(n_615),
.Y(n_4308)
);

BUFx3_ASAP7_75t_L g4309 ( 
.A(n_3882),
.Y(n_4309)
);

INVx2_ASAP7_75t_L g4310 ( 
.A(n_3612),
.Y(n_4310)
);

NAND2xp5_ASAP7_75t_L g4311 ( 
.A(n_3896),
.B(n_615),
.Y(n_4311)
);

AOI22xp33_ASAP7_75t_L g4312 ( 
.A1(n_3666),
.A2(n_618),
.B1(n_619),
.B2(n_616),
.Y(n_4312)
);

AND2x2_ASAP7_75t_L g4313 ( 
.A(n_4020),
.B(n_1104),
.Y(n_4313)
);

INVx1_ASAP7_75t_SL g4314 ( 
.A(n_3527),
.Y(n_4314)
);

NAND2xp5_ASAP7_75t_SL g4315 ( 
.A(n_3527),
.B(n_618),
.Y(n_4315)
);

NAND2xp5_ASAP7_75t_SL g4316 ( 
.A(n_3527),
.B(n_619),
.Y(n_4316)
);

INVx2_ASAP7_75t_SL g4317 ( 
.A(n_3882),
.Y(n_4317)
);

OAI22xp5_ASAP7_75t_L g4318 ( 
.A1(n_3998),
.A2(n_620),
.B1(n_622),
.B2(n_619),
.Y(n_4318)
);

INVx3_ASAP7_75t_L g4319 ( 
.A(n_3581),
.Y(n_4319)
);

INVx2_ASAP7_75t_L g4320 ( 
.A(n_3619),
.Y(n_4320)
);

INVx4_ASAP7_75t_L g4321 ( 
.A(n_3581),
.Y(n_4321)
);

NAND2xp5_ASAP7_75t_L g4322 ( 
.A(n_3899),
.B(n_620),
.Y(n_4322)
);

AOI21xp5_ASAP7_75t_L g4323 ( 
.A1(n_4002),
.A2(n_623),
.B(n_622),
.Y(n_4323)
);

NAND2xp5_ASAP7_75t_L g4324 ( 
.A(n_3910),
.B(n_623),
.Y(n_4324)
);

AOI21xp5_ASAP7_75t_L g4325 ( 
.A1(n_4003),
.A2(n_625),
.B(n_623),
.Y(n_4325)
);

INVx2_ASAP7_75t_L g4326 ( 
.A(n_3635),
.Y(n_4326)
);

INVx2_ASAP7_75t_L g4327 ( 
.A(n_3656),
.Y(n_4327)
);

CKINVDCx20_ASAP7_75t_R g4328 ( 
.A(n_3491),
.Y(n_4328)
);

O2A1O1Ixp33_ASAP7_75t_L g4329 ( 
.A1(n_3874),
.A2(n_3783),
.B(n_3830),
.C(n_3811),
.Y(n_4329)
);

O2A1O1Ixp5_ASAP7_75t_L g4330 ( 
.A1(n_3630),
.A2(n_627),
.B(n_628),
.C(n_625),
.Y(n_4330)
);

BUFx6f_ASAP7_75t_L g4331 ( 
.A(n_3581),
.Y(n_4331)
);

AOI21xp5_ASAP7_75t_L g4332 ( 
.A1(n_4010),
.A2(n_627),
.B(n_625),
.Y(n_4332)
);

NAND2xp5_ASAP7_75t_SL g4333 ( 
.A(n_3620),
.B(n_627),
.Y(n_4333)
);

AOI21xp5_ASAP7_75t_L g4334 ( 
.A1(n_4013),
.A2(n_629),
.B(n_628),
.Y(n_4334)
);

INVx2_ASAP7_75t_L g4335 ( 
.A(n_3697),
.Y(n_4335)
);

O2A1O1Ixp33_ASAP7_75t_L g4336 ( 
.A1(n_3840),
.A2(n_3849),
.B(n_3837),
.C(n_3916),
.Y(n_4336)
);

AND2x2_ASAP7_75t_L g4337 ( 
.A(n_3557),
.B(n_1115),
.Y(n_4337)
);

INVx2_ASAP7_75t_SL g4338 ( 
.A(n_3907),
.Y(n_4338)
);

AOI21xp5_ASAP7_75t_L g4339 ( 
.A1(n_3469),
.A2(n_630),
.B(n_628),
.Y(n_4339)
);

NAND2x1_ASAP7_75t_L g4340 ( 
.A(n_3620),
.B(n_630),
.Y(n_4340)
);

OAI22xp5_ASAP7_75t_L g4341 ( 
.A1(n_3850),
.A2(n_632),
.B1(n_633),
.B2(n_630),
.Y(n_4341)
);

INVx1_ASAP7_75t_L g4342 ( 
.A(n_3510),
.Y(n_4342)
);

NAND2xp5_ASAP7_75t_SL g4343 ( 
.A(n_3620),
.B(n_632),
.Y(n_4343)
);

NAND2x1p5_ASAP7_75t_L g4344 ( 
.A(n_3629),
.B(n_636),
.Y(n_4344)
);

O2A1O1Ixp33_ASAP7_75t_L g4345 ( 
.A1(n_3917),
.A2(n_633),
.B(n_634),
.C(n_632),
.Y(n_4345)
);

NAND2xp5_ASAP7_75t_L g4346 ( 
.A(n_3716),
.B(n_3734),
.Y(n_4346)
);

INVx5_ASAP7_75t_L g4347 ( 
.A(n_3629),
.Y(n_4347)
);

INVxp67_ASAP7_75t_SL g4348 ( 
.A(n_3629),
.Y(n_4348)
);

BUFx6f_ASAP7_75t_L g4349 ( 
.A(n_3639),
.Y(n_4349)
);

CKINVDCx5p33_ASAP7_75t_R g4350 ( 
.A(n_3525),
.Y(n_4350)
);

AOI21xp5_ASAP7_75t_L g4351 ( 
.A1(n_3471),
.A2(n_634),
.B(n_633),
.Y(n_4351)
);

OAI22xp5_ASAP7_75t_L g4352 ( 
.A1(n_3865),
.A2(n_635),
.B1(n_636),
.B2(n_634),
.Y(n_4352)
);

OR2x6_ASAP7_75t_L g4353 ( 
.A(n_3588),
.B(n_3540),
.Y(n_4353)
);

OAI22xp5_ASAP7_75t_L g4354 ( 
.A1(n_3866),
.A2(n_637),
.B1(n_638),
.B2(n_635),
.Y(n_4354)
);

NOR2xp67_ASAP7_75t_R g4355 ( 
.A(n_3495),
.B(n_638),
.Y(n_4355)
);

INVx2_ASAP7_75t_SL g4356 ( 
.A(n_3907),
.Y(n_4356)
);

NAND3xp33_ASAP7_75t_SL g4357 ( 
.A(n_3559),
.B(n_66),
.C(n_67),
.Y(n_4357)
);

NAND2xp5_ASAP7_75t_L g4358 ( 
.A(n_3809),
.B(n_639),
.Y(n_4358)
);

INVxp67_ASAP7_75t_L g4359 ( 
.A(n_3546),
.Y(n_4359)
);

A2O1A1Ixp33_ASAP7_75t_L g4360 ( 
.A1(n_3875),
.A2(n_640),
.B(n_641),
.C(n_639),
.Y(n_4360)
);

BUFx6f_ASAP7_75t_L g4361 ( 
.A(n_3639),
.Y(n_4361)
);

OAI22xp5_ASAP7_75t_L g4362 ( 
.A1(n_3934),
.A2(n_640),
.B1(n_641),
.B2(n_639),
.Y(n_4362)
);

OAI22xp5_ASAP7_75t_L g4363 ( 
.A1(n_3954),
.A2(n_642),
.B1(n_643),
.B2(n_640),
.Y(n_4363)
);

INVx2_ASAP7_75t_L g4364 ( 
.A(n_3721),
.Y(n_4364)
);

A2O1A1Ixp33_ASAP7_75t_L g4365 ( 
.A1(n_3971),
.A2(n_644),
.B(n_645),
.C(n_643),
.Y(n_4365)
);

OAI21x1_ASAP7_75t_L g4366 ( 
.A1(n_4023),
.A2(n_644),
.B(n_643),
.Y(n_4366)
);

AOI21xp5_ASAP7_75t_L g4367 ( 
.A1(n_3478),
.A2(n_645),
.B(n_644),
.Y(n_4367)
);

NOR2xp33_ASAP7_75t_R g4368 ( 
.A(n_3919),
.B(n_645),
.Y(n_4368)
);

NOR2xp33_ASAP7_75t_L g4369 ( 
.A(n_3826),
.B(n_646),
.Y(n_4369)
);

NAND2xp33_ASAP7_75t_SL g4370 ( 
.A(n_3565),
.B(n_1115),
.Y(n_4370)
);

INVx1_ASAP7_75t_L g4371 ( 
.A(n_3512),
.Y(n_4371)
);

OAI22xp5_ASAP7_75t_L g4372 ( 
.A1(n_3987),
.A2(n_647),
.B1(n_648),
.B2(n_646),
.Y(n_4372)
);

AOI21xp5_ASAP7_75t_L g4373 ( 
.A1(n_3752),
.A2(n_647),
.B(n_646),
.Y(n_4373)
);

INVx2_ASAP7_75t_SL g4374 ( 
.A(n_3919),
.Y(n_4374)
);

HB1xp67_ASAP7_75t_L g4375 ( 
.A(n_3745),
.Y(n_4375)
);

CKINVDCx5p33_ASAP7_75t_R g4376 ( 
.A(n_3914),
.Y(n_4376)
);

AND2x4_ASAP7_75t_L g4377 ( 
.A(n_3933),
.B(n_647),
.Y(n_4377)
);

INVx2_ASAP7_75t_L g4378 ( 
.A(n_3761),
.Y(n_4378)
);

NAND2xp5_ASAP7_75t_SL g4379 ( 
.A(n_3639),
.B(n_649),
.Y(n_4379)
);

O2A1O1Ixp33_ASAP7_75t_L g4380 ( 
.A1(n_3939),
.A2(n_651),
.B(n_652),
.C(n_650),
.Y(n_4380)
);

O2A1O1Ixp33_ASAP7_75t_L g4381 ( 
.A1(n_3953),
.A2(n_651),
.B(n_652),
.C(n_650),
.Y(n_4381)
);

OAI22xp5_ASAP7_75t_L g4382 ( 
.A1(n_3990),
.A2(n_653),
.B1(n_654),
.B2(n_652),
.Y(n_4382)
);

NAND2xp5_ASAP7_75t_L g4383 ( 
.A(n_3819),
.B(n_653),
.Y(n_4383)
);

AND2x4_ASAP7_75t_L g4384 ( 
.A(n_3933),
.B(n_653),
.Y(n_4384)
);

INVxp33_ASAP7_75t_SL g4385 ( 
.A(n_4009),
.Y(n_4385)
);

NAND2xp5_ASAP7_75t_L g4386 ( 
.A(n_3832),
.B(n_654),
.Y(n_4386)
);

AND2x2_ASAP7_75t_L g4387 ( 
.A(n_3781),
.B(n_1104),
.Y(n_4387)
);

NOR2xp67_ASAP7_75t_L g4388 ( 
.A(n_3951),
.B(n_654),
.Y(n_4388)
);

AND2x2_ASAP7_75t_L g4389 ( 
.A(n_3827),
.B(n_3780),
.Y(n_4389)
);

NOR3xp33_ASAP7_75t_L g4390 ( 
.A(n_3643),
.B(n_656),
.C(n_655),
.Y(n_4390)
);

AND2x2_ASAP7_75t_L g4391 ( 
.A(n_3784),
.B(n_1108),
.Y(n_4391)
);

A2O1A1Ixp33_ASAP7_75t_L g4392 ( 
.A1(n_3995),
.A2(n_3785),
.B(n_3758),
.C(n_3646),
.Y(n_4392)
);

INVx3_ASAP7_75t_L g4393 ( 
.A(n_3739),
.Y(n_4393)
);

NAND3xp33_ASAP7_75t_L g4394 ( 
.A(n_3818),
.B(n_1109),
.C(n_1108),
.Y(n_4394)
);

HB1xp67_ASAP7_75t_L g4395 ( 
.A(n_3798),
.Y(n_4395)
);

O2A1O1Ixp33_ASAP7_75t_L g4396 ( 
.A1(n_3973),
.A2(n_656),
.B(n_657),
.C(n_655),
.Y(n_4396)
);

OAI22xp5_ASAP7_75t_L g4397 ( 
.A1(n_3925),
.A2(n_3820),
.B1(n_3918),
.B2(n_3464),
.Y(n_4397)
);

NAND2xp5_ASAP7_75t_L g4398 ( 
.A(n_3836),
.B(n_655),
.Y(n_4398)
);

BUFx2_ASAP7_75t_L g4399 ( 
.A(n_3951),
.Y(n_4399)
);

O2A1O1Ixp5_ASAP7_75t_SL g4400 ( 
.A1(n_3729),
.A2(n_657),
.B(n_658),
.C(n_656),
.Y(n_4400)
);

AO22x1_ASAP7_75t_L g4401 ( 
.A1(n_3964),
.A2(n_3652),
.B1(n_3655),
.B2(n_3753),
.Y(n_4401)
);

BUFx8_ASAP7_75t_SL g4402 ( 
.A(n_3964),
.Y(n_4402)
);

OAI21x1_ASAP7_75t_L g4403 ( 
.A1(n_3751),
.A2(n_658),
.B(n_657),
.Y(n_4403)
);

NAND2xp5_ASAP7_75t_L g4404 ( 
.A(n_3461),
.B(n_658),
.Y(n_4404)
);

NAND2xp5_ASAP7_75t_L g4405 ( 
.A(n_3778),
.B(n_659),
.Y(n_4405)
);

A2O1A1Ixp33_ASAP7_75t_SL g4406 ( 
.A1(n_3682),
.A2(n_68),
.B(n_66),
.C(n_67),
.Y(n_4406)
);

AOI21xp5_ASAP7_75t_L g4407 ( 
.A1(n_3645),
.A2(n_660),
.B(n_659),
.Y(n_4407)
);

NAND2xp5_ASAP7_75t_SL g4408 ( 
.A(n_3739),
.B(n_660),
.Y(n_4408)
);

NAND2xp5_ASAP7_75t_L g4409 ( 
.A(n_3872),
.B(n_660),
.Y(n_4409)
);

NOR3xp33_ASAP7_75t_L g4410 ( 
.A(n_4026),
.B(n_662),
.C(n_661),
.Y(n_4410)
);

INVx2_ASAP7_75t_L g4411 ( 
.A(n_3812),
.Y(n_4411)
);

NOR3xp33_ASAP7_75t_L g4412 ( 
.A(n_3989),
.B(n_663),
.C(n_661),
.Y(n_4412)
);

INVx2_ASAP7_75t_L g4413 ( 
.A(n_3845),
.Y(n_4413)
);

NAND2x1p5_ASAP7_75t_L g4414 ( 
.A(n_3739),
.B(n_668),
.Y(n_4414)
);

AOI21xp5_ASAP7_75t_L g4415 ( 
.A1(n_3958),
.A2(n_663),
.B(n_661),
.Y(n_4415)
);

AOI21xp5_ASAP7_75t_L g4416 ( 
.A1(n_3738),
.A2(n_664),
.B(n_663),
.Y(n_4416)
);

AND2x2_ASAP7_75t_L g4417 ( 
.A(n_3928),
.B(n_1098),
.Y(n_4417)
);

O2A1O1Ixp33_ASAP7_75t_L g4418 ( 
.A1(n_3726),
.A2(n_665),
.B(n_666),
.C(n_664),
.Y(n_4418)
);

INVx1_ASAP7_75t_L g4419 ( 
.A(n_3518),
.Y(n_4419)
);

O2A1O1Ixp5_ASAP7_75t_L g4420 ( 
.A1(n_4018),
.A2(n_665),
.B(n_666),
.C(n_664),
.Y(n_4420)
);

NAND2xp5_ASAP7_75t_SL g4421 ( 
.A(n_3766),
.B(n_665),
.Y(n_4421)
);

OAI22xp5_ASAP7_75t_L g4422 ( 
.A1(n_3868),
.A2(n_667),
.B1(n_668),
.B2(n_666),
.Y(n_4422)
);

NAND2xp5_ASAP7_75t_SL g4423 ( 
.A(n_3766),
.B(n_667),
.Y(n_4423)
);

NOR2xp33_ASAP7_75t_L g4424 ( 
.A(n_3870),
.B(n_667),
.Y(n_4424)
);

AOI21xp5_ASAP7_75t_L g4425 ( 
.A1(n_3644),
.A2(n_3659),
.B(n_3647),
.Y(n_4425)
);

NOR2xp33_ASAP7_75t_L g4426 ( 
.A(n_3791),
.B(n_669),
.Y(n_4426)
);

INVx2_ASAP7_75t_L g4427 ( 
.A(n_3955),
.Y(n_4427)
);

OR2x6_ASAP7_75t_SL g4428 ( 
.A(n_3710),
.B(n_1110),
.Y(n_4428)
);

BUFx6f_ASAP7_75t_L g4429 ( 
.A(n_3766),
.Y(n_4429)
);

INVxp67_ASAP7_75t_L g4430 ( 
.A(n_3794),
.Y(n_4430)
);

NOR2xp33_ASAP7_75t_L g4431 ( 
.A(n_3520),
.B(n_3523),
.Y(n_4431)
);

NAND2xp5_ASAP7_75t_L g4432 ( 
.A(n_3536),
.B(n_670),
.Y(n_4432)
);

NAND2xp5_ASAP7_75t_L g4433 ( 
.A(n_3549),
.B(n_670),
.Y(n_4433)
);

NAND2xp5_ASAP7_75t_L g4434 ( 
.A(n_3552),
.B(n_670),
.Y(n_4434)
);

NOR2xp33_ASAP7_75t_L g4435 ( 
.A(n_3554),
.B(n_671),
.Y(n_4435)
);

AND2x2_ASAP7_75t_L g4436 ( 
.A(n_3556),
.B(n_1111),
.Y(n_4436)
);

NOR2xp33_ASAP7_75t_L g4437 ( 
.A(n_3566),
.B(n_3572),
.Y(n_4437)
);

NOR2xp33_ASAP7_75t_L g4438 ( 
.A(n_3579),
.B(n_671),
.Y(n_4438)
);

NOR2xp33_ASAP7_75t_L g4439 ( 
.A(n_3580),
.B(n_671),
.Y(n_4439)
);

NOR2xp33_ASAP7_75t_L g4440 ( 
.A(n_3589),
.B(n_672),
.Y(n_4440)
);

NAND2xp5_ASAP7_75t_L g4441 ( 
.A(n_3595),
.B(n_672),
.Y(n_4441)
);

NAND2xp5_ASAP7_75t_SL g4442 ( 
.A(n_3792),
.B(n_673),
.Y(n_4442)
);

NAND2xp5_ASAP7_75t_L g4443 ( 
.A(n_3596),
.B(n_673),
.Y(n_4443)
);

O2A1O1Ixp33_ASAP7_75t_L g4444 ( 
.A1(n_3626),
.A2(n_674),
.B(n_675),
.C(n_673),
.Y(n_4444)
);

INVx4_ASAP7_75t_L g4445 ( 
.A(n_3792),
.Y(n_4445)
);

NAND2xp5_ASAP7_75t_SL g4446 ( 
.A(n_3792),
.B(n_674),
.Y(n_4446)
);

AND2x4_ASAP7_75t_L g4447 ( 
.A(n_3728),
.B(n_674),
.Y(n_4447)
);

NOR2xp33_ASAP7_75t_L g4448 ( 
.A(n_3602),
.B(n_675),
.Y(n_4448)
);

O2A1O1Ixp33_ASAP7_75t_L g4449 ( 
.A1(n_3709),
.A2(n_676),
.B(n_677),
.C(n_675),
.Y(n_4449)
);

BUFx2_ASAP7_75t_L g4450 ( 
.A(n_3808),
.Y(n_4450)
);

BUFx3_ASAP7_75t_L g4451 ( 
.A(n_3808),
.Y(n_4451)
);

OAI22xp5_ASAP7_75t_L g4452 ( 
.A1(n_3476),
.A2(n_677),
.B1(n_678),
.B2(n_676),
.Y(n_4452)
);

AOI21xp5_ASAP7_75t_L g4453 ( 
.A1(n_3529),
.A2(n_678),
.B(n_677),
.Y(n_4453)
);

INVx1_ASAP7_75t_L g4454 ( 
.A(n_3618),
.Y(n_4454)
);

NAND2xp5_ASAP7_75t_SL g4455 ( 
.A(n_3808),
.B(n_4015),
.Y(n_4455)
);

INVx1_ASAP7_75t_L g4456 ( 
.A(n_3622),
.Y(n_4456)
);

AND2x2_ASAP7_75t_L g4457 ( 
.A(n_3623),
.B(n_1097),
.Y(n_4457)
);

AOI21xp5_ASAP7_75t_L g4458 ( 
.A1(n_3531),
.A2(n_3553),
.B(n_3534),
.Y(n_4458)
);

NOR2x1_ASAP7_75t_L g4459 ( 
.A(n_3855),
.B(n_679),
.Y(n_4459)
);

NOR2xp33_ASAP7_75t_L g4460 ( 
.A(n_3632),
.B(n_3633),
.Y(n_4460)
);

INVx2_ASAP7_75t_L g4461 ( 
.A(n_3955),
.Y(n_4461)
);

AND2x4_ASAP7_75t_L g4462 ( 
.A(n_3873),
.B(n_679),
.Y(n_4462)
);

NOR2xp33_ASAP7_75t_L g4463 ( 
.A(n_3641),
.B(n_679),
.Y(n_4463)
);

BUFx2_ASAP7_75t_L g4464 ( 
.A(n_3873),
.Y(n_4464)
);

O2A1O1Ixp33_ASAP7_75t_L g4465 ( 
.A1(n_3771),
.A2(n_681),
.B(n_682),
.C(n_680),
.Y(n_4465)
);

NOR2xp33_ASAP7_75t_L g4466 ( 
.A(n_3661),
.B(n_3672),
.Y(n_4466)
);

NOR2xp33_ASAP7_75t_L g4467 ( 
.A(n_3676),
.B(n_680),
.Y(n_4467)
);

INVx1_ASAP7_75t_L g4468 ( 
.A(n_3679),
.Y(n_4468)
);

AOI21xp5_ASAP7_75t_L g4469 ( 
.A1(n_3585),
.A2(n_681),
.B(n_680),
.Y(n_4469)
);

CKINVDCx5p33_ASAP7_75t_R g4470 ( 
.A(n_3755),
.Y(n_4470)
);

AOI21xp5_ASAP7_75t_L g4471 ( 
.A1(n_3593),
.A2(n_682),
.B(n_681),
.Y(n_4471)
);

INVx1_ASAP7_75t_L g4472 ( 
.A(n_3684),
.Y(n_4472)
);

BUFx2_ASAP7_75t_L g4473 ( 
.A(n_3873),
.Y(n_4473)
);

BUFx2_ASAP7_75t_L g4474 ( 
.A(n_3880),
.Y(n_4474)
);

BUFx6f_ASAP7_75t_L g4475 ( 
.A(n_3880),
.Y(n_4475)
);

OR2x2_ASAP7_75t_L g4476 ( 
.A(n_3693),
.B(n_683),
.Y(n_4476)
);

INVx2_ASAP7_75t_L g4477 ( 
.A(n_3855),
.Y(n_4477)
);

NAND2xp5_ASAP7_75t_L g4478 ( 
.A(n_3694),
.B(n_683),
.Y(n_4478)
);

INVx3_ASAP7_75t_L g4479 ( 
.A(n_3880),
.Y(n_4479)
);

O2A1O1Ixp5_ASAP7_75t_L g4480 ( 
.A1(n_3747),
.A2(n_684),
.B(n_685),
.C(n_683),
.Y(n_4480)
);

NAND2xp5_ASAP7_75t_L g4481 ( 
.A(n_3695),
.B(n_684),
.Y(n_4481)
);

HB1xp67_ASAP7_75t_L g4482 ( 
.A(n_3799),
.Y(n_4482)
);

BUFx6f_ASAP7_75t_L g4483 ( 
.A(n_3895),
.Y(n_4483)
);

AO21x1_ASAP7_75t_L g4484 ( 
.A1(n_3782),
.A2(n_686),
.B(n_685),
.Y(n_4484)
);

NAND2xp5_ASAP7_75t_L g4485 ( 
.A(n_3775),
.B(n_686),
.Y(n_4485)
);

NOR2xp33_ASAP7_75t_L g4486 ( 
.A(n_3802),
.B(n_687),
.Y(n_4486)
);

NAND2xp5_ASAP7_75t_L g4487 ( 
.A(n_3621),
.B(n_687),
.Y(n_4487)
);

HB1xp67_ASAP7_75t_L g4488 ( 
.A(n_3895),
.Y(n_4488)
);

INVx2_ASAP7_75t_L g4489 ( 
.A(n_3902),
.Y(n_4489)
);

NAND2xp5_ASAP7_75t_SL g4490 ( 
.A(n_3895),
.B(n_687),
.Y(n_4490)
);

INVx1_ASAP7_75t_SL g4491 ( 
.A(n_3931),
.Y(n_4491)
);

BUFx2_ASAP7_75t_L g4492 ( 
.A(n_3931),
.Y(n_4492)
);

NAND2xp5_ASAP7_75t_SL g4493 ( 
.A(n_3931),
.B(n_688),
.Y(n_4493)
);

O2A1O1Ixp33_ASAP7_75t_L g4494 ( 
.A1(n_3795),
.A2(n_689),
.B(n_690),
.C(n_688),
.Y(n_4494)
);

AOI21xp5_ASAP7_75t_L g4495 ( 
.A1(n_3519),
.A2(n_3524),
.B(n_3970),
.Y(n_4495)
);

A2O1A1Ixp33_ASAP7_75t_L g4496 ( 
.A1(n_3711),
.A2(n_689),
.B(n_690),
.C(n_688),
.Y(n_4496)
);

NAND2xp5_ASAP7_75t_L g4497 ( 
.A(n_3638),
.B(n_689),
.Y(n_4497)
);

AND2x2_ASAP7_75t_L g4498 ( 
.A(n_3640),
.B(n_690),
.Y(n_4498)
);

OAI21xp5_ASAP7_75t_L g4499 ( 
.A1(n_3860),
.A2(n_692),
.B(n_691),
.Y(n_4499)
);

OAI22xp5_ASAP7_75t_SL g4500 ( 
.A1(n_3776),
.A2(n_692),
.B1(n_693),
.B2(n_691),
.Y(n_4500)
);

HB1xp67_ASAP7_75t_L g4501 ( 
.A(n_3970),
.Y(n_4501)
);

INVx1_ASAP7_75t_SL g4502 ( 
.A(n_3970),
.Y(n_4502)
);

BUFx2_ASAP7_75t_L g4503 ( 
.A(n_4015),
.Y(n_4503)
);

NAND2xp5_ASAP7_75t_L g4504 ( 
.A(n_3642),
.B(n_691),
.Y(n_4504)
);

NOR2xp33_ASAP7_75t_L g4505 ( 
.A(n_3650),
.B(n_692),
.Y(n_4505)
);

INVx1_ASAP7_75t_L g4506 ( 
.A(n_3779),
.Y(n_4506)
);

NOR2xp33_ASAP7_75t_L g4507 ( 
.A(n_3654),
.B(n_693),
.Y(n_4507)
);

BUFx3_ASAP7_75t_L g4508 ( 
.A(n_4015),
.Y(n_4508)
);

OAI21xp5_ASAP7_75t_L g4509 ( 
.A1(n_3952),
.A2(n_694),
.B(n_693),
.Y(n_4509)
);

INVx2_ASAP7_75t_L g4510 ( 
.A(n_3724),
.Y(n_4510)
);

OAI22xp33_ASAP7_75t_L g4511 ( 
.A1(n_3891),
.A2(n_695),
.B1(n_696),
.B2(n_694),
.Y(n_4511)
);

NAND2xp5_ASAP7_75t_L g4512 ( 
.A(n_3658),
.B(n_694),
.Y(n_4512)
);

AOI21xp33_ASAP7_75t_L g4513 ( 
.A1(n_3649),
.A2(n_698),
.B(n_697),
.Y(n_4513)
);

A2O1A1Ixp33_ASAP7_75t_L g4514 ( 
.A1(n_3665),
.A2(n_698),
.B(n_699),
.C(n_697),
.Y(n_4514)
);

NOR2xp33_ASAP7_75t_L g4515 ( 
.A(n_3669),
.B(n_698),
.Y(n_4515)
);

NAND2xp5_ASAP7_75t_SL g4516 ( 
.A(n_3560),
.B(n_700),
.Y(n_4516)
);

O2A1O1Ixp33_ASAP7_75t_L g4517 ( 
.A1(n_3859),
.A2(n_701),
.B(n_702),
.C(n_700),
.Y(n_4517)
);

AOI21xp5_ASAP7_75t_L g4518 ( 
.A1(n_3894),
.A2(n_701),
.B(n_700),
.Y(n_4518)
);

INVx2_ASAP7_75t_L g4519 ( 
.A(n_3625),
.Y(n_4519)
);

A2O1A1Ixp33_ASAP7_75t_L g4520 ( 
.A1(n_3678),
.A2(n_703),
.B(n_704),
.C(n_702),
.Y(n_4520)
);

INVx1_ASAP7_75t_L g4521 ( 
.A(n_3915),
.Y(n_4521)
);

OAI22xp5_ASAP7_75t_L g4522 ( 
.A1(n_3824),
.A2(n_3901),
.B1(n_3920),
.B2(n_3898),
.Y(n_4522)
);

NAND2xp5_ASAP7_75t_L g4523 ( 
.A(n_3683),
.B(n_702),
.Y(n_4523)
);

INVxp67_ASAP7_75t_L g4524 ( 
.A(n_3686),
.Y(n_4524)
);

HB1xp67_ASAP7_75t_L g4525 ( 
.A(n_3945),
.Y(n_4525)
);

AOI21x1_ASAP7_75t_L g4526 ( 
.A1(n_3637),
.A2(n_704),
.B(n_703),
.Y(n_4526)
);

OR2x2_ASAP7_75t_L g4527 ( 
.A(n_3921),
.B(n_703),
.Y(n_4527)
);

AND2x4_ASAP7_75t_L g4528 ( 
.A(n_3688),
.B(n_705),
.Y(n_4528)
);

NOR2x1_ASAP7_75t_SL g4529 ( 
.A(n_3972),
.B(n_1115),
.Y(n_4529)
);

AND2x2_ASAP7_75t_L g4530 ( 
.A(n_3691),
.B(n_705),
.Y(n_4530)
);

NAND2xp5_ASAP7_75t_L g4531 ( 
.A(n_3703),
.B(n_706),
.Y(n_4531)
);

AOI33xp33_ASAP7_75t_L g4532 ( 
.A1(n_3900),
.A2(n_70),
.A3(n_72),
.B1(n_68),
.B2(n_69),
.B3(n_71),
.Y(n_4532)
);

INVx2_ASAP7_75t_L g4533 ( 
.A(n_3966),
.Y(n_4533)
);

NAND2xp5_ASAP7_75t_L g4534 ( 
.A(n_3705),
.B(n_3712),
.Y(n_4534)
);

INVx1_ASAP7_75t_L g4535 ( 
.A(n_4025),
.Y(n_4535)
);

INVx1_ASAP7_75t_L g4536 ( 
.A(n_3653),
.Y(n_4536)
);

AND2x2_ASAP7_75t_SL g4537 ( 
.A(n_3605),
.B(n_706),
.Y(n_4537)
);

NAND2xp5_ASAP7_75t_L g4538 ( 
.A(n_3718),
.B(n_706),
.Y(n_4538)
);

AOI21xp5_ASAP7_75t_L g4539 ( 
.A1(n_3923),
.A2(n_708),
.B(n_707),
.Y(n_4539)
);

BUFx2_ASAP7_75t_L g4540 ( 
.A(n_3772),
.Y(n_4540)
);

AND2x4_ASAP7_75t_L g4541 ( 
.A(n_3723),
.B(n_707),
.Y(n_4541)
);

AND2x2_ASAP7_75t_L g4542 ( 
.A(n_3730),
.B(n_3735),
.Y(n_4542)
);

NAND2xp5_ASAP7_75t_L g4543 ( 
.A(n_3736),
.B(n_707),
.Y(n_4543)
);

A2O1A1Ixp33_ASAP7_75t_L g4544 ( 
.A1(n_3737),
.A2(n_709),
.B(n_710),
.C(n_708),
.Y(n_4544)
);

AOI21xp5_ASAP7_75t_L g4545 ( 
.A1(n_3924),
.A2(n_709),
.B(n_708),
.Y(n_4545)
);

AOI222xp33_ASAP7_75t_L g4546 ( 
.A1(n_3935),
.A2(n_740),
.B1(n_724),
.B2(n_748),
.C1(n_732),
.C2(n_716),
.Y(n_4546)
);

O2A1O1Ixp33_ASAP7_75t_L g4547 ( 
.A1(n_3949),
.A2(n_710),
.B(n_711),
.C(n_709),
.Y(n_4547)
);

NAND2xp5_ASAP7_75t_SL g4548 ( 
.A(n_3611),
.B(n_3988),
.Y(n_4548)
);

BUFx8_ASAP7_75t_SL g4549 ( 
.A(n_3960),
.Y(n_4549)
);

INVx2_ASAP7_75t_SL g4550 ( 
.A(n_3927),
.Y(n_4550)
);

INVx1_ASAP7_75t_L g4551 ( 
.A(n_3929),
.Y(n_4551)
);

NOR2xp67_ASAP7_75t_SL g4552 ( 
.A(n_3930),
.B(n_710),
.Y(n_4552)
);

O2A1O1Ixp33_ASAP7_75t_L g4553 ( 
.A1(n_3992),
.A2(n_712),
.B(n_713),
.C(n_711),
.Y(n_4553)
);

AOI22xp33_ASAP7_75t_L g4554 ( 
.A1(n_3746),
.A2(n_712),
.B1(n_714),
.B2(n_711),
.Y(n_4554)
);

AOI21xp5_ASAP7_75t_L g4555 ( 
.A1(n_3932),
.A2(n_715),
.B(n_714),
.Y(n_4555)
);

CKINVDCx5p33_ASAP7_75t_R g4556 ( 
.A(n_3749),
.Y(n_4556)
);

AOI21xp5_ASAP7_75t_L g4557 ( 
.A1(n_3940),
.A2(n_715),
.B(n_714),
.Y(n_4557)
);

AO32x1_ASAP7_75t_L g4558 ( 
.A1(n_3813),
.A2(n_4024),
.A3(n_3948),
.B1(n_3956),
.B2(n_3943),
.Y(n_4558)
);

A2O1A1Ixp33_ASAP7_75t_L g4559 ( 
.A1(n_3942),
.A2(n_716),
.B(n_717),
.C(n_715),
.Y(n_4559)
);

OAI22xp5_ASAP7_75t_L g4560 ( 
.A1(n_3962),
.A2(n_717),
.B1(n_718),
.B2(n_716),
.Y(n_4560)
);

INVx1_ASAP7_75t_L g4561 ( 
.A(n_3974),
.Y(n_4561)
);

OAI22xp5_ASAP7_75t_L g4562 ( 
.A1(n_3997),
.A2(n_719),
.B1(n_720),
.B2(n_718),
.Y(n_4562)
);

NAND3xp33_ASAP7_75t_SL g4563 ( 
.A(n_3750),
.B(n_69),
.C(n_70),
.Y(n_4563)
);

BUFx2_ASAP7_75t_L g4564 ( 
.A(n_3514),
.Y(n_4564)
);

NAND2xp5_ASAP7_75t_L g4565 ( 
.A(n_3999),
.B(n_718),
.Y(n_4565)
);

AND2x6_ASAP7_75t_L g4566 ( 
.A(n_4014),
.B(n_719),
.Y(n_4566)
);

AND2x2_ASAP7_75t_L g4567 ( 
.A(n_4016),
.B(n_1092),
.Y(n_4567)
);

NOR2xp33_ASAP7_75t_L g4568 ( 
.A(n_4017),
.B(n_720),
.Y(n_4568)
);

OR2x2_ASAP7_75t_L g4569 ( 
.A(n_4021),
.B(n_720),
.Y(n_4569)
);

NAND2xp5_ASAP7_75t_L g4570 ( 
.A(n_3893),
.B(n_721),
.Y(n_4570)
);

INVx6_ASAP7_75t_L g4571 ( 
.A(n_3852),
.Y(n_4571)
);

O2A1O1Ixp33_ASAP7_75t_L g4572 ( 
.A1(n_3853),
.A2(n_722),
.B(n_723),
.C(n_721),
.Y(n_4572)
);

A2O1A1Ixp33_ASAP7_75t_L g4573 ( 
.A1(n_4022),
.A2(n_722),
.B(n_723),
.C(n_721),
.Y(n_4573)
);

NAND2xp5_ASAP7_75t_L g4574 ( 
.A(n_3854),
.B(n_723),
.Y(n_4574)
);

OAI22xp5_ASAP7_75t_L g4575 ( 
.A1(n_3479),
.A2(n_725),
.B1(n_726),
.B2(n_724),
.Y(n_4575)
);

INVx3_ASAP7_75t_SL g4576 ( 
.A(n_4027),
.Y(n_4576)
);

NAND2xp5_ASAP7_75t_SL g4577 ( 
.A(n_3486),
.B(n_3490),
.Y(n_4577)
);

INVx1_ASAP7_75t_L g4578 ( 
.A(n_3756),
.Y(n_4578)
);

NAND2xp5_ASAP7_75t_L g4579 ( 
.A(n_3869),
.B(n_725),
.Y(n_4579)
);

OAI22xp5_ASAP7_75t_L g4580 ( 
.A1(n_3493),
.A2(n_726),
.B1(n_727),
.B2(n_725),
.Y(n_4580)
);

NAND2xp5_ASAP7_75t_L g4581 ( 
.A(n_3759),
.B(n_726),
.Y(n_4581)
);

NAND2xp5_ASAP7_75t_SL g4582 ( 
.A(n_3760),
.B(n_728),
.Y(n_4582)
);

AND2x2_ASAP7_75t_SL g4583 ( 
.A(n_3762),
.B(n_728),
.Y(n_4583)
);

AOI21xp5_ASAP7_75t_L g4584 ( 
.A1(n_3879),
.A2(n_729),
.B(n_728),
.Y(n_4584)
);

BUFx3_ASAP7_75t_L g4585 ( 
.A(n_3883),
.Y(n_4585)
);

INVx1_ASAP7_75t_L g4586 ( 
.A(n_3765),
.Y(n_4586)
);

INVx2_ASAP7_75t_L g4587 ( 
.A(n_3793),
.Y(n_4587)
);

INVx4_ASAP7_75t_L g4588 ( 
.A(n_3801),
.Y(n_4588)
);

AND3x1_ASAP7_75t_SL g4589 ( 
.A(n_3817),
.B(n_730),
.C(n_729),
.Y(n_4589)
);

NOR2xp33_ASAP7_75t_L g4590 ( 
.A(n_3844),
.B(n_729),
.Y(n_4590)
);

NAND2xp5_ASAP7_75t_L g4591 ( 
.A(n_4039),
.B(n_3828),
.Y(n_4591)
);

AO31x2_ASAP7_75t_L g4592 ( 
.A1(n_4074),
.A2(n_3833),
.A3(n_3838),
.B(n_3768),
.Y(n_4592)
);

AOI21x1_ASAP7_75t_L g4593 ( 
.A1(n_4127),
.A2(n_731),
.B(n_730),
.Y(n_4593)
);

NAND2xp33_ASAP7_75t_L g4594 ( 
.A(n_4208),
.B(n_730),
.Y(n_4594)
);

OAI21x1_ASAP7_75t_SL g4595 ( 
.A1(n_4119),
.A2(n_4031),
.B(n_4266),
.Y(n_4595)
);

BUFx8_ASAP7_75t_SL g4596 ( 
.A(n_4087),
.Y(n_4596)
);

OA22x2_ASAP7_75t_L g4597 ( 
.A1(n_4067),
.A2(n_732),
.B1(n_733),
.B2(n_731),
.Y(n_4597)
);

OA21x2_ASAP7_75t_L g4598 ( 
.A1(n_4427),
.A2(n_732),
.B(n_731),
.Y(n_4598)
);

AOI21xp5_ASAP7_75t_L g4599 ( 
.A1(n_4118),
.A2(n_734),
.B(n_733),
.Y(n_4599)
);

O2A1O1Ixp33_ASAP7_75t_SL g4600 ( 
.A1(n_4406),
.A2(n_734),
.B(n_735),
.C(n_733),
.Y(n_4600)
);

BUFx6f_ASAP7_75t_L g4601 ( 
.A(n_4128),
.Y(n_4601)
);

AOI21x1_ASAP7_75t_L g4602 ( 
.A1(n_4540),
.A2(n_736),
.B(n_735),
.Y(n_4602)
);

OR2x2_ASAP7_75t_L g4603 ( 
.A(n_4073),
.B(n_735),
.Y(n_4603)
);

OAI21x1_ASAP7_75t_L g4604 ( 
.A1(n_4055),
.A2(n_737),
.B(n_736),
.Y(n_4604)
);

CKINVDCx8_ASAP7_75t_R g4605 ( 
.A(n_4069),
.Y(n_4605)
);

INVx8_ASAP7_75t_L g4606 ( 
.A(n_4097),
.Y(n_4606)
);

INVx3_ASAP7_75t_L g4607 ( 
.A(n_4304),
.Y(n_4607)
);

CKINVDCx5p33_ASAP7_75t_R g4608 ( 
.A(n_4046),
.Y(n_4608)
);

OR2x2_ASAP7_75t_L g4609 ( 
.A(n_4375),
.B(n_736),
.Y(n_4609)
);

INVx1_ASAP7_75t_SL g4610 ( 
.A(n_4163),
.Y(n_4610)
);

OAI21xp5_ASAP7_75t_L g4611 ( 
.A1(n_4052),
.A2(n_738),
.B(n_737),
.Y(n_4611)
);

OAI21x1_ASAP7_75t_SL g4612 ( 
.A1(n_4145),
.A2(n_739),
.B(n_738),
.Y(n_4612)
);

OAI21xp33_ASAP7_75t_L g4613 ( 
.A1(n_4257),
.A2(n_739),
.B(n_738),
.Y(n_4613)
);

OAI21x1_ASAP7_75t_L g4614 ( 
.A1(n_4111),
.A2(n_740),
.B(n_739),
.Y(n_4614)
);

AND2x4_ASAP7_75t_L g4615 ( 
.A(n_4067),
.B(n_742),
.Y(n_4615)
);

INVx2_ASAP7_75t_L g4616 ( 
.A(n_4220),
.Y(n_4616)
);

INVx1_ASAP7_75t_L g4617 ( 
.A(n_4071),
.Y(n_4617)
);

NAND2xp5_ASAP7_75t_L g4618 ( 
.A(n_4090),
.B(n_741),
.Y(n_4618)
);

AOI22xp5_ASAP7_75t_L g4619 ( 
.A1(n_4224),
.A2(n_1098),
.B1(n_1100),
.B2(n_1097),
.Y(n_4619)
);

NAND2xp5_ASAP7_75t_L g4620 ( 
.A(n_4103),
.B(n_741),
.Y(n_4620)
);

OAI22x1_ASAP7_75t_L g4621 ( 
.A1(n_4168),
.A2(n_742),
.B1(n_743),
.B2(n_741),
.Y(n_4621)
);

OAI21x1_ASAP7_75t_SL g4622 ( 
.A1(n_4459),
.A2(n_743),
.B(n_742),
.Y(n_4622)
);

INVx2_ASAP7_75t_L g4623 ( 
.A(n_4041),
.Y(n_4623)
);

OAI21x1_ASAP7_75t_L g4624 ( 
.A1(n_4100),
.A2(n_745),
.B(n_744),
.Y(n_4624)
);

AOI21x1_ASAP7_75t_L g4625 ( 
.A1(n_4519),
.A2(n_745),
.B(n_744),
.Y(n_4625)
);

OA22x2_ASAP7_75t_L g4626 ( 
.A1(n_4218),
.A2(n_4353),
.B1(n_4217),
.B2(n_4350),
.Y(n_4626)
);

AO31x2_ASAP7_75t_L g4627 ( 
.A1(n_4461),
.A2(n_745),
.A3(n_746),
.B(n_744),
.Y(n_4627)
);

AND2x6_ASAP7_75t_L g4628 ( 
.A(n_4084),
.B(n_746),
.Y(n_4628)
);

NAND3xp33_ASAP7_75t_L g4629 ( 
.A(n_4064),
.B(n_747),
.C(n_746),
.Y(n_4629)
);

INVx2_ASAP7_75t_L g4630 ( 
.A(n_4089),
.Y(n_4630)
);

AO31x2_ASAP7_75t_L g4631 ( 
.A1(n_4477),
.A2(n_4510),
.A3(n_4489),
.B(n_4588),
.Y(n_4631)
);

AND2x2_ASAP7_75t_L g4632 ( 
.A(n_4201),
.B(n_747),
.Y(n_4632)
);

AOI21xp5_ASAP7_75t_L g4633 ( 
.A1(n_4252),
.A2(n_748),
.B(n_747),
.Y(n_4633)
);

OAI21x1_ASAP7_75t_L g4634 ( 
.A1(n_4099),
.A2(n_749),
.B(n_748),
.Y(n_4634)
);

AOI21x1_ASAP7_75t_L g4635 ( 
.A1(n_4536),
.A2(n_4455),
.B(n_4256),
.Y(n_4635)
);

A2O1A1Ixp33_ASAP7_75t_L g4636 ( 
.A1(n_4199),
.A2(n_750),
.B(n_751),
.C(n_749),
.Y(n_4636)
);

OAI21x1_ASAP7_75t_L g4637 ( 
.A1(n_4495),
.A2(n_750),
.B(n_749),
.Y(n_4637)
);

OAI22xp5_ASAP7_75t_L g4638 ( 
.A1(n_4199),
.A2(n_4428),
.B1(n_4385),
.B2(n_4218),
.Y(n_4638)
);

BUFx3_ASAP7_75t_L g4639 ( 
.A(n_4304),
.Y(n_4639)
);

AO31x2_ASAP7_75t_L g4640 ( 
.A1(n_4588),
.A2(n_751),
.A3(n_752),
.B(n_750),
.Y(n_4640)
);

OAI22xp5_ASAP7_75t_L g4641 ( 
.A1(n_4300),
.A2(n_752),
.B1(n_753),
.B2(n_751),
.Y(n_4641)
);

OAI21x1_ASAP7_75t_L g4642 ( 
.A1(n_4084),
.A2(n_754),
.B(n_753),
.Y(n_4642)
);

OR2x2_ASAP7_75t_L g4643 ( 
.A(n_4395),
.B(n_753),
.Y(n_4643)
);

INVx1_ASAP7_75t_L g4644 ( 
.A(n_4109),
.Y(n_4644)
);

OAI21x1_ASAP7_75t_L g4645 ( 
.A1(n_4116),
.A2(n_755),
.B(n_754),
.Y(n_4645)
);

AOI21xp5_ASAP7_75t_L g4646 ( 
.A1(n_4577),
.A2(n_755),
.B(n_754),
.Y(n_4646)
);

INVx1_ASAP7_75t_L g4647 ( 
.A(n_4117),
.Y(n_4647)
);

AOI211x1_ASAP7_75t_L g4648 ( 
.A1(n_4050),
.A2(n_757),
.B(n_758),
.C(n_756),
.Y(n_4648)
);

INVxp67_ASAP7_75t_SL g4649 ( 
.A(n_4091),
.Y(n_4649)
);

NOR3xp33_ASAP7_75t_L g4650 ( 
.A(n_4303),
.B(n_4033),
.C(n_4062),
.Y(n_4650)
);

BUFx2_ASAP7_75t_L g4651 ( 
.A(n_4402),
.Y(n_4651)
);

AOI21xp5_ASAP7_75t_L g4652 ( 
.A1(n_4223),
.A2(n_757),
.B(n_756),
.Y(n_4652)
);

AOI21xp33_ASAP7_75t_L g4653 ( 
.A1(n_4038),
.A2(n_757),
.B(n_756),
.Y(n_4653)
);

INVx2_ASAP7_75t_SL g4654 ( 
.A(n_4079),
.Y(n_4654)
);

OR2x6_ASAP7_75t_L g4655 ( 
.A(n_4148),
.B(n_758),
.Y(n_4655)
);

CKINVDCx5p33_ASAP7_75t_R g4656 ( 
.A(n_4044),
.Y(n_4656)
);

AND2x4_ASAP7_75t_L g4657 ( 
.A(n_4061),
.B(n_759),
.Y(n_4657)
);

OAI21x1_ASAP7_75t_SL g4658 ( 
.A1(n_4261),
.A2(n_759),
.B(n_758),
.Y(n_4658)
);

A2O1A1Ixp33_ASAP7_75t_L g4659 ( 
.A1(n_4370),
.A2(n_760),
.B(n_761),
.C(n_759),
.Y(n_4659)
);

OAI21xp5_ASAP7_75t_L g4660 ( 
.A1(n_4034),
.A2(n_761),
.B(n_760),
.Y(n_4660)
);

AO32x2_ASAP7_75t_L g4661 ( 
.A1(n_4082),
.A2(n_763),
.A3(n_764),
.B1(n_762),
.B2(n_761),
.Y(n_4661)
);

AOI21xp5_ASAP7_75t_L g4662 ( 
.A1(n_4392),
.A2(n_763),
.B(n_762),
.Y(n_4662)
);

NAND2xp5_ASAP7_75t_L g4663 ( 
.A(n_4124),
.B(n_762),
.Y(n_4663)
);

INVx3_ASAP7_75t_L g4664 ( 
.A(n_4079),
.Y(n_4664)
);

AO22x2_ASAP7_75t_L g4665 ( 
.A1(n_4214),
.A2(n_765),
.B1(n_766),
.B2(n_763),
.Y(n_4665)
);

AOI21x1_ASAP7_75t_SL g4666 ( 
.A1(n_4447),
.A2(n_766),
.B(n_765),
.Y(n_4666)
);

OAI21x1_ASAP7_75t_L g4667 ( 
.A1(n_4587),
.A2(n_766),
.B(n_765),
.Y(n_4667)
);

INVx1_ASAP7_75t_L g4668 ( 
.A(n_4134),
.Y(n_4668)
);

A2O1A1Ixp33_ASAP7_75t_L g4669 ( 
.A1(n_4272),
.A2(n_4232),
.B(n_4240),
.C(n_4270),
.Y(n_4669)
);

CKINVDCx5p33_ASAP7_75t_R g4670 ( 
.A(n_4037),
.Y(n_4670)
);

OAI21xp5_ASAP7_75t_SL g4671 ( 
.A1(n_4198),
.A2(n_4042),
.B(n_4043),
.Y(n_4671)
);

INVx3_ASAP7_75t_L g4672 ( 
.A(n_4144),
.Y(n_4672)
);

OAI21x1_ASAP7_75t_L g4673 ( 
.A1(n_4578),
.A2(n_768),
.B(n_767),
.Y(n_4673)
);

NAND2xp5_ASAP7_75t_L g4674 ( 
.A(n_4149),
.B(n_767),
.Y(n_4674)
);

OAI21x1_ASAP7_75t_L g4675 ( 
.A1(n_4586),
.A2(n_769),
.B(n_768),
.Y(n_4675)
);

INVx2_ASAP7_75t_L g4676 ( 
.A(n_4121),
.Y(n_4676)
);

CKINVDCx5p33_ASAP7_75t_R g4677 ( 
.A(n_4138),
.Y(n_4677)
);

INVx1_ASAP7_75t_L g4678 ( 
.A(n_4153),
.Y(n_4678)
);

A2O1A1Ixp33_ASAP7_75t_L g4679 ( 
.A1(n_4345),
.A2(n_4380),
.B(n_4396),
.C(n_4381),
.Y(n_4679)
);

OR2x2_ASAP7_75t_L g4680 ( 
.A(n_4080),
.B(n_769),
.Y(n_4680)
);

OA21x2_ASAP7_75t_L g4681 ( 
.A1(n_4506),
.A2(n_4535),
.B(n_4521),
.Y(n_4681)
);

A2O1A1Ixp33_ASAP7_75t_L g4682 ( 
.A1(n_4294),
.A2(n_770),
.B(n_771),
.C(n_769),
.Y(n_4682)
);

NAND2xp5_ASAP7_75t_L g4683 ( 
.A(n_4154),
.B(n_4166),
.Y(n_4683)
);

CKINVDCx16_ASAP7_75t_R g4684 ( 
.A(n_4129),
.Y(n_4684)
);

NAND2xp5_ASAP7_75t_L g4685 ( 
.A(n_4182),
.B(n_770),
.Y(n_4685)
);

OR2x2_ASAP7_75t_SL g4686 ( 
.A(n_4253),
.B(n_771),
.Y(n_4686)
);

INVx1_ASAP7_75t_L g4687 ( 
.A(n_4183),
.Y(n_4687)
);

INVx2_ASAP7_75t_L g4688 ( 
.A(n_4132),
.Y(n_4688)
);

AOI21xp5_ASAP7_75t_L g4689 ( 
.A1(n_4028),
.A2(n_773),
.B(n_772),
.Y(n_4689)
);

NAND2xp5_ASAP7_75t_L g4690 ( 
.A(n_4187),
.B(n_772),
.Y(n_4690)
);

INVx1_ASAP7_75t_L g4691 ( 
.A(n_4192),
.Y(n_4691)
);

NAND2xp5_ASAP7_75t_L g4692 ( 
.A(n_4211),
.B(n_773),
.Y(n_4692)
);

OAI21x1_ASAP7_75t_L g4693 ( 
.A1(n_4403),
.A2(n_774),
.B(n_773),
.Y(n_4693)
);

AOI21xp5_ASAP7_75t_L g4694 ( 
.A1(n_4534),
.A2(n_775),
.B(n_774),
.Y(n_4694)
);

AND2x4_ASAP7_75t_L g4695 ( 
.A(n_4144),
.B(n_775),
.Y(n_4695)
);

AOI21xp5_ASAP7_75t_L g4696 ( 
.A1(n_4102),
.A2(n_775),
.B(n_774),
.Y(n_4696)
);

INVx4_ASAP7_75t_L g4697 ( 
.A(n_4105),
.Y(n_4697)
);

OAI21xp5_ASAP7_75t_L g4698 ( 
.A1(n_4070),
.A2(n_777),
.B(n_776),
.Y(n_4698)
);

OR2x6_ASAP7_75t_L g4699 ( 
.A(n_4179),
.B(n_4214),
.Y(n_4699)
);

AOI21x1_ASAP7_75t_SL g4700 ( 
.A1(n_4447),
.A2(n_777),
.B(n_776),
.Y(n_4700)
);

AOI21xp5_ASAP7_75t_L g4701 ( 
.A1(n_4063),
.A2(n_778),
.B(n_777),
.Y(n_4701)
);

OAI21xp5_ASAP7_75t_L g4702 ( 
.A1(n_4293),
.A2(n_779),
.B(n_778),
.Y(n_4702)
);

BUFx12f_ASAP7_75t_L g4703 ( 
.A(n_4095),
.Y(n_4703)
);

INVx1_ASAP7_75t_L g4704 ( 
.A(n_4228),
.Y(n_4704)
);

NAND2xp5_ASAP7_75t_L g4705 ( 
.A(n_4297),
.B(n_779),
.Y(n_4705)
);

OR2x2_ASAP7_75t_L g4706 ( 
.A(n_4209),
.B(n_780),
.Y(n_4706)
);

AOI21xp5_ASAP7_75t_L g4707 ( 
.A1(n_4057),
.A2(n_781),
.B(n_780),
.Y(n_4707)
);

INVx1_ASAP7_75t_L g4708 ( 
.A(n_4205),
.Y(n_4708)
);

AND2x2_ASAP7_75t_L g4709 ( 
.A(n_4212),
.B(n_781),
.Y(n_4709)
);

INVx1_ASAP7_75t_L g4710 ( 
.A(n_4221),
.Y(n_4710)
);

INVx1_ASAP7_75t_L g4711 ( 
.A(n_4142),
.Y(n_4711)
);

OAI21x1_ASAP7_75t_L g4712 ( 
.A1(n_4250),
.A2(n_783),
.B(n_782),
.Y(n_4712)
);

AO21x2_ASAP7_75t_L g4713 ( 
.A1(n_4390),
.A2(n_783),
.B(n_782),
.Y(n_4713)
);

INVx6_ASAP7_75t_L g4714 ( 
.A(n_4083),
.Y(n_4714)
);

NAND3xp33_ASAP7_75t_SL g4715 ( 
.A(n_4368),
.B(n_70),
.C(n_71),
.Y(n_4715)
);

A2O1A1Ixp33_ASAP7_75t_L g4716 ( 
.A1(n_4336),
.A2(n_783),
.B(n_784),
.C(n_782),
.Y(n_4716)
);

NAND2xp5_ASAP7_75t_L g4717 ( 
.A(n_4306),
.B(n_784),
.Y(n_4717)
);

AOI21xp5_ASAP7_75t_L g4718 ( 
.A1(n_4057),
.A2(n_785),
.B(n_784),
.Y(n_4718)
);

OR2x2_ASAP7_75t_L g4719 ( 
.A(n_4227),
.B(n_785),
.Y(n_4719)
);

CKINVDCx5p33_ASAP7_75t_R g4720 ( 
.A(n_4246),
.Y(n_4720)
);

OAI21x1_ASAP7_75t_L g4721 ( 
.A1(n_4250),
.A2(n_787),
.B(n_786),
.Y(n_4721)
);

INVxp67_ASAP7_75t_SL g4722 ( 
.A(n_4488),
.Y(n_4722)
);

NAND2xp5_ASAP7_75t_L g4723 ( 
.A(n_4342),
.B(n_786),
.Y(n_4723)
);

NAND2xp5_ASAP7_75t_L g4724 ( 
.A(n_4371),
.B(n_787),
.Y(n_4724)
);

HB1xp67_ASAP7_75t_L g4725 ( 
.A(n_4197),
.Y(n_4725)
);

INVx1_ASAP7_75t_L g4726 ( 
.A(n_4164),
.Y(n_4726)
);

AO31x2_ASAP7_75t_L g4727 ( 
.A1(n_4529),
.A2(n_789),
.A3(n_790),
.B(n_788),
.Y(n_4727)
);

AOI22xp5_ASAP7_75t_L g4728 ( 
.A1(n_4131),
.A2(n_1100),
.B1(n_1101),
.B2(n_1097),
.Y(n_4728)
);

AOI22xp5_ASAP7_75t_L g4729 ( 
.A1(n_4238),
.A2(n_1102),
.B1(n_1106),
.B2(n_1101),
.Y(n_4729)
);

AO31x2_ASAP7_75t_L g4730 ( 
.A1(n_4484),
.A2(n_789),
.A3(n_790),
.B(n_788),
.Y(n_4730)
);

NAND2xp5_ASAP7_75t_L g4731 ( 
.A(n_4419),
.B(n_788),
.Y(n_4731)
);

CKINVDCx20_ASAP7_75t_R g4732 ( 
.A(n_4295),
.Y(n_4732)
);

O2A1O1Ixp5_ASAP7_75t_L g4733 ( 
.A1(n_4548),
.A2(n_792),
.B(n_793),
.C(n_791),
.Y(n_4733)
);

AND3x4_ASAP7_75t_L g4734 ( 
.A(n_4141),
.B(n_793),
.C(n_792),
.Y(n_4734)
);

OAI21xp33_ASAP7_75t_SL g4735 ( 
.A1(n_4123),
.A2(n_794),
.B(n_792),
.Y(n_4735)
);

AOI21xp5_ASAP7_75t_L g4736 ( 
.A1(n_4524),
.A2(n_794),
.B(n_793),
.Y(n_4736)
);

NAND2xp5_ASAP7_75t_L g4737 ( 
.A(n_4454),
.B(n_795),
.Y(n_4737)
);

AOI21xp5_ASAP7_75t_L g4738 ( 
.A1(n_4550),
.A2(n_796),
.B(n_795),
.Y(n_4738)
);

AOI22xp33_ASAP7_75t_L g4739 ( 
.A1(n_4313),
.A2(n_796),
.B1(n_797),
.B2(n_795),
.Y(n_4739)
);

NAND3x1_ASAP7_75t_L g4740 ( 
.A(n_4098),
.B(n_798),
.C(n_797),
.Y(n_4740)
);

AOI21xp5_ASAP7_75t_L g4741 ( 
.A1(n_4458),
.A2(n_798),
.B(n_797),
.Y(n_4741)
);

INVxp67_ASAP7_75t_L g4742 ( 
.A(n_4259),
.Y(n_4742)
);

OAI22xp33_ASAP7_75t_L g4743 ( 
.A1(n_4470),
.A2(n_799),
.B1(n_800),
.B2(n_798),
.Y(n_4743)
);

OA21x2_ASAP7_75t_L g4744 ( 
.A1(n_4204),
.A2(n_800),
.B(n_799),
.Y(n_4744)
);

AND2x2_ASAP7_75t_L g4745 ( 
.A(n_4235),
.B(n_799),
.Y(n_4745)
);

NAND2xp5_ASAP7_75t_L g4746 ( 
.A(n_4456),
.B(n_801),
.Y(n_4746)
);

AOI21x1_ASAP7_75t_SL g4747 ( 
.A1(n_4190),
.A2(n_802),
.B(n_801),
.Y(n_4747)
);

INVx3_ASAP7_75t_L g4748 ( 
.A(n_4207),
.Y(n_4748)
);

INVx1_ASAP7_75t_L g4749 ( 
.A(n_4177),
.Y(n_4749)
);

OAI22xp5_ASAP7_75t_L g4750 ( 
.A1(n_4045),
.A2(n_803),
.B1(n_804),
.B2(n_802),
.Y(n_4750)
);

A2O1A1Ixp33_ASAP7_75t_L g4751 ( 
.A1(n_4444),
.A2(n_804),
.B(n_805),
.C(n_803),
.Y(n_4751)
);

INVx2_ASAP7_75t_SL g4752 ( 
.A(n_4114),
.Y(n_4752)
);

INVx2_ASAP7_75t_L g4753 ( 
.A(n_4181),
.Y(n_4753)
);

INVx1_ASAP7_75t_L g4754 ( 
.A(n_4267),
.Y(n_4754)
);

AOI221x1_ASAP7_75t_L g4755 ( 
.A1(n_4279),
.A2(n_807),
.B1(n_808),
.B2(n_806),
.C(n_803),
.Y(n_4755)
);

AO31x2_ASAP7_75t_L g4756 ( 
.A1(n_4564),
.A2(n_807),
.A3(n_808),
.B(n_806),
.Y(n_4756)
);

INVx1_ASAP7_75t_L g4757 ( 
.A(n_4292),
.Y(n_4757)
);

NAND3x1_ASAP7_75t_L g4758 ( 
.A(n_4036),
.B(n_808),
.C(n_807),
.Y(n_4758)
);

AND2x4_ASAP7_75t_L g4759 ( 
.A(n_4184),
.B(n_4092),
.Y(n_4759)
);

AND2x2_ASAP7_75t_L g4760 ( 
.A(n_4249),
.B(n_809),
.Y(n_4760)
);

AOI21xp5_ASAP7_75t_L g4761 ( 
.A1(n_4068),
.A2(n_810),
.B(n_809),
.Y(n_4761)
);

AOI21xp5_ASAP7_75t_L g4762 ( 
.A1(n_4551),
.A2(n_810),
.B(n_809),
.Y(n_4762)
);

OAI21xp5_ASAP7_75t_L g4763 ( 
.A1(n_4420),
.A2(n_811),
.B(n_810),
.Y(n_4763)
);

INVx1_ASAP7_75t_L g4764 ( 
.A(n_4310),
.Y(n_4764)
);

INVx1_ASAP7_75t_L g4765 ( 
.A(n_4320),
.Y(n_4765)
);

BUFx3_ASAP7_75t_L g4766 ( 
.A(n_4234),
.Y(n_4766)
);

A2O1A1Ixp33_ASAP7_75t_L g4767 ( 
.A1(n_4274),
.A2(n_812),
.B(n_814),
.C(n_811),
.Y(n_4767)
);

O2A1O1Ixp5_ASAP7_75t_L g4768 ( 
.A1(n_4516),
.A2(n_4552),
.B(n_4401),
.C(n_4582),
.Y(n_4768)
);

NAND2xp5_ASAP7_75t_L g4769 ( 
.A(n_4468),
.B(n_811),
.Y(n_4769)
);

NOR2xp33_ASAP7_75t_L g4770 ( 
.A(n_4376),
.B(n_812),
.Y(n_4770)
);

INVx1_ASAP7_75t_L g4771 ( 
.A(n_4326),
.Y(n_4771)
);

INVx1_ASAP7_75t_L g4772 ( 
.A(n_4327),
.Y(n_4772)
);

AND2x2_ASAP7_75t_L g4773 ( 
.A(n_4282),
.B(n_812),
.Y(n_4773)
);

NOR2xp33_ASAP7_75t_L g4774 ( 
.A(n_4359),
.B(n_814),
.Y(n_4774)
);

INVxp67_ASAP7_75t_L g4775 ( 
.A(n_4155),
.Y(n_4775)
);

AND2x2_ASAP7_75t_L g4776 ( 
.A(n_4107),
.B(n_814),
.Y(n_4776)
);

AND2x4_ASAP7_75t_L g4777 ( 
.A(n_4241),
.B(n_815),
.Y(n_4777)
);

INVx1_ASAP7_75t_L g4778 ( 
.A(n_4335),
.Y(n_4778)
);

OAI21xp5_ASAP7_75t_L g4779 ( 
.A1(n_4060),
.A2(n_817),
.B(n_816),
.Y(n_4779)
);

INVxp67_ASAP7_75t_SL g4780 ( 
.A(n_4501),
.Y(n_4780)
);

AND2x2_ASAP7_75t_L g4781 ( 
.A(n_4146),
.B(n_816),
.Y(n_4781)
);

BUFx3_ASAP7_75t_L g4782 ( 
.A(n_4156),
.Y(n_4782)
);

NAND2xp5_ASAP7_75t_L g4783 ( 
.A(n_4472),
.B(n_816),
.Y(n_4783)
);

OAI21x1_ASAP7_75t_SL g4784 ( 
.A1(n_4283),
.A2(n_818),
.B(n_817),
.Y(n_4784)
);

AOI21xp5_ASAP7_75t_SL g4785 ( 
.A1(n_4496),
.A2(n_820),
.B(n_818),
.Y(n_4785)
);

INVx3_ASAP7_75t_L g4786 ( 
.A(n_4156),
.Y(n_4786)
);

BUFx6f_ASAP7_75t_L g4787 ( 
.A(n_4157),
.Y(n_4787)
);

NAND3xp33_ASAP7_75t_L g4788 ( 
.A(n_4233),
.B(n_820),
.C(n_818),
.Y(n_4788)
);

CKINVDCx8_ASAP7_75t_R g4789 ( 
.A(n_4072),
.Y(n_4789)
);

AOI21xp5_ASAP7_75t_SL g4790 ( 
.A1(n_4108),
.A2(n_821),
.B(n_820),
.Y(n_4790)
);

OA21x2_ASAP7_75t_L g4791 ( 
.A1(n_4561),
.A2(n_822),
.B(n_821),
.Y(n_4791)
);

AO21x2_ASAP7_75t_L g4792 ( 
.A1(n_4357),
.A2(n_824),
.B(n_823),
.Y(n_4792)
);

NAND3x1_ASAP7_75t_L g4793 ( 
.A(n_4243),
.B(n_824),
.C(n_823),
.Y(n_4793)
);

AOI221x1_ASAP7_75t_L g4794 ( 
.A1(n_4407),
.A2(n_825),
.B1(n_826),
.B2(n_824),
.C(n_823),
.Y(n_4794)
);

NAND2xp5_ASAP7_75t_L g4795 ( 
.A(n_4029),
.B(n_826),
.Y(n_4795)
);

OAI21xp5_ASAP7_75t_L g4796 ( 
.A1(n_4330),
.A2(n_828),
.B(n_827),
.Y(n_4796)
);

AOI21xp5_ASAP7_75t_L g4797 ( 
.A1(n_4147),
.A2(n_828),
.B(n_827),
.Y(n_4797)
);

NAND3x1_ASAP7_75t_L g4798 ( 
.A(n_4265),
.B(n_829),
.C(n_827),
.Y(n_4798)
);

AOI21xp33_ASAP7_75t_L g4799 ( 
.A1(n_4329),
.A2(n_830),
.B(n_829),
.Y(n_4799)
);

AOI21xp33_ASAP7_75t_L g4800 ( 
.A1(n_4137),
.A2(n_830),
.B(n_829),
.Y(n_4800)
);

HB1xp67_ASAP7_75t_L g4801 ( 
.A(n_4081),
.Y(n_4801)
);

AOI21xp5_ASAP7_75t_L g4802 ( 
.A1(n_4150),
.A2(n_831),
.B(n_830),
.Y(n_4802)
);

OA21x2_ASAP7_75t_L g4803 ( 
.A1(n_4366),
.A2(n_832),
.B(n_831),
.Y(n_4803)
);

AND3x4_ASAP7_75t_L g4804 ( 
.A(n_4219),
.B(n_4388),
.C(n_4412),
.Y(n_4804)
);

NAND2xp5_ASAP7_75t_L g4805 ( 
.A(n_4389),
.B(n_4430),
.Y(n_4805)
);

OAI21xp5_ASAP7_75t_SL g4806 ( 
.A1(n_4546),
.A2(n_4237),
.B(n_4093),
.Y(n_4806)
);

O2A1O1Ixp33_ASAP7_75t_L g4807 ( 
.A1(n_4076),
.A2(n_832),
.B(n_833),
.C(n_831),
.Y(n_4807)
);

INVx2_ASAP7_75t_L g4808 ( 
.A(n_4364),
.Y(n_4808)
);

CKINVDCx20_ASAP7_75t_R g4809 ( 
.A(n_4328),
.Y(n_4809)
);

AO32x2_ASAP7_75t_L g4810 ( 
.A1(n_4500),
.A2(n_834),
.A3(n_835),
.B1(n_833),
.B2(n_832),
.Y(n_4810)
);

NAND2xp5_ASAP7_75t_SL g4811 ( 
.A(n_4157),
.B(n_833),
.Y(n_4811)
);

INVx1_ASAP7_75t_L g4812 ( 
.A(n_4378),
.Y(n_4812)
);

OAI21x1_ASAP7_75t_L g4813 ( 
.A1(n_4275),
.A2(n_835),
.B(n_834),
.Y(n_4813)
);

BUFx2_ASAP7_75t_L g4814 ( 
.A(n_4072),
.Y(n_4814)
);

AOI21xp33_ASAP7_75t_L g4815 ( 
.A1(n_4251),
.A2(n_836),
.B(n_835),
.Y(n_4815)
);

NAND2xp5_ASAP7_75t_L g4816 ( 
.A(n_4065),
.B(n_836),
.Y(n_4816)
);

NAND3x1_ASAP7_75t_L g4817 ( 
.A(n_4196),
.B(n_837),
.C(n_836),
.Y(n_4817)
);

OAI21x1_ASAP7_75t_L g4818 ( 
.A1(n_4275),
.A2(n_838),
.B(n_837),
.Y(n_4818)
);

OAI22xp5_ASAP7_75t_L g4819 ( 
.A1(n_4353),
.A2(n_838),
.B1(n_839),
.B2(n_837),
.Y(n_4819)
);

INVx2_ASAP7_75t_L g4820 ( 
.A(n_4411),
.Y(n_4820)
);

OAI21x1_ASAP7_75t_L g4821 ( 
.A1(n_4278),
.A2(n_839),
.B(n_838),
.Y(n_4821)
);

OAI21xp33_ASAP7_75t_L g4822 ( 
.A1(n_4075),
.A2(n_841),
.B(n_840),
.Y(n_4822)
);

OAI21x1_ASAP7_75t_L g4823 ( 
.A1(n_4278),
.A2(n_4393),
.B(n_4319),
.Y(n_4823)
);

INVx1_ASAP7_75t_L g4824 ( 
.A(n_4413),
.Y(n_4824)
);

OAI21xp33_ASAP7_75t_L g4825 ( 
.A1(n_4286),
.A2(n_842),
.B(n_840),
.Y(n_4825)
);

NOR2xp33_ASAP7_75t_L g4826 ( 
.A(n_4140),
.B(n_842),
.Y(n_4826)
);

AO31x2_ASAP7_75t_L g4827 ( 
.A1(n_4397),
.A2(n_843),
.A3(n_844),
.B(n_842),
.Y(n_4827)
);

OAI22xp5_ASAP7_75t_L g4828 ( 
.A1(n_4165),
.A2(n_844),
.B1(n_845),
.B2(n_843),
.Y(n_4828)
);

INVx1_ASAP7_75t_L g4829 ( 
.A(n_4231),
.Y(n_4829)
);

INVx1_ASAP7_75t_L g4830 ( 
.A(n_4193),
.Y(n_4830)
);

AOI221xp5_ASAP7_75t_SL g4831 ( 
.A1(n_4369),
.A2(n_73),
.B1(n_71),
.B2(n_72),
.C(n_74),
.Y(n_4831)
);

NAND2xp5_ASAP7_75t_L g4832 ( 
.A(n_4066),
.B(n_843),
.Y(n_4832)
);

NOR2xp33_ASAP7_75t_SL g4833 ( 
.A(n_4032),
.B(n_1089),
.Y(n_4833)
);

OAI21x1_ASAP7_75t_L g4834 ( 
.A1(n_4319),
.A2(n_845),
.B(n_844),
.Y(n_4834)
);

OAI22xp5_ASAP7_75t_L g4835 ( 
.A1(n_4583),
.A2(n_846),
.B1(n_847),
.B2(n_845),
.Y(n_4835)
);

NAND2xp5_ASAP7_75t_L g4836 ( 
.A(n_4482),
.B(n_848),
.Y(n_4836)
);

NAND2xp5_ASAP7_75t_L g4837 ( 
.A(n_4120),
.B(n_848),
.Y(n_4837)
);

INVxp67_ASAP7_75t_SL g4838 ( 
.A(n_4230),
.Y(n_4838)
);

INVx3_ASAP7_75t_SL g4839 ( 
.A(n_4178),
.Y(n_4839)
);

A2O1A1Ixp33_ASAP7_75t_L g4840 ( 
.A1(n_4532),
.A2(n_849),
.B(n_850),
.C(n_848),
.Y(n_4840)
);

A2O1A1Ixp33_ASAP7_75t_L g4841 ( 
.A1(n_4449),
.A2(n_850),
.B(n_851),
.C(n_849),
.Y(n_4841)
);

INVx1_ASAP7_75t_L g4842 ( 
.A(n_4088),
.Y(n_4842)
);

NAND2xp5_ASAP7_75t_L g4843 ( 
.A(n_4112),
.B(n_851),
.Y(n_4843)
);

INVx5_ASAP7_75t_L g4844 ( 
.A(n_4072),
.Y(n_4844)
);

OAI21x1_ASAP7_75t_L g4845 ( 
.A1(n_4393),
.A2(n_852),
.B(n_851),
.Y(n_4845)
);

OAI21x1_ASAP7_75t_L g4846 ( 
.A1(n_4479),
.A2(n_853),
.B(n_852),
.Y(n_4846)
);

CKINVDCx12_ASAP7_75t_R g4847 ( 
.A(n_4169),
.Y(n_4847)
);

NOR2xp33_ASAP7_75t_L g4848 ( 
.A(n_4030),
.B(n_853),
.Y(n_4848)
);

OAI21x1_ASAP7_75t_SL g4849 ( 
.A1(n_4341),
.A2(n_4354),
.B(n_4352),
.Y(n_4849)
);

OAI21x1_ASAP7_75t_L g4850 ( 
.A1(n_4479),
.A2(n_854),
.B(n_853),
.Y(n_4850)
);

AOI21xp5_ASAP7_75t_L g4851 ( 
.A1(n_4558),
.A2(n_855),
.B(n_854),
.Y(n_4851)
);

INVx2_ASAP7_75t_L g4852 ( 
.A(n_4391),
.Y(n_4852)
);

AOI21xp5_ASAP7_75t_L g4853 ( 
.A1(n_4558),
.A2(n_855),
.B(n_854),
.Y(n_4853)
);

OAI21x1_ASAP7_75t_L g4854 ( 
.A1(n_4526),
.A2(n_856),
.B(n_855),
.Y(n_4854)
);

BUFx6f_ASAP7_75t_L g4855 ( 
.A(n_4157),
.Y(n_4855)
);

AOI21xp5_ASAP7_75t_L g4856 ( 
.A1(n_4558),
.A2(n_857),
.B(n_856),
.Y(n_4856)
);

NAND2xp5_ASAP7_75t_L g4857 ( 
.A(n_4078),
.B(n_856),
.Y(n_4857)
);

AO31x2_ASAP7_75t_L g4858 ( 
.A1(n_4522),
.A2(n_858),
.A3(n_859),
.B(n_857),
.Y(n_4858)
);

INVx1_ASAP7_75t_L g4859 ( 
.A(n_4291),
.Y(n_4859)
);

OAI21xp5_ASAP7_75t_L g4860 ( 
.A1(n_4480),
.A2(n_858),
.B(n_857),
.Y(n_4860)
);

AO21x2_ASAP7_75t_L g4861 ( 
.A1(n_4499),
.A2(n_859),
.B(n_858),
.Y(n_4861)
);

NAND2xp5_ASAP7_75t_L g4862 ( 
.A(n_4106),
.B(n_860),
.Y(n_4862)
);

NAND2xp5_ASAP7_75t_L g4863 ( 
.A(n_4110),
.B(n_860),
.Y(n_4863)
);

INVx2_ASAP7_75t_L g4864 ( 
.A(n_4291),
.Y(n_4864)
);

NAND2xp5_ASAP7_75t_L g4865 ( 
.A(n_4152),
.B(n_4133),
.Y(n_4865)
);

OAI21x1_ASAP7_75t_L g4866 ( 
.A1(n_4160),
.A2(n_861),
.B(n_860),
.Y(n_4866)
);

AOI21x1_ASAP7_75t_SL g4867 ( 
.A1(n_4191),
.A2(n_862),
.B(n_861),
.Y(n_4867)
);

NOR2xp67_ASAP7_75t_L g4868 ( 
.A(n_4175),
.B(n_862),
.Y(n_4868)
);

INVx2_ASAP7_75t_L g4869 ( 
.A(n_4302),
.Y(n_4869)
);

AO21x2_ASAP7_75t_L g4870 ( 
.A1(n_4509),
.A2(n_863),
.B(n_861),
.Y(n_4870)
);

O2A1O1Ixp33_ASAP7_75t_SL g4871 ( 
.A1(n_4254),
.A2(n_864),
.B(n_865),
.C(n_863),
.Y(n_4871)
);

NOR2x1_ASAP7_75t_SL g4872 ( 
.A(n_4040),
.B(n_864),
.Y(n_4872)
);

AO31x2_ASAP7_75t_L g4873 ( 
.A1(n_4533),
.A2(n_865),
.A3(n_866),
.B(n_864),
.Y(n_4873)
);

CKINVDCx5p33_ASAP7_75t_R g4874 ( 
.A(n_4549),
.Y(n_4874)
);

INVx1_ASAP7_75t_SL g4875 ( 
.A(n_4175),
.Y(n_4875)
);

INVx2_ASAP7_75t_L g4876 ( 
.A(n_4302),
.Y(n_4876)
);

NOR2x1_ASAP7_75t_SL g4877 ( 
.A(n_4040),
.B(n_4047),
.Y(n_4877)
);

NOR2x1_ASAP7_75t_L g4878 ( 
.A(n_4263),
.B(n_865),
.Y(n_4878)
);

OAI21xp5_ASAP7_75t_L g4879 ( 
.A1(n_4367),
.A2(n_868),
.B(n_867),
.Y(n_4879)
);

NAND2xp5_ASAP7_75t_SL g4880 ( 
.A(n_4175),
.B(n_867),
.Y(n_4880)
);

AND2x2_ASAP7_75t_L g4881 ( 
.A(n_4337),
.B(n_867),
.Y(n_4881)
);

OAI22xp5_ASAP7_75t_L g4882 ( 
.A1(n_4188),
.A2(n_869),
.B1(n_870),
.B2(n_868),
.Y(n_4882)
);

NAND2xp5_ASAP7_75t_L g4883 ( 
.A(n_4431),
.B(n_868),
.Y(n_4883)
);

OAI21x1_ASAP7_75t_L g4884 ( 
.A1(n_4125),
.A2(n_870),
.B(n_869),
.Y(n_4884)
);

OAI21x1_ASAP7_75t_L g4885 ( 
.A1(n_4173),
.A2(n_871),
.B(n_869),
.Y(n_4885)
);

INVx1_ASAP7_75t_L g4886 ( 
.A(n_4377),
.Y(n_4886)
);

INVx1_ASAP7_75t_L g4887 ( 
.A(n_4377),
.Y(n_4887)
);

NAND2xp5_ASAP7_75t_L g4888 ( 
.A(n_4437),
.B(n_871),
.Y(n_4888)
);

AOI221xp5_ASAP7_75t_L g4889 ( 
.A1(n_4460),
.A2(n_873),
.B1(n_874),
.B2(n_872),
.C(n_871),
.Y(n_4889)
);

INVx1_ASAP7_75t_L g4890 ( 
.A(n_4384),
.Y(n_4890)
);

NAND2xp5_ASAP7_75t_L g4891 ( 
.A(n_4466),
.B(n_873),
.Y(n_4891)
);

INVx3_ASAP7_75t_L g4892 ( 
.A(n_4178),
.Y(n_4892)
);

BUFx4f_ASAP7_75t_L g4893 ( 
.A(n_4072),
.Y(n_4893)
);

NOR2xp33_ASAP7_75t_L g4894 ( 
.A(n_4143),
.B(n_873),
.Y(n_4894)
);

OAI21x1_ASAP7_75t_L g4895 ( 
.A1(n_4348),
.A2(n_875),
.B(n_874),
.Y(n_4895)
);

AO31x2_ASAP7_75t_L g4896 ( 
.A1(n_4139),
.A2(n_4321),
.A3(n_4445),
.B(n_4236),
.Y(n_4896)
);

INVx1_ASAP7_75t_L g4897 ( 
.A(n_4384),
.Y(n_4897)
);

OAI21x1_ASAP7_75t_L g4898 ( 
.A1(n_4425),
.A2(n_876),
.B(n_875),
.Y(n_4898)
);

OAI21x1_ASAP7_75t_L g4899 ( 
.A1(n_4085),
.A2(n_876),
.B(n_875),
.Y(n_4899)
);

INVx1_ASAP7_75t_L g4900 ( 
.A(n_4263),
.Y(n_4900)
);

OAI22xp5_ASAP7_75t_L g4901 ( 
.A1(n_4537),
.A2(n_4360),
.B1(n_4365),
.B2(n_4035),
.Y(n_4901)
);

INVx1_ASAP7_75t_SL g4902 ( 
.A(n_4347),
.Y(n_4902)
);

AOI21xp5_ASAP7_75t_L g4903 ( 
.A1(n_4159),
.A2(n_877),
.B(n_876),
.Y(n_4903)
);

NAND3xp33_ASAP7_75t_L g4904 ( 
.A(n_4298),
.B(n_878),
.C(n_877),
.Y(n_4904)
);

INVx1_ASAP7_75t_L g4905 ( 
.A(n_4462),
.Y(n_4905)
);

INVx1_ASAP7_75t_L g4906 ( 
.A(n_4462),
.Y(n_4906)
);

OAI21x1_ASAP7_75t_L g4907 ( 
.A1(n_4086),
.A2(n_879),
.B(n_878),
.Y(n_4907)
);

OAI21xp5_ASAP7_75t_L g4908 ( 
.A1(n_4373),
.A2(n_880),
.B(n_879),
.Y(n_4908)
);

NAND3x1_ASAP7_75t_L g4909 ( 
.A(n_4200),
.B(n_881),
.C(n_880),
.Y(n_4909)
);

OAI21xp5_ASAP7_75t_L g4910 ( 
.A1(n_4400),
.A2(n_4226),
.B(n_4394),
.Y(n_4910)
);

BUFx3_ASAP7_75t_L g4911 ( 
.A(n_4185),
.Y(n_4911)
);

INVx2_ASAP7_75t_SL g4912 ( 
.A(n_4185),
.Y(n_4912)
);

OAI22xp5_ASAP7_75t_L g4913 ( 
.A1(n_4556),
.A2(n_881),
.B1(n_882),
.B2(n_880),
.Y(n_4913)
);

AO31x2_ASAP7_75t_L g4914 ( 
.A1(n_4236),
.A2(n_882),
.A3(n_883),
.B(n_881),
.Y(n_4914)
);

OAI21x1_ASAP7_75t_L g4915 ( 
.A1(n_4096),
.A2(n_883),
.B(n_882),
.Y(n_4915)
);

HB1xp67_ASAP7_75t_L g4916 ( 
.A(n_4290),
.Y(n_4916)
);

OAI22xp5_ASAP7_75t_L g4917 ( 
.A1(n_4262),
.A2(n_884),
.B1(n_885),
.B2(n_883),
.Y(n_4917)
);

A2O1A1Ixp33_ASAP7_75t_L g4918 ( 
.A1(n_4465),
.A2(n_885),
.B(n_886),
.C(n_884),
.Y(n_4918)
);

AOI21xp33_ASAP7_75t_L g4919 ( 
.A1(n_4094),
.A2(n_885),
.B(n_884),
.Y(n_4919)
);

AOI21xp5_ASAP7_75t_L g4920 ( 
.A1(n_4051),
.A2(n_887),
.B(n_886),
.Y(n_4920)
);

NAND2xp5_ASAP7_75t_L g4921 ( 
.A(n_4215),
.B(n_4346),
.Y(n_4921)
);

NOR2x1_ASAP7_75t_SL g4922 ( 
.A(n_4040),
.B(n_886),
.Y(n_4922)
);

AOI21xp5_ASAP7_75t_L g4923 ( 
.A1(n_4053),
.A2(n_888),
.B(n_887),
.Y(n_4923)
);

INVx2_ASAP7_75t_L g4924 ( 
.A(n_4451),
.Y(n_4924)
);

AND2x2_ASAP7_75t_L g4925 ( 
.A(n_4387),
.B(n_888),
.Y(n_4925)
);

NAND2xp5_ASAP7_75t_L g4926 ( 
.A(n_4113),
.B(n_888),
.Y(n_4926)
);

OR2x2_ASAP7_75t_L g4927 ( 
.A(n_4299),
.B(n_889),
.Y(n_4927)
);

AO31x2_ASAP7_75t_L g4928 ( 
.A1(n_4321),
.A2(n_4445),
.A3(n_4464),
.B(n_4450),
.Y(n_4928)
);

INVx2_ASAP7_75t_L g4929 ( 
.A(n_4508),
.Y(n_4929)
);

NAND3xp33_ASAP7_75t_L g4930 ( 
.A(n_4424),
.B(n_890),
.C(n_889),
.Y(n_4930)
);

AO31x2_ASAP7_75t_L g4931 ( 
.A1(n_4473),
.A2(n_890),
.A3(n_891),
.B(n_889),
.Y(n_4931)
);

AOI21xp5_ASAP7_75t_L g4932 ( 
.A1(n_4056),
.A2(n_891),
.B(n_890),
.Y(n_4932)
);

NAND3x1_ASAP7_75t_L g4933 ( 
.A(n_4225),
.B(n_892),
.C(n_891),
.Y(n_4933)
);

NAND2xp5_ASAP7_75t_L g4934 ( 
.A(n_4436),
.B(n_4457),
.Y(n_4934)
);

OAI21x1_ASAP7_75t_L g4935 ( 
.A1(n_4172),
.A2(n_893),
.B(n_892),
.Y(n_4935)
);

OAI21x1_ASAP7_75t_L g4936 ( 
.A1(n_4281),
.A2(n_894),
.B(n_893),
.Y(n_4936)
);

AND2x4_ASAP7_75t_L g4937 ( 
.A(n_4280),
.B(n_894),
.Y(n_4937)
);

OAI22xp5_ASAP7_75t_L g4938 ( 
.A1(n_4284),
.A2(n_895),
.B1(n_896),
.B2(n_894),
.Y(n_4938)
);

AND2x2_ASAP7_75t_L g4939 ( 
.A(n_4417),
.B(n_896),
.Y(n_4939)
);

INVx3_ASAP7_75t_L g4940 ( 
.A(n_4309),
.Y(n_4940)
);

NOR2xp67_ASAP7_75t_SL g4941 ( 
.A(n_4347),
.B(n_896),
.Y(n_4941)
);

INVx3_ASAP7_75t_L g4942 ( 
.A(n_4399),
.Y(n_4942)
);

NAND2xp5_ASAP7_75t_L g4943 ( 
.A(n_4104),
.B(n_897),
.Y(n_4943)
);

NAND2xp5_ASAP7_75t_L g4944 ( 
.A(n_4048),
.B(n_897),
.Y(n_4944)
);

AOI211x1_ASAP7_75t_L g4945 ( 
.A1(n_4049),
.A2(n_898),
.B(n_899),
.C(n_897),
.Y(n_4945)
);

INVx1_ASAP7_75t_L g4946 ( 
.A(n_4527),
.Y(n_4946)
);

AO31x2_ASAP7_75t_L g4947 ( 
.A1(n_4474),
.A2(n_899),
.A3(n_900),
.B(n_898),
.Y(n_4947)
);

O2A1O1Ixp33_ASAP7_75t_L g4948 ( 
.A1(n_4115),
.A2(n_901),
.B(n_902),
.C(n_898),
.Y(n_4948)
);

INVx1_ASAP7_75t_L g4949 ( 
.A(n_4569),
.Y(n_4949)
);

NAND2xp5_ASAP7_75t_L g4950 ( 
.A(n_4242),
.B(n_901),
.Y(n_4950)
);

INVx1_ASAP7_75t_L g4951 ( 
.A(n_4476),
.Y(n_4951)
);

OAI21x1_ASAP7_75t_L g4952 ( 
.A1(n_4151),
.A2(n_903),
.B(n_902),
.Y(n_4952)
);

NAND2xp5_ASAP7_75t_L g4953 ( 
.A(n_4247),
.B(n_903),
.Y(n_4953)
);

AOI21xp5_ASAP7_75t_L g4954 ( 
.A1(n_4542),
.A2(n_904),
.B(n_903),
.Y(n_4954)
);

OAI21x1_ASAP7_75t_L g4955 ( 
.A1(n_4340),
.A2(n_905),
.B(n_904),
.Y(n_4955)
);

OA21x2_ASAP7_75t_L g4956 ( 
.A1(n_4513),
.A2(n_905),
.B(n_904),
.Y(n_4956)
);

CKINVDCx5p33_ASAP7_75t_R g4957 ( 
.A(n_4122),
.Y(n_4957)
);

INVx1_ASAP7_75t_L g4958 ( 
.A(n_4567),
.Y(n_4958)
);

INVxp67_ASAP7_75t_L g4959 ( 
.A(n_4355),
.Y(n_4959)
);

BUFx8_ASAP7_75t_L g4960 ( 
.A(n_4492),
.Y(n_4960)
);

INVx4_ASAP7_75t_L g4961 ( 
.A(n_4347),
.Y(n_4961)
);

BUFx6f_ASAP7_75t_L g4962 ( 
.A(n_4077),
.Y(n_4962)
);

AOI31xp67_ASAP7_75t_L g4963 ( 
.A1(n_4276),
.A2(n_906),
.A3(n_907),
.B(n_905),
.Y(n_4963)
);

AOI21xp5_ASAP7_75t_L g4964 ( 
.A1(n_4314),
.A2(n_907),
.B(n_906),
.Y(n_4964)
);

AO31x2_ASAP7_75t_L g4965 ( 
.A1(n_4503),
.A2(n_908),
.A3(n_909),
.B(n_907),
.Y(n_4965)
);

NAND2xp5_ASAP7_75t_L g4966 ( 
.A(n_4264),
.B(n_908),
.Y(n_4966)
);

OAI22xp5_ASAP7_75t_L g4967 ( 
.A1(n_4248),
.A2(n_910),
.B1(n_911),
.B2(n_909),
.Y(n_4967)
);

AND2x4_ASAP7_75t_L g4968 ( 
.A(n_4158),
.B(n_909),
.Y(n_4968)
);

NOR2xp67_ASAP7_75t_SL g4969 ( 
.A(n_4244),
.B(n_910),
.Y(n_4969)
);

AOI21xp5_ASAP7_75t_L g4970 ( 
.A1(n_4491),
.A2(n_911),
.B(n_910),
.Y(n_4970)
);

NAND2xp5_ASAP7_75t_L g4971 ( 
.A(n_4426),
.B(n_911),
.Y(n_4971)
);

NOR2xp33_ASAP7_75t_L g4972 ( 
.A(n_4130),
.B(n_912),
.Y(n_4972)
);

INVx4_ASAP7_75t_L g4973 ( 
.A(n_4077),
.Y(n_4973)
);

BUFx5_ASAP7_75t_L g4974 ( 
.A(n_4566),
.Y(n_4974)
);

NAND2xp5_ASAP7_75t_L g4975 ( 
.A(n_4435),
.B(n_912),
.Y(n_4975)
);

OAI21xp5_ASAP7_75t_SL g4976 ( 
.A1(n_4362),
.A2(n_914),
.B(n_913),
.Y(n_4976)
);

AO31x2_ASAP7_75t_L g4977 ( 
.A1(n_4307),
.A2(n_914),
.A3(n_915),
.B(n_913),
.Y(n_4977)
);

BUFx2_ASAP7_75t_L g4978 ( 
.A(n_4273),
.Y(n_4978)
);

AOI21xp5_ASAP7_75t_L g4979 ( 
.A1(n_4502),
.A2(n_915),
.B(n_913),
.Y(n_4979)
);

OAI21x1_ASAP7_75t_L g4980 ( 
.A1(n_4161),
.A2(n_916),
.B(n_915),
.Y(n_4980)
);

OR2x2_ASAP7_75t_L g4981 ( 
.A(n_4301),
.B(n_916),
.Y(n_4981)
);

INVx1_ASAP7_75t_L g4982 ( 
.A(n_4305),
.Y(n_4982)
);

AO21x1_ASAP7_75t_L g4983 ( 
.A1(n_4344),
.A2(n_917),
.B(n_916),
.Y(n_4983)
);

BUFx2_ASAP7_75t_L g4984 ( 
.A(n_4317),
.Y(n_4984)
);

BUFx2_ASAP7_75t_SL g4985 ( 
.A(n_4338),
.Y(n_4985)
);

AOI221xp5_ASAP7_75t_L g4986 ( 
.A1(n_4438),
.A2(n_919),
.B1(n_920),
.B2(n_918),
.C(n_917),
.Y(n_4986)
);

NAND3xp33_ASAP7_75t_L g4987 ( 
.A(n_4439),
.B(n_4448),
.C(n_4440),
.Y(n_4987)
);

OAI21x1_ASAP7_75t_L g4988 ( 
.A1(n_4174),
.A2(n_4414),
.B(n_4058),
.Y(n_4988)
);

INVx1_ASAP7_75t_L g4989 ( 
.A(n_4356),
.Y(n_4989)
);

OAI21x1_ASAP7_75t_L g4990 ( 
.A1(n_4584),
.A2(n_919),
.B(n_918),
.Y(n_4990)
);

OAI22xp5_ASAP7_75t_L g4991 ( 
.A1(n_4363),
.A2(n_920),
.B1(n_921),
.B2(n_918),
.Y(n_4991)
);

OAI21xp5_ASAP7_75t_L g4992 ( 
.A1(n_4494),
.A2(n_922),
.B(n_921),
.Y(n_4992)
);

AOI21xp33_ASAP7_75t_L g4993 ( 
.A1(n_4101),
.A2(n_923),
.B(n_922),
.Y(n_4993)
);

AND2x4_ASAP7_75t_L g4994 ( 
.A(n_4374),
.B(n_4528),
.Y(n_4994)
);

INVx1_ASAP7_75t_L g4995 ( 
.A(n_4498),
.Y(n_4995)
);

AO31x2_ASAP7_75t_L g4996 ( 
.A1(n_4135),
.A2(n_4382),
.A3(n_4372),
.B(n_4573),
.Y(n_4996)
);

AND2x6_ASAP7_75t_L g4997 ( 
.A(n_4585),
.B(n_922),
.Y(n_4997)
);

OAI21x1_ASAP7_75t_L g4998 ( 
.A1(n_4136),
.A2(n_924),
.B(n_923),
.Y(n_4998)
);

NAND2xp5_ASAP7_75t_L g4999 ( 
.A(n_4463),
.B(n_923),
.Y(n_4999)
);

INVx1_ASAP7_75t_L g5000 ( 
.A(n_4530),
.Y(n_5000)
);

OAI21x1_ASAP7_75t_L g5001 ( 
.A1(n_4176),
.A2(n_925),
.B(n_924),
.Y(n_5001)
);

AOI21xp5_ASAP7_75t_L g5002 ( 
.A1(n_4077),
.A2(n_925),
.B(n_924),
.Y(n_5002)
);

NOR2xp33_ASAP7_75t_L g5003 ( 
.A(n_4467),
.B(n_4162),
.Y(n_5003)
);

INVx5_ASAP7_75t_L g5004 ( 
.A(n_4186),
.Y(n_5004)
);

AOI21xp5_ASAP7_75t_L g5005 ( 
.A1(n_4186),
.A2(n_926),
.B(n_925),
.Y(n_5005)
);

OAI21x1_ASAP7_75t_L g5006 ( 
.A1(n_4574),
.A2(n_927),
.B(n_926),
.Y(n_5006)
);

OAI21x1_ASAP7_75t_L g5007 ( 
.A1(n_4579),
.A2(n_927),
.B(n_926),
.Y(n_5007)
);

INVx1_ASAP7_75t_L g5008 ( 
.A(n_4222),
.Y(n_5008)
);

OAI21x1_ASAP7_75t_L g5009 ( 
.A1(n_4581),
.A2(n_928),
.B(n_927),
.Y(n_5009)
);

CKINVDCx5p33_ASAP7_75t_R g5010 ( 
.A(n_4318),
.Y(n_5010)
);

INVx1_ASAP7_75t_L g5011 ( 
.A(n_4528),
.Y(n_5011)
);

O2A1O1Ixp5_ASAP7_75t_L g5012 ( 
.A1(n_4315),
.A2(n_929),
.B(n_930),
.C(n_928),
.Y(n_5012)
);

AOI21xp5_ASAP7_75t_L g5013 ( 
.A1(n_4186),
.A2(n_930),
.B(n_928),
.Y(n_5013)
);

HB1xp67_ASAP7_75t_L g5014 ( 
.A(n_4206),
.Y(n_5014)
);

BUFx10_ASAP7_75t_L g5015 ( 
.A(n_4541),
.Y(n_5015)
);

NAND2xp5_ASAP7_75t_L g5016 ( 
.A(n_4525),
.B(n_931),
.Y(n_5016)
);

OAI21x1_ASAP7_75t_L g5017 ( 
.A1(n_4453),
.A2(n_932),
.B(n_931),
.Y(n_5017)
);

INVx1_ASAP7_75t_SL g5018 ( 
.A(n_4206),
.Y(n_5018)
);

AO21x1_ASAP7_75t_L g5019 ( 
.A1(n_4511),
.A2(n_932),
.B(n_931),
.Y(n_5019)
);

NOR2x1_ASAP7_75t_R g5020 ( 
.A(n_4541),
.B(n_932),
.Y(n_5020)
);

AOI221x1_ASAP7_75t_L g5021 ( 
.A1(n_4054),
.A2(n_935),
.B1(n_936),
.B2(n_934),
.C(n_933),
.Y(n_5021)
);

OA21x2_ASAP7_75t_L g5022 ( 
.A1(n_4514),
.A2(n_934),
.B(n_933),
.Y(n_5022)
);

AND2x4_ASAP7_75t_L g5023 ( 
.A(n_4126),
.B(n_933),
.Y(n_5023)
);

NAND2xp5_ASAP7_75t_L g5024 ( 
.A(n_4213),
.B(n_4486),
.Y(n_5024)
);

INVx2_ASAP7_75t_L g5025 ( 
.A(n_4206),
.Y(n_5025)
);

NAND2xp5_ASAP7_75t_L g5026 ( 
.A(n_4568),
.B(n_935),
.Y(n_5026)
);

NOR3xp33_ASAP7_75t_L g5027 ( 
.A(n_4563),
.B(n_936),
.C(n_935),
.Y(n_5027)
);

NAND2xp5_ASAP7_75t_L g5028 ( 
.A(n_4210),
.B(n_937),
.Y(n_5028)
);

OAI21x1_ASAP7_75t_L g5029 ( 
.A1(n_4469),
.A2(n_4471),
.B(n_4333),
.Y(n_5029)
);

AOI21xp5_ASAP7_75t_L g5030 ( 
.A1(n_4277),
.A2(n_938),
.B(n_937),
.Y(n_5030)
);

OAI21x1_ASAP7_75t_L g5031 ( 
.A1(n_4316),
.A2(n_939),
.B(n_938),
.Y(n_5031)
);

INVx2_ASAP7_75t_L g5032 ( 
.A(n_4277),
.Y(n_5032)
);

BUFx10_ASAP7_75t_L g5033 ( 
.A(n_4277),
.Y(n_5033)
);

NAND2xp5_ASAP7_75t_L g5034 ( 
.A(n_4505),
.B(n_938),
.Y(n_5034)
);

OAI21x1_ASAP7_75t_L g5035 ( 
.A1(n_4343),
.A2(n_4408),
.B(n_4379),
.Y(n_5035)
);

NAND2xp5_ASAP7_75t_SL g5036 ( 
.A(n_4296),
.B(n_4331),
.Y(n_5036)
);

OAI21x1_ASAP7_75t_L g5037 ( 
.A1(n_4421),
.A2(n_940),
.B(n_939),
.Y(n_5037)
);

AOI21xp5_ASAP7_75t_L g5038 ( 
.A1(n_4296),
.A2(n_4349),
.B(n_4331),
.Y(n_5038)
);

AOI21xp5_ASAP7_75t_L g5039 ( 
.A1(n_4296),
.A2(n_941),
.B(n_939),
.Y(n_5039)
);

NAND2xp5_ASAP7_75t_L g5040 ( 
.A(n_4507),
.B(n_941),
.Y(n_5040)
);

AO31x2_ASAP7_75t_L g5041 ( 
.A1(n_4575),
.A2(n_943),
.A3(n_944),
.B(n_942),
.Y(n_5041)
);

O2A1O1Ixp5_ASAP7_75t_SL g5042 ( 
.A1(n_4423),
.A2(n_944),
.B(n_945),
.C(n_942),
.Y(n_5042)
);

A2O1A1Ixp33_ASAP7_75t_L g5043 ( 
.A1(n_4517),
.A2(n_4553),
.B(n_4547),
.C(n_4189),
.Y(n_5043)
);

BUFx12f_ASAP7_75t_L g5044 ( 
.A(n_4566),
.Y(n_5044)
);

INVx1_ASAP7_75t_L g5045 ( 
.A(n_4432),
.Y(n_5045)
);

OR2x2_ASAP7_75t_L g5046 ( 
.A(n_4409),
.B(n_944),
.Y(n_5046)
);

AOI31xp67_ASAP7_75t_L g5047 ( 
.A1(n_4442),
.A2(n_946),
.A3(n_947),
.B(n_945),
.Y(n_5047)
);

AOI21xp5_ASAP7_75t_L g5048 ( 
.A1(n_4331),
.A2(n_946),
.B(n_945),
.Y(n_5048)
);

HB1xp67_ASAP7_75t_L g5049 ( 
.A(n_4349),
.Y(n_5049)
);

OAI21xp5_ASAP7_75t_SL g5050 ( 
.A1(n_4410),
.A2(n_947),
.B(n_946),
.Y(n_5050)
);

NOR2xp33_ASAP7_75t_L g5051 ( 
.A(n_4271),
.B(n_947),
.Y(n_5051)
);

INVx2_ASAP7_75t_L g5052 ( 
.A(n_4349),
.Y(n_5052)
);

NAND3x1_ASAP7_75t_L g5053 ( 
.A(n_4515),
.B(n_949),
.C(n_948),
.Y(n_5053)
);

OAI21x1_ASAP7_75t_L g5054 ( 
.A1(n_4446),
.A2(n_949),
.B(n_948),
.Y(n_5054)
);

OAI21x1_ASAP7_75t_L g5055 ( 
.A1(n_4490),
.A2(n_950),
.B(n_948),
.Y(n_5055)
);

NAND2xp5_ASAP7_75t_L g5056 ( 
.A(n_4287),
.B(n_950),
.Y(n_5056)
);

AOI21x1_ASAP7_75t_L g5057 ( 
.A1(n_4170),
.A2(n_952),
.B(n_951),
.Y(n_5057)
);

INVx1_ASAP7_75t_L g5058 ( 
.A(n_4433),
.Y(n_5058)
);

OR2x6_ASAP7_75t_L g5059 ( 
.A(n_4245),
.B(n_951),
.Y(n_5059)
);

AOI21x1_ASAP7_75t_SL g5060 ( 
.A1(n_4268),
.A2(n_952),
.B(n_951),
.Y(n_5060)
);

NAND2xp5_ASAP7_75t_L g5061 ( 
.A(n_4358),
.B(n_952),
.Y(n_5061)
);

INVx1_ASAP7_75t_L g5062 ( 
.A(n_4434),
.Y(n_5062)
);

A2O1A1Ixp33_ASAP7_75t_L g5063 ( 
.A1(n_4418),
.A2(n_954),
.B(n_955),
.C(n_953),
.Y(n_5063)
);

AOI21xp5_ASAP7_75t_L g5064 ( 
.A1(n_4361),
.A2(n_954),
.B(n_953),
.Y(n_5064)
);

OAI22xp5_ASAP7_75t_L g5065 ( 
.A1(n_4312),
.A2(n_956),
.B1(n_957),
.B2(n_954),
.Y(n_5065)
);

INVx2_ASAP7_75t_L g5066 ( 
.A(n_4361),
.Y(n_5066)
);

INVx1_ASAP7_75t_L g5067 ( 
.A(n_4617),
.Y(n_5067)
);

INVx4_ASAP7_75t_SL g5068 ( 
.A(n_4639),
.Y(n_5068)
);

OAI21x1_ASAP7_75t_L g5069 ( 
.A1(n_4635),
.A2(n_4493),
.B(n_4415),
.Y(n_5069)
);

INVx6_ASAP7_75t_L g5070 ( 
.A(n_4606),
.Y(n_5070)
);

INVx2_ASAP7_75t_SL g5071 ( 
.A(n_4606),
.Y(n_5071)
);

OAI21xp5_ASAP7_75t_L g5072 ( 
.A1(n_4594),
.A2(n_4255),
.B(n_4239),
.Y(n_5072)
);

AOI221xp5_ASAP7_75t_L g5073 ( 
.A1(n_4750),
.A2(n_4195),
.B1(n_4194),
.B2(n_4260),
.C(n_4229),
.Y(n_5073)
);

INVx1_ASAP7_75t_L g5074 ( 
.A(n_4644),
.Y(n_5074)
);

AO21x2_ASAP7_75t_L g5075 ( 
.A1(n_4851),
.A2(n_4322),
.B(n_4311),
.Y(n_5075)
);

INVx1_ASAP7_75t_L g5076 ( 
.A(n_4647),
.Y(n_5076)
);

AOI21xp5_ASAP7_75t_L g5077 ( 
.A1(n_4893),
.A2(n_4203),
.B(n_4361),
.Y(n_5077)
);

INVx1_ASAP7_75t_SL g5078 ( 
.A(n_4714),
.Y(n_5078)
);

OAI21x1_ASAP7_75t_L g5079 ( 
.A1(n_4988),
.A2(n_4416),
.B(n_4572),
.Y(n_5079)
);

AOI22xp33_ASAP7_75t_L g5080 ( 
.A1(n_4626),
.A2(n_4566),
.B1(n_4285),
.B2(n_4571),
.Y(n_5080)
);

BUFx6f_ASAP7_75t_L g5081 ( 
.A(n_4787),
.Y(n_5081)
);

BUFx10_ASAP7_75t_L g5082 ( 
.A(n_4608),
.Y(n_5082)
);

NAND2xp5_ASAP7_75t_L g5083 ( 
.A(n_4842),
.B(n_4566),
.Y(n_5083)
);

A2O1A1Ixp33_ASAP7_75t_L g5084 ( 
.A1(n_4671),
.A2(n_4613),
.B(n_4976),
.C(n_5050),
.Y(n_5084)
);

AND2x4_ASAP7_75t_L g5085 ( 
.A(n_4844),
.B(n_4429),
.Y(n_5085)
);

BUFx3_ASAP7_75t_L g5086 ( 
.A(n_4607),
.Y(n_5086)
);

OA21x2_ASAP7_75t_L g5087 ( 
.A1(n_4900),
.A2(n_4544),
.B(n_4520),
.Y(n_5087)
);

OA21x2_ASAP7_75t_L g5088 ( 
.A1(n_4707),
.A2(n_4559),
.B(n_4497),
.Y(n_5088)
);

OAI21x1_ASAP7_75t_L g5089 ( 
.A1(n_5038),
.A2(n_4539),
.B(n_4518),
.Y(n_5089)
);

INVx2_ASAP7_75t_L g5090 ( 
.A(n_4623),
.Y(n_5090)
);

INVx1_ASAP7_75t_L g5091 ( 
.A(n_4668),
.Y(n_5091)
);

AND2x2_ASAP7_75t_L g5092 ( 
.A(n_4775),
.B(n_4781),
.Y(n_5092)
);

AO21x2_ASAP7_75t_L g5093 ( 
.A1(n_4853),
.A2(n_4324),
.B(n_4405),
.Y(n_5093)
);

INVx1_ASAP7_75t_SL g5094 ( 
.A(n_4714),
.Y(n_5094)
);

OAI21x1_ASAP7_75t_L g5095 ( 
.A1(n_4614),
.A2(n_4555),
.B(n_4545),
.Y(n_5095)
);

INVx2_ASAP7_75t_L g5096 ( 
.A(n_4630),
.Y(n_5096)
);

BUFx6f_ASAP7_75t_L g5097 ( 
.A(n_4787),
.Y(n_5097)
);

AOI22xp33_ASAP7_75t_L g5098 ( 
.A1(n_4595),
.A2(n_5044),
.B1(n_4650),
.B2(n_5003),
.Y(n_5098)
);

INVx2_ASAP7_75t_L g5099 ( 
.A(n_4676),
.Y(n_5099)
);

AOI21xp5_ASAP7_75t_L g5100 ( 
.A1(n_5036),
.A2(n_4475),
.B(n_4429),
.Y(n_5100)
);

OR2x2_ASAP7_75t_L g5101 ( 
.A(n_4649),
.B(n_4441),
.Y(n_5101)
);

AND2x2_ASAP7_75t_L g5102 ( 
.A(n_4776),
.B(n_4429),
.Y(n_5102)
);

A2O1A1Ixp33_ASAP7_75t_L g5103 ( 
.A1(n_4638),
.A2(n_4590),
.B(n_4059),
.C(n_4557),
.Y(n_5103)
);

AOI21xp5_ASAP7_75t_L g5104 ( 
.A1(n_4844),
.A2(n_4483),
.B(n_4475),
.Y(n_5104)
);

OR2x2_ASAP7_75t_L g5105 ( 
.A(n_4838),
.B(n_4443),
.Y(n_5105)
);

INVx2_ASAP7_75t_L g5106 ( 
.A(n_4688),
.Y(n_5106)
);

INVx1_ASAP7_75t_L g5107 ( 
.A(n_4678),
.Y(n_5107)
);

AOI21xp5_ASAP7_75t_L g5108 ( 
.A1(n_4844),
.A2(n_4483),
.B(n_4475),
.Y(n_5108)
);

INVx1_ASAP7_75t_L g5109 ( 
.A(n_4687),
.Y(n_5109)
);

OAI21x1_ASAP7_75t_L g5110 ( 
.A1(n_4604),
.A2(n_4288),
.B(n_4258),
.Y(n_5110)
);

OAI21x1_ASAP7_75t_L g5111 ( 
.A1(n_4823),
.A2(n_4308),
.B(n_4289),
.Y(n_5111)
);

OAI21x1_ASAP7_75t_L g5112 ( 
.A1(n_4637),
.A2(n_4325),
.B(n_4323),
.Y(n_5112)
);

INVx2_ASAP7_75t_L g5113 ( 
.A(n_4753),
.Y(n_5113)
);

OAI21x1_ASAP7_75t_L g5114 ( 
.A1(n_4624),
.A2(n_4334),
.B(n_4332),
.Y(n_5114)
);

OA21x2_ASAP7_75t_L g5115 ( 
.A1(n_4718),
.A2(n_4504),
.B(n_4487),
.Y(n_5115)
);

OAI21x1_ASAP7_75t_L g5116 ( 
.A1(n_4667),
.A2(n_4351),
.B(n_4339),
.Y(n_5116)
);

INVx1_ASAP7_75t_L g5117 ( 
.A(n_4691),
.Y(n_5117)
);

BUFx10_ASAP7_75t_L g5118 ( 
.A(n_4656),
.Y(n_5118)
);

INVx1_ASAP7_75t_L g5119 ( 
.A(n_4683),
.Y(n_5119)
);

AOI21xp33_ASAP7_75t_L g5120 ( 
.A1(n_4959),
.A2(n_4386),
.B(n_4383),
.Y(n_5120)
);

NAND3xp33_ASAP7_75t_L g5121 ( 
.A(n_4987),
.B(n_4806),
.C(n_4972),
.Y(n_5121)
);

INVx1_ASAP7_75t_L g5122 ( 
.A(n_4704),
.Y(n_5122)
);

INVx3_ASAP7_75t_L g5123 ( 
.A(n_4782),
.Y(n_5123)
);

OAI21x1_ASAP7_75t_L g5124 ( 
.A1(n_4768),
.A2(n_4565),
.B(n_4523),
.Y(n_5124)
);

OA21x2_ASAP7_75t_L g5125 ( 
.A1(n_4935),
.A2(n_4531),
.B(n_4512),
.Y(n_5125)
);

OAI21x1_ASAP7_75t_L g5126 ( 
.A1(n_5035),
.A2(n_4543),
.B(n_4538),
.Y(n_5126)
);

INVx1_ASAP7_75t_L g5127 ( 
.A(n_4725),
.Y(n_5127)
);

A2O1A1Ixp33_ASAP7_75t_L g5128 ( 
.A1(n_4948),
.A2(n_4562),
.B(n_4560),
.C(n_4202),
.Y(n_5128)
);

INVx2_ASAP7_75t_SL g5129 ( 
.A(n_4703),
.Y(n_5129)
);

INVx1_ASAP7_75t_L g5130 ( 
.A(n_4708),
.Y(n_5130)
);

OR2x2_ASAP7_75t_L g5131 ( 
.A(n_4805),
.B(n_4478),
.Y(n_5131)
);

O2A1O1Ixp33_ASAP7_75t_SL g5132 ( 
.A1(n_4654),
.A2(n_4216),
.B(n_4422),
.C(n_4452),
.Y(n_5132)
);

OAI21x1_ASAP7_75t_SL g5133 ( 
.A1(n_4872),
.A2(n_4570),
.B(n_4485),
.Y(n_5133)
);

INVx2_ASAP7_75t_L g5134 ( 
.A(n_4808),
.Y(n_5134)
);

OAI21x1_ASAP7_75t_L g5135 ( 
.A1(n_4634),
.A2(n_4580),
.B(n_4180),
.Y(n_5135)
);

OAI21x1_ASAP7_75t_L g5136 ( 
.A1(n_5060),
.A2(n_4167),
.B(n_4554),
.Y(n_5136)
);

AOI22xp5_ASAP7_75t_L g5137 ( 
.A1(n_4734),
.A2(n_4589),
.B1(n_4576),
.B2(n_4269),
.Y(n_5137)
);

OAI21x1_ASAP7_75t_L g5138 ( 
.A1(n_4625),
.A2(n_4867),
.B(n_4747),
.Y(n_5138)
);

NAND2xp5_ASAP7_75t_L g5139 ( 
.A(n_4829),
.B(n_4398),
.Y(n_5139)
);

A2O1A1Ixp33_ASAP7_75t_L g5140 ( 
.A1(n_4735),
.A2(n_4404),
.B(n_4481),
.C(n_4171),
.Y(n_5140)
);

OA21x2_ASAP7_75t_L g5141 ( 
.A1(n_4910),
.A2(n_4571),
.B(n_4483),
.Y(n_5141)
);

INVx6_ASAP7_75t_L g5142 ( 
.A(n_4960),
.Y(n_5142)
);

INVx2_ASAP7_75t_L g5143 ( 
.A(n_4820),
.Y(n_5143)
);

AO21x2_ASAP7_75t_L g5144 ( 
.A1(n_4856),
.A2(n_958),
.B(n_956),
.Y(n_5144)
);

OAI21x1_ASAP7_75t_L g5145 ( 
.A1(n_4878),
.A2(n_958),
.B(n_956),
.Y(n_5145)
);

INVx2_ASAP7_75t_L g5146 ( 
.A(n_4616),
.Y(n_5146)
);

OAI221xp5_ASAP7_75t_SL g5147 ( 
.A1(n_4729),
.A2(n_960),
.B1(n_961),
.B2(n_959),
.C(n_958),
.Y(n_5147)
);

OAI21x1_ASAP7_75t_L g5148 ( 
.A1(n_4666),
.A2(n_960),
.B(n_959),
.Y(n_5148)
);

NAND2xp5_ASAP7_75t_L g5149 ( 
.A(n_4830),
.B(n_1114),
.Y(n_5149)
);

AND2x4_ASAP7_75t_L g5150 ( 
.A(n_4911),
.B(n_960),
.Y(n_5150)
);

INVx2_ASAP7_75t_L g5151 ( 
.A(n_4710),
.Y(n_5151)
);

CKINVDCx20_ASAP7_75t_R g5152 ( 
.A(n_4596),
.Y(n_5152)
);

NAND2xp5_ASAP7_75t_L g5153 ( 
.A(n_4946),
.B(n_961),
.Y(n_5153)
);

OA21x2_ASAP7_75t_L g5154 ( 
.A1(n_4854),
.A2(n_962),
.B(n_961),
.Y(n_5154)
);

INVx2_ASAP7_75t_SL g5155 ( 
.A(n_4664),
.Y(n_5155)
);

INVx1_ASAP7_75t_L g5156 ( 
.A(n_4801),
.Y(n_5156)
);

NAND2xp5_ASAP7_75t_L g5157 ( 
.A(n_4949),
.B(n_1114),
.Y(n_5157)
);

INVx2_ASAP7_75t_L g5158 ( 
.A(n_4711),
.Y(n_5158)
);

NAND2xp5_ASAP7_75t_L g5159 ( 
.A(n_4958),
.B(n_962),
.Y(n_5159)
);

AO31x2_ASAP7_75t_L g5160 ( 
.A1(n_4983),
.A2(n_5021),
.A3(n_4794),
.B(n_5025),
.Y(n_5160)
);

AND2x2_ASAP7_75t_L g5161 ( 
.A(n_4632),
.B(n_4709),
.Y(n_5161)
);

A2O1A1Ixp33_ASAP7_75t_L g5162 ( 
.A1(n_4825),
.A2(n_964),
.B(n_965),
.C(n_963),
.Y(n_5162)
);

NAND2xp5_ASAP7_75t_L g5163 ( 
.A(n_4995),
.B(n_1113),
.Y(n_5163)
);

OAI21x1_ASAP7_75t_L g5164 ( 
.A1(n_4700),
.A2(n_4675),
.B(n_4673),
.Y(n_5164)
);

AO31x2_ASAP7_75t_L g5165 ( 
.A1(n_5032),
.A2(n_1113),
.A3(n_964),
.B(n_965),
.Y(n_5165)
);

NAND2xp5_ASAP7_75t_L g5166 ( 
.A(n_5000),
.B(n_1113),
.Y(n_5166)
);

INVx2_ASAP7_75t_L g5167 ( 
.A(n_4726),
.Y(n_5167)
);

OAI21x1_ASAP7_75t_L g5168 ( 
.A1(n_5029),
.A2(n_964),
.B(n_963),
.Y(n_5168)
);

NAND2xp5_ASAP7_75t_L g5169 ( 
.A(n_4951),
.B(n_965),
.Y(n_5169)
);

OAI22xp5_ASAP7_75t_L g5170 ( 
.A1(n_4686),
.A2(n_967),
.B1(n_968),
.B2(n_966),
.Y(n_5170)
);

AO21x2_ASAP7_75t_L g5171 ( 
.A1(n_4602),
.A2(n_967),
.B(n_966),
.Y(n_5171)
);

AOI22xp33_ASAP7_75t_L g5172 ( 
.A1(n_4715),
.A2(n_968),
.B1(n_969),
.B2(n_967),
.Y(n_5172)
);

INVx1_ASAP7_75t_L g5173 ( 
.A(n_4749),
.Y(n_5173)
);

NOR2xp33_ASAP7_75t_L g5174 ( 
.A(n_4732),
.B(n_71),
.Y(n_5174)
);

OA21x2_ASAP7_75t_L g5175 ( 
.A1(n_4660),
.A2(n_970),
.B(n_969),
.Y(n_5175)
);

OR2x2_ASAP7_75t_L g5176 ( 
.A(n_4742),
.B(n_1110),
.Y(n_5176)
);

INVx1_ASAP7_75t_L g5177 ( 
.A(n_4754),
.Y(n_5177)
);

NOR2x1_ASAP7_75t_L g5178 ( 
.A(n_4699),
.B(n_4655),
.Y(n_5178)
);

INVx2_ASAP7_75t_L g5179 ( 
.A(n_4757),
.Y(n_5179)
);

OAI21x1_ASAP7_75t_L g5180 ( 
.A1(n_4645),
.A2(n_970),
.B(n_969),
.Y(n_5180)
);

AND2x2_ASAP7_75t_L g5181 ( 
.A(n_4745),
.B(n_4760),
.Y(n_5181)
);

O2A1O1Ixp33_ASAP7_75t_L g5182 ( 
.A1(n_4819),
.A2(n_972),
.B(n_973),
.C(n_971),
.Y(n_5182)
);

INVx1_ASAP7_75t_L g5183 ( 
.A(n_4764),
.Y(n_5183)
);

OAI21x1_ASAP7_75t_SL g5184 ( 
.A1(n_4922),
.A2(n_972),
.B(n_971),
.Y(n_5184)
);

INVx1_ASAP7_75t_L g5185 ( 
.A(n_4765),
.Y(n_5185)
);

OAI22xp5_ASAP7_75t_L g5186 ( 
.A1(n_4789),
.A2(n_972),
.B1(n_973),
.B2(n_971),
.Y(n_5186)
);

BUFx2_ASAP7_75t_L g5187 ( 
.A(n_4722),
.Y(n_5187)
);

OAI21x1_ASAP7_75t_L g5188 ( 
.A1(n_4885),
.A2(n_975),
.B(n_974),
.Y(n_5188)
);

INVx2_ASAP7_75t_L g5189 ( 
.A(n_4771),
.Y(n_5189)
);

NAND2xp5_ASAP7_75t_L g5190 ( 
.A(n_4865),
.B(n_974),
.Y(n_5190)
);

BUFx8_ASAP7_75t_L g5191 ( 
.A(n_4601),
.Y(n_5191)
);

INVx1_ASAP7_75t_L g5192 ( 
.A(n_4772),
.Y(n_5192)
);

NOR2xp67_ASAP7_75t_L g5193 ( 
.A(n_4748),
.B(n_974),
.Y(n_5193)
);

INVx2_ASAP7_75t_L g5194 ( 
.A(n_4778),
.Y(n_5194)
);

INVx2_ASAP7_75t_L g5195 ( 
.A(n_4812),
.Y(n_5195)
);

NAND2xp5_ASAP7_75t_L g5196 ( 
.A(n_4852),
.B(n_1110),
.Y(n_5196)
);

OAI21x1_ASAP7_75t_L g5197 ( 
.A1(n_4952),
.A2(n_976),
.B(n_975),
.Y(n_5197)
);

BUFx4f_ASAP7_75t_L g5198 ( 
.A(n_4655),
.Y(n_5198)
);

AOI22xp33_ASAP7_75t_L g5199 ( 
.A1(n_4901),
.A2(n_976),
.B1(n_977),
.B2(n_975),
.Y(n_5199)
);

CKINVDCx11_ASAP7_75t_R g5200 ( 
.A(n_4605),
.Y(n_5200)
);

NOR2xp33_ASAP7_75t_L g5201 ( 
.A(n_4610),
.B(n_72),
.Y(n_5201)
);

NAND2x1p5_ASAP7_75t_L g5202 ( 
.A(n_4697),
.B(n_977),
.Y(n_5202)
);

NAND2xp5_ASAP7_75t_L g5203 ( 
.A(n_4824),
.B(n_978),
.Y(n_5203)
);

INVx2_ASAP7_75t_L g5204 ( 
.A(n_5011),
.Y(n_5204)
);

OAI21x1_ASAP7_75t_L g5205 ( 
.A1(n_4936),
.A2(n_979),
.B(n_978),
.Y(n_5205)
);

AOI221xp5_ASAP7_75t_L g5206 ( 
.A1(n_4743),
.A2(n_75),
.B1(n_73),
.B2(n_74),
.C(n_76),
.Y(n_5206)
);

AOI22xp33_ASAP7_75t_L g5207 ( 
.A1(n_4849),
.A2(n_979),
.B1(n_980),
.B2(n_978),
.Y(n_5207)
);

NAND2x1p5_ASAP7_75t_L g5208 ( 
.A(n_4601),
.B(n_979),
.Y(n_5208)
);

OR2x2_ASAP7_75t_L g5209 ( 
.A(n_4916),
.B(n_980),
.Y(n_5209)
);

OAI21x1_ASAP7_75t_L g5210 ( 
.A1(n_4866),
.A2(n_981),
.B(n_980),
.Y(n_5210)
);

AO31x2_ASAP7_75t_L g5211 ( 
.A1(n_5052),
.A2(n_1109),
.A3(n_982),
.B(n_983),
.Y(n_5211)
);

O2A1O1Ixp33_ASAP7_75t_SL g5212 ( 
.A1(n_4636),
.A2(n_983),
.B(n_984),
.C(n_981),
.Y(n_5212)
);

AOI22xp33_ASAP7_75t_L g5213 ( 
.A1(n_5059),
.A2(n_983),
.B1(n_984),
.B2(n_981),
.Y(n_5213)
);

BUFx3_ASAP7_75t_L g5214 ( 
.A(n_4766),
.Y(n_5214)
);

CKINVDCx20_ASAP7_75t_R g5215 ( 
.A(n_4670),
.Y(n_5215)
);

NAND2xp5_ASAP7_75t_L g5216 ( 
.A(n_5008),
.B(n_5045),
.Y(n_5216)
);

INVx2_ASAP7_75t_L g5217 ( 
.A(n_4598),
.Y(n_5217)
);

INVx4_ASAP7_75t_L g5218 ( 
.A(n_4699),
.Y(n_5218)
);

OAI21x1_ASAP7_75t_L g5219 ( 
.A1(n_4693),
.A2(n_985),
.B(n_984),
.Y(n_5219)
);

AND2x2_ASAP7_75t_L g5220 ( 
.A(n_4773),
.B(n_73),
.Y(n_5220)
);

INVx2_ASAP7_75t_SL g5221 ( 
.A(n_4759),
.Y(n_5221)
);

AND2x4_ASAP7_75t_L g5222 ( 
.A(n_4814),
.B(n_986),
.Y(n_5222)
);

INVx1_ASAP7_75t_L g5223 ( 
.A(n_4680),
.Y(n_5223)
);

OAI21x1_ASAP7_75t_L g5224 ( 
.A1(n_4672),
.A2(n_987),
.B(n_986),
.Y(n_5224)
);

AND2x2_ASAP7_75t_L g5225 ( 
.A(n_4752),
.B(n_73),
.Y(n_5225)
);

O2A1O1Ixp33_ASAP7_75t_SL g5226 ( 
.A1(n_4809),
.A2(n_4659),
.B(n_4840),
.C(n_4716),
.Y(n_5226)
);

AOI22xp33_ASAP7_75t_L g5227 ( 
.A1(n_5059),
.A2(n_987),
.B1(n_988),
.B2(n_986),
.Y(n_5227)
);

OAI21x1_ASAP7_75t_L g5228 ( 
.A1(n_4884),
.A2(n_4980),
.B(n_5001),
.Y(n_5228)
);

AOI22xp5_ASAP7_75t_L g5229 ( 
.A1(n_5010),
.A2(n_988),
.B1(n_989),
.B2(n_987),
.Y(n_5229)
);

CKINVDCx5p33_ASAP7_75t_R g5230 ( 
.A(n_4720),
.Y(n_5230)
);

INVx1_ASAP7_75t_L g5231 ( 
.A(n_4609),
.Y(n_5231)
);

NAND2xp5_ASAP7_75t_L g5232 ( 
.A(n_5058),
.B(n_5062),
.Y(n_5232)
);

INVx2_ASAP7_75t_L g5233 ( 
.A(n_4598),
.Y(n_5233)
);

INVx2_ASAP7_75t_L g5234 ( 
.A(n_5014),
.Y(n_5234)
);

AO21x2_ASAP7_75t_L g5235 ( 
.A1(n_4622),
.A2(n_989),
.B(n_988),
.Y(n_5235)
);

INVx2_ASAP7_75t_L g5236 ( 
.A(n_5049),
.Y(n_5236)
);

INVx2_ASAP7_75t_L g5237 ( 
.A(n_5066),
.Y(n_5237)
);

NAND2xp5_ASAP7_75t_L g5238 ( 
.A(n_4921),
.B(n_989),
.Y(n_5238)
);

OA21x2_ASAP7_75t_L g5239 ( 
.A1(n_4599),
.A2(n_991),
.B(n_990),
.Y(n_5239)
);

OAI21xp5_ASAP7_75t_L g5240 ( 
.A1(n_4817),
.A2(n_4798),
.B(n_4933),
.Y(n_5240)
);

AND2x2_ASAP7_75t_SL g5241 ( 
.A(n_4651),
.B(n_1109),
.Y(n_5241)
);

INVx2_ASAP7_75t_L g5242 ( 
.A(n_4974),
.Y(n_5242)
);

AOI21xp5_ASAP7_75t_L g5243 ( 
.A1(n_4600),
.A2(n_991),
.B(n_990),
.Y(n_5243)
);

OAI21x1_ASAP7_75t_L g5244 ( 
.A1(n_5042),
.A2(n_4895),
.B(n_4998),
.Y(n_5244)
);

BUFx3_ASAP7_75t_L g5245 ( 
.A(n_4940),
.Y(n_5245)
);

OAI21x1_ASAP7_75t_L g5246 ( 
.A1(n_5042),
.A2(n_991),
.B(n_990),
.Y(n_5246)
);

NAND2xp5_ASAP7_75t_L g5247 ( 
.A(n_5016),
.B(n_992),
.Y(n_5247)
);

INVx1_ASAP7_75t_L g5248 ( 
.A(n_4643),
.Y(n_5248)
);

CKINVDCx20_ASAP7_75t_R g5249 ( 
.A(n_4677),
.Y(n_5249)
);

NAND2xp5_ASAP7_75t_L g5250 ( 
.A(n_4786),
.B(n_992),
.Y(n_5250)
);

OAI21x1_ASAP7_75t_L g5251 ( 
.A1(n_4642),
.A2(n_994),
.B(n_993),
.Y(n_5251)
);

AOI21xp33_ASAP7_75t_L g5252 ( 
.A1(n_5020),
.A2(n_994),
.B(n_993),
.Y(n_5252)
);

OAI21x1_ASAP7_75t_L g5253 ( 
.A1(n_4712),
.A2(n_995),
.B(n_993),
.Y(n_5253)
);

OA21x2_ASAP7_75t_L g5254 ( 
.A1(n_4779),
.A2(n_996),
.B(n_995),
.Y(n_5254)
);

AND2x2_ASAP7_75t_L g5255 ( 
.A(n_4881),
.B(n_4925),
.Y(n_5255)
);

INVx2_ASAP7_75t_L g5256 ( 
.A(n_4974),
.Y(n_5256)
);

OAI21x1_ASAP7_75t_L g5257 ( 
.A1(n_4721),
.A2(n_997),
.B(n_996),
.Y(n_5257)
);

OAI222xp33_ASAP7_75t_L g5258 ( 
.A1(n_4597),
.A2(n_1000),
.B1(n_998),
.B2(n_1001),
.C1(n_999),
.C2(n_996),
.Y(n_5258)
);

AND2x4_ASAP7_75t_L g5259 ( 
.A(n_4780),
.B(n_998),
.Y(n_5259)
);

OA21x2_ASAP7_75t_L g5260 ( 
.A1(n_4591),
.A2(n_999),
.B(n_998),
.Y(n_5260)
);

AOI221xp5_ASAP7_75t_L g5261 ( 
.A1(n_4665),
.A2(n_4641),
.B1(n_4835),
.B2(n_4882),
.C(n_4913),
.Y(n_5261)
);

NAND2x1p5_ASAP7_75t_L g5262 ( 
.A(n_4941),
.B(n_1000),
.Y(n_5262)
);

NOR2xp33_ASAP7_75t_L g5263 ( 
.A(n_4957),
.B(n_74),
.Y(n_5263)
);

OAI21x1_ASAP7_75t_L g5264 ( 
.A1(n_4813),
.A2(n_1001),
.B(n_1000),
.Y(n_5264)
);

INVx2_ASAP7_75t_L g5265 ( 
.A(n_4974),
.Y(n_5265)
);

NOR2xp33_ASAP7_75t_L g5266 ( 
.A(n_4770),
.B(n_74),
.Y(n_5266)
);

AND2x2_ASAP7_75t_L g5267 ( 
.A(n_4934),
.B(n_75),
.Y(n_5267)
);

INVx2_ASAP7_75t_L g5268 ( 
.A(n_4974),
.Y(n_5268)
);

BUFx3_ASAP7_75t_L g5269 ( 
.A(n_4855),
.Y(n_5269)
);

O2A1O1Ixp33_ASAP7_75t_L g5270 ( 
.A1(n_5024),
.A2(n_1002),
.B(n_1003),
.C(n_1001),
.Y(n_5270)
);

O2A1O1Ixp33_ASAP7_75t_SL g5271 ( 
.A1(n_4919),
.A2(n_1004),
.B(n_1005),
.C(n_1002),
.Y(n_5271)
);

HB1xp67_ASAP7_75t_L g5272 ( 
.A(n_4994),
.Y(n_5272)
);

NAND3xp33_ASAP7_75t_L g5273 ( 
.A(n_4648),
.B(n_1006),
.C(n_1005),
.Y(n_5273)
);

AOI22x1_ASAP7_75t_L g5274 ( 
.A1(n_4684),
.A2(n_1006),
.B1(n_1007),
.B2(n_1005),
.Y(n_5274)
);

INVx2_ASAP7_75t_SL g5275 ( 
.A(n_4855),
.Y(n_5275)
);

INVx2_ASAP7_75t_L g5276 ( 
.A(n_4928),
.Y(n_5276)
);

CKINVDCx11_ASAP7_75t_R g5277 ( 
.A(n_4839),
.Y(n_5277)
);

INVx2_ASAP7_75t_L g5278 ( 
.A(n_4928),
.Y(n_5278)
);

OAI21x1_ASAP7_75t_L g5279 ( 
.A1(n_4818),
.A2(n_4834),
.B(n_4821),
.Y(n_5279)
);

NAND2x1p5_ASAP7_75t_L g5280 ( 
.A(n_4961),
.B(n_1006),
.Y(n_5280)
);

OAI21x1_ASAP7_75t_L g5281 ( 
.A1(n_4845),
.A2(n_1008),
.B(n_1007),
.Y(n_5281)
);

BUFx12f_ASAP7_75t_L g5282 ( 
.A(n_4874),
.Y(n_5282)
);

AO22x2_ASAP7_75t_L g5283 ( 
.A1(n_4942),
.A2(n_1008),
.B1(n_1009),
.B2(n_1007),
.Y(n_5283)
);

OAI21x1_ASAP7_75t_L g5284 ( 
.A1(n_4846),
.A2(n_1010),
.B(n_1008),
.Y(n_5284)
);

INVx1_ASAP7_75t_L g5285 ( 
.A(n_4982),
.Y(n_5285)
);

AOI22xp33_ASAP7_75t_L g5286 ( 
.A1(n_4997),
.A2(n_1012),
.B1(n_1013),
.B2(n_1010),
.Y(n_5286)
);

BUFx2_ASAP7_75t_L g5287 ( 
.A(n_4896),
.Y(n_5287)
);

BUFx4_ASAP7_75t_SL g5288 ( 
.A(n_4978),
.Y(n_5288)
);

AND2x4_ASAP7_75t_L g5289 ( 
.A(n_4859),
.B(n_1012),
.Y(n_5289)
);

AOI21xp5_ASAP7_75t_L g5290 ( 
.A1(n_4679),
.A2(n_1014),
.B(n_1013),
.Y(n_5290)
);

NAND2x1p5_ASAP7_75t_L g5291 ( 
.A(n_4615),
.B(n_4695),
.Y(n_5291)
);

OA21x2_ASAP7_75t_L g5292 ( 
.A1(n_4800),
.A2(n_1014),
.B(n_1013),
.Y(n_5292)
);

INVx3_ASAP7_75t_L g5293 ( 
.A(n_5015),
.Y(n_5293)
);

OAI21x1_ASAP7_75t_L g5294 ( 
.A1(n_4850),
.A2(n_1016),
.B(n_1015),
.Y(n_5294)
);

INVx4_ASAP7_75t_SL g5295 ( 
.A(n_4628),
.Y(n_5295)
);

INVx2_ASAP7_75t_L g5296 ( 
.A(n_4681),
.Y(n_5296)
);

OAI21x1_ASAP7_75t_L g5297 ( 
.A1(n_4593),
.A2(n_1016),
.B(n_1015),
.Y(n_5297)
);

AND2x2_ASAP7_75t_L g5298 ( 
.A(n_4939),
.B(n_75),
.Y(n_5298)
);

OA21x2_ASAP7_75t_L g5299 ( 
.A1(n_4698),
.A2(n_1016),
.B(n_1015),
.Y(n_5299)
);

AOI221xp5_ASAP7_75t_L g5300 ( 
.A1(n_4665),
.A2(n_78),
.B1(n_76),
.B2(n_77),
.C(n_79),
.Y(n_5300)
);

OR2x6_ASAP7_75t_L g5301 ( 
.A(n_4985),
.B(n_1017),
.Y(n_5301)
);

BUFx3_ASAP7_75t_L g5302 ( 
.A(n_4984),
.Y(n_5302)
);

OAI21xp5_ASAP7_75t_L g5303 ( 
.A1(n_4930),
.A2(n_1019),
.B(n_1018),
.Y(n_5303)
);

OAI21x1_ASAP7_75t_L g5304 ( 
.A1(n_4898),
.A2(n_1019),
.B(n_1018),
.Y(n_5304)
);

AO32x2_ASAP7_75t_L g5305 ( 
.A1(n_4828),
.A2(n_1021),
.A3(n_1022),
.B1(n_1020),
.B2(n_1018),
.Y(n_5305)
);

AND2x4_ASAP7_75t_L g5306 ( 
.A(n_4886),
.B(n_1020),
.Y(n_5306)
);

O2A1O1Ixp33_ASAP7_75t_L g5307 ( 
.A1(n_5026),
.A2(n_5040),
.B(n_5034),
.C(n_4944),
.Y(n_5307)
);

CKINVDCx5p33_ASAP7_75t_R g5308 ( 
.A(n_4847),
.Y(n_5308)
);

AOI21x1_ASAP7_75t_L g5309 ( 
.A1(n_4791),
.A2(n_4802),
.B(n_4797),
.Y(n_5309)
);

INVx1_ASAP7_75t_L g5310 ( 
.A(n_4989),
.Y(n_5310)
);

INVx1_ASAP7_75t_L g5311 ( 
.A(n_4681),
.Y(n_5311)
);

INVx2_ASAP7_75t_SL g5312 ( 
.A(n_4912),
.Y(n_5312)
);

AOI22x1_ASAP7_75t_L g5313 ( 
.A1(n_4621),
.A2(n_1021),
.B1(n_1023),
.B2(n_1020),
.Y(n_5313)
);

OAI21x1_ASAP7_75t_SL g5314 ( 
.A1(n_4612),
.A2(n_5019),
.B(n_4611),
.Y(n_5314)
);

NOR2xp33_ASAP7_75t_L g5315 ( 
.A(n_4857),
.B(n_76),
.Y(n_5315)
);

AO21x2_ASAP7_75t_L g5316 ( 
.A1(n_4868),
.A2(n_1024),
.B(n_1023),
.Y(n_5316)
);

INVx1_ASAP7_75t_L g5317 ( 
.A(n_4603),
.Y(n_5317)
);

O2A1O1Ixp33_ASAP7_75t_L g5318 ( 
.A1(n_4883),
.A2(n_1024),
.B(n_1025),
.C(n_1023),
.Y(n_5318)
);

OR2x2_ASAP7_75t_L g5319 ( 
.A(n_4706),
.B(n_4719),
.Y(n_5319)
);

NAND2x1p5_ASAP7_75t_L g5320 ( 
.A(n_4875),
.B(n_1024),
.Y(n_5320)
);

OAI21x1_ASAP7_75t_L g5321 ( 
.A1(n_4955),
.A2(n_1026),
.B(n_1025),
.Y(n_5321)
);

BUFx3_ASAP7_75t_L g5322 ( 
.A(n_4777),
.Y(n_5322)
);

OAI21x1_ASAP7_75t_L g5323 ( 
.A1(n_4899),
.A2(n_1026),
.B(n_1025),
.Y(n_5323)
);

OAI21x1_ASAP7_75t_L g5324 ( 
.A1(n_4907),
.A2(n_1028),
.B(n_1027),
.Y(n_5324)
);

OAI21x1_ASAP7_75t_L g5325 ( 
.A1(n_4915),
.A2(n_1028),
.B(n_1027),
.Y(n_5325)
);

AOI332xp33_ASAP7_75t_L g5326 ( 
.A1(n_4739),
.A2(n_1101),
.A3(n_1096),
.B1(n_1095),
.B2(n_1094),
.B3(n_1093),
.C1(n_1092),
.C2(n_1091),
.Y(n_5326)
);

AND2x2_ASAP7_75t_L g5327 ( 
.A(n_4887),
.B(n_77),
.Y(n_5327)
);

O2A1O1Ixp33_ASAP7_75t_SL g5328 ( 
.A1(n_4811),
.A2(n_1028),
.B(n_1029),
.C(n_1027),
.Y(n_5328)
);

AND2x2_ASAP7_75t_L g5329 ( 
.A(n_4890),
.B(n_77),
.Y(n_5329)
);

OAI21x1_ASAP7_75t_L g5330 ( 
.A1(n_4741),
.A2(n_1030),
.B(n_1029),
.Y(n_5330)
);

O2A1O1Ixp33_ASAP7_75t_L g5331 ( 
.A1(n_4888),
.A2(n_1030),
.B(n_1032),
.C(n_1029),
.Y(n_5331)
);

NOR2xp33_ASAP7_75t_L g5332 ( 
.A(n_4894),
.B(n_77),
.Y(n_5332)
);

OAI221xp5_ASAP7_75t_L g5333 ( 
.A1(n_4619),
.A2(n_1034),
.B1(n_1035),
.B2(n_1033),
.C(n_1030),
.Y(n_5333)
);

CKINVDCx5p33_ASAP7_75t_R g5334 ( 
.A(n_4657),
.Y(n_5334)
);

INVx1_ASAP7_75t_L g5335 ( 
.A(n_4897),
.Y(n_5335)
);

AOI221xp5_ASAP7_75t_SL g5336 ( 
.A1(n_4826),
.A2(n_80),
.B1(n_78),
.B2(n_79),
.C(n_81),
.Y(n_5336)
);

NAND3xp33_ASAP7_75t_L g5337 ( 
.A(n_4831),
.B(n_1034),
.C(n_1033),
.Y(n_5337)
);

BUFx6f_ASAP7_75t_L g5338 ( 
.A(n_5033),
.Y(n_5338)
);

INVx1_ASAP7_75t_L g5339 ( 
.A(n_4627),
.Y(n_5339)
);

OAI21x1_ASAP7_75t_L g5340 ( 
.A1(n_5006),
.A2(n_1036),
.B(n_1034),
.Y(n_5340)
);

OAI21x1_ASAP7_75t_L g5341 ( 
.A1(n_5007),
.A2(n_1038),
.B(n_1037),
.Y(n_5341)
);

HB1xp67_ASAP7_75t_L g5342 ( 
.A(n_4927),
.Y(n_5342)
);

OAI21x1_ASAP7_75t_L g5343 ( 
.A1(n_5009),
.A2(n_1038),
.B(n_1037),
.Y(n_5343)
);

OR2x2_ASAP7_75t_L g5344 ( 
.A(n_4836),
.B(n_1038),
.Y(n_5344)
);

INVx8_ASAP7_75t_L g5345 ( 
.A(n_4628),
.Y(n_5345)
);

OAI21x1_ASAP7_75t_L g5346 ( 
.A1(n_5031),
.A2(n_1040),
.B(n_1039),
.Y(n_5346)
);

INVx1_ASAP7_75t_L g5347 ( 
.A(n_4627),
.Y(n_5347)
);

OR2x6_ASAP7_75t_L g5348 ( 
.A(n_4945),
.B(n_1039),
.Y(n_5348)
);

NAND2xp5_ASAP7_75t_SL g5349 ( 
.A(n_4902),
.B(n_1039),
.Y(n_5349)
);

BUFx3_ASAP7_75t_L g5350 ( 
.A(n_4892),
.Y(n_5350)
);

INVx1_ASAP7_75t_L g5351 ( 
.A(n_4618),
.Y(n_5351)
);

OAI21x1_ASAP7_75t_L g5352 ( 
.A1(n_5037),
.A2(n_1041),
.B(n_1040),
.Y(n_5352)
);

INVx1_ASAP7_75t_SL g5353 ( 
.A(n_4937),
.Y(n_5353)
);

NOR2x1_ASAP7_75t_L g5354 ( 
.A(n_4713),
.B(n_1040),
.Y(n_5354)
);

INVx1_ASAP7_75t_L g5355 ( 
.A(n_4620),
.Y(n_5355)
);

AOI21xp5_ASAP7_75t_L g5356 ( 
.A1(n_4669),
.A2(n_1042),
.B(n_1041),
.Y(n_5356)
);

NOR2xp33_ASAP7_75t_L g5357 ( 
.A(n_4891),
.B(n_78),
.Y(n_5357)
);

INVx1_ASAP7_75t_L g5358 ( 
.A(n_4663),
.Y(n_5358)
);

NAND2x1p5_ASAP7_75t_L g5359 ( 
.A(n_5004),
.B(n_1041),
.Y(n_5359)
);

INVx2_ASAP7_75t_L g5360 ( 
.A(n_4864),
.Y(n_5360)
);

OAI21x1_ASAP7_75t_L g5361 ( 
.A1(n_5054),
.A2(n_1043),
.B(n_1042),
.Y(n_5361)
);

OAI22xp5_ASAP7_75t_SL g5362 ( 
.A1(n_4804),
.A2(n_1043),
.B1(n_1044),
.B2(n_1042),
.Y(n_5362)
);

OAI21x1_ASAP7_75t_L g5363 ( 
.A1(n_5055),
.A2(n_1045),
.B(n_1044),
.Y(n_5363)
);

NOR2xp67_ASAP7_75t_L g5364 ( 
.A(n_4788),
.B(n_1044),
.Y(n_5364)
);

OAI21x1_ASAP7_75t_L g5365 ( 
.A1(n_4689),
.A2(n_1046),
.B(n_1045),
.Y(n_5365)
);

OAI21x1_ASAP7_75t_L g5366 ( 
.A1(n_4738),
.A2(n_4696),
.B(n_5057),
.Y(n_5366)
);

INVx1_ASAP7_75t_L g5367 ( 
.A(n_4674),
.Y(n_5367)
);

OAI21x1_ASAP7_75t_L g5368 ( 
.A1(n_4646),
.A2(n_1046),
.B(n_1045),
.Y(n_5368)
);

NOR2xp33_ASAP7_75t_L g5369 ( 
.A(n_4774),
.B(n_78),
.Y(n_5369)
);

CKINVDCx20_ASAP7_75t_R g5370 ( 
.A(n_4848),
.Y(n_5370)
);

OAI21x1_ASAP7_75t_L g5371 ( 
.A1(n_4791),
.A2(n_1047),
.B(n_1046),
.Y(n_5371)
);

NAND2xp5_ASAP7_75t_SL g5372 ( 
.A(n_5004),
.B(n_1047),
.Y(n_5372)
);

INVx3_ASAP7_75t_L g5373 ( 
.A(n_4628),
.Y(n_5373)
);

INVx1_ASAP7_75t_L g5374 ( 
.A(n_4685),
.Y(n_5374)
);

OA21x2_ASAP7_75t_L g5375 ( 
.A1(n_4905),
.A2(n_1048),
.B(n_1047),
.Y(n_5375)
);

AND2x4_ASAP7_75t_L g5376 ( 
.A(n_4869),
.B(n_1048),
.Y(n_5376)
);

OAI21x1_ASAP7_75t_L g5377 ( 
.A1(n_4860),
.A2(n_1050),
.B(n_1049),
.Y(n_5377)
);

OAI21xp5_ASAP7_75t_L g5378 ( 
.A1(n_4904),
.A2(n_1050),
.B(n_1049),
.Y(n_5378)
);

OAI21x1_ASAP7_75t_L g5379 ( 
.A1(n_4694),
.A2(n_1051),
.B(n_1050),
.Y(n_5379)
);

INVx1_ASAP7_75t_L g5380 ( 
.A(n_4690),
.Y(n_5380)
);

AOI22xp5_ASAP7_75t_L g5381 ( 
.A1(n_4833),
.A2(n_1052),
.B1(n_1053),
.B2(n_1051),
.Y(n_5381)
);

BUFx8_ASAP7_75t_SL g5382 ( 
.A(n_4924),
.Y(n_5382)
);

AOI22xp33_ASAP7_75t_L g5383 ( 
.A1(n_5362),
.A2(n_5121),
.B1(n_5261),
.B2(n_4997),
.Y(n_5383)
);

NAND2xp5_ASAP7_75t_L g5384 ( 
.A(n_5119),
.B(n_4795),
.Y(n_5384)
);

AOI21x1_ASAP7_75t_L g5385 ( 
.A1(n_5178),
.A2(n_4969),
.B(n_4880),
.Y(n_5385)
);

AOI22xp33_ASAP7_75t_L g5386 ( 
.A1(n_5080),
.A2(n_4997),
.B1(n_5027),
.B2(n_5023),
.Y(n_5386)
);

NOR2xp33_ASAP7_75t_L g5387 ( 
.A(n_5078),
.B(n_4971),
.Y(n_5387)
);

INVx3_ASAP7_75t_L g5388 ( 
.A(n_5070),
.Y(n_5388)
);

NAND2xp5_ASAP7_75t_L g5389 ( 
.A(n_5231),
.B(n_4906),
.Y(n_5389)
);

AOI21xp5_ASAP7_75t_L g5390 ( 
.A1(n_5084),
.A2(n_5132),
.B(n_5077),
.Y(n_5390)
);

OR2x6_ASAP7_75t_L g5391 ( 
.A(n_5345),
.B(n_4790),
.Y(n_5391)
);

AOI21x1_ASAP7_75t_L g5392 ( 
.A1(n_5193),
.A2(n_4903),
.B(n_4755),
.Y(n_5392)
);

AND2x2_ASAP7_75t_L g5393 ( 
.A(n_5272),
.B(n_4876),
.Y(n_5393)
);

OA21x2_ASAP7_75t_L g5394 ( 
.A1(n_5276),
.A2(n_4929),
.B(n_4717),
.Y(n_5394)
);

NAND2x1p5_ASAP7_75t_L g5395 ( 
.A(n_5198),
.B(n_5004),
.Y(n_5395)
);

CKINVDCx5p33_ASAP7_75t_R g5396 ( 
.A(n_5200),
.Y(n_5396)
);

INVx2_ASAP7_75t_L g5397 ( 
.A(n_5187),
.Y(n_5397)
);

AND2x2_ASAP7_75t_L g5398 ( 
.A(n_5092),
.B(n_5018),
.Y(n_5398)
);

OAI21x1_ASAP7_75t_L g5399 ( 
.A1(n_5141),
.A2(n_5138),
.B(n_5278),
.Y(n_5399)
);

AO31x2_ASAP7_75t_L g5400 ( 
.A1(n_5287),
.A2(n_4973),
.A3(n_4877),
.B(n_5043),
.Y(n_5400)
);

AOI21xp5_ASAP7_75t_L g5401 ( 
.A1(n_5100),
.A2(n_4871),
.B(n_4785),
.Y(n_5401)
);

INVx2_ASAP7_75t_L g5402 ( 
.A(n_5187),
.Y(n_5402)
);

AOI21xp5_ASAP7_75t_L g5403 ( 
.A1(n_5345),
.A2(n_4993),
.B(n_4822),
.Y(n_5403)
);

AO21x2_ASAP7_75t_L g5404 ( 
.A1(n_5311),
.A2(n_4799),
.B(n_4653),
.Y(n_5404)
);

NOR2xp33_ASAP7_75t_L g5405 ( 
.A(n_5094),
.B(n_4975),
.Y(n_5405)
);

BUFx6f_ASAP7_75t_L g5406 ( 
.A(n_5338),
.Y(n_5406)
);

AOI21xp5_ASAP7_75t_L g5407 ( 
.A1(n_5104),
.A2(n_4992),
.B(n_4954),
.Y(n_5407)
);

INVx1_ASAP7_75t_L g5408 ( 
.A(n_5067),
.Y(n_5408)
);

BUFx12f_ASAP7_75t_L g5409 ( 
.A(n_5070),
.Y(n_5409)
);

OAI22xp5_ASAP7_75t_L g5410 ( 
.A1(n_5098),
.A2(n_4758),
.B1(n_4740),
.B2(n_5053),
.Y(n_5410)
);

A2O1A1Ixp33_ASAP7_75t_L g5411 ( 
.A1(n_5252),
.A2(n_5240),
.B(n_5373),
.C(n_5364),
.Y(n_5411)
);

AOI31xp33_ASAP7_75t_SL g5412 ( 
.A1(n_5300),
.A2(n_4943),
.A3(n_4815),
.B(n_4986),
.Y(n_5412)
);

INVx1_ASAP7_75t_SL g5413 ( 
.A(n_5288),
.Y(n_5413)
);

AO31x2_ASAP7_75t_L g5414 ( 
.A1(n_5287),
.A2(n_5051),
.A3(n_4692),
.B(n_4926),
.Y(n_5414)
);

AND2x2_ASAP7_75t_L g5415 ( 
.A(n_5161),
.B(n_4631),
.Y(n_5415)
);

AOI21xp5_ASAP7_75t_L g5416 ( 
.A1(n_5108),
.A2(n_4918),
.B(n_4841),
.Y(n_5416)
);

INVx2_ASAP7_75t_L g5417 ( 
.A(n_5090),
.Y(n_5417)
);

OAI21xp5_ASAP7_75t_L g5418 ( 
.A1(n_5170),
.A2(n_4793),
.B(n_4909),
.Y(n_5418)
);

OA21x2_ASAP7_75t_L g5419 ( 
.A1(n_5296),
.A2(n_4723),
.B(n_4705),
.Y(n_5419)
);

OAI21x1_ASAP7_75t_L g5420 ( 
.A1(n_5141),
.A2(n_4733),
.B(n_4762),
.Y(n_5420)
);

NAND2xp5_ASAP7_75t_L g5421 ( 
.A(n_5248),
.B(n_4858),
.Y(n_5421)
);

BUFx2_ASAP7_75t_L g5422 ( 
.A(n_5214),
.Y(n_5422)
);

NAND2xp5_ASAP7_75t_L g5423 ( 
.A(n_5127),
.B(n_4858),
.Y(n_5423)
);

OAI21x1_ASAP7_75t_SL g5424 ( 
.A1(n_5218),
.A2(n_4784),
.B(n_4658),
.Y(n_5424)
);

INVx1_ASAP7_75t_L g5425 ( 
.A(n_5074),
.Y(n_5425)
);

INVx1_ASAP7_75t_L g5426 ( 
.A(n_5076),
.Y(n_5426)
);

NAND2x1_ASAP7_75t_L g5427 ( 
.A(n_5301),
.B(n_4744),
.Y(n_5427)
);

AND2x4_ASAP7_75t_L g5428 ( 
.A(n_5295),
.B(n_4896),
.Y(n_5428)
);

OA21x2_ASAP7_75t_L g5429 ( 
.A1(n_5339),
.A2(n_4731),
.B(n_4724),
.Y(n_5429)
);

OAI22xp33_ASAP7_75t_L g5430 ( 
.A1(n_5301),
.A2(n_4629),
.B1(n_4728),
.B2(n_5022),
.Y(n_5430)
);

AND2x4_ASAP7_75t_L g5431 ( 
.A(n_5295),
.B(n_4962),
.Y(n_5431)
);

OAI21x1_ASAP7_75t_L g5432 ( 
.A1(n_5126),
.A2(n_4744),
.B(n_5012),
.Y(n_5432)
);

AO21x2_ASAP7_75t_L g5433 ( 
.A1(n_5347),
.A2(n_4746),
.B(n_4737),
.Y(n_5433)
);

OR2x6_ASAP7_75t_L g5434 ( 
.A(n_5142),
.B(n_4968),
.Y(n_5434)
);

INVx1_ASAP7_75t_L g5435 ( 
.A(n_5091),
.Y(n_5435)
);

AOI21xp5_ASAP7_75t_L g5436 ( 
.A1(n_5133),
.A2(n_5063),
.B(n_4767),
.Y(n_5436)
);

NAND2xp5_ASAP7_75t_L g5437 ( 
.A(n_5156),
.B(n_4756),
.Y(n_5437)
);

INVx2_ASAP7_75t_L g5438 ( 
.A(n_5096),
.Y(n_5438)
);

AND2x2_ASAP7_75t_L g5439 ( 
.A(n_5181),
.B(n_4631),
.Y(n_5439)
);

INVx2_ASAP7_75t_L g5440 ( 
.A(n_5099),
.Y(n_5440)
);

HB1xp67_ASAP7_75t_L g5441 ( 
.A(n_5302),
.Y(n_5441)
);

NOR2xp33_ASAP7_75t_L g5442 ( 
.A(n_5155),
.B(n_4999),
.Y(n_5442)
);

AOI21xp5_ASAP7_75t_L g5443 ( 
.A1(n_5133),
.A2(n_4751),
.B(n_4682),
.Y(n_5443)
);

AOI21xp5_ASAP7_75t_L g5444 ( 
.A1(n_5103),
.A2(n_5260),
.B(n_5072),
.Y(n_5444)
);

NAND2xp5_ASAP7_75t_L g5445 ( 
.A(n_5223),
.B(n_4756),
.Y(n_5445)
);

OAI21x1_ASAP7_75t_SL g5446 ( 
.A1(n_5184),
.A2(n_5314),
.B(n_5071),
.Y(n_5446)
);

INVx3_ASAP7_75t_L g5447 ( 
.A(n_5086),
.Y(n_5447)
);

NAND2xp5_ASAP7_75t_L g5448 ( 
.A(n_5317),
.B(n_4827),
.Y(n_5448)
);

BUFx2_ASAP7_75t_R g5449 ( 
.A(n_5308),
.Y(n_5449)
);

OA21x2_ASAP7_75t_L g5450 ( 
.A1(n_5217),
.A2(n_4783),
.B(n_4769),
.Y(n_5450)
);

OAI21x1_ASAP7_75t_SL g5451 ( 
.A1(n_5184),
.A2(n_4807),
.B(n_4702),
.Y(n_5451)
);

NAND2xp5_ASAP7_75t_L g5452 ( 
.A(n_5351),
.B(n_4827),
.Y(n_5452)
);

BUFx8_ASAP7_75t_L g5453 ( 
.A(n_5282),
.Y(n_5453)
);

AOI21xp5_ASAP7_75t_L g5454 ( 
.A1(n_5260),
.A2(n_5022),
.B(n_4763),
.Y(n_5454)
);

AOI21xp5_ASAP7_75t_L g5455 ( 
.A1(n_5271),
.A2(n_4796),
.B(n_4662),
.Y(n_5455)
);

AOI21xp5_ASAP7_75t_L g5456 ( 
.A1(n_5212),
.A2(n_4736),
.B(n_4956),
.Y(n_5456)
);

AND2x2_ASAP7_75t_L g5457 ( 
.A(n_5255),
.B(n_5102),
.Y(n_5457)
);

NAND2xp5_ASAP7_75t_L g5458 ( 
.A(n_5355),
.B(n_4640),
.Y(n_5458)
);

AND2x2_ASAP7_75t_L g5459 ( 
.A(n_5234),
.B(n_4640),
.Y(n_5459)
);

AOI21xp5_ASAP7_75t_L g5460 ( 
.A1(n_5128),
.A2(n_4956),
.B(n_4633),
.Y(n_5460)
);

HB1xp67_ASAP7_75t_L g5461 ( 
.A(n_5236),
.Y(n_5461)
);

OA21x2_ASAP7_75t_L g5462 ( 
.A1(n_5233),
.A2(n_4652),
.B(n_4920),
.Y(n_5462)
);

NAND2xp5_ASAP7_75t_L g5463 ( 
.A(n_5358),
.B(n_5380),
.Y(n_5463)
);

AND2x4_ASAP7_75t_L g5464 ( 
.A(n_5068),
.B(n_4962),
.Y(n_5464)
);

AOI22x1_ASAP7_75t_L g5465 ( 
.A1(n_5202),
.A2(n_4964),
.B1(n_4979),
.B2(n_4970),
.Y(n_5465)
);

NAND2xp5_ASAP7_75t_L g5466 ( 
.A(n_5367),
.B(n_4837),
.Y(n_5466)
);

INVxp67_ASAP7_75t_L g5467 ( 
.A(n_5245),
.Y(n_5467)
);

AO21x2_ASAP7_75t_L g5468 ( 
.A1(n_5120),
.A2(n_4953),
.B(n_4950),
.Y(n_5468)
);

BUFx6f_ASAP7_75t_L g5469 ( 
.A(n_5338),
.Y(n_5469)
);

AND2x4_ASAP7_75t_L g5470 ( 
.A(n_5068),
.B(n_4981),
.Y(n_5470)
);

INVx1_ASAP7_75t_L g5471 ( 
.A(n_5107),
.Y(n_5471)
);

AO31x2_ASAP7_75t_L g5472 ( 
.A1(n_5242),
.A2(n_4991),
.A3(n_4843),
.B(n_4966),
.Y(n_5472)
);

OAI21x1_ASAP7_75t_L g5473 ( 
.A1(n_5279),
.A2(n_4932),
.B(n_4923),
.Y(n_5473)
);

OAI21x1_ASAP7_75t_L g5474 ( 
.A1(n_5069),
.A2(n_4803),
.B(n_4761),
.Y(n_5474)
);

INVx2_ASAP7_75t_L g5475 ( 
.A(n_5106),
.Y(n_5475)
);

INVx1_ASAP7_75t_L g5476 ( 
.A(n_5109),
.Y(n_5476)
);

BUFx2_ASAP7_75t_L g5477 ( 
.A(n_5269),
.Y(n_5477)
);

OAI21x1_ASAP7_75t_L g5478 ( 
.A1(n_5164),
.A2(n_4803),
.B(n_4990),
.Y(n_5478)
);

AOI21xp5_ASAP7_75t_L g5479 ( 
.A1(n_5075),
.A2(n_4792),
.B(n_4879),
.Y(n_5479)
);

NOR2x1_ASAP7_75t_L g5480 ( 
.A(n_5322),
.B(n_4861),
.Y(n_5480)
);

INVx3_ASAP7_75t_L g5481 ( 
.A(n_5142),
.Y(n_5481)
);

INVx1_ASAP7_75t_L g5482 ( 
.A(n_5117),
.Y(n_5482)
);

OAI21x1_ASAP7_75t_L g5483 ( 
.A1(n_5228),
.A2(n_5017),
.B(n_4701),
.Y(n_5483)
);

INVx1_ASAP7_75t_L g5484 ( 
.A(n_5122),
.Y(n_5484)
);

INVx1_ASAP7_75t_L g5485 ( 
.A(n_5285),
.Y(n_5485)
);

AOI21xp5_ASAP7_75t_L g5486 ( 
.A1(n_5093),
.A2(n_4908),
.B(n_4870),
.Y(n_5486)
);

INVx2_ASAP7_75t_L g5487 ( 
.A(n_5113),
.Y(n_5487)
);

OA21x2_ASAP7_75t_L g5488 ( 
.A1(n_5256),
.A2(n_5061),
.B(n_5056),
.Y(n_5488)
);

OAI21xp5_ASAP7_75t_L g5489 ( 
.A1(n_5274),
.A2(n_5047),
.B(n_4963),
.Y(n_5489)
);

AND2x4_ASAP7_75t_L g5490 ( 
.A(n_5123),
.B(n_5221),
.Y(n_5490)
);

NAND2xp5_ASAP7_75t_L g5491 ( 
.A(n_5374),
.B(n_5046),
.Y(n_5491)
);

OR2x4_ASAP7_75t_L g5492 ( 
.A(n_5174),
.B(n_5028),
.Y(n_5492)
);

INVx2_ASAP7_75t_L g5493 ( 
.A(n_5134),
.Y(n_5493)
);

OAI22xp5_ASAP7_75t_L g5494 ( 
.A1(n_5137),
.A2(n_4889),
.B1(n_4863),
.B2(n_4862),
.Y(n_5494)
);

AND2x2_ASAP7_75t_L g5495 ( 
.A(n_5310),
.B(n_4914),
.Y(n_5495)
);

A2O1A1Ixp33_ASAP7_75t_L g5496 ( 
.A1(n_5326),
.A2(n_5005),
.B(n_5013),
.C(n_5002),
.Y(n_5496)
);

INVx4_ASAP7_75t_SL g5497 ( 
.A(n_5222),
.Y(n_5497)
);

INVx1_ASAP7_75t_L g5498 ( 
.A(n_5130),
.Y(n_5498)
);

NAND2xp5_ASAP7_75t_L g5499 ( 
.A(n_5151),
.B(n_4816),
.Y(n_5499)
);

NAND2xp5_ASAP7_75t_L g5500 ( 
.A(n_5158),
.B(n_5167),
.Y(n_5500)
);

OAI21x1_ASAP7_75t_L g5501 ( 
.A1(n_5371),
.A2(n_5039),
.B(n_5030),
.Y(n_5501)
);

HB1xp67_ASAP7_75t_L g5502 ( 
.A(n_5179),
.Y(n_5502)
);

AOI21xp5_ASAP7_75t_L g5503 ( 
.A1(n_5162),
.A2(n_4832),
.B(n_4967),
.Y(n_5503)
);

NAND2xp5_ASAP7_75t_L g5504 ( 
.A(n_5189),
.B(n_4931),
.Y(n_5504)
);

AOI21x1_ASAP7_75t_L g5505 ( 
.A1(n_5283),
.A2(n_5259),
.B(n_5354),
.Y(n_5505)
);

AND2x4_ASAP7_75t_L g5506 ( 
.A(n_5312),
.B(n_4727),
.Y(n_5506)
);

NOR2xp33_ASAP7_75t_L g5507 ( 
.A(n_5382),
.B(n_1052),
.Y(n_5507)
);

AO21x2_ASAP7_75t_L g5508 ( 
.A1(n_5314),
.A2(n_5064),
.B(n_5048),
.Y(n_5508)
);

AND2x2_ASAP7_75t_L g5509 ( 
.A(n_5204),
.B(n_4914),
.Y(n_5509)
);

INVx2_ASAP7_75t_L g5510 ( 
.A(n_5143),
.Y(n_5510)
);

AOI21xp5_ASAP7_75t_L g5511 ( 
.A1(n_5140),
.A2(n_4938),
.B(n_4917),
.Y(n_5511)
);

AND2x2_ASAP7_75t_L g5512 ( 
.A(n_5335),
.B(n_4931),
.Y(n_5512)
);

NAND2xp5_ASAP7_75t_L g5513 ( 
.A(n_5194),
.B(n_4947),
.Y(n_5513)
);

OAI21x1_ASAP7_75t_L g5514 ( 
.A1(n_5244),
.A2(n_5065),
.B(n_4873),
.Y(n_5514)
);

NAND2xp5_ASAP7_75t_L g5515 ( 
.A(n_5195),
.B(n_4947),
.Y(n_5515)
);

INVx1_ASAP7_75t_L g5516 ( 
.A(n_5173),
.Y(n_5516)
);

INVx1_ASAP7_75t_L g5517 ( 
.A(n_5177),
.Y(n_5517)
);

NAND2x1p5_ASAP7_75t_L g5518 ( 
.A(n_5150),
.B(n_4810),
.Y(n_5518)
);

OR2x2_ASAP7_75t_L g5519 ( 
.A(n_5319),
.B(n_4965),
.Y(n_5519)
);

AOI21xp5_ASAP7_75t_L g5520 ( 
.A1(n_5254),
.A2(n_4996),
.B(n_4661),
.Y(n_5520)
);

AO21x2_ASAP7_75t_L g5521 ( 
.A1(n_5203),
.A2(n_4661),
.B(n_4965),
.Y(n_5521)
);

AOI21xp5_ASAP7_75t_L g5522 ( 
.A1(n_5254),
.A2(n_4996),
.B(n_4810),
.Y(n_5522)
);

AO21x2_ASAP7_75t_L g5523 ( 
.A1(n_5303),
.A2(n_4873),
.B(n_4730),
.Y(n_5523)
);

OAI21x1_ASAP7_75t_L g5524 ( 
.A1(n_5124),
.A2(n_4727),
.B(n_4730),
.Y(n_5524)
);

OAI21x1_ASAP7_75t_L g5525 ( 
.A1(n_5366),
.A2(n_4592),
.B(n_4977),
.Y(n_5525)
);

A2O1A1Ixp33_ASAP7_75t_L g5526 ( 
.A1(n_5270),
.A2(n_4977),
.B(n_5041),
.C(n_1053),
.Y(n_5526)
);

INVx3_ASAP7_75t_L g5527 ( 
.A(n_5277),
.Y(n_5527)
);

AOI21xp5_ASAP7_75t_SL g5528 ( 
.A1(n_5222),
.A2(n_5041),
.B(n_1054),
.Y(n_5528)
);

OR2x2_ASAP7_75t_L g5529 ( 
.A(n_5101),
.B(n_4592),
.Y(n_5529)
);

INVx6_ASAP7_75t_L g5530 ( 
.A(n_5191),
.Y(n_5530)
);

OAI21xp33_ASAP7_75t_L g5531 ( 
.A1(n_5241),
.A2(n_79),
.B(n_80),
.Y(n_5531)
);

AO21x2_ASAP7_75t_L g5532 ( 
.A1(n_5153),
.A2(n_1055),
.B(n_1052),
.Y(n_5532)
);

AND2x2_ASAP7_75t_L g5533 ( 
.A(n_5360),
.B(n_5342),
.Y(n_5533)
);

AO21x2_ASAP7_75t_L g5534 ( 
.A1(n_5157),
.A2(n_1056),
.B(n_1055),
.Y(n_5534)
);

A2O1A1Ixp33_ASAP7_75t_L g5535 ( 
.A1(n_5318),
.A2(n_1056),
.B(n_1057),
.C(n_1055),
.Y(n_5535)
);

NAND2xp5_ASAP7_75t_L g5536 ( 
.A(n_5183),
.B(n_1056),
.Y(n_5536)
);

INVx4_ASAP7_75t_SL g5537 ( 
.A(n_5081),
.Y(n_5537)
);

BUFx2_ASAP7_75t_L g5538 ( 
.A(n_5081),
.Y(n_5538)
);

INVx2_ASAP7_75t_L g5539 ( 
.A(n_5146),
.Y(n_5539)
);

AOI21xp5_ASAP7_75t_L g5540 ( 
.A1(n_5328),
.A2(n_1058),
.B(n_1057),
.Y(n_5540)
);

INVx1_ASAP7_75t_L g5541 ( 
.A(n_5185),
.Y(n_5541)
);

INVx2_ASAP7_75t_L g5542 ( 
.A(n_5237),
.Y(n_5542)
);

AO31x2_ASAP7_75t_L g5543 ( 
.A1(n_5265),
.A2(n_5268),
.A3(n_5083),
.B(n_5192),
.Y(n_5543)
);

NOR2xp33_ASAP7_75t_L g5544 ( 
.A(n_5353),
.B(n_1057),
.Y(n_5544)
);

OAI22xp33_ASAP7_75t_SL g5545 ( 
.A1(n_5291),
.A2(n_5320),
.B1(n_5259),
.B2(n_5209),
.Y(n_5545)
);

OAI21x1_ASAP7_75t_L g5546 ( 
.A1(n_5309),
.A2(n_1059),
.B(n_1058),
.Y(n_5546)
);

AOI21xp5_ASAP7_75t_L g5547 ( 
.A1(n_5226),
.A2(n_1059),
.B(n_1058),
.Y(n_5547)
);

A2O1A1Ixp33_ASAP7_75t_L g5548 ( 
.A1(n_5331),
.A2(n_1060),
.B(n_1061),
.C(n_1059),
.Y(n_5548)
);

INVx1_ASAP7_75t_L g5549 ( 
.A(n_5485),
.Y(n_5549)
);

INVx1_ASAP7_75t_L g5550 ( 
.A(n_5408),
.Y(n_5550)
);

INVx2_ASAP7_75t_L g5551 ( 
.A(n_5502),
.Y(n_5551)
);

INVx2_ASAP7_75t_L g5552 ( 
.A(n_5461),
.Y(n_5552)
);

BUFx6f_ASAP7_75t_L g5553 ( 
.A(n_5409),
.Y(n_5553)
);

OAI21xp5_ASAP7_75t_L g5554 ( 
.A1(n_5390),
.A2(n_5336),
.B(n_5258),
.Y(n_5554)
);

NAND2xp5_ASAP7_75t_L g5555 ( 
.A(n_5519),
.B(n_5216),
.Y(n_5555)
);

INVx1_ASAP7_75t_L g5556 ( 
.A(n_5425),
.Y(n_5556)
);

INVx1_ASAP7_75t_L g5557 ( 
.A(n_5426),
.Y(n_5557)
);

INVx1_ASAP7_75t_L g5558 ( 
.A(n_5435),
.Y(n_5558)
);

OAI21x1_ASAP7_75t_L g5559 ( 
.A1(n_5399),
.A2(n_5293),
.B(n_5309),
.Y(n_5559)
);

INVx1_ASAP7_75t_L g5560 ( 
.A(n_5471),
.Y(n_5560)
);

INVx2_ASAP7_75t_L g5561 ( 
.A(n_5397),
.Y(n_5561)
);

BUFx2_ASAP7_75t_L g5562 ( 
.A(n_5422),
.Y(n_5562)
);

BUFx3_ASAP7_75t_L g5563 ( 
.A(n_5530),
.Y(n_5563)
);

INVx2_ASAP7_75t_L g5564 ( 
.A(n_5402),
.Y(n_5564)
);

INVx1_ASAP7_75t_L g5565 ( 
.A(n_5476),
.Y(n_5565)
);

INVx3_ASAP7_75t_L g5566 ( 
.A(n_5428),
.Y(n_5566)
);

NAND2x1p5_ASAP7_75t_L g5567 ( 
.A(n_5413),
.B(n_5097),
.Y(n_5567)
);

INVx2_ASAP7_75t_L g5568 ( 
.A(n_5417),
.Y(n_5568)
);

INVx1_ASAP7_75t_L g5569 ( 
.A(n_5482),
.Y(n_5569)
);

AOI21xp5_ASAP7_75t_SL g5570 ( 
.A1(n_5411),
.A2(n_5375),
.B(n_5299),
.Y(n_5570)
);

INVx2_ASAP7_75t_L g5571 ( 
.A(n_5438),
.Y(n_5571)
);

INVx2_ASAP7_75t_L g5572 ( 
.A(n_5440),
.Y(n_5572)
);

HB1xp67_ASAP7_75t_L g5573 ( 
.A(n_5441),
.Y(n_5573)
);

INVx5_ASAP7_75t_L g5574 ( 
.A(n_5530),
.Y(n_5574)
);

INVx1_ASAP7_75t_L g5575 ( 
.A(n_5484),
.Y(n_5575)
);

INVx1_ASAP7_75t_L g5576 ( 
.A(n_5500),
.Y(n_5576)
);

INVx2_ASAP7_75t_L g5577 ( 
.A(n_5475),
.Y(n_5577)
);

BUFx3_ASAP7_75t_L g5578 ( 
.A(n_5447),
.Y(n_5578)
);

OR2x6_ASAP7_75t_L g5579 ( 
.A(n_5434),
.B(n_5208),
.Y(n_5579)
);

INVx1_ASAP7_75t_L g5580 ( 
.A(n_5498),
.Y(n_5580)
);

BUFx2_ASAP7_75t_L g5581 ( 
.A(n_5477),
.Y(n_5581)
);

OA21x2_ASAP7_75t_L g5582 ( 
.A1(n_5444),
.A2(n_5232),
.B(n_5139),
.Y(n_5582)
);

OR2x2_ASAP7_75t_L g5583 ( 
.A(n_5529),
.B(n_5415),
.Y(n_5583)
);

INVx1_ASAP7_75t_SL g5584 ( 
.A(n_5406),
.Y(n_5584)
);

INVx2_ASAP7_75t_L g5585 ( 
.A(n_5487),
.Y(n_5585)
);

AND2x2_ASAP7_75t_L g5586 ( 
.A(n_5457),
.B(n_5350),
.Y(n_5586)
);

AO21x2_ASAP7_75t_L g5587 ( 
.A1(n_5479),
.A2(n_5149),
.B(n_5378),
.Y(n_5587)
);

NOR2xp33_ASAP7_75t_L g5588 ( 
.A(n_5481),
.B(n_5129),
.Y(n_5588)
);

INVx1_ASAP7_75t_L g5589 ( 
.A(n_5516),
.Y(n_5589)
);

INVx2_ASAP7_75t_L g5590 ( 
.A(n_5493),
.Y(n_5590)
);

INVx1_ASAP7_75t_L g5591 ( 
.A(n_5517),
.Y(n_5591)
);

INVx1_ASAP7_75t_L g5592 ( 
.A(n_5541),
.Y(n_5592)
);

NAND2xp5_ASAP7_75t_L g5593 ( 
.A(n_5519),
.B(n_5105),
.Y(n_5593)
);

AND2x2_ASAP7_75t_L g5594 ( 
.A(n_5439),
.B(n_5334),
.Y(n_5594)
);

BUFx2_ASAP7_75t_L g5595 ( 
.A(n_5497),
.Y(n_5595)
);

INVx1_ASAP7_75t_L g5596 ( 
.A(n_5463),
.Y(n_5596)
);

OA21x2_ASAP7_75t_L g5597 ( 
.A1(n_5520),
.A2(n_5168),
.B(n_5079),
.Y(n_5597)
);

INVx1_ASAP7_75t_L g5598 ( 
.A(n_5533),
.Y(n_5598)
);

INVxp67_ASAP7_75t_L g5599 ( 
.A(n_5387),
.Y(n_5599)
);

INVx1_ASAP7_75t_L g5600 ( 
.A(n_5389),
.Y(n_5600)
);

NAND2xp5_ASAP7_75t_L g5601 ( 
.A(n_5529),
.B(n_5131),
.Y(n_5601)
);

BUFx12f_ASAP7_75t_L g5602 ( 
.A(n_5453),
.Y(n_5602)
);

NAND2xp5_ASAP7_75t_L g5603 ( 
.A(n_5448),
.B(n_5421),
.Y(n_5603)
);

INVx1_ASAP7_75t_L g5604 ( 
.A(n_5510),
.Y(n_5604)
);

INVx1_ASAP7_75t_L g5605 ( 
.A(n_5539),
.Y(n_5605)
);

BUFx3_ASAP7_75t_L g5606 ( 
.A(n_5406),
.Y(n_5606)
);

INVx4_ASAP7_75t_SL g5607 ( 
.A(n_5434),
.Y(n_5607)
);

AOI21x1_ASAP7_75t_L g5608 ( 
.A1(n_5427),
.A2(n_5505),
.B(n_5385),
.Y(n_5608)
);

AND2x2_ASAP7_75t_L g5609 ( 
.A(n_5398),
.B(n_5275),
.Y(n_5609)
);

INVx2_ASAP7_75t_L g5610 ( 
.A(n_5542),
.Y(n_5610)
);

INVx1_ASAP7_75t_L g5611 ( 
.A(n_5499),
.Y(n_5611)
);

INVx2_ASAP7_75t_L g5612 ( 
.A(n_5506),
.Y(n_5612)
);

HB1xp67_ASAP7_75t_L g5613 ( 
.A(n_5394),
.Y(n_5613)
);

AO21x2_ASAP7_75t_L g5614 ( 
.A1(n_5446),
.A2(n_5169),
.B(n_5201),
.Y(n_5614)
);

BUFx2_ASAP7_75t_L g5615 ( 
.A(n_5497),
.Y(n_5615)
);

INVx3_ASAP7_75t_L g5616 ( 
.A(n_5464),
.Y(n_5616)
);

OAI21x1_ASAP7_75t_L g5617 ( 
.A1(n_5480),
.A2(n_5280),
.B(n_5135),
.Y(n_5617)
);

HB1xp67_ASAP7_75t_L g5618 ( 
.A(n_5543),
.Y(n_5618)
);

AND2x2_ASAP7_75t_L g5619 ( 
.A(n_5393),
.B(n_5225),
.Y(n_5619)
);

NOR2xp33_ASAP7_75t_R g5620 ( 
.A(n_5396),
.B(n_5152),
.Y(n_5620)
);

BUFx2_ASAP7_75t_L g5621 ( 
.A(n_5469),
.Y(n_5621)
);

INVx1_ASAP7_75t_L g5622 ( 
.A(n_5495),
.Y(n_5622)
);

INVx2_ASAP7_75t_L g5623 ( 
.A(n_5543),
.Y(n_5623)
);

INVx1_ASAP7_75t_L g5624 ( 
.A(n_5437),
.Y(n_5624)
);

INVx2_ASAP7_75t_SL g5625 ( 
.A(n_5469),
.Y(n_5625)
);

AND2x2_ASAP7_75t_L g5626 ( 
.A(n_5490),
.B(n_5220),
.Y(n_5626)
);

INVx2_ASAP7_75t_L g5627 ( 
.A(n_5459),
.Y(n_5627)
);

BUFx2_ASAP7_75t_L g5628 ( 
.A(n_5467),
.Y(n_5628)
);

INVx1_ASAP7_75t_L g5629 ( 
.A(n_5423),
.Y(n_5629)
);

OA21x2_ASAP7_75t_L g5630 ( 
.A1(n_5522),
.A2(n_5111),
.B(n_5247),
.Y(n_5630)
);

AND2x2_ASAP7_75t_L g5631 ( 
.A(n_5509),
.B(n_5298),
.Y(n_5631)
);

INVx2_ASAP7_75t_L g5632 ( 
.A(n_5429),
.Y(n_5632)
);

HB1xp67_ASAP7_75t_L g5633 ( 
.A(n_5488),
.Y(n_5633)
);

INVx1_ASAP7_75t_L g5634 ( 
.A(n_5512),
.Y(n_5634)
);

BUFx2_ASAP7_75t_L g5635 ( 
.A(n_5538),
.Y(n_5635)
);

AND2x2_ASAP7_75t_L g5636 ( 
.A(n_5405),
.B(n_5327),
.Y(n_5636)
);

INVx1_ASAP7_75t_L g5637 ( 
.A(n_5504),
.Y(n_5637)
);

HB1xp67_ASAP7_75t_L g5638 ( 
.A(n_5419),
.Y(n_5638)
);

AOI21x1_ASAP7_75t_L g5639 ( 
.A1(n_5391),
.A2(n_5283),
.B(n_5349),
.Y(n_5639)
);

HB1xp67_ASAP7_75t_L g5640 ( 
.A(n_5450),
.Y(n_5640)
);

OAI21x1_ASAP7_75t_L g5641 ( 
.A1(n_5525),
.A2(n_5148),
.B(n_5313),
.Y(n_5641)
);

INVx1_ASAP7_75t_L g5642 ( 
.A(n_5513),
.Y(n_5642)
);

HB1xp67_ASAP7_75t_L g5643 ( 
.A(n_5433),
.Y(n_5643)
);

INVx1_ASAP7_75t_L g5644 ( 
.A(n_5515),
.Y(n_5644)
);

INVx3_ASAP7_75t_L g5645 ( 
.A(n_5400),
.Y(n_5645)
);

INVx3_ASAP7_75t_L g5646 ( 
.A(n_5400),
.Y(n_5646)
);

INVx2_ASAP7_75t_L g5647 ( 
.A(n_5458),
.Y(n_5647)
);

INVx1_ASAP7_75t_L g5648 ( 
.A(n_5445),
.Y(n_5648)
);

HB1xp67_ASAP7_75t_L g5649 ( 
.A(n_5414),
.Y(n_5649)
);

INVx1_ASAP7_75t_L g5650 ( 
.A(n_5452),
.Y(n_5650)
);

INVx2_ASAP7_75t_L g5651 ( 
.A(n_5414),
.Y(n_5651)
);

INVx2_ASAP7_75t_L g5652 ( 
.A(n_5524),
.Y(n_5652)
);

CKINVDCx5p33_ASAP7_75t_R g5653 ( 
.A(n_5449),
.Y(n_5653)
);

OR2x2_ASAP7_75t_L g5654 ( 
.A(n_5491),
.B(n_5176),
.Y(n_5654)
);

INVx1_ASAP7_75t_L g5655 ( 
.A(n_5384),
.Y(n_5655)
);

BUFx3_ASAP7_75t_L g5656 ( 
.A(n_5388),
.Y(n_5656)
);

BUFx4f_ASAP7_75t_L g5657 ( 
.A(n_5395),
.Y(n_5657)
);

AND2x2_ASAP7_75t_L g5658 ( 
.A(n_5442),
.B(n_5329),
.Y(n_5658)
);

INVx2_ASAP7_75t_L g5659 ( 
.A(n_5518),
.Y(n_5659)
);

CKINVDCx5p33_ASAP7_75t_R g5660 ( 
.A(n_5527),
.Y(n_5660)
);

AND2x2_ASAP7_75t_L g5661 ( 
.A(n_5470),
.B(n_5267),
.Y(n_5661)
);

BUFx2_ASAP7_75t_L g5662 ( 
.A(n_5537),
.Y(n_5662)
);

AND2x2_ASAP7_75t_L g5663 ( 
.A(n_5468),
.B(n_5376),
.Y(n_5663)
);

INVx2_ASAP7_75t_L g5664 ( 
.A(n_5478),
.Y(n_5664)
);

BUFx2_ASAP7_75t_L g5665 ( 
.A(n_5537),
.Y(n_5665)
);

INVx1_ASAP7_75t_L g5666 ( 
.A(n_5536),
.Y(n_5666)
);

INVx1_ASAP7_75t_L g5667 ( 
.A(n_5466),
.Y(n_5667)
);

INVx1_ASAP7_75t_L g5668 ( 
.A(n_5521),
.Y(n_5668)
);

INVx2_ASAP7_75t_L g5669 ( 
.A(n_5546),
.Y(n_5669)
);

INVx1_ASAP7_75t_L g5670 ( 
.A(n_5523),
.Y(n_5670)
);

INVx1_ASAP7_75t_L g5671 ( 
.A(n_5432),
.Y(n_5671)
);

INVx1_ASAP7_75t_L g5672 ( 
.A(n_5472),
.Y(n_5672)
);

AOI22xp33_ASAP7_75t_L g5673 ( 
.A1(n_5659),
.A2(n_5383),
.B1(n_5410),
.B2(n_5386),
.Y(n_5673)
);

INVx3_ASAP7_75t_L g5674 ( 
.A(n_5574),
.Y(n_5674)
);

INVx1_ASAP7_75t_L g5675 ( 
.A(n_5549),
.Y(n_5675)
);

AOI21xp33_ASAP7_75t_L g5676 ( 
.A1(n_5614),
.A2(n_5587),
.B(n_5545),
.Y(n_5676)
);

AOI222xp33_ASAP7_75t_L g5677 ( 
.A1(n_5554),
.A2(n_5531),
.B1(n_5418),
.B2(n_5544),
.C1(n_5494),
.C2(n_5369),
.Y(n_5677)
);

BUFx12f_ASAP7_75t_L g5678 ( 
.A(n_5602),
.Y(n_5678)
);

NOR2xp33_ASAP7_75t_L g5679 ( 
.A(n_5574),
.B(n_5492),
.Y(n_5679)
);

INVx1_ASAP7_75t_L g5680 ( 
.A(n_5549),
.Y(n_5680)
);

BUFx4f_ASAP7_75t_L g5681 ( 
.A(n_5553),
.Y(n_5681)
);

AND2x4_ASAP7_75t_L g5682 ( 
.A(n_5607),
.B(n_5431),
.Y(n_5682)
);

NAND2xp5_ASAP7_75t_L g5683 ( 
.A(n_5629),
.B(n_5486),
.Y(n_5683)
);

INVx2_ASAP7_75t_L g5684 ( 
.A(n_5562),
.Y(n_5684)
);

OAI22xp33_ASAP7_75t_L g5685 ( 
.A1(n_5595),
.A2(n_5391),
.B1(n_5403),
.B2(n_5454),
.Y(n_5685)
);

AND2x4_ASAP7_75t_SL g5686 ( 
.A(n_5553),
.B(n_5118),
.Y(n_5686)
);

AOI22xp33_ASAP7_75t_L g5687 ( 
.A1(n_5663),
.A2(n_5465),
.B1(n_5508),
.B2(n_5451),
.Y(n_5687)
);

INVx1_ASAP7_75t_L g5688 ( 
.A(n_5550),
.Y(n_5688)
);

INVx3_ASAP7_75t_L g5689 ( 
.A(n_5574),
.Y(n_5689)
);

INVx1_ASAP7_75t_L g5690 ( 
.A(n_5550),
.Y(n_5690)
);

INVx3_ASAP7_75t_L g5691 ( 
.A(n_5563),
.Y(n_5691)
);

OAI22xp33_ASAP7_75t_L g5692 ( 
.A1(n_5615),
.A2(n_5348),
.B1(n_5547),
.B2(n_5460),
.Y(n_5692)
);

OAI221xp5_ASAP7_75t_L g5693 ( 
.A1(n_5639),
.A2(n_5207),
.B1(n_5507),
.B2(n_5526),
.C(n_5511),
.Y(n_5693)
);

INVx2_ASAP7_75t_L g5694 ( 
.A(n_5551),
.Y(n_5694)
);

AOI22xp33_ASAP7_75t_SL g5695 ( 
.A1(n_5581),
.A2(n_5578),
.B1(n_5628),
.B2(n_5582),
.Y(n_5695)
);

INVx2_ASAP7_75t_L g5696 ( 
.A(n_5552),
.Y(n_5696)
);

AOI21xp33_ASAP7_75t_L g5697 ( 
.A1(n_5630),
.A2(n_5307),
.B(n_5532),
.Y(n_5697)
);

BUFx2_ASAP7_75t_L g5698 ( 
.A(n_5607),
.Y(n_5698)
);

CKINVDCx5p33_ASAP7_75t_R g5699 ( 
.A(n_5620),
.Y(n_5699)
);

AOI22xp33_ASAP7_75t_L g5700 ( 
.A1(n_5631),
.A2(n_5430),
.B1(n_5404),
.B2(n_5424),
.Y(n_5700)
);

AOI22xp33_ASAP7_75t_SL g5701 ( 
.A1(n_5582),
.A2(n_5306),
.B1(n_5289),
.B2(n_5534),
.Y(n_5701)
);

NOR2xp33_ASAP7_75t_L g5702 ( 
.A(n_5553),
.B(n_5082),
.Y(n_5702)
);

AOI22xp33_ASAP7_75t_SL g5703 ( 
.A1(n_5657),
.A2(n_5289),
.B1(n_5306),
.B2(n_5376),
.Y(n_5703)
);

INVx4_ASAP7_75t_L g5704 ( 
.A(n_5657),
.Y(n_5704)
);

OAI22xp5_ASAP7_75t_SL g5705 ( 
.A1(n_5653),
.A2(n_5249),
.B1(n_5215),
.B2(n_5370),
.Y(n_5705)
);

AOI22xp33_ASAP7_75t_L g5706 ( 
.A1(n_5598),
.A2(n_5348),
.B1(n_5407),
.B2(n_5503),
.Y(n_5706)
);

NAND2xp5_ASAP7_75t_L g5707 ( 
.A(n_5624),
.B(n_5648),
.Y(n_5707)
);

AOI22xp33_ASAP7_75t_SL g5708 ( 
.A1(n_5573),
.A2(n_5332),
.B1(n_5263),
.B2(n_5266),
.Y(n_5708)
);

NAND2xp5_ASAP7_75t_L g5709 ( 
.A(n_5648),
.B(n_5472),
.Y(n_5709)
);

AOI22xp33_ASAP7_75t_L g5710 ( 
.A1(n_5601),
.A2(n_5436),
.B1(n_5443),
.B2(n_5462),
.Y(n_5710)
);

INVxp67_ASAP7_75t_L g5711 ( 
.A(n_5635),
.Y(n_5711)
);

AOI22xp5_ASAP7_75t_L g5712 ( 
.A1(n_5579),
.A2(n_5357),
.B1(n_5315),
.B2(n_5227),
.Y(n_5712)
);

INVx1_ASAP7_75t_L g5713 ( 
.A(n_5556),
.Y(n_5713)
);

OAI21x1_ASAP7_75t_SL g5714 ( 
.A1(n_5608),
.A2(n_5392),
.B(n_5401),
.Y(n_5714)
);

AOI22xp33_ASAP7_75t_L g5715 ( 
.A1(n_5593),
.A2(n_5462),
.B1(n_5235),
.B2(n_5213),
.Y(n_5715)
);

INVx1_ASAP7_75t_L g5716 ( 
.A(n_5556),
.Y(n_5716)
);

AOI221xp5_ASAP7_75t_L g5717 ( 
.A1(n_5649),
.A2(n_5528),
.B1(n_5186),
.B2(n_5147),
.C(n_5333),
.Y(n_5717)
);

AND2x2_ASAP7_75t_L g5718 ( 
.A(n_5594),
.B(n_5583),
.Y(n_5718)
);

AOI22xp33_ASAP7_75t_SL g5719 ( 
.A1(n_5586),
.A2(n_5175),
.B1(n_5299),
.B2(n_5097),
.Y(n_5719)
);

AOI22xp33_ASAP7_75t_L g5720 ( 
.A1(n_5599),
.A2(n_5473),
.B1(n_5489),
.B2(n_5175),
.Y(n_5720)
);

OA21x2_ASAP7_75t_L g5721 ( 
.A1(n_5632),
.A2(n_5474),
.B(n_5514),
.Y(n_5721)
);

BUFx2_ASAP7_75t_L g5722 ( 
.A(n_5662),
.Y(n_5722)
);

INVx1_ASAP7_75t_L g5723 ( 
.A(n_5557),
.Y(n_5723)
);

AOI21xp5_ASAP7_75t_L g5724 ( 
.A1(n_5570),
.A2(n_5456),
.B(n_5372),
.Y(n_5724)
);

INVx1_ASAP7_75t_SL g5725 ( 
.A(n_5584),
.Y(n_5725)
);

OAI221xp5_ASAP7_75t_L g5726 ( 
.A1(n_5579),
.A2(n_5496),
.B1(n_5229),
.B2(n_5548),
.C(n_5535),
.Y(n_5726)
);

NAND2xp5_ASAP7_75t_L g5727 ( 
.A(n_5650),
.B(n_5087),
.Y(n_5727)
);

BUFx8_ASAP7_75t_L g5728 ( 
.A(n_5621),
.Y(n_5728)
);

NAND2xp5_ASAP7_75t_L g5729 ( 
.A(n_5650),
.B(n_5087),
.Y(n_5729)
);

OAI221xp5_ASAP7_75t_L g5730 ( 
.A1(n_5603),
.A2(n_5286),
.B1(n_5199),
.B2(n_5412),
.C(n_5381),
.Y(n_5730)
);

AOI22xp5_ASAP7_75t_L g5731 ( 
.A1(n_5666),
.A2(n_5416),
.B1(n_5316),
.B2(n_5190),
.Y(n_5731)
);

OAI21xp33_ASAP7_75t_L g5732 ( 
.A1(n_5668),
.A2(n_5238),
.B(n_5344),
.Y(n_5732)
);

AND2x2_ASAP7_75t_SL g5733 ( 
.A(n_5665),
.B(n_5375),
.Y(n_5733)
);

AOI22xp33_ASAP7_75t_L g5734 ( 
.A1(n_5666),
.A2(n_5337),
.B1(n_5273),
.B2(n_5171),
.Y(n_5734)
);

AOI22xp33_ASAP7_75t_L g5735 ( 
.A1(n_5655),
.A2(n_5667),
.B1(n_5669),
.B2(n_5611),
.Y(n_5735)
);

AND2x2_ASAP7_75t_L g5736 ( 
.A(n_5609),
.B(n_5483),
.Y(n_5736)
);

BUFx6f_ASAP7_75t_L g5737 ( 
.A(n_5606),
.Y(n_5737)
);

NAND2xp5_ASAP7_75t_L g5738 ( 
.A(n_5637),
.B(n_5115),
.Y(n_5738)
);

CKINVDCx5p33_ASAP7_75t_R g5739 ( 
.A(n_5660),
.Y(n_5739)
);

OAI211xp5_ASAP7_75t_SL g5740 ( 
.A1(n_5668),
.A2(n_5206),
.B(n_5073),
.C(n_5172),
.Y(n_5740)
);

AOI211xp5_ASAP7_75t_L g5741 ( 
.A1(n_5588),
.A2(n_5290),
.B(n_5356),
.C(n_5455),
.Y(n_5741)
);

CKINVDCx5p33_ASAP7_75t_R g5742 ( 
.A(n_5656),
.Y(n_5742)
);

AOI22xp33_ASAP7_75t_L g5743 ( 
.A1(n_5655),
.A2(n_5115),
.B1(n_5239),
.B2(n_5292),
.Y(n_5743)
);

AOI221xp5_ASAP7_75t_L g5744 ( 
.A1(n_5667),
.A2(n_5596),
.B1(n_5651),
.B2(n_5670),
.C(n_5643),
.Y(n_5744)
);

OAI221xp5_ASAP7_75t_L g5745 ( 
.A1(n_5633),
.A2(n_5359),
.B1(n_5262),
.B2(n_5540),
.C(n_5163),
.Y(n_5745)
);

AOI222xp33_ASAP7_75t_L g5746 ( 
.A1(n_5600),
.A2(n_5159),
.B1(n_5166),
.B2(n_5196),
.C1(n_5250),
.C2(n_5136),
.Y(n_5746)
);

AOI22xp33_ASAP7_75t_SL g5747 ( 
.A1(n_5645),
.A2(n_5239),
.B1(n_5085),
.B2(n_5154),
.Y(n_5747)
);

OAI22xp5_ASAP7_75t_L g5748 ( 
.A1(n_5567),
.A2(n_5230),
.B1(n_5085),
.B2(n_5154),
.Y(n_5748)
);

INVx1_ASAP7_75t_L g5749 ( 
.A(n_5557),
.Y(n_5749)
);

AND2x2_ASAP7_75t_L g5750 ( 
.A(n_5619),
.B(n_5420),
.Y(n_5750)
);

OAI211xp5_ASAP7_75t_SL g5751 ( 
.A1(n_5670),
.A2(n_5182),
.B(n_5243),
.C(n_83),
.Y(n_5751)
);

INVx2_ASAP7_75t_L g5752 ( 
.A(n_5613),
.Y(n_5752)
);

INVx2_ASAP7_75t_L g5753 ( 
.A(n_5568),
.Y(n_5753)
);

OAI211xp5_ASAP7_75t_SL g5754 ( 
.A1(n_5654),
.A2(n_83),
.B(n_81),
.C(n_82),
.Y(n_5754)
);

OAI22xp33_ASAP7_75t_L g5755 ( 
.A1(n_5616),
.A2(n_5292),
.B1(n_5088),
.B2(n_5125),
.Y(n_5755)
);

OA21x2_ASAP7_75t_L g5756 ( 
.A1(n_5559),
.A2(n_5501),
.B(n_5089),
.Y(n_5756)
);

INVx2_ASAP7_75t_L g5757 ( 
.A(n_5571),
.Y(n_5757)
);

AOI221xp5_ASAP7_75t_L g5758 ( 
.A1(n_5642),
.A2(n_5144),
.B1(n_5305),
.B2(n_1062),
.C(n_1063),
.Y(n_5758)
);

AOI22xp33_ASAP7_75t_L g5759 ( 
.A1(n_5636),
.A2(n_5088),
.B1(n_5125),
.B2(n_5365),
.Y(n_5759)
);

AO31x2_ASAP7_75t_L g5760 ( 
.A1(n_5623),
.A2(n_5305),
.A3(n_5165),
.B(n_5211),
.Y(n_5760)
);

CKINVDCx5p33_ASAP7_75t_R g5761 ( 
.A(n_5625),
.Y(n_5761)
);

INVx3_ASAP7_75t_L g5762 ( 
.A(n_5616),
.Y(n_5762)
);

AOI22xp33_ASAP7_75t_SL g5763 ( 
.A1(n_5645),
.A2(n_5145),
.B1(n_5224),
.B2(n_5379),
.Y(n_5763)
);

OA21x2_ASAP7_75t_L g5764 ( 
.A1(n_5638),
.A2(n_5246),
.B(n_5112),
.Y(n_5764)
);

HB1xp67_ASAP7_75t_L g5765 ( 
.A(n_5640),
.Y(n_5765)
);

NAND2xp5_ASAP7_75t_L g5766 ( 
.A(n_5644),
.B(n_5634),
.Y(n_5766)
);

BUFx3_ASAP7_75t_L g5767 ( 
.A(n_5626),
.Y(n_5767)
);

AOI22xp33_ASAP7_75t_SL g5768 ( 
.A1(n_5646),
.A2(n_5377),
.B1(n_5251),
.B2(n_5341),
.Y(n_5768)
);

AOI21xp33_ASAP7_75t_L g5769 ( 
.A1(n_5630),
.A2(n_5368),
.B(n_5330),
.Y(n_5769)
);

OAI211xp5_ASAP7_75t_L g5770 ( 
.A1(n_5646),
.A2(n_5114),
.B(n_5343),
.C(n_5340),
.Y(n_5770)
);

AOI22xp33_ASAP7_75t_L g5771 ( 
.A1(n_5612),
.A2(n_5110),
.B1(n_5297),
.B2(n_5321),
.Y(n_5771)
);

AND2x2_ASAP7_75t_L g5772 ( 
.A(n_5627),
.B(n_5566),
.Y(n_5772)
);

INVxp67_ASAP7_75t_SL g5773 ( 
.A(n_5618),
.Y(n_5773)
);

BUFx10_ASAP7_75t_L g5774 ( 
.A(n_5576),
.Y(n_5774)
);

INVx3_ASAP7_75t_L g5775 ( 
.A(n_5566),
.Y(n_5775)
);

INVx1_ASAP7_75t_L g5776 ( 
.A(n_5558),
.Y(n_5776)
);

AOI21xp5_ASAP7_75t_L g5777 ( 
.A1(n_5617),
.A2(n_5257),
.B(n_5253),
.Y(n_5777)
);

AOI22xp33_ASAP7_75t_SL g5778 ( 
.A1(n_5661),
.A2(n_5281),
.B1(n_5284),
.B2(n_5264),
.Y(n_5778)
);

OAI22xp33_ASAP7_75t_L g5779 ( 
.A1(n_5555),
.A2(n_5160),
.B1(n_5211),
.B2(n_5165),
.Y(n_5779)
);

BUFx6f_ASAP7_75t_L g5780 ( 
.A(n_5678),
.Y(n_5780)
);

HB1xp67_ASAP7_75t_L g5781 ( 
.A(n_5765),
.Y(n_5781)
);

INVx2_ASAP7_75t_L g5782 ( 
.A(n_5752),
.Y(n_5782)
);

INVx2_ASAP7_75t_SL g5783 ( 
.A(n_5681),
.Y(n_5783)
);

NAND2xp5_ASAP7_75t_SL g5784 ( 
.A(n_5695),
.B(n_5672),
.Y(n_5784)
);

INVx1_ASAP7_75t_L g5785 ( 
.A(n_5707),
.Y(n_5785)
);

OR2x2_ASAP7_75t_L g5786 ( 
.A(n_5738),
.B(n_5622),
.Y(n_5786)
);

INVx1_ASAP7_75t_L g5787 ( 
.A(n_5766),
.Y(n_5787)
);

BUFx6f_ASAP7_75t_L g5788 ( 
.A(n_5704),
.Y(n_5788)
);

INVx1_ASAP7_75t_L g5789 ( 
.A(n_5675),
.Y(n_5789)
);

AND2x2_ASAP7_75t_L g5790 ( 
.A(n_5750),
.B(n_5658),
.Y(n_5790)
);

AND2x2_ASAP7_75t_L g5791 ( 
.A(n_5736),
.B(n_5647),
.Y(n_5791)
);

INVx1_ASAP7_75t_L g5792 ( 
.A(n_5680),
.Y(n_5792)
);

NOR2xp33_ASAP7_75t_L g5793 ( 
.A(n_5699),
.B(n_5565),
.Y(n_5793)
);

AND2x2_ASAP7_75t_L g5794 ( 
.A(n_5722),
.B(n_5672),
.Y(n_5794)
);

INVx3_ASAP7_75t_L g5795 ( 
.A(n_5682),
.Y(n_5795)
);

INVx2_ASAP7_75t_L g5796 ( 
.A(n_5774),
.Y(n_5796)
);

NAND2xp5_ASAP7_75t_L g5797 ( 
.A(n_5683),
.B(n_5558),
.Y(n_5797)
);

NAND2xp5_ASAP7_75t_SL g5798 ( 
.A(n_5685),
.B(n_5572),
.Y(n_5798)
);

BUFx3_ASAP7_75t_L g5799 ( 
.A(n_5686),
.Y(n_5799)
);

OR2x2_ASAP7_75t_L g5800 ( 
.A(n_5727),
.B(n_5561),
.Y(n_5800)
);

AND2x2_ASAP7_75t_L g5801 ( 
.A(n_5775),
.B(n_5564),
.Y(n_5801)
);

AND2x2_ASAP7_75t_L g5802 ( 
.A(n_5762),
.B(n_5569),
.Y(n_5802)
);

INVx1_ASAP7_75t_L g5803 ( 
.A(n_5688),
.Y(n_5803)
);

AND2x2_ASAP7_75t_L g5804 ( 
.A(n_5772),
.B(n_5575),
.Y(n_5804)
);

AND2x2_ASAP7_75t_L g5805 ( 
.A(n_5718),
.B(n_5580),
.Y(n_5805)
);

BUFx2_ASAP7_75t_L g5806 ( 
.A(n_5728),
.Y(n_5806)
);

INVx2_ASAP7_75t_L g5807 ( 
.A(n_5753),
.Y(n_5807)
);

INVx1_ASAP7_75t_L g5808 ( 
.A(n_5690),
.Y(n_5808)
);

AOI22xp33_ASAP7_75t_SL g5809 ( 
.A1(n_5698),
.A2(n_5597),
.B1(n_5671),
.B2(n_5664),
.Y(n_5809)
);

INVx2_ASAP7_75t_L g5810 ( 
.A(n_5757),
.Y(n_5810)
);

INVx1_ASAP7_75t_L g5811 ( 
.A(n_5713),
.Y(n_5811)
);

INVx1_ASAP7_75t_L g5812 ( 
.A(n_5716),
.Y(n_5812)
);

INVx2_ASAP7_75t_L g5813 ( 
.A(n_5723),
.Y(n_5813)
);

AND2x4_ASAP7_75t_L g5814 ( 
.A(n_5682),
.B(n_5671),
.Y(n_5814)
);

AND2x2_ASAP7_75t_L g5815 ( 
.A(n_5725),
.B(n_5589),
.Y(n_5815)
);

OAI221xp5_ASAP7_75t_L g5816 ( 
.A1(n_5700),
.A2(n_5560),
.B1(n_5592),
.B2(n_5591),
.C(n_5652),
.Y(n_5816)
);

AND2x2_ASAP7_75t_L g5817 ( 
.A(n_5684),
.B(n_5560),
.Y(n_5817)
);

AND2x2_ASAP7_75t_L g5818 ( 
.A(n_5711),
.B(n_5767),
.Y(n_5818)
);

INVx1_ASAP7_75t_L g5819 ( 
.A(n_5749),
.Y(n_5819)
);

NAND2xp5_ASAP7_75t_L g5820 ( 
.A(n_5735),
.B(n_5604),
.Y(n_5820)
);

INVx1_ASAP7_75t_L g5821 ( 
.A(n_5776),
.Y(n_5821)
);

NAND2xp5_ASAP7_75t_L g5822 ( 
.A(n_5710),
.B(n_5605),
.Y(n_5822)
);

OR2x2_ASAP7_75t_L g5823 ( 
.A(n_5729),
.B(n_5577),
.Y(n_5823)
);

INVx1_ASAP7_75t_L g5824 ( 
.A(n_5709),
.Y(n_5824)
);

INVx2_ASAP7_75t_L g5825 ( 
.A(n_5694),
.Y(n_5825)
);

AND2x2_ASAP7_75t_L g5826 ( 
.A(n_5691),
.B(n_5585),
.Y(n_5826)
);

INVx1_ASAP7_75t_L g5827 ( 
.A(n_5696),
.Y(n_5827)
);

INVx2_ASAP7_75t_L g5828 ( 
.A(n_5721),
.Y(n_5828)
);

OR2x2_ASAP7_75t_L g5829 ( 
.A(n_5773),
.B(n_5590),
.Y(n_5829)
);

INVx1_ASAP7_75t_L g5830 ( 
.A(n_5721),
.Y(n_5830)
);

AND2x2_ASAP7_75t_L g5831 ( 
.A(n_5737),
.B(n_5610),
.Y(n_5831)
);

HB1xp67_ASAP7_75t_L g5832 ( 
.A(n_5737),
.Y(n_5832)
);

NAND2xp5_ASAP7_75t_L g5833 ( 
.A(n_5687),
.B(n_5597),
.Y(n_5833)
);

NOR2x1_ASAP7_75t_SL g5834 ( 
.A(n_5748),
.B(n_5641),
.Y(n_5834)
);

INVx1_ASAP7_75t_L g5835 ( 
.A(n_5732),
.Y(n_5835)
);

AND2x2_ASAP7_75t_L g5836 ( 
.A(n_5737),
.B(n_5679),
.Y(n_5836)
);

NAND2x1_ASAP7_75t_L g5837 ( 
.A(n_5674),
.B(n_5689),
.Y(n_5837)
);

INVxp67_ASAP7_75t_L g5838 ( 
.A(n_5728),
.Y(n_5838)
);

NAND2xp5_ASAP7_75t_L g5839 ( 
.A(n_5759),
.B(n_5160),
.Y(n_5839)
);

INVx1_ASAP7_75t_L g5840 ( 
.A(n_5760),
.Y(n_5840)
);

INVx2_ASAP7_75t_L g5841 ( 
.A(n_5733),
.Y(n_5841)
);

OAI22xp5_ASAP7_75t_L g5842 ( 
.A1(n_5701),
.A2(n_5294),
.B1(n_5188),
.B2(n_5304),
.Y(n_5842)
);

INVx1_ASAP7_75t_L g5843 ( 
.A(n_5760),
.Y(n_5843)
);

AND2x4_ASAP7_75t_L g5844 ( 
.A(n_5720),
.B(n_5095),
.Y(n_5844)
);

HB1xp67_ASAP7_75t_L g5845 ( 
.A(n_5742),
.Y(n_5845)
);

INVx1_ASAP7_75t_L g5846 ( 
.A(n_5760),
.Y(n_5846)
);

AND2x4_ASAP7_75t_L g5847 ( 
.A(n_5724),
.B(n_5731),
.Y(n_5847)
);

HB1xp67_ASAP7_75t_L g5848 ( 
.A(n_5761),
.Y(n_5848)
);

INVx1_ASAP7_75t_L g5849 ( 
.A(n_5764),
.Y(n_5849)
);

AND2x4_ASAP7_75t_L g5850 ( 
.A(n_5777),
.B(n_5116),
.Y(n_5850)
);

NOR2xp33_ASAP7_75t_SL g5851 ( 
.A(n_5702),
.B(n_5705),
.Y(n_5851)
);

AND2x2_ASAP7_75t_L g5852 ( 
.A(n_5673),
.B(n_5180),
.Y(n_5852)
);

BUFx2_ASAP7_75t_L g5853 ( 
.A(n_5739),
.Y(n_5853)
);

INVx6_ASAP7_75t_L g5854 ( 
.A(n_5703),
.Y(n_5854)
);

AND2x2_ASAP7_75t_L g5855 ( 
.A(n_5744),
.B(n_5210),
.Y(n_5855)
);

NAND2xp5_ASAP7_75t_SL g5856 ( 
.A(n_5676),
.B(n_5219),
.Y(n_5856)
);

NAND2xp5_ASAP7_75t_L g5857 ( 
.A(n_5697),
.B(n_5715),
.Y(n_5857)
);

INVx1_ASAP7_75t_L g5858 ( 
.A(n_5764),
.Y(n_5858)
);

INVx1_ASAP7_75t_L g5859 ( 
.A(n_5813),
.Y(n_5859)
);

INVx2_ASAP7_75t_L g5860 ( 
.A(n_5829),
.Y(n_5860)
);

AND2x2_ASAP7_75t_L g5861 ( 
.A(n_5795),
.B(n_5706),
.Y(n_5861)
);

HB1xp67_ASAP7_75t_L g5862 ( 
.A(n_5781),
.Y(n_5862)
);

AND2x2_ASAP7_75t_L g5863 ( 
.A(n_5795),
.B(n_5836),
.Y(n_5863)
);

AND2x2_ASAP7_75t_L g5864 ( 
.A(n_5832),
.B(n_5719),
.Y(n_5864)
);

NAND2xp5_ASAP7_75t_L g5865 ( 
.A(n_5852),
.B(n_5835),
.Y(n_5865)
);

AOI221xp5_ASAP7_75t_L g5866 ( 
.A1(n_5857),
.A2(n_5693),
.B1(n_5726),
.B2(n_5730),
.C(n_5692),
.Y(n_5866)
);

INVx1_ASAP7_75t_L g5867 ( 
.A(n_5797),
.Y(n_5867)
);

INVx1_ASAP7_75t_L g5868 ( 
.A(n_5787),
.Y(n_5868)
);

INVx1_ASAP7_75t_L g5869 ( 
.A(n_5785),
.Y(n_5869)
);

INVx2_ASAP7_75t_L g5870 ( 
.A(n_5782),
.Y(n_5870)
);

OR2x2_ASAP7_75t_L g5871 ( 
.A(n_5786),
.B(n_5743),
.Y(n_5871)
);

AND2x2_ASAP7_75t_L g5872 ( 
.A(n_5790),
.B(n_5747),
.Y(n_5872)
);

OAI221xp5_ASAP7_75t_SL g5873 ( 
.A1(n_5816),
.A2(n_5677),
.B1(n_5712),
.B2(n_5717),
.C(n_5741),
.Y(n_5873)
);

AND2x4_ASAP7_75t_L g5874 ( 
.A(n_5799),
.B(n_5771),
.Y(n_5874)
);

NAND2xp5_ASAP7_75t_L g5875 ( 
.A(n_5855),
.B(n_5779),
.Y(n_5875)
);

AND2x2_ASAP7_75t_L g5876 ( 
.A(n_5814),
.B(n_5756),
.Y(n_5876)
);

AND2x2_ASAP7_75t_L g5877 ( 
.A(n_5814),
.B(n_5756),
.Y(n_5877)
);

AND2x2_ASAP7_75t_L g5878 ( 
.A(n_5791),
.B(n_5746),
.Y(n_5878)
);

HB1xp67_ASAP7_75t_L g5879 ( 
.A(n_5840),
.Y(n_5879)
);

INVx2_ASAP7_75t_L g5880 ( 
.A(n_5807),
.Y(n_5880)
);

AND2x4_ASAP7_75t_L g5881 ( 
.A(n_5796),
.B(n_5734),
.Y(n_5881)
);

INVx1_ASAP7_75t_L g5882 ( 
.A(n_5789),
.Y(n_5882)
);

AND2x4_ASAP7_75t_L g5883 ( 
.A(n_5818),
.B(n_5197),
.Y(n_5883)
);

AND2x2_ASAP7_75t_L g5884 ( 
.A(n_5831),
.B(n_5769),
.Y(n_5884)
);

AND2x4_ASAP7_75t_L g5885 ( 
.A(n_5788),
.B(n_5346),
.Y(n_5885)
);

INVx1_ASAP7_75t_L g5886 ( 
.A(n_5792),
.Y(n_5886)
);

NAND2xp5_ASAP7_75t_L g5887 ( 
.A(n_5839),
.B(n_5755),
.Y(n_5887)
);

INVx1_ASAP7_75t_L g5888 ( 
.A(n_5803),
.Y(n_5888)
);

BUFx2_ASAP7_75t_L g5889 ( 
.A(n_5848),
.Y(n_5889)
);

INVx2_ASAP7_75t_L g5890 ( 
.A(n_5810),
.Y(n_5890)
);

INVx1_ASAP7_75t_L g5891 ( 
.A(n_5808),
.Y(n_5891)
);

INVx1_ASAP7_75t_L g5892 ( 
.A(n_5811),
.Y(n_5892)
);

NAND2xp5_ASAP7_75t_L g5893 ( 
.A(n_5847),
.B(n_5778),
.Y(n_5893)
);

AND2x4_ASAP7_75t_L g5894 ( 
.A(n_5788),
.B(n_5352),
.Y(n_5894)
);

INVx1_ASAP7_75t_L g5895 ( 
.A(n_5812),
.Y(n_5895)
);

AND2x2_ASAP7_75t_L g5896 ( 
.A(n_5834),
.B(n_5708),
.Y(n_5896)
);

NAND2xp5_ASAP7_75t_L g5897 ( 
.A(n_5847),
.B(n_5768),
.Y(n_5897)
);

OR2x2_ASAP7_75t_L g5898 ( 
.A(n_5822),
.B(n_5770),
.Y(n_5898)
);

AND2x2_ASAP7_75t_L g5899 ( 
.A(n_5834),
.B(n_5763),
.Y(n_5899)
);

NAND2xp5_ASAP7_75t_L g5900 ( 
.A(n_5824),
.B(n_5758),
.Y(n_5900)
);

OR2x2_ASAP7_75t_L g5901 ( 
.A(n_5823),
.B(n_5745),
.Y(n_5901)
);

INVx2_ASAP7_75t_L g5902 ( 
.A(n_5825),
.Y(n_5902)
);

NAND2xp5_ASAP7_75t_L g5903 ( 
.A(n_5856),
.B(n_5714),
.Y(n_5903)
);

INVx2_ASAP7_75t_L g5904 ( 
.A(n_5800),
.Y(n_5904)
);

NAND2x1p5_ASAP7_75t_L g5905 ( 
.A(n_5806),
.B(n_5788),
.Y(n_5905)
);

NOR2xp33_ASAP7_75t_R g5906 ( 
.A(n_5780),
.B(n_81),
.Y(n_5906)
);

OR2x2_ASAP7_75t_L g5907 ( 
.A(n_5820),
.B(n_81),
.Y(n_5907)
);

NOR2xp67_ASAP7_75t_L g5908 ( 
.A(n_5841),
.B(n_82),
.Y(n_5908)
);

INVx1_ASAP7_75t_L g5909 ( 
.A(n_5819),
.Y(n_5909)
);

AND2x2_ASAP7_75t_L g5910 ( 
.A(n_5794),
.B(n_5205),
.Y(n_5910)
);

AND2x2_ASAP7_75t_L g5911 ( 
.A(n_5815),
.B(n_5802),
.Y(n_5911)
);

NAND2xp5_ASAP7_75t_L g5912 ( 
.A(n_5805),
.B(n_5361),
.Y(n_5912)
);

NAND2xp5_ASAP7_75t_L g5913 ( 
.A(n_5833),
.B(n_5363),
.Y(n_5913)
);

INVx2_ASAP7_75t_L g5914 ( 
.A(n_5828),
.Y(n_5914)
);

INVx1_ASAP7_75t_L g5915 ( 
.A(n_5821),
.Y(n_5915)
);

OR2x2_ASAP7_75t_L g5916 ( 
.A(n_5798),
.B(n_82),
.Y(n_5916)
);

INVx2_ASAP7_75t_L g5917 ( 
.A(n_5817),
.Y(n_5917)
);

HB1xp67_ASAP7_75t_L g5918 ( 
.A(n_5843),
.Y(n_5918)
);

INVx1_ASAP7_75t_L g5919 ( 
.A(n_5821),
.Y(n_5919)
);

NAND2xp5_ASAP7_75t_L g5920 ( 
.A(n_5844),
.B(n_5323),
.Y(n_5920)
);

INVx1_ASAP7_75t_SL g5921 ( 
.A(n_5853),
.Y(n_5921)
);

INVx1_ASAP7_75t_L g5922 ( 
.A(n_5846),
.Y(n_5922)
);

NAND2xp5_ASAP7_75t_L g5923 ( 
.A(n_5844),
.B(n_5324),
.Y(n_5923)
);

INVxp67_ASAP7_75t_L g5924 ( 
.A(n_5851),
.Y(n_5924)
);

OR2x6_ASAP7_75t_L g5925 ( 
.A(n_5780),
.B(n_5325),
.Y(n_5925)
);

NOR2xp33_ASAP7_75t_L g5926 ( 
.A(n_5838),
.B(n_5740),
.Y(n_5926)
);

AND2x4_ASAP7_75t_L g5927 ( 
.A(n_5783),
.B(n_1060),
.Y(n_5927)
);

OAI22xp5_ASAP7_75t_L g5928 ( 
.A1(n_5854),
.A2(n_5754),
.B1(n_5751),
.B2(n_84),
.Y(n_5928)
);

AND2x2_ASAP7_75t_L g5929 ( 
.A(n_5889),
.B(n_5854),
.Y(n_5929)
);

NOR3xp33_ASAP7_75t_L g5930 ( 
.A(n_5873),
.B(n_5842),
.C(n_5784),
.Y(n_5930)
);

INVx2_ASAP7_75t_SL g5931 ( 
.A(n_5905),
.Y(n_5931)
);

INVx1_ASAP7_75t_L g5932 ( 
.A(n_5862),
.Y(n_5932)
);

NAND2x1_ASAP7_75t_L g5933 ( 
.A(n_5899),
.B(n_5830),
.Y(n_5933)
);

NOR2xp33_ASAP7_75t_L g5934 ( 
.A(n_5924),
.B(n_5780),
.Y(n_5934)
);

OAI33xp33_ASAP7_75t_L g5935 ( 
.A1(n_5875),
.A2(n_5858),
.A3(n_5849),
.B1(n_5827),
.B2(n_5809),
.B3(n_5793),
.Y(n_5935)
);

INVx1_ASAP7_75t_L g5936 ( 
.A(n_5879),
.Y(n_5936)
);

AND2x4_ASAP7_75t_L g5937 ( 
.A(n_5921),
.B(n_5845),
.Y(n_5937)
);

HB1xp67_ASAP7_75t_L g5938 ( 
.A(n_5918),
.Y(n_5938)
);

INVx3_ASAP7_75t_L g5939 ( 
.A(n_5927),
.Y(n_5939)
);

AND2x4_ASAP7_75t_L g5940 ( 
.A(n_5863),
.B(n_5837),
.Y(n_5940)
);

NAND3xp33_ASAP7_75t_L g5941 ( 
.A(n_5926),
.B(n_5858),
.C(n_5850),
.Y(n_5941)
);

INVx1_ASAP7_75t_L g5942 ( 
.A(n_5916),
.Y(n_5942)
);

OR2x2_ASAP7_75t_L g5943 ( 
.A(n_5900),
.B(n_5850),
.Y(n_5943)
);

INVx2_ASAP7_75t_SL g5944 ( 
.A(n_5927),
.Y(n_5944)
);

NAND3xp33_ASAP7_75t_L g5945 ( 
.A(n_5866),
.B(n_5826),
.C(n_5801),
.Y(n_5945)
);

AND2x2_ASAP7_75t_L g5946 ( 
.A(n_5864),
.B(n_5804),
.Y(n_5946)
);

INVx1_ASAP7_75t_SL g5947 ( 
.A(n_5906),
.Y(n_5947)
);

AND2x4_ASAP7_75t_SL g5948 ( 
.A(n_5874),
.B(n_82),
.Y(n_5948)
);

NAND2xp5_ASAP7_75t_L g5949 ( 
.A(n_5881),
.B(n_83),
.Y(n_5949)
);

OAI221xp5_ASAP7_75t_L g5950 ( 
.A1(n_5893),
.A2(n_86),
.B1(n_84),
.B2(n_85),
.C(n_87),
.Y(n_5950)
);

AND2x2_ASAP7_75t_L g5951 ( 
.A(n_5874),
.B(n_84),
.Y(n_5951)
);

INVx3_ASAP7_75t_L g5952 ( 
.A(n_5860),
.Y(n_5952)
);

OAI33xp33_ASAP7_75t_L g5953 ( 
.A1(n_5887),
.A2(n_87),
.A3(n_89),
.B1(n_85),
.B2(n_86),
.B3(n_88),
.Y(n_5953)
);

NOR3xp33_ASAP7_75t_SL g5954 ( 
.A(n_5928),
.B(n_85),
.C(n_86),
.Y(n_5954)
);

OAI22xp5_ASAP7_75t_L g5955 ( 
.A1(n_5897),
.A2(n_87),
.B1(n_85),
.B2(n_86),
.Y(n_5955)
);

AND2x2_ASAP7_75t_L g5956 ( 
.A(n_5861),
.B(n_87),
.Y(n_5956)
);

AND2x2_ASAP7_75t_L g5957 ( 
.A(n_5896),
.B(n_88),
.Y(n_5957)
);

AND2x4_ASAP7_75t_L g5958 ( 
.A(n_5881),
.B(n_1060),
.Y(n_5958)
);

AND2x2_ASAP7_75t_L g5959 ( 
.A(n_5911),
.B(n_88),
.Y(n_5959)
);

AOI322xp5_ASAP7_75t_L g5960 ( 
.A1(n_5865),
.A2(n_1096),
.A3(n_1095),
.B1(n_1094),
.B2(n_1093),
.C1(n_1091),
.C2(n_1090),
.Y(n_5960)
);

AND2x2_ASAP7_75t_L g5961 ( 
.A(n_5884),
.B(n_88),
.Y(n_5961)
);

HB1xp67_ASAP7_75t_L g5962 ( 
.A(n_5914),
.Y(n_5962)
);

AND2x2_ASAP7_75t_L g5963 ( 
.A(n_5910),
.B(n_89),
.Y(n_5963)
);

AND2x2_ASAP7_75t_L g5964 ( 
.A(n_5872),
.B(n_90),
.Y(n_5964)
);

OR2x2_ASAP7_75t_L g5965 ( 
.A(n_5913),
.B(n_90),
.Y(n_5965)
);

NAND3xp33_ASAP7_75t_L g5966 ( 
.A(n_5903),
.B(n_90),
.C(n_91),
.Y(n_5966)
);

NAND2xp33_ASAP7_75t_L g5967 ( 
.A(n_5907),
.B(n_91),
.Y(n_5967)
);

AND2x2_ASAP7_75t_L g5968 ( 
.A(n_5904),
.B(n_91),
.Y(n_5968)
);

OR2x2_ASAP7_75t_L g5969 ( 
.A(n_5867),
.B(n_91),
.Y(n_5969)
);

INVx1_ASAP7_75t_L g5970 ( 
.A(n_5868),
.Y(n_5970)
);

AND2x2_ASAP7_75t_L g5971 ( 
.A(n_5883),
.B(n_92),
.Y(n_5971)
);

INVx2_ASAP7_75t_L g5972 ( 
.A(n_5880),
.Y(n_5972)
);

NOR3xp33_ASAP7_75t_L g5973 ( 
.A(n_5898),
.B(n_5923),
.C(n_5920),
.Y(n_5973)
);

NAND2xp5_ASAP7_75t_L g5974 ( 
.A(n_5964),
.B(n_5869),
.Y(n_5974)
);

AND2x4_ASAP7_75t_L g5975 ( 
.A(n_5937),
.B(n_5925),
.Y(n_5975)
);

NAND2xp5_ASAP7_75t_L g5976 ( 
.A(n_5951),
.B(n_5878),
.Y(n_5976)
);

AND2x2_ASAP7_75t_L g5977 ( 
.A(n_5934),
.B(n_5883),
.Y(n_5977)
);

INVxp67_ASAP7_75t_L g5978 ( 
.A(n_5937),
.Y(n_5978)
);

AND2x2_ASAP7_75t_L g5979 ( 
.A(n_5929),
.B(n_5901),
.Y(n_5979)
);

INVx1_ASAP7_75t_L g5980 ( 
.A(n_5938),
.Y(n_5980)
);

AND2x4_ASAP7_75t_L g5981 ( 
.A(n_5944),
.B(n_5925),
.Y(n_5981)
);

HB1xp67_ASAP7_75t_L g5982 ( 
.A(n_5932),
.Y(n_5982)
);

NOR2xp67_ASAP7_75t_SL g5983 ( 
.A(n_5939),
.B(n_5912),
.Y(n_5983)
);

NAND2xp5_ASAP7_75t_L g5984 ( 
.A(n_5930),
.B(n_5956),
.Y(n_5984)
);

INVxp67_ASAP7_75t_L g5985 ( 
.A(n_5949),
.Y(n_5985)
);

AND2x2_ASAP7_75t_L g5986 ( 
.A(n_5948),
.B(n_5871),
.Y(n_5986)
);

NAND2xp5_ASAP7_75t_L g5987 ( 
.A(n_5963),
.B(n_5882),
.Y(n_5987)
);

OR2x2_ASAP7_75t_L g5988 ( 
.A(n_5965),
.B(n_5886),
.Y(n_5988)
);

NAND2xp5_ASAP7_75t_L g5989 ( 
.A(n_5961),
.B(n_5888),
.Y(n_5989)
);

NAND2xp5_ASAP7_75t_L g5990 ( 
.A(n_5957),
.B(n_5891),
.Y(n_5990)
);

AND2x4_ASAP7_75t_L g5991 ( 
.A(n_5939),
.B(n_5885),
.Y(n_5991)
);

NAND2xp5_ASAP7_75t_L g5992 ( 
.A(n_5958),
.B(n_5892),
.Y(n_5992)
);

AND3x2_ASAP7_75t_L g5993 ( 
.A(n_5958),
.B(n_5894),
.C(n_5885),
.Y(n_5993)
);

AOI22xp33_ASAP7_75t_L g5994 ( 
.A1(n_5973),
.A2(n_5935),
.B1(n_5931),
.B2(n_5945),
.Y(n_5994)
);

NAND3xp33_ASAP7_75t_L g5995 ( 
.A(n_5960),
.B(n_5922),
.C(n_5894),
.Y(n_5995)
);

NOR2xp67_ASAP7_75t_L g5996 ( 
.A(n_5941),
.B(n_5876),
.Y(n_5996)
);

NOR2x1_ASAP7_75t_L g5997 ( 
.A(n_5966),
.B(n_5908),
.Y(n_5997)
);

AOI22xp5_ASAP7_75t_L g5998 ( 
.A1(n_5955),
.A2(n_5895),
.B1(n_5909),
.B2(n_5877),
.Y(n_5998)
);

AND2x2_ASAP7_75t_L g5999 ( 
.A(n_5940),
.B(n_5917),
.Y(n_5999)
);

OR2x2_ASAP7_75t_L g6000 ( 
.A(n_5942),
.B(n_5870),
.Y(n_6000)
);

INVx1_ASAP7_75t_L g6001 ( 
.A(n_5971),
.Y(n_6001)
);

AND2x2_ASAP7_75t_L g6002 ( 
.A(n_5940),
.B(n_5890),
.Y(n_6002)
);

HB1xp67_ASAP7_75t_L g6003 ( 
.A(n_5962),
.Y(n_6003)
);

INVx1_ASAP7_75t_L g6004 ( 
.A(n_5968),
.Y(n_6004)
);

NAND2xp5_ASAP7_75t_L g6005 ( 
.A(n_5936),
.B(n_5959),
.Y(n_6005)
);

INVx1_ASAP7_75t_L g6006 ( 
.A(n_5969),
.Y(n_6006)
);

INVx2_ASAP7_75t_L g6007 ( 
.A(n_5952),
.Y(n_6007)
);

AND2x2_ASAP7_75t_L g6008 ( 
.A(n_5946),
.B(n_5902),
.Y(n_6008)
);

NAND2xp5_ASAP7_75t_L g6009 ( 
.A(n_5970),
.B(n_5859),
.Y(n_6009)
);

AND2x4_ASAP7_75t_L g6010 ( 
.A(n_5947),
.B(n_5859),
.Y(n_6010)
);

OR2x2_ASAP7_75t_L g6011 ( 
.A(n_5980),
.B(n_5933),
.Y(n_6011)
);

INVx1_ASAP7_75t_L g6012 ( 
.A(n_6003),
.Y(n_6012)
);

INVx1_ASAP7_75t_SL g6013 ( 
.A(n_6010),
.Y(n_6013)
);

INVx1_ASAP7_75t_L g6014 ( 
.A(n_5982),
.Y(n_6014)
);

AND2x2_ASAP7_75t_L g6015 ( 
.A(n_5979),
.B(n_5978),
.Y(n_6015)
);

NAND2xp5_ASAP7_75t_L g6016 ( 
.A(n_6010),
.B(n_5954),
.Y(n_6016)
);

AND2x4_ASAP7_75t_L g6017 ( 
.A(n_5975),
.B(n_5972),
.Y(n_6017)
);

AND2x2_ASAP7_75t_L g6018 ( 
.A(n_5986),
.B(n_5943),
.Y(n_6018)
);

INVx2_ASAP7_75t_SL g6019 ( 
.A(n_5975),
.Y(n_6019)
);

INVx1_ASAP7_75t_L g6020 ( 
.A(n_6000),
.Y(n_6020)
);

INVx1_ASAP7_75t_L g6021 ( 
.A(n_6004),
.Y(n_6021)
);

INVx1_ASAP7_75t_L g6022 ( 
.A(n_6001),
.Y(n_6022)
);

AND2x2_ASAP7_75t_L g6023 ( 
.A(n_5977),
.B(n_5933),
.Y(n_6023)
);

AND2x2_ASAP7_75t_L g6024 ( 
.A(n_6002),
.B(n_5967),
.Y(n_6024)
);

AND2x2_ASAP7_75t_L g6025 ( 
.A(n_6008),
.B(n_5915),
.Y(n_6025)
);

INVx1_ASAP7_75t_L g6026 ( 
.A(n_6009),
.Y(n_6026)
);

INVx1_ASAP7_75t_SL g6027 ( 
.A(n_5981),
.Y(n_6027)
);

AND2x2_ASAP7_75t_L g6028 ( 
.A(n_6007),
.B(n_5919),
.Y(n_6028)
);

NAND2xp5_ASAP7_75t_L g6029 ( 
.A(n_5994),
.B(n_5950),
.Y(n_6029)
);

AND2x2_ASAP7_75t_L g6030 ( 
.A(n_5999),
.B(n_92),
.Y(n_6030)
);

OR2x2_ASAP7_75t_L g6031 ( 
.A(n_6006),
.B(n_92),
.Y(n_6031)
);

OR2x2_ASAP7_75t_L g6032 ( 
.A(n_6005),
.B(n_92),
.Y(n_6032)
);

INVx1_ASAP7_75t_L g6033 ( 
.A(n_5988),
.Y(n_6033)
);

AND2x2_ASAP7_75t_L g6034 ( 
.A(n_5981),
.B(n_93),
.Y(n_6034)
);

OR2x2_ASAP7_75t_L g6035 ( 
.A(n_5974),
.B(n_93),
.Y(n_6035)
);

NAND2xp5_ASAP7_75t_L g6036 ( 
.A(n_5984),
.B(n_5953),
.Y(n_6036)
);

INVx1_ASAP7_75t_L g6037 ( 
.A(n_5992),
.Y(n_6037)
);

OR2x2_ASAP7_75t_L g6038 ( 
.A(n_5989),
.B(n_93),
.Y(n_6038)
);

AND2x2_ASAP7_75t_L g6039 ( 
.A(n_5996),
.B(n_94),
.Y(n_6039)
);

NOR2xp33_ASAP7_75t_L g6040 ( 
.A(n_5976),
.B(n_94),
.Y(n_6040)
);

OAI21xp33_ASAP7_75t_L g6041 ( 
.A1(n_5998),
.A2(n_94),
.B(n_95),
.Y(n_6041)
);

INVx1_ASAP7_75t_L g6042 ( 
.A(n_5990),
.Y(n_6042)
);

INVx1_ASAP7_75t_L g6043 ( 
.A(n_5987),
.Y(n_6043)
);

INVx2_ASAP7_75t_L g6044 ( 
.A(n_5991),
.Y(n_6044)
);

NAND2xp5_ASAP7_75t_L g6045 ( 
.A(n_5985),
.B(n_95),
.Y(n_6045)
);

OR2x2_ASAP7_75t_L g6046 ( 
.A(n_5995),
.B(n_95),
.Y(n_6046)
);

AND2x2_ASAP7_75t_L g6047 ( 
.A(n_5997),
.B(n_5991),
.Y(n_6047)
);

OR2x2_ASAP7_75t_L g6048 ( 
.A(n_5983),
.B(n_95),
.Y(n_6048)
);

OR2x2_ASAP7_75t_L g6049 ( 
.A(n_5993),
.B(n_96),
.Y(n_6049)
);

AOI22xp33_ASAP7_75t_L g6050 ( 
.A1(n_5979),
.A2(n_1062),
.B1(n_1063),
.B2(n_1061),
.Y(n_6050)
);

INVx1_ASAP7_75t_L g6051 ( 
.A(n_6012),
.Y(n_6051)
);

AOI22xp5_ASAP7_75t_L g6052 ( 
.A1(n_6027),
.A2(n_98),
.B1(n_96),
.B2(n_97),
.Y(n_6052)
);

NAND2xp5_ASAP7_75t_L g6053 ( 
.A(n_6013),
.B(n_96),
.Y(n_6053)
);

INVx1_ASAP7_75t_L g6054 ( 
.A(n_6034),
.Y(n_6054)
);

INVx2_ASAP7_75t_SL g6055 ( 
.A(n_6017),
.Y(n_6055)
);

INVx2_ASAP7_75t_L g6056 ( 
.A(n_6044),
.Y(n_6056)
);

INVx3_ASAP7_75t_SL g6057 ( 
.A(n_6019),
.Y(n_6057)
);

AOI21xp5_ASAP7_75t_L g6058 ( 
.A1(n_6016),
.A2(n_97),
.B(n_98),
.Y(n_6058)
);

NAND2xp5_ASAP7_75t_L g6059 ( 
.A(n_6015),
.B(n_97),
.Y(n_6059)
);

AND2x2_ASAP7_75t_L g6060 ( 
.A(n_6023),
.B(n_97),
.Y(n_6060)
);

INVx2_ASAP7_75t_L g6061 ( 
.A(n_6017),
.Y(n_6061)
);

BUFx2_ASAP7_75t_L g6062 ( 
.A(n_6018),
.Y(n_6062)
);

INVx2_ASAP7_75t_L g6063 ( 
.A(n_6012),
.Y(n_6063)
);

AOI21xp33_ASAP7_75t_SL g6064 ( 
.A1(n_6049),
.A2(n_98),
.B(n_99),
.Y(n_6064)
);

NOR2xp33_ASAP7_75t_L g6065 ( 
.A(n_6046),
.B(n_98),
.Y(n_6065)
);

NAND2xp5_ASAP7_75t_L g6066 ( 
.A(n_6039),
.B(n_99),
.Y(n_6066)
);

AOI22xp33_ASAP7_75t_SL g6067 ( 
.A1(n_6047),
.A2(n_101),
.B1(n_99),
.B2(n_100),
.Y(n_6067)
);

NOR2xp33_ASAP7_75t_L g6068 ( 
.A(n_6048),
.B(n_6041),
.Y(n_6068)
);

BUFx3_ASAP7_75t_L g6069 ( 
.A(n_6014),
.Y(n_6069)
);

AOI22xp5_ASAP7_75t_L g6070 ( 
.A1(n_6024),
.A2(n_102),
.B1(n_100),
.B2(n_101),
.Y(n_6070)
);

AOI32xp33_ASAP7_75t_L g6071 ( 
.A1(n_6029),
.A2(n_103),
.A3(n_100),
.B1(n_102),
.B2(n_104),
.Y(n_6071)
);

INVx1_ASAP7_75t_L g6072 ( 
.A(n_6030),
.Y(n_6072)
);

AND2x4_ASAP7_75t_L g6073 ( 
.A(n_6020),
.B(n_100),
.Y(n_6073)
);

AOI222xp33_ASAP7_75t_L g6074 ( 
.A1(n_6036),
.A2(n_105),
.B1(n_107),
.B2(n_103),
.C1(n_104),
.C2(n_106),
.Y(n_6074)
);

INVx2_ASAP7_75t_L g6075 ( 
.A(n_6028),
.Y(n_6075)
);

INVxp67_ASAP7_75t_SL g6076 ( 
.A(n_6045),
.Y(n_6076)
);

INVx1_ASAP7_75t_L g6077 ( 
.A(n_6031),
.Y(n_6077)
);

AND2x2_ASAP7_75t_L g6078 ( 
.A(n_6025),
.B(n_103),
.Y(n_6078)
);

HB1xp67_ASAP7_75t_L g6079 ( 
.A(n_6033),
.Y(n_6079)
);

INVx1_ASAP7_75t_L g6080 ( 
.A(n_6032),
.Y(n_6080)
);

INVx1_ASAP7_75t_L g6081 ( 
.A(n_6011),
.Y(n_6081)
);

INVx2_ASAP7_75t_L g6082 ( 
.A(n_6035),
.Y(n_6082)
);

INVx1_ASAP7_75t_L g6083 ( 
.A(n_6038),
.Y(n_6083)
);

INVx2_ASAP7_75t_SL g6084 ( 
.A(n_6021),
.Y(n_6084)
);

NAND2xp5_ASAP7_75t_L g6085 ( 
.A(n_6040),
.B(n_103),
.Y(n_6085)
);

INVx1_ASAP7_75t_L g6086 ( 
.A(n_6037),
.Y(n_6086)
);

AO22x1_ASAP7_75t_L g6087 ( 
.A1(n_6042),
.A2(n_106),
.B1(n_104),
.B2(n_105),
.Y(n_6087)
);

OR2x2_ASAP7_75t_L g6088 ( 
.A(n_6042),
.B(n_104),
.Y(n_6088)
);

INVx1_ASAP7_75t_L g6089 ( 
.A(n_6022),
.Y(n_6089)
);

INVx1_ASAP7_75t_L g6090 ( 
.A(n_6026),
.Y(n_6090)
);

INVx2_ASAP7_75t_L g6091 ( 
.A(n_6026),
.Y(n_6091)
);

INVxp67_ASAP7_75t_L g6092 ( 
.A(n_6043),
.Y(n_6092)
);

INVx1_ASAP7_75t_L g6093 ( 
.A(n_6050),
.Y(n_6093)
);

NAND2xp5_ASAP7_75t_L g6094 ( 
.A(n_6057),
.B(n_106),
.Y(n_6094)
);

NAND2xp5_ASAP7_75t_L g6095 ( 
.A(n_6062),
.B(n_107),
.Y(n_6095)
);

NAND2xp5_ASAP7_75t_L g6096 ( 
.A(n_6055),
.B(n_107),
.Y(n_6096)
);

OR2x2_ASAP7_75t_L g6097 ( 
.A(n_6059),
.B(n_6053),
.Y(n_6097)
);

NAND2xp33_ASAP7_75t_L g6098 ( 
.A(n_6061),
.B(n_107),
.Y(n_6098)
);

NOR2xp33_ASAP7_75t_L g6099 ( 
.A(n_6064),
.B(n_108),
.Y(n_6099)
);

NAND2xp5_ASAP7_75t_L g6100 ( 
.A(n_6087),
.B(n_108),
.Y(n_6100)
);

INVx1_ASAP7_75t_L g6101 ( 
.A(n_6056),
.Y(n_6101)
);

NAND2xp5_ASAP7_75t_SL g6102 ( 
.A(n_6074),
.B(n_108),
.Y(n_6102)
);

INVx1_ASAP7_75t_L g6103 ( 
.A(n_6073),
.Y(n_6103)
);

OAI22xp5_ASAP7_75t_L g6104 ( 
.A1(n_6093),
.A2(n_111),
.B1(n_109),
.B2(n_110),
.Y(n_6104)
);

NAND3xp33_ASAP7_75t_L g6105 ( 
.A(n_6071),
.B(n_109),
.C(n_110),
.Y(n_6105)
);

NAND2xp5_ASAP7_75t_L g6106 ( 
.A(n_6060),
.B(n_109),
.Y(n_6106)
);

OAI22xp5_ASAP7_75t_L g6107 ( 
.A1(n_6093),
.A2(n_111),
.B1(n_109),
.B2(n_110),
.Y(n_6107)
);

NAND2xp5_ASAP7_75t_L g6108 ( 
.A(n_6067),
.B(n_6073),
.Y(n_6108)
);

INVx1_ASAP7_75t_L g6109 ( 
.A(n_6079),
.Y(n_6109)
);

O2A1O1Ixp33_ASAP7_75t_L g6110 ( 
.A1(n_6092),
.A2(n_113),
.B(n_111),
.C(n_112),
.Y(n_6110)
);

INVx1_ASAP7_75t_L g6111 ( 
.A(n_6081),
.Y(n_6111)
);

OAI21xp5_ASAP7_75t_L g6112 ( 
.A1(n_6058),
.A2(n_111),
.B(n_112),
.Y(n_6112)
);

NOR2xp33_ASAP7_75t_L g6113 ( 
.A(n_6072),
.B(n_112),
.Y(n_6113)
);

AOI22xp5_ASAP7_75t_L g6114 ( 
.A1(n_6065),
.A2(n_115),
.B1(n_113),
.B2(n_114),
.Y(n_6114)
);

NAND2xp5_ASAP7_75t_L g6115 ( 
.A(n_6078),
.B(n_113),
.Y(n_6115)
);

NAND2xp5_ASAP7_75t_L g6116 ( 
.A(n_6052),
.B(n_113),
.Y(n_6116)
);

OR2x2_ASAP7_75t_L g6117 ( 
.A(n_6088),
.B(n_114),
.Y(n_6117)
);

AOI22xp5_ASAP7_75t_L g6118 ( 
.A1(n_6068),
.A2(n_116),
.B1(n_114),
.B2(n_115),
.Y(n_6118)
);

NOR3xp33_ASAP7_75t_SL g6119 ( 
.A(n_6086),
.B(n_114),
.C(n_115),
.Y(n_6119)
);

INVx1_ASAP7_75t_L g6120 ( 
.A(n_6069),
.Y(n_6120)
);

OAI321xp33_ASAP7_75t_L g6121 ( 
.A1(n_6051),
.A2(n_115),
.A3(n_116),
.B1(n_117),
.B2(n_118),
.C(n_119),
.Y(n_6121)
);

INVxp67_ASAP7_75t_SL g6122 ( 
.A(n_6066),
.Y(n_6122)
);

O2A1O1Ixp33_ASAP7_75t_SL g6123 ( 
.A1(n_6054),
.A2(n_6084),
.B(n_6077),
.C(n_6080),
.Y(n_6123)
);

AO32x1_ASAP7_75t_L g6124 ( 
.A1(n_6082),
.A2(n_118),
.A3(n_116),
.B1(n_117),
.B2(n_119),
.Y(n_6124)
);

AOI22xp5_ASAP7_75t_L g6125 ( 
.A1(n_6070),
.A2(n_119),
.B1(n_117),
.B2(n_118),
.Y(n_6125)
);

HB1xp67_ASAP7_75t_L g6126 ( 
.A(n_6063),
.Y(n_6126)
);

INVx1_ASAP7_75t_L g6127 ( 
.A(n_6051),
.Y(n_6127)
);

INVx2_ASAP7_75t_L g6128 ( 
.A(n_6075),
.Y(n_6128)
);

NAND2xp5_ASAP7_75t_SL g6129 ( 
.A(n_6091),
.B(n_117),
.Y(n_6129)
);

INVx2_ASAP7_75t_L g6130 ( 
.A(n_6083),
.Y(n_6130)
);

INVx1_ASAP7_75t_L g6131 ( 
.A(n_6085),
.Y(n_6131)
);

INVxp67_ASAP7_75t_L g6132 ( 
.A(n_6076),
.Y(n_6132)
);

NAND2xp5_ASAP7_75t_L g6133 ( 
.A(n_6090),
.B(n_118),
.Y(n_6133)
);

INVx1_ASAP7_75t_L g6134 ( 
.A(n_6089),
.Y(n_6134)
);

INVxp67_ASAP7_75t_L g6135 ( 
.A(n_6062),
.Y(n_6135)
);

NAND3xp33_ASAP7_75t_L g6136 ( 
.A(n_6074),
.B(n_119),
.C(n_120),
.Y(n_6136)
);

NOR2xp67_ASAP7_75t_L g6137 ( 
.A(n_6055),
.B(n_120),
.Y(n_6137)
);

INVx2_ASAP7_75t_SL g6138 ( 
.A(n_6057),
.Y(n_6138)
);

NAND2xp5_ASAP7_75t_L g6139 ( 
.A(n_6057),
.B(n_120),
.Y(n_6139)
);

INVx1_ASAP7_75t_L g6140 ( 
.A(n_6053),
.Y(n_6140)
);

NAND2xp5_ASAP7_75t_L g6141 ( 
.A(n_6057),
.B(n_121),
.Y(n_6141)
);

A2O1A1Ixp33_ASAP7_75t_L g6142 ( 
.A1(n_6068),
.A2(n_123),
.B(n_121),
.C(n_122),
.Y(n_6142)
);

INVx1_ASAP7_75t_L g6143 ( 
.A(n_6053),
.Y(n_6143)
);

AOI22xp5_ASAP7_75t_L g6144 ( 
.A1(n_6057),
.A2(n_123),
.B1(n_121),
.B2(n_122),
.Y(n_6144)
);

OR2x2_ASAP7_75t_L g6145 ( 
.A(n_6062),
.B(n_122),
.Y(n_6145)
);

NAND4xp25_ASAP7_75t_L g6146 ( 
.A(n_6062),
.B(n_125),
.C(n_123),
.D(n_124),
.Y(n_6146)
);

HB1xp67_ASAP7_75t_L g6147 ( 
.A(n_6056),
.Y(n_6147)
);

OAI21xp33_ASAP7_75t_L g6148 ( 
.A1(n_6055),
.A2(n_123),
.B(n_124),
.Y(n_6148)
);

INVx1_ASAP7_75t_L g6149 ( 
.A(n_6053),
.Y(n_6149)
);

INVx1_ASAP7_75t_L g6150 ( 
.A(n_6053),
.Y(n_6150)
);

O2A1O1Ixp33_ASAP7_75t_L g6151 ( 
.A1(n_6057),
.A2(n_128),
.B(n_126),
.C(n_127),
.Y(n_6151)
);

AOI22xp5_ASAP7_75t_L g6152 ( 
.A1(n_6057),
.A2(n_128),
.B1(n_126),
.B2(n_127),
.Y(n_6152)
);

INVx1_ASAP7_75t_L g6153 ( 
.A(n_6053),
.Y(n_6153)
);

NAND2xp5_ASAP7_75t_L g6154 ( 
.A(n_6057),
.B(n_126),
.Y(n_6154)
);

NOR2xp33_ASAP7_75t_L g6155 ( 
.A(n_6057),
.B(n_126),
.Y(n_6155)
);

OAI322xp33_ASAP7_75t_L g6156 ( 
.A1(n_6081),
.A2(n_127),
.A3(n_128),
.B1(n_129),
.B2(n_130),
.C1(n_131),
.C2(n_132),
.Y(n_6156)
);

AOI22xp5_ASAP7_75t_L g6157 ( 
.A1(n_6138),
.A2(n_129),
.B1(n_127),
.B2(n_128),
.Y(n_6157)
);

NAND2xp33_ASAP7_75t_R g6158 ( 
.A(n_6119),
.B(n_129),
.Y(n_6158)
);

INVx1_ASAP7_75t_SL g6159 ( 
.A(n_6147),
.Y(n_6159)
);

XNOR2x1_ASAP7_75t_L g6160 ( 
.A(n_6104),
.B(n_130),
.Y(n_6160)
);

NAND2xp5_ASAP7_75t_L g6161 ( 
.A(n_6155),
.B(n_130),
.Y(n_6161)
);

HB1xp67_ASAP7_75t_L g6162 ( 
.A(n_6094),
.Y(n_6162)
);

INVx1_ASAP7_75t_L g6163 ( 
.A(n_6139),
.Y(n_6163)
);

NAND2xp5_ASAP7_75t_L g6164 ( 
.A(n_6137),
.B(n_130),
.Y(n_6164)
);

INVx2_ASAP7_75t_L g6165 ( 
.A(n_6101),
.Y(n_6165)
);

OAI21xp33_ASAP7_75t_L g6166 ( 
.A1(n_6120),
.A2(n_131),
.B(n_132),
.Y(n_6166)
);

NAND3xp33_ASAP7_75t_L g6167 ( 
.A(n_6136),
.B(n_131),
.C(n_132),
.Y(n_6167)
);

INVx1_ASAP7_75t_L g6168 ( 
.A(n_6141),
.Y(n_6168)
);

INVx1_ASAP7_75t_SL g6169 ( 
.A(n_6154),
.Y(n_6169)
);

NAND4xp25_ASAP7_75t_L g6170 ( 
.A(n_6108),
.B(n_133),
.C(n_131),
.D(n_132),
.Y(n_6170)
);

AND2x2_ASAP7_75t_L g6171 ( 
.A(n_6135),
.B(n_133),
.Y(n_6171)
);

NAND2xp5_ASAP7_75t_L g6172 ( 
.A(n_6099),
.B(n_133),
.Y(n_6172)
);

OAI322xp33_ASAP7_75t_L g6173 ( 
.A1(n_6132),
.A2(n_133),
.A3(n_134),
.B1(n_135),
.B2(n_136),
.C1(n_137),
.C2(n_138),
.Y(n_6173)
);

NAND2xp5_ASAP7_75t_L g6174 ( 
.A(n_6148),
.B(n_134),
.Y(n_6174)
);

OAI21xp33_ASAP7_75t_SL g6175 ( 
.A1(n_6109),
.A2(n_134),
.B(n_135),
.Y(n_6175)
);

OR2x2_ASAP7_75t_L g6176 ( 
.A(n_6100),
.B(n_134),
.Y(n_6176)
);

OR4x1_ASAP7_75t_L g6177 ( 
.A(n_6103),
.B(n_137),
.C(n_135),
.D(n_136),
.Y(n_6177)
);

INVx1_ASAP7_75t_SL g6178 ( 
.A(n_6096),
.Y(n_6178)
);

INVx1_ASAP7_75t_L g6179 ( 
.A(n_6124),
.Y(n_6179)
);

AOI22xp5_ASAP7_75t_L g6180 ( 
.A1(n_6107),
.A2(n_138),
.B1(n_135),
.B2(n_137),
.Y(n_6180)
);

AOI22xp5_ASAP7_75t_L g6181 ( 
.A1(n_6146),
.A2(n_139),
.B1(n_137),
.B2(n_138),
.Y(n_6181)
);

OR2x2_ASAP7_75t_L g6182 ( 
.A(n_6095),
.B(n_138),
.Y(n_6182)
);

NOR2xp33_ASAP7_75t_L g6183 ( 
.A(n_6102),
.B(n_139),
.Y(n_6183)
);

INVx2_ASAP7_75t_L g6184 ( 
.A(n_6128),
.Y(n_6184)
);

NAND2xp5_ASAP7_75t_L g6185 ( 
.A(n_6144),
.B(n_139),
.Y(n_6185)
);

OAI22xp5_ASAP7_75t_L g6186 ( 
.A1(n_6145),
.A2(n_141),
.B1(n_139),
.B2(n_140),
.Y(n_6186)
);

NAND2xp5_ASAP7_75t_L g6187 ( 
.A(n_6152),
.B(n_140),
.Y(n_6187)
);

XOR2xp5_ASAP7_75t_L g6188 ( 
.A(n_6105),
.B(n_140),
.Y(n_6188)
);

NOR3xp33_ASAP7_75t_L g6189 ( 
.A(n_6151),
.B(n_140),
.C(n_141),
.Y(n_6189)
);

NOR2x1_ASAP7_75t_L g6190 ( 
.A(n_6133),
.B(n_141),
.Y(n_6190)
);

AND2x2_ASAP7_75t_L g6191 ( 
.A(n_6112),
.B(n_141),
.Y(n_6191)
);

NAND2xp5_ASAP7_75t_L g6192 ( 
.A(n_6126),
.B(n_142),
.Y(n_6192)
);

NOR3xp33_ASAP7_75t_L g6193 ( 
.A(n_6121),
.B(n_142),
.C(n_143),
.Y(n_6193)
);

INVxp67_ASAP7_75t_SL g6194 ( 
.A(n_6116),
.Y(n_6194)
);

NAND4xp25_ASAP7_75t_SL g6195 ( 
.A(n_6140),
.B(n_6149),
.C(n_6150),
.D(n_6143),
.Y(n_6195)
);

OR2x2_ASAP7_75t_L g6196 ( 
.A(n_6117),
.B(n_142),
.Y(n_6196)
);

INVx2_ASAP7_75t_L g6197 ( 
.A(n_6130),
.Y(n_6197)
);

INVx1_ASAP7_75t_L g6198 ( 
.A(n_6124),
.Y(n_6198)
);

NAND2xp5_ASAP7_75t_L g6199 ( 
.A(n_6142),
.B(n_142),
.Y(n_6199)
);

OAI21xp5_ASAP7_75t_L g6200 ( 
.A1(n_6113),
.A2(n_143),
.B(n_144),
.Y(n_6200)
);

OAI22xp5_ASAP7_75t_L g6201 ( 
.A1(n_6111),
.A2(n_145),
.B1(n_143),
.B2(n_144),
.Y(n_6201)
);

NAND2xp5_ASAP7_75t_L g6202 ( 
.A(n_6122),
.B(n_143),
.Y(n_6202)
);

OAI22xp5_ASAP7_75t_SL g6203 ( 
.A1(n_6153),
.A2(n_146),
.B1(n_144),
.B2(n_145),
.Y(n_6203)
);

NOR2x1_ASAP7_75t_L g6204 ( 
.A(n_6098),
.B(n_145),
.Y(n_6204)
);

INVx1_ASAP7_75t_L g6205 ( 
.A(n_6124),
.Y(n_6205)
);

INVx1_ASAP7_75t_L g6206 ( 
.A(n_6106),
.Y(n_6206)
);

AOI221x1_ASAP7_75t_L g6207 ( 
.A1(n_6127),
.A2(n_147),
.B1(n_145),
.B2(n_146),
.C(n_148),
.Y(n_6207)
);

AO22x1_ASAP7_75t_L g6208 ( 
.A1(n_6131),
.A2(n_148),
.B1(n_146),
.B2(n_147),
.Y(n_6208)
);

AND2x4_ASAP7_75t_L g6209 ( 
.A(n_6129),
.B(n_146),
.Y(n_6209)
);

INVx1_ASAP7_75t_L g6210 ( 
.A(n_6115),
.Y(n_6210)
);

OAI221xp5_ASAP7_75t_L g6211 ( 
.A1(n_6181),
.A2(n_6118),
.B1(n_6125),
.B2(n_6110),
.C(n_6114),
.Y(n_6211)
);

AOI211x1_ASAP7_75t_L g6212 ( 
.A1(n_6167),
.A2(n_6134),
.B(n_6123),
.C(n_6097),
.Y(n_6212)
);

NAND4xp25_ASAP7_75t_L g6213 ( 
.A(n_6189),
.B(n_6156),
.C(n_149),
.D(n_147),
.Y(n_6213)
);

AOI221xp5_ASAP7_75t_L g6214 ( 
.A1(n_6175),
.A2(n_149),
.B1(n_147),
.B2(n_148),
.C(n_150),
.Y(n_6214)
);

NAND2xp5_ASAP7_75t_SL g6215 ( 
.A(n_6184),
.B(n_149),
.Y(n_6215)
);

AOI211xp5_ASAP7_75t_L g6216 ( 
.A1(n_6183),
.A2(n_151),
.B(n_149),
.C(n_150),
.Y(n_6216)
);

AOI21xp5_ASAP7_75t_L g6217 ( 
.A1(n_6179),
.A2(n_150),
.B(n_151),
.Y(n_6217)
);

AOI221xp5_ASAP7_75t_L g6218 ( 
.A1(n_6159),
.A2(n_152),
.B1(n_150),
.B2(n_151),
.C(n_153),
.Y(n_6218)
);

INVx1_ASAP7_75t_L g6219 ( 
.A(n_6198),
.Y(n_6219)
);

AOI221xp5_ASAP7_75t_L g6220 ( 
.A1(n_6177),
.A2(n_153),
.B1(n_151),
.B2(n_152),
.C(n_154),
.Y(n_6220)
);

AOI221xp5_ASAP7_75t_L g6221 ( 
.A1(n_6170),
.A2(n_6165),
.B1(n_6205),
.B2(n_6186),
.C(n_6197),
.Y(n_6221)
);

AOI211xp5_ASAP7_75t_SL g6222 ( 
.A1(n_6192),
.A2(n_154),
.B(n_152),
.C(n_153),
.Y(n_6222)
);

OAI21xp33_ASAP7_75t_L g6223 ( 
.A1(n_6171),
.A2(n_152),
.B(n_154),
.Y(n_6223)
);

AOI221x1_ASAP7_75t_L g6224 ( 
.A1(n_6193),
.A2(n_6202),
.B1(n_6166),
.B2(n_6163),
.C(n_6168),
.Y(n_6224)
);

NOR3xp33_ASAP7_75t_L g6225 ( 
.A(n_6173),
.B(n_154),
.C(n_155),
.Y(n_6225)
);

AOI21xp5_ASAP7_75t_L g6226 ( 
.A1(n_6164),
.A2(n_6188),
.B(n_6174),
.Y(n_6226)
);

NOR3xp33_ASAP7_75t_L g6227 ( 
.A(n_6201),
.B(n_6203),
.C(n_6208),
.Y(n_6227)
);

INVx1_ASAP7_75t_L g6228 ( 
.A(n_6191),
.Y(n_6228)
);

OAI22xp5_ASAP7_75t_L g6229 ( 
.A1(n_6172),
.A2(n_6176),
.B1(n_6161),
.B2(n_6185),
.Y(n_6229)
);

INVx1_ASAP7_75t_L g6230 ( 
.A(n_6196),
.Y(n_6230)
);

AOI21xp5_ASAP7_75t_L g6231 ( 
.A1(n_6199),
.A2(n_155),
.B(n_156),
.Y(n_6231)
);

INVx1_ASAP7_75t_L g6232 ( 
.A(n_6209),
.Y(n_6232)
);

NAND4xp25_ASAP7_75t_SL g6233 ( 
.A(n_6169),
.B(n_157),
.C(n_155),
.D(n_156),
.Y(n_6233)
);

NOR2xp33_ASAP7_75t_L g6234 ( 
.A(n_6160),
.B(n_6187),
.Y(n_6234)
);

NOR3xp33_ASAP7_75t_L g6235 ( 
.A(n_6195),
.B(n_155),
.C(n_156),
.Y(n_6235)
);

OAI21xp5_ASAP7_75t_L g6236 ( 
.A1(n_6204),
.A2(n_157),
.B(n_158),
.Y(n_6236)
);

AOI21xp5_ASAP7_75t_L g6237 ( 
.A1(n_6200),
.A2(n_158),
.B(n_159),
.Y(n_6237)
);

OAI22xp5_ASAP7_75t_L g6238 ( 
.A1(n_6182),
.A2(n_160),
.B1(n_158),
.B2(n_159),
.Y(n_6238)
);

OAI211xp5_ASAP7_75t_L g6239 ( 
.A1(n_6180),
.A2(n_161),
.B(n_159),
.C(n_160),
.Y(n_6239)
);

OAI21xp5_ASAP7_75t_L g6240 ( 
.A1(n_6190),
.A2(n_159),
.B(n_160),
.Y(n_6240)
);

INVx1_ASAP7_75t_L g6241 ( 
.A(n_6209),
.Y(n_6241)
);

OAI221xp5_ASAP7_75t_SL g6242 ( 
.A1(n_6178),
.A2(n_163),
.B1(n_161),
.B2(n_162),
.C(n_164),
.Y(n_6242)
);

CKINVDCx20_ASAP7_75t_L g6243 ( 
.A(n_6158),
.Y(n_6243)
);

AOI221xp5_ASAP7_75t_L g6244 ( 
.A1(n_6194),
.A2(n_163),
.B1(n_161),
.B2(n_162),
.C(n_164),
.Y(n_6244)
);

OAI311xp33_ASAP7_75t_L g6245 ( 
.A1(n_6210),
.A2(n_163),
.A3(n_161),
.B1(n_162),
.C1(n_164),
.Y(n_6245)
);

AOI222xp33_ASAP7_75t_L g6246 ( 
.A1(n_6206),
.A2(n_162),
.B1(n_163),
.B2(n_164),
.C1(n_165),
.C2(n_166),
.Y(n_6246)
);

AOI22xp5_ASAP7_75t_L g6247 ( 
.A1(n_6157),
.A2(n_6162),
.B1(n_6207),
.B2(n_167),
.Y(n_6247)
);

NAND2xp5_ASAP7_75t_L g6248 ( 
.A(n_6179),
.B(n_165),
.Y(n_6248)
);

NOR2xp33_ASAP7_75t_L g6249 ( 
.A(n_6175),
.B(n_165),
.Y(n_6249)
);

XNOR2x1_ASAP7_75t_L g6250 ( 
.A(n_6160),
.B(n_166),
.Y(n_6250)
);

NAND3xp33_ASAP7_75t_SL g6251 ( 
.A(n_6159),
.B(n_166),
.C(n_167),
.Y(n_6251)
);

AOI211xp5_ASAP7_75t_L g6252 ( 
.A1(n_6189),
.A2(n_168),
.B(n_166),
.C(n_167),
.Y(n_6252)
);

AOI321xp33_ASAP7_75t_L g6253 ( 
.A1(n_6194),
.A2(n_167),
.A3(n_168),
.B1(n_169),
.B2(n_170),
.C(n_171),
.Y(n_6253)
);

INVx1_ASAP7_75t_L g6254 ( 
.A(n_6179),
.Y(n_6254)
);

OAI21xp5_ASAP7_75t_L g6255 ( 
.A1(n_6175),
.A2(n_168),
.B(n_169),
.Y(n_6255)
);

OAI21xp5_ASAP7_75t_SL g6256 ( 
.A1(n_6181),
.A2(n_168),
.B(n_169),
.Y(n_6256)
);

NOR2xp33_ASAP7_75t_L g6257 ( 
.A(n_6175),
.B(n_170),
.Y(n_6257)
);

AOI221xp5_ASAP7_75t_L g6258 ( 
.A1(n_6175),
.A2(n_170),
.B1(n_171),
.B2(n_172),
.C(n_173),
.Y(n_6258)
);

NAND2xp5_ASAP7_75t_L g6259 ( 
.A(n_6179),
.B(n_171),
.Y(n_6259)
);

NAND2xp5_ASAP7_75t_L g6260 ( 
.A(n_6179),
.B(n_171),
.Y(n_6260)
);

AOI22xp5_ASAP7_75t_L g6261 ( 
.A1(n_6158),
.A2(n_174),
.B1(n_172),
.B2(n_173),
.Y(n_6261)
);

AOI321xp33_ASAP7_75t_L g6262 ( 
.A1(n_6194),
.A2(n_172),
.A3(n_173),
.B1(n_174),
.B2(n_175),
.C(n_176),
.Y(n_6262)
);

NOR2xp33_ASAP7_75t_SL g6263 ( 
.A(n_6232),
.B(n_173),
.Y(n_6263)
);

OR2x2_ASAP7_75t_L g6264 ( 
.A(n_6219),
.B(n_6254),
.Y(n_6264)
);

AOI22xp5_ASAP7_75t_L g6265 ( 
.A1(n_6243),
.A2(n_176),
.B1(n_174),
.B2(n_175),
.Y(n_6265)
);

INVx1_ASAP7_75t_L g6266 ( 
.A(n_6248),
.Y(n_6266)
);

AOI322xp5_ASAP7_75t_L g6267 ( 
.A1(n_6235),
.A2(n_174),
.A3(n_175),
.B1(n_176),
.B2(n_177),
.C1(n_178),
.C2(n_179),
.Y(n_6267)
);

AND2x2_ASAP7_75t_L g6268 ( 
.A(n_6225),
.B(n_177),
.Y(n_6268)
);

AOI322xp5_ASAP7_75t_L g6269 ( 
.A1(n_6221),
.A2(n_6234),
.A3(n_6241),
.B1(n_6227),
.B2(n_6228),
.C1(n_6251),
.C2(n_6230),
.Y(n_6269)
);

AOI222xp33_ASAP7_75t_L g6270 ( 
.A1(n_6220),
.A2(n_177),
.B1(n_178),
.B2(n_179),
.C1(n_180),
.C2(n_181),
.Y(n_6270)
);

O2A1O1Ixp33_ASAP7_75t_SL g6271 ( 
.A1(n_6259),
.A2(n_180),
.B(n_178),
.C(n_179),
.Y(n_6271)
);

AOI221xp5_ASAP7_75t_L g6272 ( 
.A1(n_6217),
.A2(n_178),
.B1(n_179),
.B2(n_180),
.C(n_181),
.Y(n_6272)
);

AOI21xp33_ASAP7_75t_SL g6273 ( 
.A1(n_6250),
.A2(n_181),
.B(n_182),
.Y(n_6273)
);

AOI221xp5_ASAP7_75t_L g6274 ( 
.A1(n_6249),
.A2(n_181),
.B1(n_182),
.B2(n_183),
.C(n_184),
.Y(n_6274)
);

INVx1_ASAP7_75t_L g6275 ( 
.A(n_6260),
.Y(n_6275)
);

INVxp67_ASAP7_75t_SL g6276 ( 
.A(n_6215),
.Y(n_6276)
);

INVx2_ASAP7_75t_L g6277 ( 
.A(n_6212),
.Y(n_6277)
);

OAI22xp5_ASAP7_75t_L g6278 ( 
.A1(n_6261),
.A2(n_184),
.B1(n_182),
.B2(n_183),
.Y(n_6278)
);

INVx1_ASAP7_75t_L g6279 ( 
.A(n_6255),
.Y(n_6279)
);

XNOR2x1_ASAP7_75t_L g6280 ( 
.A(n_6238),
.B(n_182),
.Y(n_6280)
);

AOI22xp33_ASAP7_75t_L g6281 ( 
.A1(n_6213),
.A2(n_6257),
.B1(n_6233),
.B2(n_6223),
.Y(n_6281)
);

O2A1O1Ixp33_ASAP7_75t_L g6282 ( 
.A1(n_6245),
.A2(n_185),
.B(n_183),
.C(n_184),
.Y(n_6282)
);

OAI321xp33_ASAP7_75t_L g6283 ( 
.A1(n_6229),
.A2(n_185),
.A3(n_186),
.B1(n_187),
.B2(n_188),
.C(n_189),
.Y(n_6283)
);

OAI21xp33_ASAP7_75t_L g6284 ( 
.A1(n_6256),
.A2(n_185),
.B(n_187),
.Y(n_6284)
);

NAND2xp5_ASAP7_75t_L g6285 ( 
.A(n_6222),
.B(n_187),
.Y(n_6285)
);

INVx1_ASAP7_75t_SL g6286 ( 
.A(n_6237),
.Y(n_6286)
);

OAI21x1_ASAP7_75t_SL g6287 ( 
.A1(n_6226),
.A2(n_188),
.B(n_189),
.Y(n_6287)
);

INVx1_ASAP7_75t_L g6288 ( 
.A(n_6247),
.Y(n_6288)
);

NOR2xp33_ASAP7_75t_L g6289 ( 
.A(n_6211),
.B(n_188),
.Y(n_6289)
);

AOI21xp5_ASAP7_75t_L g6290 ( 
.A1(n_6231),
.A2(n_188),
.B(n_189),
.Y(n_6290)
);

AOI321xp33_ASAP7_75t_L g6291 ( 
.A1(n_6252),
.A2(n_189),
.A3(n_190),
.B1(n_191),
.B2(n_192),
.C(n_193),
.Y(n_6291)
);

INVx1_ASAP7_75t_L g6292 ( 
.A(n_6236),
.Y(n_6292)
);

OAI22xp5_ASAP7_75t_L g6293 ( 
.A1(n_6242),
.A2(n_192),
.B1(n_190),
.B2(n_191),
.Y(n_6293)
);

AOI22xp5_ASAP7_75t_L g6294 ( 
.A1(n_6218),
.A2(n_192),
.B1(n_190),
.B2(n_191),
.Y(n_6294)
);

AND2x2_ASAP7_75t_L g6295 ( 
.A(n_6216),
.B(n_190),
.Y(n_6295)
);

INVxp67_ASAP7_75t_L g6296 ( 
.A(n_6246),
.Y(n_6296)
);

OAI21xp33_ASAP7_75t_L g6297 ( 
.A1(n_6214),
.A2(n_193),
.B(n_194),
.Y(n_6297)
);

INVx1_ASAP7_75t_L g6298 ( 
.A(n_6262),
.Y(n_6298)
);

AOI22xp5_ASAP7_75t_L g6299 ( 
.A1(n_6239),
.A2(n_195),
.B1(n_193),
.B2(n_194),
.Y(n_6299)
);

AOI22xp5_ASAP7_75t_L g6300 ( 
.A1(n_6258),
.A2(n_196),
.B1(n_194),
.B2(n_195),
.Y(n_6300)
);

NOR3xp33_ASAP7_75t_L g6301 ( 
.A(n_6244),
.B(n_194),
.C(n_195),
.Y(n_6301)
);

OAI21xp33_ASAP7_75t_SL g6302 ( 
.A1(n_6240),
.A2(n_195),
.B(n_196),
.Y(n_6302)
);

OAI21xp5_ASAP7_75t_L g6303 ( 
.A1(n_6224),
.A2(n_196),
.B(n_197),
.Y(n_6303)
);

NAND2xp5_ASAP7_75t_L g6304 ( 
.A(n_6253),
.B(n_197),
.Y(n_6304)
);

AOI221xp5_ASAP7_75t_L g6305 ( 
.A1(n_6219),
.A2(n_197),
.B1(n_198),
.B2(n_199),
.C(n_200),
.Y(n_6305)
);

NAND2xp5_ASAP7_75t_SL g6306 ( 
.A(n_6220),
.B(n_197),
.Y(n_6306)
);

NOR2x1_ASAP7_75t_L g6307 ( 
.A(n_6219),
.B(n_198),
.Y(n_6307)
);

OAI21xp5_ASAP7_75t_L g6308 ( 
.A1(n_6217),
.A2(n_198),
.B(n_199),
.Y(n_6308)
);

INVx1_ASAP7_75t_L g6309 ( 
.A(n_6264),
.Y(n_6309)
);

AOI22xp5_ASAP7_75t_L g6310 ( 
.A1(n_6289),
.A2(n_201),
.B1(n_199),
.B2(n_200),
.Y(n_6310)
);

AND4x1_ASAP7_75t_L g6311 ( 
.A(n_6263),
.B(n_202),
.C(n_200),
.D(n_201),
.Y(n_6311)
);

AOI221xp5_ASAP7_75t_L g6312 ( 
.A1(n_6293),
.A2(n_200),
.B1(n_201),
.B2(n_202),
.C(n_203),
.Y(n_6312)
);

AND2x2_ASAP7_75t_L g6313 ( 
.A(n_6268),
.B(n_201),
.Y(n_6313)
);

A2O1A1Ixp33_ASAP7_75t_L g6314 ( 
.A1(n_6282),
.A2(n_204),
.B(n_202),
.C(n_203),
.Y(n_6314)
);

INVx1_ASAP7_75t_L g6315 ( 
.A(n_6285),
.Y(n_6315)
);

NOR3xp33_ASAP7_75t_SL g6316 ( 
.A(n_6306),
.B(n_203),
.C(n_204),
.Y(n_6316)
);

NAND2xp5_ASAP7_75t_L g6317 ( 
.A(n_6267),
.B(n_203),
.Y(n_6317)
);

INVx2_ASAP7_75t_L g6318 ( 
.A(n_6287),
.Y(n_6318)
);

OAI211xp5_ASAP7_75t_L g6319 ( 
.A1(n_6269),
.A2(n_206),
.B(n_204),
.C(n_205),
.Y(n_6319)
);

OAI31xp33_ASAP7_75t_L g6320 ( 
.A1(n_6284),
.A2(n_206),
.A3(n_204),
.B(n_205),
.Y(n_6320)
);

OAI22xp5_ASAP7_75t_L g6321 ( 
.A1(n_6281),
.A2(n_207),
.B1(n_205),
.B2(n_206),
.Y(n_6321)
);

AOI22xp33_ASAP7_75t_L g6322 ( 
.A1(n_6298),
.A2(n_208),
.B1(n_206),
.B2(n_207),
.Y(n_6322)
);

AOI21xp33_ASAP7_75t_L g6323 ( 
.A1(n_6270),
.A2(n_6304),
.B(n_6296),
.Y(n_6323)
);

AOI221xp5_ASAP7_75t_L g6324 ( 
.A1(n_6283),
.A2(n_207),
.B1(n_208),
.B2(n_209),
.C(n_210),
.Y(n_6324)
);

OAI211xp5_ASAP7_75t_L g6325 ( 
.A1(n_6274),
.A2(n_209),
.B(n_207),
.C(n_208),
.Y(n_6325)
);

AOI21xp5_ASAP7_75t_L g6326 ( 
.A1(n_6271),
.A2(n_208),
.B(n_209),
.Y(n_6326)
);

NOR2x1_ASAP7_75t_L g6327 ( 
.A(n_6303),
.B(n_209),
.Y(n_6327)
);

BUFx2_ASAP7_75t_L g6328 ( 
.A(n_6302),
.Y(n_6328)
);

NOR3xp33_ASAP7_75t_L g6329 ( 
.A(n_6305),
.B(n_210),
.C(n_211),
.Y(n_6329)
);

OAI211xp5_ASAP7_75t_SL g6330 ( 
.A1(n_6297),
.A2(n_6294),
.B(n_6300),
.C(n_6286),
.Y(n_6330)
);

OAI22xp5_ASAP7_75t_L g6331 ( 
.A1(n_6277),
.A2(n_212),
.B1(n_210),
.B2(n_211),
.Y(n_6331)
);

AOI321xp33_ASAP7_75t_L g6332 ( 
.A1(n_6276),
.A2(n_211),
.A3(n_212),
.B1(n_213),
.B2(n_214),
.C(n_215),
.Y(n_6332)
);

NAND2xp5_ASAP7_75t_L g6333 ( 
.A(n_6299),
.B(n_211),
.Y(n_6333)
);

AOI221xp5_ASAP7_75t_L g6334 ( 
.A1(n_6273),
.A2(n_212),
.B1(n_213),
.B2(n_214),
.C(n_215),
.Y(n_6334)
);

AOI211x1_ASAP7_75t_L g6335 ( 
.A1(n_6308),
.A2(n_214),
.B(n_212),
.C(n_213),
.Y(n_6335)
);

NAND2xp5_ASAP7_75t_L g6336 ( 
.A(n_6295),
.B(n_213),
.Y(n_6336)
);

XOR2x2_ASAP7_75t_L g6337 ( 
.A(n_6280),
.B(n_215),
.Y(n_6337)
);

BUFx2_ASAP7_75t_L g6338 ( 
.A(n_6307),
.Y(n_6338)
);

NAND2xp5_ASAP7_75t_L g6339 ( 
.A(n_6272),
.B(n_216),
.Y(n_6339)
);

INVxp67_ASAP7_75t_L g6340 ( 
.A(n_6288),
.Y(n_6340)
);

OAI21xp5_ASAP7_75t_SL g6341 ( 
.A1(n_6265),
.A2(n_216),
.B(n_217),
.Y(n_6341)
);

OAI22xp33_ASAP7_75t_L g6342 ( 
.A1(n_6279),
.A2(n_6275),
.B1(n_6266),
.B2(n_6292),
.Y(n_6342)
);

AOI221xp5_ASAP7_75t_L g6343 ( 
.A1(n_6278),
.A2(n_216),
.B1(n_217),
.B2(n_218),
.C(n_219),
.Y(n_6343)
);

XNOR2xp5_ASAP7_75t_L g6344 ( 
.A(n_6290),
.B(n_217),
.Y(n_6344)
);

OAI21xp5_ASAP7_75t_L g6345 ( 
.A1(n_6301),
.A2(n_218),
.B(n_219),
.Y(n_6345)
);

INVx2_ASAP7_75t_SL g6346 ( 
.A(n_6291),
.Y(n_6346)
);

OAI21xp33_ASAP7_75t_L g6347 ( 
.A1(n_6289),
.A2(n_218),
.B(n_220),
.Y(n_6347)
);

A2O1A1Ixp33_ASAP7_75t_L g6348 ( 
.A1(n_6289),
.A2(n_222),
.B(n_220),
.C(n_221),
.Y(n_6348)
);

OAI21xp33_ASAP7_75t_L g6349 ( 
.A1(n_6289),
.A2(n_220),
.B(n_221),
.Y(n_6349)
);

OAI211xp5_ASAP7_75t_SL g6350 ( 
.A1(n_6269),
.A2(n_222),
.B(n_220),
.C(n_221),
.Y(n_6350)
);

AOI321xp33_ASAP7_75t_L g6351 ( 
.A1(n_6329),
.A2(n_222),
.A3(n_223),
.B1(n_224),
.B2(n_225),
.C(n_226),
.Y(n_6351)
);

NOR2x1_ASAP7_75t_L g6352 ( 
.A(n_6319),
.B(n_223),
.Y(n_6352)
);

XOR2x2_ASAP7_75t_L g6353 ( 
.A(n_6344),
.B(n_223),
.Y(n_6353)
);

NAND4xp25_ASAP7_75t_L g6354 ( 
.A(n_6323),
.B(n_225),
.C(n_223),
.D(n_224),
.Y(n_6354)
);

NOR2x1_ASAP7_75t_SL g6355 ( 
.A(n_6318),
.B(n_224),
.Y(n_6355)
);

INVxp67_ASAP7_75t_L g6356 ( 
.A(n_6327),
.Y(n_6356)
);

INVx2_ASAP7_75t_SL g6357 ( 
.A(n_6309),
.Y(n_6357)
);

INVx1_ASAP7_75t_L g6358 ( 
.A(n_6336),
.Y(n_6358)
);

OAI211xp5_ASAP7_75t_L g6359 ( 
.A1(n_6322),
.A2(n_6332),
.B(n_6312),
.C(n_6314),
.Y(n_6359)
);

O2A1O1Ixp5_ASAP7_75t_SL g6360 ( 
.A1(n_6340),
.A2(n_226),
.B(n_224),
.C(n_225),
.Y(n_6360)
);

XNOR2x2_ASAP7_75t_L g6361 ( 
.A(n_6337),
.B(n_225),
.Y(n_6361)
);

XNOR2xp5_ASAP7_75t_L g6362 ( 
.A(n_6311),
.B(n_226),
.Y(n_6362)
);

AO22x2_ASAP7_75t_L g6363 ( 
.A1(n_6346),
.A2(n_228),
.B1(n_226),
.B2(n_227),
.Y(n_6363)
);

BUFx8_ASAP7_75t_SL g6364 ( 
.A(n_6328),
.Y(n_6364)
);

INVx1_ASAP7_75t_L g6365 ( 
.A(n_6333),
.Y(n_6365)
);

AOI221xp5_ASAP7_75t_L g6366 ( 
.A1(n_6321),
.A2(n_227),
.B1(n_228),
.B2(n_229),
.C(n_230),
.Y(n_6366)
);

BUFx4f_ASAP7_75t_SL g6367 ( 
.A(n_6315),
.Y(n_6367)
);

INVxp33_ASAP7_75t_SL g6368 ( 
.A(n_6331),
.Y(n_6368)
);

O2A1O1Ixp33_ASAP7_75t_L g6369 ( 
.A1(n_6348),
.A2(n_229),
.B(n_227),
.C(n_228),
.Y(n_6369)
);

INVx1_ASAP7_75t_L g6370 ( 
.A(n_6313),
.Y(n_6370)
);

INVxp67_ASAP7_75t_L g6371 ( 
.A(n_6326),
.Y(n_6371)
);

OAI22xp5_ASAP7_75t_L g6372 ( 
.A1(n_6310),
.A2(n_230),
.B1(n_228),
.B2(n_229),
.Y(n_6372)
);

AOI221xp5_ASAP7_75t_SL g6373 ( 
.A1(n_6347),
.A2(n_229),
.B1(n_230),
.B2(n_231),
.C(n_232),
.Y(n_6373)
);

AOI22xp5_ASAP7_75t_L g6374 ( 
.A1(n_6350),
.A2(n_6349),
.B1(n_6330),
.B2(n_6317),
.Y(n_6374)
);

AOI211xp5_ASAP7_75t_L g6375 ( 
.A1(n_6342),
.A2(n_233),
.B(n_231),
.C(n_232),
.Y(n_6375)
);

AND2x2_ASAP7_75t_L g6376 ( 
.A(n_6316),
.B(n_231),
.Y(n_6376)
);

XNOR2xp5_ASAP7_75t_L g6377 ( 
.A(n_6335),
.B(n_231),
.Y(n_6377)
);

OAI22xp5_ASAP7_75t_L g6378 ( 
.A1(n_6339),
.A2(n_234),
.B1(n_232),
.B2(n_233),
.Y(n_6378)
);

INVxp67_ASAP7_75t_SL g6379 ( 
.A(n_6345),
.Y(n_6379)
);

NAND5xp2_ASAP7_75t_L g6380 ( 
.A(n_6324),
.B(n_232),
.C(n_233),
.D(n_234),
.E(n_235),
.Y(n_6380)
);

INVx1_ASAP7_75t_L g6381 ( 
.A(n_6363),
.Y(n_6381)
);

NOR2x1_ASAP7_75t_L g6382 ( 
.A(n_6354),
.B(n_6338),
.Y(n_6382)
);

NOR2x1_ASAP7_75t_L g6383 ( 
.A(n_6352),
.B(n_6359),
.Y(n_6383)
);

AOI22xp5_ASAP7_75t_L g6384 ( 
.A1(n_6376),
.A2(n_6325),
.B1(n_6341),
.B2(n_6334),
.Y(n_6384)
);

AND2x4_ASAP7_75t_L g6385 ( 
.A(n_6357),
.B(n_6320),
.Y(n_6385)
);

INVx1_ASAP7_75t_L g6386 ( 
.A(n_6363),
.Y(n_6386)
);

NOR2x1_ASAP7_75t_L g6387 ( 
.A(n_6378),
.B(n_6343),
.Y(n_6387)
);

NOR2xp67_ASAP7_75t_SL g6388 ( 
.A(n_6365),
.B(n_6358),
.Y(n_6388)
);

INVx1_ASAP7_75t_L g6389 ( 
.A(n_6355),
.Y(n_6389)
);

AND2x2_ASAP7_75t_L g6390 ( 
.A(n_6370),
.B(n_233),
.Y(n_6390)
);

INVx1_ASAP7_75t_L g6391 ( 
.A(n_6362),
.Y(n_6391)
);

INVx1_ASAP7_75t_L g6392 ( 
.A(n_6364),
.Y(n_6392)
);

HB1xp67_ASAP7_75t_L g6393 ( 
.A(n_6371),
.Y(n_6393)
);

OAI22xp5_ASAP7_75t_SL g6394 ( 
.A1(n_6377),
.A2(n_234),
.B1(n_235),
.B2(n_236),
.Y(n_6394)
);

INVx1_ASAP7_75t_L g6395 ( 
.A(n_6361),
.Y(n_6395)
);

INVx1_ASAP7_75t_L g6396 ( 
.A(n_6369),
.Y(n_6396)
);

NOR2xp33_ASAP7_75t_L g6397 ( 
.A(n_6368),
.B(n_234),
.Y(n_6397)
);

NOR2x1_ASAP7_75t_L g6398 ( 
.A(n_6380),
.B(n_235),
.Y(n_6398)
);

NAND2xp5_ASAP7_75t_L g6399 ( 
.A(n_6375),
.B(n_235),
.Y(n_6399)
);

NOR2x1_ASAP7_75t_L g6400 ( 
.A(n_6372),
.B(n_237),
.Y(n_6400)
);

INVx1_ASAP7_75t_L g6401 ( 
.A(n_6374),
.Y(n_6401)
);

INVx1_ASAP7_75t_L g6402 ( 
.A(n_6351),
.Y(n_6402)
);

AOI22xp33_ASAP7_75t_L g6403 ( 
.A1(n_6367),
.A2(n_237),
.B1(n_238),
.B2(n_239),
.Y(n_6403)
);

AOI22xp5_ASAP7_75t_L g6404 ( 
.A1(n_6379),
.A2(n_238),
.B1(n_239),
.B2(n_240),
.Y(n_6404)
);

INVx2_ASAP7_75t_L g6405 ( 
.A(n_6356),
.Y(n_6405)
);

AND3x4_ASAP7_75t_L g6406 ( 
.A(n_6353),
.B(n_238),
.C(n_239),
.Y(n_6406)
);

INVx1_ASAP7_75t_L g6407 ( 
.A(n_6366),
.Y(n_6407)
);

AOI22xp5_ASAP7_75t_L g6408 ( 
.A1(n_6373),
.A2(n_6360),
.B1(n_240),
.B2(n_241),
.Y(n_6408)
);

NOR2xp33_ASAP7_75t_L g6409 ( 
.A(n_6354),
.B(n_238),
.Y(n_6409)
);

INVx1_ASAP7_75t_L g6410 ( 
.A(n_6389),
.Y(n_6410)
);

AO22x2_ASAP7_75t_L g6411 ( 
.A1(n_6406),
.A2(n_240),
.B1(n_241),
.B2(n_242),
.Y(n_6411)
);

AND2x4_ASAP7_75t_L g6412 ( 
.A(n_6392),
.B(n_241),
.Y(n_6412)
);

INVxp33_ASAP7_75t_L g6413 ( 
.A(n_6397),
.Y(n_6413)
);

INVx1_ASAP7_75t_L g6414 ( 
.A(n_6390),
.Y(n_6414)
);

INVx2_ASAP7_75t_L g6415 ( 
.A(n_6385),
.Y(n_6415)
);

OR2x2_ASAP7_75t_L g6416 ( 
.A(n_6399),
.B(n_242),
.Y(n_6416)
);

OR2x2_ASAP7_75t_L g6417 ( 
.A(n_6402),
.B(n_6395),
.Y(n_6417)
);

AND3x4_ASAP7_75t_L g6418 ( 
.A(n_6398),
.B(n_243),
.C(n_244),
.Y(n_6418)
);

AOI22x1_ASAP7_75t_SL g6419 ( 
.A1(n_6401),
.A2(n_243),
.B1(n_244),
.B2(n_245),
.Y(n_6419)
);

NOR3xp33_ASAP7_75t_L g6420 ( 
.A(n_6394),
.B(n_244),
.C(n_245),
.Y(n_6420)
);

OR2x2_ASAP7_75t_L g6421 ( 
.A(n_6381),
.B(n_245),
.Y(n_6421)
);

NAND4xp75_ASAP7_75t_L g6422 ( 
.A(n_6383),
.B(n_6382),
.C(n_6387),
.D(n_6400),
.Y(n_6422)
);

INVx1_ASAP7_75t_L g6423 ( 
.A(n_6404),
.Y(n_6423)
);

NAND5xp2_ASAP7_75t_L g6424 ( 
.A(n_6384),
.B(n_245),
.C(n_246),
.D(n_247),
.E(n_248),
.Y(n_6424)
);

AND2x4_ASAP7_75t_L g6425 ( 
.A(n_6405),
.B(n_246),
.Y(n_6425)
);

INVx1_ASAP7_75t_L g6426 ( 
.A(n_6408),
.Y(n_6426)
);

INVx1_ASAP7_75t_L g6427 ( 
.A(n_6386),
.Y(n_6427)
);

INVx1_ASAP7_75t_L g6428 ( 
.A(n_6385),
.Y(n_6428)
);

NAND4xp75_ASAP7_75t_L g6429 ( 
.A(n_6409),
.B(n_246),
.C(n_247),
.D(n_248),
.Y(n_6429)
);

HB1xp67_ASAP7_75t_L g6430 ( 
.A(n_6393),
.Y(n_6430)
);

INVxp33_ASAP7_75t_L g6431 ( 
.A(n_6388),
.Y(n_6431)
);

OAI211xp5_ASAP7_75t_L g6432 ( 
.A1(n_6410),
.A2(n_6403),
.B(n_6396),
.C(n_6407),
.Y(n_6432)
);

A2O1A1Ixp33_ASAP7_75t_L g6433 ( 
.A1(n_6431),
.A2(n_6391),
.B(n_247),
.C(n_248),
.Y(n_6433)
);

AOI222xp33_ASAP7_75t_L g6434 ( 
.A1(n_6428),
.A2(n_246),
.B1(n_247),
.B2(n_248),
.C1(n_249),
.C2(n_250),
.Y(n_6434)
);

AOI22xp5_ASAP7_75t_L g6435 ( 
.A1(n_6415),
.A2(n_249),
.B1(n_250),
.B2(n_251),
.Y(n_6435)
);

INVx1_ASAP7_75t_L g6436 ( 
.A(n_6419),
.Y(n_6436)
);

AOI21xp5_ASAP7_75t_L g6437 ( 
.A1(n_6417),
.A2(n_249),
.B(n_250),
.Y(n_6437)
);

OAI22xp5_ASAP7_75t_SL g6438 ( 
.A1(n_6418),
.A2(n_6426),
.B1(n_6414),
.B2(n_6427),
.Y(n_6438)
);

AOI22xp5_ASAP7_75t_SL g6439 ( 
.A1(n_6412),
.A2(n_249),
.B1(n_251),
.B2(n_252),
.Y(n_6439)
);

NAND2xp5_ASAP7_75t_L g6440 ( 
.A(n_6425),
.B(n_251),
.Y(n_6440)
);

OAI221xp5_ASAP7_75t_L g6441 ( 
.A1(n_6420),
.A2(n_252),
.B1(n_253),
.B2(n_254),
.C(n_255),
.Y(n_6441)
);

OAI22xp5_ASAP7_75t_L g6442 ( 
.A1(n_6421),
.A2(n_6430),
.B1(n_6416),
.B2(n_6423),
.Y(n_6442)
);

NAND2xp5_ASAP7_75t_SL g6443 ( 
.A(n_6413),
.B(n_252),
.Y(n_6443)
);

AOI22x1_ASAP7_75t_L g6444 ( 
.A1(n_6411),
.A2(n_252),
.B1(n_253),
.B2(n_254),
.Y(n_6444)
);

AOI22xp5_ASAP7_75t_L g6445 ( 
.A1(n_6422),
.A2(n_253),
.B1(n_254),
.B2(n_255),
.Y(n_6445)
);

NAND2xp5_ASAP7_75t_SL g6446 ( 
.A(n_6429),
.B(n_253),
.Y(n_6446)
);

INVx1_ASAP7_75t_SL g6447 ( 
.A(n_6440),
.Y(n_6447)
);

AND3x4_ASAP7_75t_L g6448 ( 
.A(n_6432),
.B(n_6424),
.C(n_6411),
.Y(n_6448)
);

INVx1_ASAP7_75t_L g6449 ( 
.A(n_6445),
.Y(n_6449)
);

AND3x2_ASAP7_75t_L g6450 ( 
.A(n_6436),
.B(n_254),
.C(n_255),
.Y(n_6450)
);

AND3x4_ASAP7_75t_L g6451 ( 
.A(n_6438),
.B(n_255),
.C(n_256),
.Y(n_6451)
);

INVx3_ASAP7_75t_L g6452 ( 
.A(n_6439),
.Y(n_6452)
);

NOR2x1_ASAP7_75t_L g6453 ( 
.A(n_6433),
.B(n_256),
.Y(n_6453)
);

INVx1_ASAP7_75t_L g6454 ( 
.A(n_6435),
.Y(n_6454)
);

AND3x4_ASAP7_75t_L g6455 ( 
.A(n_6434),
.B(n_256),
.C(n_257),
.Y(n_6455)
);

AND2x4_ASAP7_75t_L g6456 ( 
.A(n_6443),
.B(n_256),
.Y(n_6456)
);

XNOR2xp5_ASAP7_75t_L g6457 ( 
.A(n_6442),
.B(n_257),
.Y(n_6457)
);

BUFx2_ASAP7_75t_L g6458 ( 
.A(n_6450),
.Y(n_6458)
);

INVx2_ASAP7_75t_L g6459 ( 
.A(n_6456),
.Y(n_6459)
);

INVx1_ASAP7_75t_L g6460 ( 
.A(n_6457),
.Y(n_6460)
);

INVx2_ASAP7_75t_L g6461 ( 
.A(n_6452),
.Y(n_6461)
);

INVx2_ASAP7_75t_L g6462 ( 
.A(n_6449),
.Y(n_6462)
);

INVx1_ASAP7_75t_L g6463 ( 
.A(n_6451),
.Y(n_6463)
);

OAI22x1_ASAP7_75t_L g6464 ( 
.A1(n_6462),
.A2(n_6448),
.B1(n_6461),
.B2(n_6444),
.Y(n_6464)
);

AOI22xp33_ASAP7_75t_L g6465 ( 
.A1(n_6458),
.A2(n_6454),
.B1(n_6441),
.B2(n_6447),
.Y(n_6465)
);

XNOR2xp5_ASAP7_75t_L g6466 ( 
.A(n_6464),
.B(n_6455),
.Y(n_6466)
);

INVx2_ASAP7_75t_L g6467 ( 
.A(n_6465),
.Y(n_6467)
);

HB1xp67_ASAP7_75t_L g6468 ( 
.A(n_6467),
.Y(n_6468)
);

AND2x4_ASAP7_75t_L g6469 ( 
.A(n_6466),
.B(n_6460),
.Y(n_6469)
);

NAND2xp5_ASAP7_75t_L g6470 ( 
.A(n_6468),
.B(n_6463),
.Y(n_6470)
);

AOI22xp33_ASAP7_75t_L g6471 ( 
.A1(n_6470),
.A2(n_6469),
.B1(n_6459),
.B2(n_6453),
.Y(n_6471)
);

OAI21x1_ASAP7_75t_L g6472 ( 
.A1(n_6471),
.A2(n_6437),
.B(n_6446),
.Y(n_6472)
);

AOI22xp5_ASAP7_75t_L g6473 ( 
.A1(n_6472),
.A2(n_257),
.B1(n_258),
.B2(n_259),
.Y(n_6473)
);

AOI22xp33_ASAP7_75t_L g6474 ( 
.A1(n_6472),
.A2(n_257),
.B1(n_258),
.B2(n_259),
.Y(n_6474)
);

OR2x6_ASAP7_75t_L g6475 ( 
.A(n_6473),
.B(n_1061),
.Y(n_6475)
);

NAND2xp5_ASAP7_75t_L g6476 ( 
.A(n_6474),
.B(n_258),
.Y(n_6476)
);

AOI21xp5_ASAP7_75t_L g6477 ( 
.A1(n_6476),
.A2(n_259),
.B(n_260),
.Y(n_6477)
);

AOI211xp5_ASAP7_75t_L g6478 ( 
.A1(n_6477),
.A2(n_6475),
.B(n_261),
.C(n_262),
.Y(n_6478)
);


endmodule