module fake_netlist_1_9531_n_17 (n_1, n_2, n_6, n_4, n_3, n_5, n_0, n_17);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_0;
output n_17;
wire n_11;
wire n_13;
wire n_16;
wire n_12;
wire n_9;
wire n_14;
wire n_10;
wire n_15;
wire n_7;
wire n_8;
NAND2xp5_ASAP7_75t_SL g7 ( .A(n_4), .B(n_5), .Y(n_7) );
NAND2xp5_ASAP7_75t_L g8 ( .A(n_1), .B(n_6), .Y(n_8) );
INVx1_ASAP7_75t_L g9 ( .A(n_0), .Y(n_9) );
INVx2_ASAP7_75t_L g10 ( .A(n_2), .Y(n_10) );
BUFx6f_ASAP7_75t_L g11 ( .A(n_3), .Y(n_11) );
OAI21x1_ASAP7_75t_L g12 ( .A1(n_10), .A2(n_8), .B(n_7), .Y(n_12) );
INVxp67_ASAP7_75t_L g13 ( .A(n_9), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_13), .Y(n_14) );
NAND4xp25_ASAP7_75t_L g15 ( .A(n_14), .B(n_0), .C(n_12), .D(n_11), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_15), .Y(n_16) );
NAND2xp5_ASAP7_75t_L g17 ( .A(n_16), .B(n_11), .Y(n_17) );
endmodule