module fake_jpeg_20528_n_163 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_163);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_163;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_93;
wire n_91;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_10),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_31),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_38),
.Y(n_51)
);

BUFx10_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_33),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_22),
.Y(n_55)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_9),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_6),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_36),
.Y(n_60)
);

INVx2_ASAP7_75t_R g61 ( 
.A(n_29),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_24),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_4),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_17),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_23),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_16),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_6),
.Y(n_69)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_3),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_40),
.B(n_44),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_20),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_1),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_75),
.Y(n_87)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_76),
.Y(n_85)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_70),
.B(n_0),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_79),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_59),
.B(n_61),
.C(n_53),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_81),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_0),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_74),
.Y(n_93)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_78),
.Y(n_84)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_81),
.Y(n_88)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_82),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_92),
.B(n_94),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_93),
.B(n_90),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_82),
.B(n_69),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_78),
.A2(n_61),
.B(n_68),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_95),
.A2(n_60),
.B1(n_71),
.B2(n_65),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_96),
.B(n_105),
.Y(n_120)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_97),
.A2(n_101),
.B1(n_73),
.B2(n_64),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_93),
.B(n_58),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_99),
.B(n_104),
.Y(n_121)
);

INVx2_ASAP7_75t_SL g100 ( 
.A(n_85),
.Y(n_100)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_100),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_89),
.A2(n_56),
.B1(n_52),
.B2(n_49),
.Y(n_101)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_83),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_91),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_88),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_107),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_108),
.A2(n_71),
.B1(n_67),
.B2(n_48),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_104),
.A2(n_87),
.B1(n_90),
.B2(n_52),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_109),
.A2(n_111),
.B1(n_116),
.B2(n_119),
.Y(n_126)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_106),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_115),
.Y(n_128)
);

AOI21xp33_ASAP7_75t_SL g113 ( 
.A1(n_96),
.A2(n_52),
.B(n_73),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_113),
.B(n_118),
.Y(n_125)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_97),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_102),
.A2(n_62),
.B1(n_72),
.B2(n_51),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_117),
.A2(n_50),
.B1(n_66),
.B2(n_55),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_108),
.B(n_98),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_101),
.A2(n_103),
.B1(n_100),
.B2(n_54),
.Y(n_119)
);

INVx2_ASAP7_75t_SL g143 ( 
.A(n_122),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_117),
.A2(n_59),
.B1(n_70),
.B2(n_3),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_123),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_112),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_124),
.B(n_127),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_118),
.B(n_1),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_114),
.Y(n_129)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_129),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_120),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_130),
.B(n_131),
.Y(n_136)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_121),
.Y(n_131)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_109),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_132),
.B(n_133),
.Y(n_141)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_112),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_125),
.B(n_19),
.C(n_46),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_135),
.B(n_15),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g137 ( 
.A(n_126),
.B(n_2),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_137),
.A2(n_139),
.B(n_140),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_128),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_122),
.B(n_2),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_132),
.B(n_4),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_142),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_138),
.A2(n_123),
.B(n_26),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_145),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_136),
.A2(n_25),
.B(n_45),
.Y(n_147)
);

NOR2xp67_ASAP7_75t_L g152 ( 
.A(n_147),
.B(n_148),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_SL g148 ( 
.A(n_135),
.B(n_5),
.Y(n_148)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_152),
.Y(n_153)
);

NOR3xp33_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_134),
.C(n_150),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_146),
.Y(n_155)
);

OR2x2_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_141),
.Y(n_156)
);

AOI322xp5_ASAP7_75t_L g157 ( 
.A1(n_156),
.A2(n_151),
.A3(n_144),
.B1(n_137),
.B2(n_143),
.C1(n_149),
.C2(n_5),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_157),
.A2(n_143),
.B1(n_27),
.B2(n_28),
.Y(n_158)
);

A2O1A1Ixp33_ASAP7_75t_L g159 ( 
.A1(n_158),
.A2(n_14),
.B(n_43),
.C(n_35),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_159),
.A2(n_11),
.B(n_34),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_160),
.A2(n_13),
.B1(n_32),
.B2(n_47),
.Y(n_161)
);

MAJx2_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_7),
.C(n_8),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_7),
.Y(n_163)
);


endmodule