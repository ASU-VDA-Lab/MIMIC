module fake_jpeg_23296_n_265 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_265);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_265;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_139;
wire n_45;
wire n_61;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_155;
wire n_118;
wire n_258;
wire n_96;

BUFx5_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

INVx11_ASAP7_75t_SL g21 ( 
.A(n_15),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_2),
.B(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_18),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_47),
.Y(n_53)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx3_ASAP7_75t_SL g86 ( 
.A(n_42),
.Y(n_86)
);

BUFx4f_ASAP7_75t_SL g43 ( 
.A(n_25),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx3_ASAP7_75t_SL g45 ( 
.A(n_26),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_45),
.A2(n_19),
.B1(n_34),
.B2(n_17),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_29),
.B(n_1),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_46),
.B(n_29),
.Y(n_58)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

INVx2_ASAP7_75t_R g49 ( 
.A(n_43),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_49),
.B(n_58),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_50),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_L g51 ( 
.A1(n_39),
.A2(n_45),
.B1(n_34),
.B2(n_43),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_51),
.A2(n_82),
.B1(n_41),
.B2(n_38),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_22),
.Y(n_54)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_27),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_55),
.B(n_84),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_40),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_57),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_62),
.A2(n_72),
.B1(n_33),
.B2(n_23),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_22),
.Y(n_63)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

A2O1A1Ixp33_ASAP7_75t_L g64 ( 
.A1(n_43),
.A2(n_27),
.B(n_20),
.C(n_32),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_64),
.B(n_1),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_65),
.Y(n_109)
);

CKINVDCx12_ASAP7_75t_R g66 ( 
.A(n_48),
.Y(n_66)
);

INVx6_ASAP7_75t_SL g95 ( 
.A(n_66),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_67),
.Y(n_116)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_68),
.B(n_71),
.Y(n_89)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_69),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_31),
.Y(n_70)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_70),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_37),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_45),
.A2(n_19),
.B1(n_21),
.B2(n_17),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_42),
.A2(n_19),
.B1(n_36),
.B2(n_18),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_75),
.A2(n_81),
.B1(n_23),
.B2(n_33),
.Y(n_101)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_39),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_76),
.B(n_77),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_41),
.B(n_31),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_39),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_78),
.B(n_83),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_80),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_47),
.A2(n_36),
.B1(n_20),
.B2(n_32),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_47),
.A2(n_36),
.B1(n_27),
.B2(n_24),
.Y(n_82)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_41),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_45),
.B(n_27),
.C(n_44),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_38),
.B(n_1),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_35),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_93),
.A2(n_107),
.B1(n_65),
.B2(n_5),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_101),
.A2(n_104),
.B1(n_117),
.B2(n_86),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_51),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_53),
.B(n_24),
.Y(n_103)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_103),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_64),
.B(n_74),
.Y(n_106)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_106),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_85),
.A2(n_35),
.B1(n_30),
.B2(n_28),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_74),
.B(n_16),
.Y(n_108)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_108),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_49),
.B(n_14),
.Y(n_110)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_110),
.Y(n_146)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_65),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_113),
.B(n_60),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_114),
.B(n_115),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_60),
.B(n_26),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_84),
.A2(n_35),
.B1(n_30),
.B2(n_44),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_100),
.B(n_59),
.C(n_68),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_119),
.B(n_124),
.C(n_89),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_109),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_120),
.B(n_123),
.Y(n_154)
);

FAx1_ASAP7_75t_SL g121 ( 
.A(n_100),
.B(n_55),
.CI(n_82),
.CON(n_121),
.SN(n_121)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_121),
.B(n_127),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_122),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_94),
.A2(n_86),
.B1(n_69),
.B2(n_83),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_85),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_125),
.A2(n_132),
.B1(n_99),
.B2(n_111),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_90),
.B(n_56),
.Y(n_126)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_126),
.Y(n_159)
);

A2O1A1Ixp33_ASAP7_75t_L g127 ( 
.A1(n_106),
.A2(n_55),
.B(n_56),
.C(n_50),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_133),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_93),
.A2(n_76),
.B1(n_73),
.B2(n_78),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_130),
.A2(n_131),
.B1(n_138),
.B2(n_110),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_104),
.A2(n_73),
.B1(n_59),
.B2(n_52),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_101),
.A2(n_52),
.B1(n_80),
.B2(n_79),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_105),
.B(n_4),
.Y(n_133)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_96),
.Y(n_134)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_134),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_105),
.B(n_67),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_135),
.B(n_136),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_91),
.B(n_67),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_114),
.B(n_30),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_137),
.B(n_141),
.Y(n_150)
);

INVx1_ASAP7_75t_SL g139 ( 
.A(n_109),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_139),
.B(n_142),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_94),
.B(n_87),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_92),
.B(n_61),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_91),
.B(n_4),
.Y(n_143)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_143),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_90),
.B(n_5),
.Y(n_144)
);

INVxp33_ASAP7_75t_L g163 ( 
.A(n_144),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_88),
.B(n_6),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_147),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_117),
.B(n_97),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_148),
.B(n_95),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_140),
.A2(n_92),
.B(n_115),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_149),
.A2(n_151),
.B(n_165),
.Y(n_187)
);

OA21x2_ASAP7_75t_L g151 ( 
.A1(n_130),
.A2(n_98),
.B(n_97),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_152),
.A2(n_171),
.B1(n_145),
.B2(n_134),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_155),
.A2(n_158),
.B1(n_162),
.B2(n_174),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_124),
.B(n_89),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_156),
.B(n_160),
.C(n_175),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_140),
.A2(n_98),
.B1(n_111),
.B2(n_99),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_131),
.A2(n_112),
.B1(n_108),
.B2(n_116),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_127),
.A2(n_103),
.B(n_112),
.Y(n_165)
);

AO22x1_ASAP7_75t_L g167 ( 
.A1(n_125),
.A2(n_61),
.B1(n_116),
.B2(n_96),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_167),
.A2(n_7),
.B(n_8),
.Y(n_194)
);

INVx13_ASAP7_75t_L g168 ( 
.A(n_139),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_168),
.B(n_7),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_170),
.B(n_176),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_132),
.A2(n_113),
.B1(n_88),
.B2(n_8),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_119),
.A2(n_121),
.B1(n_129),
.B2(n_148),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_142),
.B(n_95),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_121),
.B(n_6),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_158),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_177),
.B(n_180),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_175),
.B(n_150),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_178),
.A2(n_194),
.B(n_195),
.Y(n_199)
);

AOI322xp5_ASAP7_75t_L g179 ( 
.A1(n_161),
.A2(n_129),
.A3(n_118),
.B1(n_137),
.B2(n_146),
.C1(n_128),
.C2(n_141),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_179),
.B(n_174),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_169),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_173),
.B(n_128),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_181),
.B(n_166),
.Y(n_200)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_150),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_182),
.B(n_184),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_156),
.B(n_145),
.Y(n_183)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_183),
.Y(n_214)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_162),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_159),
.B(n_146),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_185),
.B(n_189),
.Y(n_205)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_152),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_171),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_190),
.B(n_192),
.Y(n_198)
);

CKINVDCx14_ASAP7_75t_R g203 ( 
.A(n_191),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_170),
.B(n_120),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_157),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_193),
.B(n_197),
.Y(n_207)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_167),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_200),
.B(n_193),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_201),
.B(n_188),
.C(n_209),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_187),
.A2(n_149),
.B(n_153),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_202),
.A2(n_213),
.B(n_194),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_187),
.A2(n_154),
.B(n_151),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_204),
.A2(n_208),
.B(n_9),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_197),
.A2(n_165),
.B(n_151),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_189),
.A2(n_155),
.B1(n_167),
.B2(n_160),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_209),
.A2(n_184),
.B1(n_190),
.B2(n_183),
.Y(n_224)
);

OA21x2_ASAP7_75t_SL g210 ( 
.A1(n_178),
.A2(n_176),
.B(n_163),
.Y(n_210)
);

MAJx2_ASAP7_75t_L g216 ( 
.A(n_210),
.B(n_178),
.C(n_196),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_188),
.A2(n_172),
.B1(n_164),
.B2(n_168),
.Y(n_211)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_211),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_192),
.A2(n_163),
.B(n_10),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_216),
.B(n_217),
.Y(n_238)
);

MAJx2_ASAP7_75t_L g217 ( 
.A(n_210),
.B(n_196),
.C(n_186),
.Y(n_217)
);

XNOR2x1_ASAP7_75t_L g218 ( 
.A(n_204),
.B(n_186),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_218),
.B(n_205),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_219),
.A2(n_227),
.B(n_228),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_207),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_220),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_207),
.B(n_182),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_221),
.B(n_222),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_223),
.B(n_201),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_224),
.A2(n_211),
.B1(n_206),
.B2(n_199),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_214),
.B(n_180),
.C(n_191),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_225),
.B(n_226),
.C(n_213),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_214),
.B(n_13),
.C(n_10),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_212),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_215),
.A2(n_203),
.B1(n_198),
.B2(n_212),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_230),
.A2(n_234),
.B1(n_9),
.B2(n_10),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_228),
.A2(n_208),
.B(n_199),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_232),
.B(n_233),
.Y(n_244)
);

XOR2x2_ASAP7_75t_L g234 ( 
.A(n_218),
.B(n_198),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_235),
.A2(n_215),
.B1(n_221),
.B2(n_205),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_236),
.B(n_237),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_225),
.B(n_202),
.C(n_206),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_239),
.B(n_200),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_241),
.A2(n_242),
.B1(n_243),
.B2(n_230),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_229),
.A2(n_224),
.B1(n_219),
.B2(n_223),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_237),
.A2(n_216),
.B1(n_217),
.B2(n_226),
.Y(n_243)
);

INVxp33_ASAP7_75t_L g245 ( 
.A(n_240),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_245),
.B(n_239),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_246),
.B(n_247),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_244),
.A2(n_231),
.B(n_234),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_249),
.B(n_251),
.C(n_238),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_245),
.B(n_233),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_250),
.B(n_254),
.Y(n_258)
);

AO21x2_ASAP7_75t_L g255 ( 
.A1(n_253),
.A2(n_241),
.B(n_242),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_248),
.B(n_243),
.Y(n_254)
);

O2A1O1Ixp33_ASAP7_75t_L g261 ( 
.A1(n_255),
.A2(n_256),
.B(n_9),
.C(n_11),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_253),
.A2(n_238),
.B(n_248),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_257),
.A2(n_252),
.B1(n_236),
.B2(n_12),
.Y(n_259)
);

BUFx24_ASAP7_75t_SL g263 ( 
.A(n_259),
.Y(n_263)
);

NOR3xp33_ASAP7_75t_L g260 ( 
.A(n_255),
.B(n_252),
.C(n_11),
.Y(n_260)
);

A2O1A1Ixp33_ASAP7_75t_L g262 ( 
.A1(n_260),
.A2(n_261),
.B(n_11),
.C(n_12),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_262),
.B(n_258),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_264),
.B(n_263),
.Y(n_265)
);


endmodule