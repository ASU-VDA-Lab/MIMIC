module fake_jpeg_30250_n_95 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_95);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_95;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

BUFx12_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_23),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

BUFx16f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_39),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_29),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_40),
.B(n_43),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx3_ASAP7_75t_SL g48 ( 
.A(n_41),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_28),
.B(n_1),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_51),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_36),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_56),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_43),
.Y(n_51)
);

AND2x6_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_32),
.Y(n_52)
);

NOR2xp67_ASAP7_75t_L g63 ( 
.A(n_52),
.B(n_1),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_39),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_57),
.B(n_58),
.Y(n_69)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_61),
.Y(n_73)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_63),
.A2(n_64),
.B(n_65),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_53),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

OA22x2_ASAP7_75t_L g78 ( 
.A1(n_66),
.A2(n_67),
.B1(n_68),
.B2(n_33),
.Y(n_78)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_62),
.A2(n_18),
.B(n_27),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_70),
.A2(n_76),
.B(n_8),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_SL g71 ( 
.A(n_59),
.B(n_62),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_71),
.B(n_75),
.C(n_77),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_63),
.A2(n_31),
.B1(n_3),
.B2(n_4),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_74),
.B(n_78),
.Y(n_84)
);

MAJx2_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_35),
.C(n_33),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_65),
.A2(n_19),
.B(n_25),
.Y(n_76)
);

XNOR2x1_ASAP7_75t_L g77 ( 
.A(n_59),
.B(n_35),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_78),
.A2(n_31),
.B1(n_4),
.B2(n_2),
.Y(n_79)
);

AO21x2_ASAP7_75t_L g87 ( 
.A1(n_79),
.A2(n_70),
.B(n_12),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_72),
.A2(n_2),
.B(n_7),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_80),
.B(n_82),
.Y(n_85)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_83),
.B(n_9),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_86),
.B(n_87),
.C(n_84),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_88),
.A2(n_89),
.B(n_87),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_85),
.B(n_81),
.C(n_69),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_90),
.B(n_10),
.C(n_13),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_91),
.B(n_14),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_92),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_93),
.A2(n_16),
.B(n_17),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_20),
.Y(n_95)
);


endmodule