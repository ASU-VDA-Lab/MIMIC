module fake_jpeg_16025_n_43 (n_3, n_2, n_1, n_0, n_4, n_5, n_43);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_43;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx3_ASAP7_75t_L g6 ( 
.A(n_5),
.Y(n_6)
);

INVx1_ASAP7_75t_L g7 ( 
.A(n_0),
.Y(n_7)
);

NOR2xp33_ASAP7_75t_L g8 ( 
.A(n_1),
.B(n_3),
.Y(n_8)
);

INVx4_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

INVx4_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_14),
.B(n_12),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_8),
.B(n_0),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_15),
.B(n_18),
.Y(n_24)
);

INVxp33_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_16),
.B(n_20),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_9),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_17)
);

XOR2xp5_ASAP7_75t_L g25 ( 
.A(n_17),
.B(n_18),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_13),
.B(n_2),
.Y(n_18)
);

AOI22xp33_ASAP7_75t_SL g19 ( 
.A1(n_9),
.A2(n_2),
.B1(n_3),
.B2(n_11),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_19),
.A2(n_21),
.B(n_6),
.Y(n_23)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

OAI21xp33_ASAP7_75t_L g21 ( 
.A1(n_11),
.A2(n_10),
.B(n_12),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_22),
.B(n_26),
.Y(n_30)
);

XNOR2x1_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_25),
.Y(n_34)
);

XNOR2xp5_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_23),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_15),
.B(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_17),
.B(n_15),
.Y(n_29)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

FAx1_ASAP7_75t_SL g36 ( 
.A(n_31),
.B(n_34),
.CI(n_24),
.CON(n_36),
.SN(n_36)
);

BUFx4f_ASAP7_75t_SL g35 ( 
.A(n_27),
.Y(n_35)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

OAI21x1_ASAP7_75t_L g39 ( 
.A1(n_36),
.A2(n_38),
.B(n_30),
.Y(n_39)
);

AO22x1_ASAP7_75t_L g38 ( 
.A1(n_34),
.A2(n_27),
.B1(n_33),
.B2(n_35),
.Y(n_38)
);

HB1xp67_ASAP7_75t_L g41 ( 
.A(n_39),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_38),
.A2(n_36),
.B1(n_32),
.B2(n_37),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_41),
.B(n_38),
.Y(n_42)
);

MAJx2_ASAP7_75t_L g43 ( 
.A(n_42),
.B(n_40),
.C(n_36),
.Y(n_43)
);


endmodule