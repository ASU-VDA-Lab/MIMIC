module fake_jpeg_458_n_62 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_62);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_62;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_47;
wire n_22;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx1_ASAP7_75t_L g7 ( 
.A(n_1),
.Y(n_7)
);

AND2x2_ASAP7_75t_L g8 ( 
.A(n_2),
.B(n_4),
.Y(n_8)
);

BUFx10_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

BUFx10_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_16),
.B(n_19),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_8),
.B(n_0),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_17),
.B(n_8),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_18),
.B(n_20),
.Y(n_21)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_8),
.B(n_3),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_23),
.B(n_24),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_17),
.B(n_14),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_20),
.B(n_12),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_26),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_16),
.Y(n_26)
);

INVx2_ASAP7_75t_SL g27 ( 
.A(n_22),
.Y(n_27)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

NAND2x1_ASAP7_75t_SL g28 ( 
.A(n_22),
.B(n_19),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_28),
.B(n_29),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_21),
.A2(n_16),
.B1(n_13),
.B2(n_7),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_21),
.A2(n_15),
.B1(n_10),
.B2(n_12),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_33),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_22),
.A2(n_15),
.B1(n_10),
.B2(n_9),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

OAI21xp33_ASAP7_75t_L g33 ( 
.A1(n_21),
.A2(n_0),
.B(n_2),
.Y(n_33)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_22),
.B(n_18),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_18),
.C(n_9),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_32),
.B(n_5),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_37),
.B(n_38),
.Y(n_47)
);

XOR2xp5_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_18),
.Y(n_38)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g45 ( 
.A1(n_42),
.A2(n_27),
.B(n_35),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_38),
.C(n_40),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_39),
.Y(n_46)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_43),
.A2(n_27),
.B1(n_29),
.B2(n_30),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_49),
.A2(n_41),
.B1(n_34),
.B2(n_36),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_48),
.C(n_45),
.Y(n_55)
);

OAI22x1_ASAP7_75t_L g52 ( 
.A1(n_49),
.A2(n_43),
.B1(n_44),
.B2(n_42),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_52),
.B(n_53),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_55),
.B(n_47),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g58 ( 
.A(n_56),
.B(n_57),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_54),
.B(n_50),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g59 ( 
.A1(n_58),
.A2(n_52),
.B(n_36),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_59),
.B(n_39),
.C(n_11),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_60),
.B(n_6),
.Y(n_61)
);

XOR2xp5_ASAP7_75t_L g62 ( 
.A(n_61),
.B(n_6),
.Y(n_62)
);


endmodule