module real_jpeg_26162_n_29 (n_17, n_8, n_0, n_21, n_2, n_132, n_139, n_10, n_137, n_9, n_12, n_135, n_24, n_134, n_6, n_136, n_28, n_133, n_23, n_11, n_14, n_131, n_138, n_25, n_7, n_22, n_18, n_3, n_5, n_4, n_1, n_26, n_27, n_20, n_19, n_140, n_16, n_15, n_13, n_29);

input n_17;
input n_8;
input n_0;
input n_21;
input n_2;
input n_132;
input n_139;
input n_10;
input n_137;
input n_9;
input n_12;
input n_135;
input n_24;
input n_134;
input n_6;
input n_136;
input n_28;
input n_133;
input n_23;
input n_11;
input n_14;
input n_131;
input n_138;
input n_25;
input n_7;
input n_22;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_26;
input n_27;
input n_20;
input n_19;
input n_140;
input n_16;
input n_15;
input n_13;

output n_29;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_56;
wire n_48;
wire n_126;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_118;
wire n_123;
wire n_116;
wire n_50;
wire n_69;
wire n_31;
wire n_129;
wire n_72;
wire n_100;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_30;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

BUFx10_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

INVx6_ASAP7_75t_SL g57 ( 
.A(n_0),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_0),
.Y(n_60)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_1),
.Y(n_91)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_3),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_4),
.B(n_39),
.C(n_90),
.Y(n_38)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_5),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_6),
.B(n_47),
.C(n_58),
.Y(n_46)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_7),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_8),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_9),
.B(n_41),
.C(n_82),
.Y(n_40)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_10),
.Y(n_112)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_11),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_12),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_13),
.B(n_37),
.C(n_99),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_14),
.Y(n_118)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_15),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_16),
.Y(n_115)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_17),
.Y(n_104)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_18),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_19),
.B(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_20),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_21),
.B(n_45),
.C(n_65),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_35),
.C(n_110),
.Y(n_34)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_23),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_24),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_25),
.B(n_43),
.C(n_74),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_33),
.C(n_117),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_27),
.B(n_31),
.C(n_124),
.Y(n_30)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_27),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_27),
.A2(n_119),
.B1(n_127),
.B2(n_128),
.Y(n_126)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_28),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_126),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_119),
.C(n_120),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_112),
.C(n_113),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_101),
.C(n_102),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_93),
.C(n_94),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_85),
.C(n_86),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_77),
.C(n_78),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_68),
.C(n_69),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_61),
.C(n_62),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_52),
.C(n_53),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_51),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_64),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g73 ( 
.A(n_51),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

BUFx12_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_56),
.Y(n_54)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g67 ( 
.A(n_57),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_60),
.Y(n_58)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_67),
.Y(n_65)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_72),
.Y(n_70)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_73),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_76),
.Y(n_74)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_81),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_84),
.Y(n_82)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_89),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_89),
.B(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_111),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_92),
.Y(n_90)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_97),
.Y(n_95)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_105),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_105),
.B(n_129),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_106),
.B(n_118),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_125),
.Y(n_124)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_107),
.Y(n_116)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_116),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_116),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_123),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_131),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_132),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_133),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_134),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_135),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_136),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_137),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_138),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_139),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_140),
.Y(n_88)
);


endmodule