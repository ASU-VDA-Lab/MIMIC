module fake_jpeg_30728_n_422 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_422);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_422;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g22 ( 
.A(n_20),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_12),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_20),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

BUFx16f_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

BUFx10_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

BUFx4f_ASAP7_75t_SL g43 ( 
.A(n_12),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_11),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_1),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_2),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_51),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_52),
.Y(n_128)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_53),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_22),
.B(n_0),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_54),
.B(n_62),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_55),
.Y(n_107)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_56),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_57),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_58),
.Y(n_126)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_59),
.Y(n_100)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_60),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_61),
.Y(n_96)
);

INVx4_ASAP7_75t_SL g62 ( 
.A(n_49),
.Y(n_62)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_63),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_64),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_65),
.Y(n_106)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_66),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_26),
.B(n_0),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_67),
.B(n_72),
.Y(n_115)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_68),
.Y(n_92)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_69),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_70),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_71),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_26),
.B(n_0),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_24),
.Y(n_73)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_73),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_74),
.Y(n_117)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_24),
.Y(n_75)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_75),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

CKINVDCx6p67_ASAP7_75t_R g93 ( 
.A(n_76),
.Y(n_93)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_34),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_78),
.Y(n_120)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_79),
.B(n_80),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_38),
.B(n_1),
.Y(n_80)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_41),
.Y(n_81)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_81),
.Y(n_130)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_24),
.Y(n_82)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_82),
.Y(n_131)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_29),
.Y(n_83)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_83),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_39),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_84),
.Y(n_109)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_39),
.Y(n_85)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_39),
.Y(n_86)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_33),
.Y(n_87)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_87),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_42),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_89),
.Y(n_112)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_34),
.Y(n_89)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_43),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_90),
.B(n_32),
.Y(n_116)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_33),
.Y(n_91)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_91),
.Y(n_122)
);

INVx6_ASAP7_75t_SL g95 ( 
.A(n_55),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_95),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_80),
.A2(n_50),
.B1(n_47),
.B2(n_45),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_101),
.A2(n_104),
.B1(n_111),
.B2(n_32),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_54),
.A2(n_50),
.B1(n_47),
.B2(n_45),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_62),
.A2(n_32),
.B1(n_30),
.B2(n_50),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_116),
.B(n_81),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_76),
.B(n_44),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_124),
.B(n_132),
.Y(n_139)
);

A2O1A1Ixp33_ASAP7_75t_L g127 ( 
.A1(n_90),
.A2(n_48),
.B(n_31),
.C(n_35),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_127),
.B(n_1),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_56),
.B(n_44),
.Y(n_132)
);

BUFx10_ASAP7_75t_L g133 ( 
.A(n_66),
.Y(n_133)
);

INVx3_ASAP7_75t_SL g138 ( 
.A(n_133),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_89),
.B(n_38),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_135),
.B(n_32),
.Y(n_143)
);

HB1xp67_ASAP7_75t_L g140 ( 
.A(n_113),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_140),
.Y(n_195)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_125),
.Y(n_141)
);

INVx4_ASAP7_75t_SL g193 ( 
.A(n_141),
.Y(n_193)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_92),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_142),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_143),
.B(n_145),
.Y(n_173)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_110),
.Y(n_144)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_144),
.Y(n_190)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_122),
.Y(n_146)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_146),
.Y(n_177)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_100),
.Y(n_147)
);

INVx6_ASAP7_75t_L g180 ( 
.A(n_147),
.Y(n_180)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_136),
.Y(n_148)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_148),
.Y(n_178)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_130),
.Y(n_149)
);

INVx8_ASAP7_75t_L g182 ( 
.A(n_149),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_150),
.B(n_157),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_115),
.B(n_42),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_151),
.B(n_152),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_98),
.B(n_42),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_117),
.Y(n_153)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_153),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_106),
.Y(n_154)
);

INVx3_ASAP7_75t_SL g188 ( 
.A(n_154),
.Y(n_188)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_129),
.Y(n_155)
);

INVx8_ASAP7_75t_L g186 ( 
.A(n_155),
.Y(n_186)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_109),
.Y(n_156)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_156),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_112),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_102),
.A2(n_53),
.B1(n_60),
.B2(n_78),
.Y(n_158)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_158),
.Y(n_184)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_120),
.Y(n_159)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_159),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_98),
.A2(n_105),
.B1(n_71),
.B2(n_74),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_160),
.B(n_168),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_137),
.A2(n_27),
.B1(n_48),
.B2(n_40),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_161),
.Y(n_194)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_112),
.Y(n_162)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_162),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_105),
.A2(n_40),
.B(n_35),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_164),
.A2(n_169),
.B(n_116),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_124),
.B(n_31),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_165),
.Y(n_172)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_103),
.Y(n_166)
);

BUFx6f_ASAP7_75t_SL g175 ( 
.A(n_166),
.Y(n_175)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_100),
.Y(n_167)
);

BUFx12_ASAP7_75t_L g181 ( 
.A(n_167),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_106),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_114),
.A2(n_27),
.B1(n_59),
.B2(n_42),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_133),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_170),
.B(n_133),
.Y(n_187)
);

AOI21xp33_ASAP7_75t_L g174 ( 
.A1(n_171),
.A2(n_139),
.B(n_132),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_174),
.B(n_164),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_183),
.B(n_169),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_187),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_151),
.B(n_118),
.C(n_131),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_196),
.B(n_152),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_187),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_199),
.B(n_218),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_200),
.A2(n_217),
.B(n_195),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_201),
.B(n_198),
.Y(n_239)
);

OAI21xp33_ASAP7_75t_SL g202 ( 
.A1(n_185),
.A2(n_194),
.B(n_176),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_202),
.A2(n_213),
.B(n_185),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_203),
.B(n_216),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_172),
.B(n_139),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_204),
.B(n_205),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_176),
.B(n_143),
.Y(n_205)
);

A2O1A1Ixp33_ASAP7_75t_SL g206 ( 
.A1(n_183),
.A2(n_93),
.B(n_163),
.C(n_111),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_206),
.A2(n_208),
.B(n_180),
.Y(n_231)
);

NOR2x1_ASAP7_75t_L g207 ( 
.A(n_173),
.B(n_93),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_207),
.B(n_219),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_173),
.A2(n_138),
.B(n_167),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_177),
.Y(n_209)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_209),
.Y(n_222)
);

BUFx5_ASAP7_75t_L g210 ( 
.A(n_186),
.Y(n_210)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_210),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_173),
.B(n_146),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_211),
.B(n_220),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_192),
.A2(n_138),
.B(n_142),
.Y(n_213)
);

OAI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_194),
.A2(n_141),
.B1(n_147),
.B2(n_121),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g238 ( 
.A1(n_214),
.A2(n_193),
.B1(n_155),
.B2(n_107),
.Y(n_238)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_177),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_215),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_172),
.B(n_2),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_193),
.A2(n_184),
.B1(n_180),
.B2(n_186),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_189),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_175),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_196),
.B(n_144),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_221),
.A2(n_232),
.B(n_206),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_212),
.A2(n_184),
.B1(n_191),
.B2(n_188),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_227),
.A2(n_233),
.B1(n_242),
.B2(n_214),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_212),
.B(n_191),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_230),
.B(n_235),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_231),
.A2(n_234),
.B(n_179),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_206),
.A2(n_193),
.B1(n_188),
.B2(n_182),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_211),
.A2(n_178),
.B1(n_188),
.B2(n_97),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_205),
.B(n_178),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_220),
.B(n_197),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_236),
.B(n_237),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_201),
.B(n_197),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_238),
.A2(n_217),
.B1(n_219),
.B2(n_195),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_239),
.B(n_201),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_200),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_241),
.B(n_200),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_202),
.A2(n_97),
.B1(n_148),
.B2(n_198),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_SL g243 ( 
.A(n_234),
.B(n_206),
.C(n_203),
.Y(n_243)
);

NAND3xp33_ASAP7_75t_L g287 ( 
.A(n_243),
.B(n_253),
.C(n_262),
.Y(n_287)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_222),
.Y(n_244)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_244),
.Y(n_268)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_222),
.Y(n_245)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_245),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_246),
.B(n_237),
.Y(n_279)
);

AO22x1_ASAP7_75t_L g247 ( 
.A1(n_231),
.A2(n_207),
.B1(n_206),
.B2(n_200),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_247),
.B(n_248),
.Y(n_269)
);

XNOR2x2_ASAP7_75t_SL g248 ( 
.A(n_228),
.B(n_208),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_229),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_249),
.B(n_240),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_251),
.A2(n_223),
.B1(n_210),
.B2(n_238),
.Y(n_289)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_225),
.Y(n_252)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_252),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_226),
.B(n_204),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_254),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_231),
.A2(n_207),
.B(n_208),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_255),
.A2(n_258),
.B(n_263),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_240),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_256),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_257),
.A2(n_242),
.B1(n_227),
.B2(n_233),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_239),
.B(n_213),
.C(n_215),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_260),
.B(n_236),
.C(n_228),
.Y(n_282)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_225),
.Y(n_261)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_261),
.Y(n_277)
);

AOI32xp33_ASAP7_75t_L g262 ( 
.A1(n_229),
.A2(n_206),
.A3(n_209),
.B1(n_218),
.B2(n_216),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_221),
.A2(n_206),
.B(n_179),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_264),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_224),
.B(n_189),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_265),
.Y(n_275)
);

BUFx2_ASAP7_75t_L g266 ( 
.A(n_223),
.Y(n_266)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_266),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_224),
.B(n_190),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_267),
.Y(n_288)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_272),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_246),
.B(n_239),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_273),
.B(n_279),
.Y(n_295)
);

OAI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_249),
.A2(n_232),
.B1(n_230),
.B2(n_225),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_274),
.A2(n_264),
.B1(n_247),
.B2(n_252),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_282),
.B(n_285),
.C(n_263),
.Y(n_293)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_244),
.Y(n_283)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_283),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_250),
.B(n_235),
.Y(n_284)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_284),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_260),
.B(n_242),
.C(n_233),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_286),
.B(n_255),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_289),
.A2(n_257),
.B1(n_251),
.B2(n_261),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_259),
.B(n_226),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_290),
.B(n_259),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_278),
.B(n_253),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_292),
.B(n_302),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_293),
.B(n_310),
.C(n_282),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_294),
.A2(n_304),
.B1(n_307),
.B2(n_271),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_296),
.A2(n_65),
.B1(n_84),
.B2(n_86),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_272),
.B(n_250),
.Y(n_297)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_297),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_SL g298 ( 
.A(n_279),
.B(n_243),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_298),
.B(n_300),
.Y(n_319)
);

CKINVDCx14_ASAP7_75t_R g302 ( 
.A(n_287),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_290),
.B(n_245),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_303),
.B(n_309),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_291),
.A2(n_247),
.B1(n_258),
.B2(n_248),
.Y(n_304)
);

BUFx12_ASAP7_75t_L g305 ( 
.A(n_281),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_305),
.B(n_308),
.Y(n_329)
);

BUFx12_ASAP7_75t_L g308 ( 
.A(n_281),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_284),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_SL g310 ( 
.A(n_273),
.B(n_248),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_276),
.B(n_266),
.Y(n_311)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_311),
.Y(n_335)
);

BUFx2_ASAP7_75t_L g312 ( 
.A(n_280),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_312),
.B(n_317),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_291),
.A2(n_266),
.B(n_93),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g323 ( 
.A(n_313),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_269),
.A2(n_210),
.B(n_156),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g332 ( 
.A(n_314),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_269),
.A2(n_128),
.B(n_99),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_315),
.B(n_316),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_275),
.B(n_182),
.Y(n_316)
);

XOR2x1_ASAP7_75t_L g317 ( 
.A(n_271),
.B(n_175),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_318),
.A2(n_320),
.B1(n_325),
.B2(n_336),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_294),
.A2(n_276),
.B1(n_277),
.B2(n_288),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_321),
.B(n_308),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_301),
.A2(n_289),
.B1(n_285),
.B2(n_283),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_322),
.A2(n_313),
.B1(n_317),
.B2(n_299),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_293),
.B(n_277),
.C(n_270),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_324),
.B(n_326),
.C(n_330),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_304),
.A2(n_270),
.B1(n_268),
.B2(n_280),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_295),
.B(n_268),
.C(n_190),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_295),
.B(n_197),
.C(n_149),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_298),
.B(n_310),
.C(n_300),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_333),
.B(n_337),
.C(n_305),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_314),
.A2(n_168),
.B1(n_154),
.B2(n_107),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_296),
.B(n_315),
.C(n_306),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_338),
.A2(n_299),
.B1(n_153),
.B2(n_159),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_306),
.A2(n_123),
.B1(n_126),
.B2(n_166),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_340),
.B(n_126),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_341),
.A2(n_342),
.B1(n_343),
.B2(n_351),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_328),
.A2(n_312),
.B1(n_297),
.B2(n_311),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_326),
.B(n_308),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_346),
.B(n_348),
.Y(n_370)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_327),
.Y(n_347)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_347),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_324),
.B(n_3),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_349),
.B(n_353),
.C(n_354),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_334),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_350),
.B(n_352),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_321),
.B(n_305),
.C(n_181),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_330),
.B(n_181),
.C(n_134),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_335),
.Y(n_355)
);

HB1xp67_ASAP7_75t_L g371 ( 
.A(n_355),
.Y(n_371)
);

HB1xp67_ASAP7_75t_L g356 ( 
.A(n_339),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_356),
.A2(n_96),
.B1(n_119),
.B2(n_58),
.Y(n_369)
);

BUFx24_ASAP7_75t_SL g357 ( 
.A(n_331),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_357),
.A2(n_358),
.B1(n_325),
.B2(n_340),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_320),
.B(n_3),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_345),
.A2(n_332),
.B1(n_323),
.B2(n_337),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g374 ( 
.A(n_360),
.B(n_362),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_352),
.A2(n_318),
.B1(n_329),
.B2(n_333),
.Y(n_362)
);

OR2x2_ASAP7_75t_L g363 ( 
.A(n_342),
.B(n_339),
.Y(n_363)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_363),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_365),
.B(n_366),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_344),
.A2(n_336),
.B1(n_338),
.B2(n_319),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_344),
.B(n_319),
.C(n_181),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_367),
.B(n_368),
.C(n_353),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_349),
.B(n_181),
.C(n_123),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_369),
.B(n_354),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_373),
.B(n_381),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_375),
.B(n_377),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_361),
.A2(n_3),
.B1(n_5),
.B2(n_7),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_360),
.A2(n_108),
.B1(n_57),
.B2(n_11),
.Y(n_378)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_378),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_359),
.B(n_109),
.C(n_94),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_379),
.B(n_383),
.C(n_368),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_372),
.A2(n_5),
.B(n_8),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_380),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_SL g381 ( 
.A1(n_359),
.A2(n_8),
.B(n_11),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_363),
.B(n_13),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_SL g393 ( 
.A1(n_382),
.A2(n_379),
.B(n_383),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_367),
.B(n_94),
.C(n_43),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_385),
.B(n_389),
.Y(n_404)
);

AOI22xp33_ASAP7_75t_SL g388 ( 
.A1(n_376),
.A2(n_371),
.B1(n_364),
.B2(n_362),
.Y(n_388)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_388),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_L g389 ( 
.A1(n_374),
.A2(n_370),
.B1(n_14),
.B2(n_15),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_374),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_390),
.B(n_395),
.Y(n_405)
);

AOI22xp33_ASAP7_75t_L g391 ( 
.A1(n_373),
.A2(n_43),
.B1(n_14),
.B2(n_15),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_391),
.B(n_393),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_384),
.A2(n_13),
.B1(n_16),
.B2(n_17),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_392),
.A2(n_18),
.B1(n_19),
.B2(n_21),
.Y(n_400)
);

HB1xp67_ASAP7_75t_L g395 ( 
.A(n_375),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_L g397 ( 
.A1(n_386),
.A2(n_16),
.B(n_17),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_SL g410 ( 
.A1(n_397),
.A2(n_399),
.B(n_402),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_L g399 ( 
.A1(n_387),
.A2(n_16),
.B(n_18),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g407 ( 
.A1(n_400),
.A2(n_385),
.B1(n_392),
.B2(n_43),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_L g402 ( 
.A1(n_390),
.A2(n_18),
.B(n_19),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_SL g403 ( 
.A(n_394),
.B(n_21),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_403),
.B(n_37),
.Y(n_409)
);

MAJx2_ASAP7_75t_L g406 ( 
.A(n_401),
.B(n_388),
.C(n_396),
.Y(n_406)
);

AO21x1_ASAP7_75t_L g412 ( 
.A1(n_406),
.A2(n_411),
.B(n_410),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_407),
.B(n_409),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_404),
.B(n_405),
.C(n_398),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_408),
.B(n_28),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_SL g411 ( 
.A1(n_401),
.A2(n_42),
.B(n_28),
.Y(n_411)
);

OR2x2_ASAP7_75t_L g417 ( 
.A(n_412),
.B(n_28),
.Y(n_417)
);

AOI21xp5_ASAP7_75t_L g416 ( 
.A1(n_414),
.A2(n_415),
.B(n_413),
.Y(n_416)
);

INVxp67_ASAP7_75t_L g415 ( 
.A(n_408),
.Y(n_415)
);

HB1xp67_ASAP7_75t_L g418 ( 
.A(n_416),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_418),
.B(n_417),
.Y(n_419)
);

BUFx24_ASAP7_75t_SL g420 ( 
.A(n_419),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_420),
.A2(n_28),
.B1(n_37),
.B2(n_415),
.Y(n_421)
);

BUFx24_ASAP7_75t_SL g422 ( 
.A(n_421),
.Y(n_422)
);


endmodule