module fake_netlist_5_2108_n_781 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_781);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_781;

wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_194;
wire n_316;
wire n_389;
wire n_549;
wire n_684;
wire n_418;
wire n_248;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_235;
wire n_226;
wire n_605;
wire n_776;
wire n_667;
wire n_515;
wire n_353;
wire n_351;
wire n_367;
wire n_620;
wire n_643;
wire n_452;
wire n_397;
wire n_493;
wire n_525;
wire n_703;
wire n_698;
wire n_483;
wire n_544;
wire n_683;
wire n_780;
wire n_649;
wire n_552;
wire n_547;
wire n_721;
wire n_467;
wire n_564;
wire n_423;
wire n_284;
wire n_245;
wire n_501;
wire n_725;
wire n_280;
wire n_744;
wire n_590;
wire n_629;
wire n_672;
wire n_378;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_254;
wire n_690;
wire n_583;
wire n_671;
wire n_718;
wire n_302;
wire n_265;
wire n_526;
wire n_719;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_677;
wire n_173;
wire n_198;
wire n_714;
wire n_447;
wire n_247;
wire n_368;
wire n_314;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_625;
wire n_621;
wire n_753;
wire n_455;
wire n_674;
wire n_417;
wire n_612;
wire n_212;
wire n_385;
wire n_498;
wire n_516;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_252;
wire n_624;
wire n_295;
wire n_330;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_692;
wire n_755;
wire n_509;
wire n_568;
wire n_373;
wire n_757;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_556;
wire n_209;
wire n_259;
wire n_448;
wire n_758;
wire n_668;
wire n_733;
wire n_375;
wire n_301;
wire n_779;
wire n_576;
wire n_186;
wire n_537;
wire n_191;
wire n_587;
wire n_659;
wire n_492;
wire n_563;
wire n_171;
wire n_756;
wire n_524;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_741;
wire n_548;
wire n_543;
wire n_260;
wire n_298;
wire n_650;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_282;
wire n_752;
wire n_331;
wire n_406;
wire n_519;
wire n_470;
wire n_325;
wire n_449;
wire n_724;
wire n_546;
wire n_760;
wire n_658;
wire n_281;
wire n_240;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_323;
wire n_569;
wire n_769;
wire n_195;
wire n_356;
wire n_227;
wire n_592;
wire n_271;
wire n_335;
wire n_654;
wire n_370;
wire n_167;
wire n_234;
wire n_343;
wire n_428;
wire n_379;
wire n_308;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_297;
wire n_603;
wire n_225;
wire n_377;
wire n_751;
wire n_484;
wire n_775;
wire n_219;
wire n_442;
wire n_157;
wire n_192;
wire n_636;
wire n_600;
wire n_660;
wire n_223;
wire n_392;
wire n_158;
wire n_655;
wire n_704;
wire n_264;
wire n_669;
wire n_472;
wire n_742;
wire n_750;
wire n_454;
wire n_387;
wire n_771;
wire n_374;
wire n_163;
wire n_276;
wire n_339;
wire n_183;
wire n_185;
wire n_243;
wire n_398;
wire n_396;
wire n_635;
wire n_347;
wire n_763;
wire n_169;
wire n_522;
wire n_550;
wire n_255;
wire n_696;
wire n_215;
wire n_350;
wire n_196;
wire n_662;
wire n_459;
wire n_646;
wire n_211;
wire n_218;
wire n_400;
wire n_181;
wire n_436;
wire n_290;
wire n_580;
wire n_221;
wire n_178;
wire n_622;
wire n_723;
wire n_386;
wire n_578;
wire n_287;
wire n_344;
wire n_555;
wire n_473;
wire n_422;
wire n_475;
wire n_777;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_496;
wire n_355;
wire n_486;
wire n_670;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_521;
wire n_614;
wire n_663;
wire n_337;
wire n_430;
wire n_313;
wire n_631;
wire n_673;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_680;
wire n_168;
wire n_395;
wire n_164;
wire n_432;
wire n_553;
wire n_727;
wire n_311;
wire n_773;
wire n_208;
wire n_743;
wire n_214;
wire n_328;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_296;
wire n_613;
wire n_241;
wire n_637;
wire n_357;
wire n_598;
wire n_685;
wire n_608;
wire n_184;
wire n_446;
wire n_445;
wire n_749;
wire n_772;
wire n_691;
wire n_717;
wire n_165;
wire n_468;
wire n_499;
wire n_213;
wire n_342;
wire n_482;
wire n_517;
wire n_588;
wire n_361;
wire n_464;
wire n_363;
wire n_402;
wire n_413;
wire n_734;
wire n_638;
wire n_700;
wire n_197;
wire n_573;
wire n_236;
wire n_388;
wire n_761;
wire n_249;
wire n_740;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_277;
wire n_338;
wire n_477;
wire n_461;
wire n_333;
wire n_571;
wire n_693;
wire n_309;
wire n_512;
wire n_462;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_778;
wire n_306;
wire n_722;
wire n_458;
wire n_288;
wire n_770;
wire n_188;
wire n_190;
wire n_201;
wire n_263;
wire n_471;
wire n_609;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_711;
wire n_474;
wire n_765;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_736;
wire n_502;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_465;
wire n_358;
wire n_362;
wire n_170;
wire n_332;
wire n_161;
wire n_273;
wire n_349;
wire n_585;
wire n_270;
wire n_616;
wire n_230;
wire n_601;
wire n_279;
wire n_253;
wire n_261;
wire n_174;
wire n_289;
wire n_745;
wire n_627;
wire n_767;
wire n_172;
wire n_206;
wire n_217;
wire n_440;
wire n_726;
wire n_478;
wire n_545;
wire n_441;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_429;
wire n_534;
wire n_345;
wire n_210;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_730;
wire n_729;
wire n_176;
wire n_557;
wire n_182;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_647;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_710;
wire n_679;
wire n_707;
wire n_695;
wire n_180;
wire n_560;
wire n_656;
wire n_340;
wire n_207;
wire n_561;
wire n_346;
wire n_393;
wire n_229;
wire n_495;
wire n_487;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_177;
wire n_403;
wire n_453;
wire n_421;
wire n_720;
wire n_623;
wire n_405;
wire n_359;
wire n_490;
wire n_326;
wire n_768;
wire n_233;
wire n_404;
wire n_686;
wire n_205;
wire n_366;
wire n_572;
wire n_754;
wire n_712;
wire n_246;
wire n_596;
wire n_179;
wire n_410;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_412;
wire n_232;
wire n_327;
wire n_657;
wire n_728;
wire n_644;
wire n_202;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_732;
wire n_193;
wire n_251;
wire n_352;
wire n_160;
wire n_566;
wire n_426;
wire n_520;
wire n_565;
wire n_409;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_300;
wire n_651;
wire n_435;
wire n_159;
wire n_334;
wire n_599;
wire n_766;
wire n_541;
wire n_391;
wire n_701;
wire n_434;
wire n_645;
wire n_539;
wire n_175;
wire n_538;
wire n_666;
wire n_262;
wire n_238;
wire n_639;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_536;
wire n_531;
wire n_242;
wire n_360;
wire n_594;
wire n_764;
wire n_200;
wire n_162;
wire n_759;
wire n_222;
wire n_438;
wire n_713;
wire n_324;
wire n_634;
wire n_416;
wire n_199;
wire n_187;
wire n_401;
wire n_348;
wire n_166;
wire n_626;
wire n_424;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_747;
wire n_278;

INVx1_ASAP7_75t_L g157 ( 
.A(n_55),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_102),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_155),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_97),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_96),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_90),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_156),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_95),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_80),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_76),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_24),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_74),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_23),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_14),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_8),
.Y(n_171)
);

INVx2_ASAP7_75t_SL g172 ( 
.A(n_139),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_121),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_101),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_147),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_150),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_149),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_143),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_28),
.Y(n_179)
);

OR2x2_ASAP7_75t_L g180 ( 
.A(n_57),
.B(n_135),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_31),
.Y(n_181)
);

CKINVDCx14_ASAP7_75t_R g182 ( 
.A(n_59),
.Y(n_182)
);

BUFx10_ASAP7_75t_L g183 ( 
.A(n_153),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_54),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_83),
.Y(n_185)
);

BUFx10_ASAP7_75t_L g186 ( 
.A(n_33),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_58),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_13),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_20),
.Y(n_189)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_138),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_51),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_29),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_110),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_91),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_53),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_25),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_18),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_60),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_88),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_10),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_104),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_62),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_146),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_64),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_86),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_109),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_47),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_141),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_34),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_82),
.Y(n_210)
);

INVx2_ASAP7_75t_SL g211 ( 
.A(n_7),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_40),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_45),
.Y(n_213)
);

INVx5_ASAP7_75t_L g214 ( 
.A(n_166),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_200),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_182),
.B(n_0),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_190),
.B(n_0),
.Y(n_217)
);

INVx5_ASAP7_75t_L g218 ( 
.A(n_166),
.Y(n_218)
);

BUFx12f_ASAP7_75t_L g219 ( 
.A(n_183),
.Y(n_219)
);

BUFx8_ASAP7_75t_L g220 ( 
.A(n_211),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_210),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_200),
.Y(n_222)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_166),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_161),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_170),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_166),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_161),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_162),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_190),
.B(n_1),
.Y(n_229)
);

INVx2_ASAP7_75t_SL g230 ( 
.A(n_183),
.Y(n_230)
);

BUFx2_ASAP7_75t_L g231 ( 
.A(n_171),
.Y(n_231)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_183),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_188),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_157),
.Y(n_234)
);

AND2x4_ASAP7_75t_L g235 ( 
.A(n_162),
.B(n_2),
.Y(n_235)
);

NAND2x1p5_ASAP7_75t_L g236 ( 
.A(n_180),
.B(n_19),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_173),
.Y(n_237)
);

BUFx12f_ASAP7_75t_L g238 ( 
.A(n_186),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_210),
.Y(n_239)
);

BUFx12f_ASAP7_75t_L g240 ( 
.A(n_186),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_186),
.Y(n_241)
);

INVx5_ASAP7_75t_L g242 ( 
.A(n_172),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_173),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_158),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_198),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_163),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_182),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_247)
);

AND2x4_ASAP7_75t_L g248 ( 
.A(n_198),
.B(n_4),
.Y(n_248)
);

INVx5_ASAP7_75t_L g249 ( 
.A(n_189),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_164),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_165),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_212),
.B(n_5),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_212),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_175),
.Y(n_254)
);

INVx2_ASAP7_75t_SL g255 ( 
.A(n_159),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_176),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_219),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_226),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_238),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_228),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_240),
.Y(n_261)
);

INVxp33_ASAP7_75t_SL g262 ( 
.A(n_225),
.Y(n_262)
);

INVx2_ASAP7_75t_SL g263 ( 
.A(n_225),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_255),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_221),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_228),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_221),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_239),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_239),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_231),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_241),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_228),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_228),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_241),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_237),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_249),
.B(n_177),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_249),
.B(n_181),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_249),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_249),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_220),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_224),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_220),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_232),
.Y(n_283)
);

AOI21x1_ASAP7_75t_L g284 ( 
.A1(n_245),
.A2(n_196),
.B(n_184),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_230),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_242),
.B(n_232),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_227),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_237),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_242),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_242),
.B(n_185),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_237),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_237),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_243),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_242),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_243),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_216),
.B(n_160),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_243),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_256),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_256),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_256),
.Y(n_300)
);

HB1xp67_ASAP7_75t_L g301 ( 
.A(n_215),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_243),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_256),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_245),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_222),
.Y(n_305)
);

NOR3xp33_ASAP7_75t_L g306 ( 
.A(n_263),
.B(n_233),
.C(n_229),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_266),
.B(n_253),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_260),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_275),
.B(n_253),
.Y(n_309)
);

NAND3xp33_ASAP7_75t_L g310 ( 
.A(n_296),
.B(n_229),
.C(n_217),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_283),
.B(n_217),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_264),
.B(n_236),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_260),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_271),
.B(n_236),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_281),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_298),
.B(n_214),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_262),
.A2(n_247),
.B1(n_235),
.B2(n_248),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_258),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_299),
.B(n_300),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_287),
.B(n_252),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_258),
.Y(n_321)
);

OR2x2_ASAP7_75t_L g322 ( 
.A(n_301),
.B(n_252),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_305),
.B(n_234),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_272),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_270),
.A2(n_235),
.B1(n_248),
.B2(n_167),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_281),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_274),
.B(n_168),
.Y(n_327)
);

NOR3xp33_ASAP7_75t_L g328 ( 
.A(n_265),
.B(n_233),
.C(n_244),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_288),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_303),
.B(n_214),
.Y(n_330)
);

NOR3xp33_ASAP7_75t_L g331 ( 
.A(n_267),
.B(n_254),
.C(n_251),
.Y(n_331)
);

NAND2xp33_ASAP7_75t_L g332 ( 
.A(n_278),
.B(n_169),
.Y(n_332)
);

NOR3xp33_ASAP7_75t_L g333 ( 
.A(n_276),
.B(n_250),
.C(n_246),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_286),
.B(n_291),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_279),
.B(n_174),
.Y(n_335)
);

BUFx5_ASAP7_75t_L g336 ( 
.A(n_292),
.Y(n_336)
);

INVx2_ASAP7_75t_SL g337 ( 
.A(n_277),
.Y(n_337)
);

OR2x2_ASAP7_75t_L g338 ( 
.A(n_304),
.B(n_223),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_293),
.B(n_214),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_295),
.B(n_214),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_280),
.B(n_178),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_282),
.B(n_179),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_289),
.B(n_294),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_272),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_273),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_297),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_257),
.B(n_187),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_302),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_290),
.B(n_223),
.Y(n_349)
);

AO221x1_ASAP7_75t_L g350 ( 
.A1(n_273),
.A2(n_208),
.B1(n_202),
.B2(n_201),
.C(n_199),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_258),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_259),
.B(n_191),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_258),
.B(n_218),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_285),
.B(n_193),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_285),
.A2(n_205),
.B1(n_194),
.B2(n_213),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_261),
.B(n_195),
.Y(n_356)
);

INVx4_ASAP7_75t_L g357 ( 
.A(n_284),
.Y(n_357)
);

NAND2xp33_ASAP7_75t_L g358 ( 
.A(n_268),
.B(n_203),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_268),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_269),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_269),
.B(n_204),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_260),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_298),
.B(n_218),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_298),
.B(n_218),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_298),
.B(n_218),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_283),
.B(n_206),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_281),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_266),
.B(n_226),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_283),
.B(n_207),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_266),
.B(n_226),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_318),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_307),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_307),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_354),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_318),
.Y(n_375)
);

AOI22xp33_ASAP7_75t_L g376 ( 
.A1(n_310),
.A2(n_197),
.B1(n_192),
.B2(n_209),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_311),
.B(n_226),
.Y(n_377)
);

AND2x4_ASAP7_75t_SL g378 ( 
.A(n_360),
.B(n_21),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_320),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_323),
.B(n_6),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_308),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_313),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_309),
.Y(n_383)
);

INVx4_ASAP7_75t_L g384 ( 
.A(n_318),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_322),
.B(n_6),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_310),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_319),
.B(n_9),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_349),
.B(n_22),
.Y(n_388)
);

INVx3_ASAP7_75t_L g389 ( 
.A(n_324),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_309),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_315),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_321),
.Y(n_392)
);

AOI22xp33_ASAP7_75t_L g393 ( 
.A1(n_306),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_367),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_344),
.Y(n_395)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_359),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_317),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_355),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_398)
);

INVx5_ASAP7_75t_L g399 ( 
.A(n_321),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_337),
.B(n_15),
.Y(n_400)
);

INVx3_ASAP7_75t_L g401 ( 
.A(n_345),
.Y(n_401)
);

BUFx3_ASAP7_75t_L g402 ( 
.A(n_329),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_368),
.Y(n_403)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_334),
.A2(n_93),
.B(n_152),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_361),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_368),
.Y(n_406)
);

INVx4_ASAP7_75t_L g407 ( 
.A(n_321),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_370),
.Y(n_408)
);

NOR2x1p5_ASAP7_75t_L g409 ( 
.A(n_358),
.B(n_16),
.Y(n_409)
);

AOI21xp33_ASAP7_75t_L g410 ( 
.A1(n_312),
.A2(n_314),
.B(n_325),
.Y(n_410)
);

INVx3_ASAP7_75t_L g411 ( 
.A(n_362),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_346),
.B(n_26),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_351),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_348),
.B(n_27),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_336),
.B(n_30),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_326),
.B(n_17),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_370),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_328),
.A2(n_17),
.B1(n_32),
.B2(n_35),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_338),
.Y(n_419)
);

HB1xp67_ASAP7_75t_L g420 ( 
.A(n_331),
.Y(n_420)
);

AND2x4_ASAP7_75t_L g421 ( 
.A(n_333),
.B(n_36),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_336),
.B(n_37),
.Y(n_422)
);

NOR3xp33_ASAP7_75t_SL g423 ( 
.A(n_366),
.B(n_38),
.C(n_39),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_336),
.B(n_41),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_327),
.Y(n_425)
);

INVx4_ASAP7_75t_L g426 ( 
.A(n_357),
.Y(n_426)
);

BUFx2_ASAP7_75t_L g427 ( 
.A(n_343),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_357),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_369),
.B(n_42),
.Y(n_429)
);

AND2x4_ASAP7_75t_L g430 ( 
.A(n_335),
.B(n_43),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_336),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_347),
.B(n_44),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_336),
.Y(n_433)
);

OR2x4_ASAP7_75t_L g434 ( 
.A(n_341),
.B(n_342),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_350),
.A2(n_46),
.B1(n_48),
.B2(n_49),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_353),
.Y(n_436)
);

AOI22xp33_ASAP7_75t_L g437 ( 
.A1(n_332),
.A2(n_50),
.B1(n_52),
.B2(n_56),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_339),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_340),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_316),
.Y(n_440)
);

INVx4_ASAP7_75t_L g441 ( 
.A(n_440),
.Y(n_441)
);

NOR2xp67_ASAP7_75t_SL g442 ( 
.A(n_428),
.B(n_399),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_L g443 ( 
.A1(n_379),
.A2(n_365),
.B1(n_364),
.B2(n_363),
.Y(n_443)
);

AOI21xp5_ASAP7_75t_L g444 ( 
.A1(n_388),
.A2(n_330),
.B(n_356),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_391),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_410),
.B(n_352),
.Y(n_446)
);

AOI222xp33_ASAP7_75t_L g447 ( 
.A1(n_397),
.A2(n_61),
.B1(n_63),
.B2(n_65),
.C1(n_66),
.C2(n_67),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_374),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_430),
.B(n_68),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_394),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_430),
.B(n_69),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_L g452 ( 
.A1(n_405),
.A2(n_70),
.B1(n_71),
.B2(n_72),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_371),
.Y(n_453)
);

O2A1O1Ixp33_ASAP7_75t_L g454 ( 
.A1(n_387),
.A2(n_73),
.B(n_75),
.C(n_77),
.Y(n_454)
);

INVx1_ASAP7_75t_SL g455 ( 
.A(n_396),
.Y(n_455)
);

BUFx4f_ASAP7_75t_L g456 ( 
.A(n_421),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_427),
.B(n_78),
.Y(n_457)
);

AOI21xp5_ASAP7_75t_L g458 ( 
.A1(n_428),
.A2(n_79),
.B(n_81),
.Y(n_458)
);

OAI21x1_ASAP7_75t_L g459 ( 
.A1(n_431),
.A2(n_84),
.B(n_85),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_381),
.Y(n_460)
);

O2A1O1Ixp33_ASAP7_75t_L g461 ( 
.A1(n_400),
.A2(n_373),
.B(n_372),
.C(n_390),
.Y(n_461)
);

INVx3_ASAP7_75t_L g462 ( 
.A(n_402),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_383),
.B(n_87),
.Y(n_463)
);

AOI21xp5_ASAP7_75t_L g464 ( 
.A1(n_428),
.A2(n_89),
.B(n_92),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_385),
.B(n_380),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_371),
.Y(n_466)
);

OAI21xp5_ASAP7_75t_L g467 ( 
.A1(n_403),
.A2(n_94),
.B(n_98),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_419),
.B(n_99),
.Y(n_468)
);

AND2x4_ASAP7_75t_L g469 ( 
.A(n_378),
.B(n_100),
.Y(n_469)
);

A2O1A1Ixp33_ASAP7_75t_L g470 ( 
.A1(n_376),
.A2(n_406),
.B(n_408),
.C(n_416),
.Y(n_470)
);

NAND2x1p5_ASAP7_75t_L g471 ( 
.A(n_399),
.B(n_103),
.Y(n_471)
);

A2O1A1Ixp33_ASAP7_75t_L g472 ( 
.A1(n_438),
.A2(n_105),
.B(n_106),
.C(n_107),
.Y(n_472)
);

AOI221xp5_ASAP7_75t_L g473 ( 
.A1(n_393),
.A2(n_108),
.B1(n_111),
.B2(n_112),
.C(n_113),
.Y(n_473)
);

AOI21xp5_ASAP7_75t_L g474 ( 
.A1(n_436),
.A2(n_114),
.B(n_115),
.Y(n_474)
);

AO21x1_ASAP7_75t_L g475 ( 
.A1(n_415),
.A2(n_116),
.B(n_117),
.Y(n_475)
);

INVx4_ASAP7_75t_L g476 ( 
.A(n_371),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_377),
.B(n_118),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_420),
.B(n_119),
.Y(n_478)
);

BUFx2_ASAP7_75t_L g479 ( 
.A(n_421),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_417),
.B(n_120),
.Y(n_480)
);

AND3x1_ASAP7_75t_SL g481 ( 
.A(n_409),
.B(n_397),
.C(n_398),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_382),
.Y(n_482)
);

AND2x4_ASAP7_75t_L g483 ( 
.A(n_440),
.B(n_122),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_425),
.Y(n_484)
);

AOI221xp5_ASAP7_75t_L g485 ( 
.A1(n_386),
.A2(n_123),
.B1(n_124),
.B2(n_125),
.C(n_126),
.Y(n_485)
);

INVx4_ASAP7_75t_L g486 ( 
.A(n_375),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_L g487 ( 
.A1(n_434),
.A2(n_127),
.B1(n_128),
.B2(n_129),
.Y(n_487)
);

AOI21xp5_ASAP7_75t_L g488 ( 
.A1(n_399),
.A2(n_130),
.B(n_131),
.Y(n_488)
);

INVxp67_ASAP7_75t_SL g489 ( 
.A(n_375),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_395),
.Y(n_490)
);

OR2x6_ASAP7_75t_L g491 ( 
.A(n_409),
.B(n_132),
.Y(n_491)
);

INVx1_ASAP7_75t_SL g492 ( 
.A(n_386),
.Y(n_492)
);

O2A1O1Ixp33_ASAP7_75t_L g493 ( 
.A1(n_429),
.A2(n_133),
.B(n_134),
.C(n_136),
.Y(n_493)
);

INVx4_ASAP7_75t_L g494 ( 
.A(n_440),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_389),
.Y(n_495)
);

AOI21xp5_ASAP7_75t_L g496 ( 
.A1(n_439),
.A2(n_137),
.B(n_140),
.Y(n_496)
);

O2A1O1Ixp33_ASAP7_75t_L g497 ( 
.A1(n_432),
.A2(n_142),
.B(n_144),
.C(n_145),
.Y(n_497)
);

INVx1_ASAP7_75t_SL g498 ( 
.A(n_455),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_445),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_465),
.B(n_417),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_450),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_459),
.Y(n_502)
);

AND2x4_ASAP7_75t_L g503 ( 
.A(n_479),
.B(n_417),
.Y(n_503)
);

OAI21x1_ASAP7_75t_L g504 ( 
.A1(n_480),
.A2(n_422),
.B(n_424),
.Y(n_504)
);

HB1xp67_ASAP7_75t_L g505 ( 
.A(n_462),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_448),
.Y(n_506)
);

NOR2xp67_ASAP7_75t_SL g507 ( 
.A(n_453),
.B(n_392),
.Y(n_507)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_453),
.Y(n_508)
);

INVx6_ASAP7_75t_L g509 ( 
.A(n_441),
.Y(n_509)
);

BUFx4f_ASAP7_75t_SL g510 ( 
.A(n_469),
.Y(n_510)
);

CKINVDCx14_ASAP7_75t_R g511 ( 
.A(n_484),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_460),
.Y(n_512)
);

NAND2x1p5_ASAP7_75t_L g513 ( 
.A(n_442),
.B(n_426),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_482),
.Y(n_514)
);

AO21x2_ASAP7_75t_L g515 ( 
.A1(n_467),
.A2(n_412),
.B(n_414),
.Y(n_515)
);

INVx1_ASAP7_75t_SL g516 ( 
.A(n_468),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_490),
.Y(n_517)
);

BUFx3_ASAP7_75t_L g518 ( 
.A(n_483),
.Y(n_518)
);

NAND2x1p5_ASAP7_75t_L g519 ( 
.A(n_494),
.B(n_426),
.Y(n_519)
);

BUFx2_ASAP7_75t_SL g520 ( 
.A(n_483),
.Y(n_520)
);

CKINVDCx16_ASAP7_75t_R g521 ( 
.A(n_491),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_453),
.Y(n_522)
);

BUFx12f_ASAP7_75t_L g523 ( 
.A(n_491),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_495),
.Y(n_524)
);

BUFx12f_ASAP7_75t_L g525 ( 
.A(n_469),
.Y(n_525)
);

OAI21x1_ASAP7_75t_L g526 ( 
.A1(n_477),
.A2(n_433),
.B(n_404),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_466),
.Y(n_527)
);

OAI21x1_ASAP7_75t_SL g528 ( 
.A1(n_475),
.A2(n_418),
.B(n_437),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_466),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_456),
.B(n_418),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_466),
.Y(n_531)
);

OAI21x1_ASAP7_75t_L g532 ( 
.A1(n_444),
.A2(n_411),
.B(n_389),
.Y(n_532)
);

CKINVDCx11_ASAP7_75t_R g533 ( 
.A(n_492),
.Y(n_533)
);

INVx8_ASAP7_75t_L g534 ( 
.A(n_476),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_476),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_486),
.Y(n_536)
);

OAI21x1_ASAP7_75t_L g537 ( 
.A1(n_463),
.A2(n_474),
.B(n_496),
.Y(n_537)
);

OAI21x1_ASAP7_75t_L g538 ( 
.A1(n_461),
.A2(n_401),
.B(n_411),
.Y(n_538)
);

BUFx6f_ASAP7_75t_L g539 ( 
.A(n_486),
.Y(n_539)
);

INVx2_ASAP7_75t_SL g540 ( 
.A(n_449),
.Y(n_540)
);

OAI21x1_ASAP7_75t_L g541 ( 
.A1(n_458),
.A2(n_401),
.B(n_435),
.Y(n_541)
);

AO21x2_ASAP7_75t_L g542 ( 
.A1(n_470),
.A2(n_435),
.B(n_423),
.Y(n_542)
);

OAI21x1_ASAP7_75t_L g543 ( 
.A1(n_464),
.A2(n_413),
.B(n_384),
.Y(n_543)
);

AO21x2_ASAP7_75t_L g544 ( 
.A1(n_446),
.A2(n_413),
.B(n_392),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_489),
.Y(n_545)
);

INVx2_ASAP7_75t_SL g546 ( 
.A(n_451),
.Y(n_546)
);

OAI21x1_ASAP7_75t_L g547 ( 
.A1(n_488),
.A2(n_413),
.B(n_384),
.Y(n_547)
);

AOI22xp33_ASAP7_75t_L g548 ( 
.A1(n_530),
.A2(n_447),
.B1(n_473),
.B2(n_485),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_524),
.Y(n_549)
);

INVx3_ASAP7_75t_L g550 ( 
.A(n_536),
.Y(n_550)
);

AOI22xp33_ASAP7_75t_SL g551 ( 
.A1(n_521),
.A2(n_457),
.B1(n_478),
.B2(n_481),
.Y(n_551)
);

BUFx2_ASAP7_75t_L g552 ( 
.A(n_498),
.Y(n_552)
);

AND2x4_ASAP7_75t_L g553 ( 
.A(n_518),
.B(n_472),
.Y(n_553)
);

OAI21x1_ASAP7_75t_L g554 ( 
.A1(n_502),
.A2(n_497),
.B(n_493),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_524),
.Y(n_555)
);

AOI21x1_ASAP7_75t_L g556 ( 
.A1(n_530),
.A2(n_443),
.B(n_487),
.Y(n_556)
);

BUFx2_ASAP7_75t_L g557 ( 
.A(n_500),
.Y(n_557)
);

AOI22xp33_ASAP7_75t_SL g558 ( 
.A1(n_523),
.A2(n_452),
.B1(n_471),
.B2(n_454),
.Y(n_558)
);

OA21x2_ASAP7_75t_L g559 ( 
.A1(n_504),
.A2(n_407),
.B(n_375),
.Y(n_559)
);

HB1xp67_ASAP7_75t_L g560 ( 
.A(n_500),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_520),
.B(n_407),
.Y(n_561)
);

NOR2x1_ASAP7_75t_R g562 ( 
.A(n_506),
.B(n_392),
.Y(n_562)
);

INVx5_ASAP7_75t_L g563 ( 
.A(n_522),
.Y(n_563)
);

NAND2x1p5_ASAP7_75t_L g564 ( 
.A(n_518),
.B(n_148),
.Y(n_564)
);

BUFx2_ASAP7_75t_R g565 ( 
.A(n_506),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_516),
.B(n_503),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_499),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_533),
.B(n_151),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_503),
.B(n_154),
.Y(n_569)
);

BUFx2_ASAP7_75t_R g570 ( 
.A(n_542),
.Y(n_570)
);

OAI22xp5_ASAP7_75t_L g571 ( 
.A1(n_540),
.A2(n_546),
.B1(n_503),
.B2(n_501),
.Y(n_571)
);

AOI22xp33_ASAP7_75t_L g572 ( 
.A1(n_540),
.A2(n_546),
.B1(n_533),
.B2(n_528),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_538),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_538),
.Y(n_574)
);

BUFx6f_ASAP7_75t_L g575 ( 
.A(n_522),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_512),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_511),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_514),
.Y(n_578)
);

BUFx2_ASAP7_75t_L g579 ( 
.A(n_525),
.Y(n_579)
);

CKINVDCx11_ASAP7_75t_R g580 ( 
.A(n_523),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_517),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_545),
.Y(n_582)
);

AOI22xp33_ASAP7_75t_L g583 ( 
.A1(n_542),
.A2(n_510),
.B1(n_525),
.B2(n_505),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_532),
.Y(n_584)
);

AOI21x1_ASAP7_75t_L g585 ( 
.A1(n_526),
.A2(n_532),
.B(n_504),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_527),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_527),
.Y(n_587)
);

CKINVDCx11_ASAP7_75t_R g588 ( 
.A(n_536),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_535),
.B(n_531),
.Y(n_589)
);

BUFx10_ASAP7_75t_L g590 ( 
.A(n_509),
.Y(n_590)
);

AND3x2_ASAP7_75t_L g591 ( 
.A(n_553),
.B(n_535),
.C(n_529),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_R g592 ( 
.A(n_588),
.B(n_511),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_560),
.B(n_557),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_557),
.B(n_508),
.Y(n_594)
);

CKINVDCx20_ASAP7_75t_R g595 ( 
.A(n_588),
.Y(n_595)
);

OAI22xp5_ASAP7_75t_L g596 ( 
.A1(n_548),
.A2(n_509),
.B1(n_513),
.B2(n_519),
.Y(n_596)
);

OR2x2_ASAP7_75t_L g597 ( 
.A(n_566),
.B(n_508),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_569),
.B(n_508),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_569),
.B(n_522),
.Y(n_599)
);

HB1xp67_ASAP7_75t_L g600 ( 
.A(n_549),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_576),
.Y(n_601)
);

CKINVDCx16_ASAP7_75t_R g602 ( 
.A(n_552),
.Y(n_602)
);

CKINVDCx16_ASAP7_75t_R g603 ( 
.A(n_552),
.Y(n_603)
);

INVx2_ASAP7_75t_SL g604 ( 
.A(n_590),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_551),
.B(n_509),
.Y(n_605)
);

NAND2xp33_ASAP7_75t_R g606 ( 
.A(n_577),
.B(n_502),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_576),
.Y(n_607)
);

HB1xp67_ASAP7_75t_L g608 ( 
.A(n_549),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_565),
.Y(n_609)
);

BUFx3_ASAP7_75t_L g610 ( 
.A(n_579),
.Y(n_610)
);

INVxp67_ASAP7_75t_L g611 ( 
.A(n_562),
.Y(n_611)
);

A2O1A1Ixp33_ASAP7_75t_L g612 ( 
.A1(n_572),
.A2(n_541),
.B(n_537),
.C(n_526),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_578),
.B(n_539),
.Y(n_613)
);

XOR2xp5_ASAP7_75t_L g614 ( 
.A(n_577),
.B(n_564),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_580),
.Y(n_615)
);

AOI22xp33_ASAP7_75t_L g616 ( 
.A1(n_558),
.A2(n_583),
.B1(n_553),
.B2(n_581),
.Y(n_616)
);

NAND2xp33_ASAP7_75t_R g617 ( 
.A(n_579),
.B(n_502),
.Y(n_617)
);

AND2x2_ASAP7_75t_L g618 ( 
.A(n_586),
.B(n_522),
.Y(n_618)
);

AOI22xp33_ASAP7_75t_L g619 ( 
.A1(n_553),
.A2(n_515),
.B1(n_544),
.B2(n_541),
.Y(n_619)
);

HB1xp67_ASAP7_75t_L g620 ( 
.A(n_555),
.Y(n_620)
);

HB1xp67_ASAP7_75t_L g621 ( 
.A(n_555),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_567),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_582),
.B(n_539),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_587),
.Y(n_624)
);

AOI22xp33_ASAP7_75t_L g625 ( 
.A1(n_571),
.A2(n_515),
.B1(n_536),
.B2(n_539),
.Y(n_625)
);

NOR3xp33_ASAP7_75t_SL g626 ( 
.A(n_568),
.B(n_507),
.C(n_534),
.Y(n_626)
);

AND2x4_ASAP7_75t_L g627 ( 
.A(n_550),
.B(n_536),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_570),
.B(n_539),
.Y(n_628)
);

AOI22xp33_ASAP7_75t_L g629 ( 
.A1(n_580),
.A2(n_564),
.B1(n_589),
.B2(n_561),
.Y(n_629)
);

NAND2xp33_ASAP7_75t_SL g630 ( 
.A(n_575),
.B(n_534),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_575),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_575),
.Y(n_632)
);

INVx4_ASAP7_75t_L g633 ( 
.A(n_590),
.Y(n_633)
);

OR2x4_ASAP7_75t_L g634 ( 
.A(n_575),
.B(n_534),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_550),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_575),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_600),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_607),
.Y(n_638)
);

BUFx3_ASAP7_75t_L g639 ( 
.A(n_634),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_601),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_600),
.Y(n_641)
);

OR2x2_ASAP7_75t_L g642 ( 
.A(n_593),
.B(n_573),
.Y(n_642)
);

OAI21xp5_ASAP7_75t_L g643 ( 
.A1(n_596),
.A2(n_556),
.B(n_629),
.Y(n_643)
);

INVx2_ASAP7_75t_SL g644 ( 
.A(n_634),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_608),
.Y(n_645)
);

HB1xp67_ASAP7_75t_L g646 ( 
.A(n_608),
.Y(n_646)
);

AOI22xp33_ASAP7_75t_SL g647 ( 
.A1(n_628),
.A2(n_605),
.B1(n_603),
.B2(n_602),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_620),
.B(n_574),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_620),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_621),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_597),
.B(n_564),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_621),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_594),
.B(n_584),
.Y(n_653)
);

INVxp67_ASAP7_75t_SL g654 ( 
.A(n_613),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_622),
.Y(n_655)
);

HB1xp67_ASAP7_75t_L g656 ( 
.A(n_631),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_599),
.B(n_563),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_598),
.B(n_623),
.Y(n_658)
);

NOR2x1_ASAP7_75t_L g659 ( 
.A(n_633),
.B(n_559),
.Y(n_659)
);

HB1xp67_ASAP7_75t_L g660 ( 
.A(n_632),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_624),
.B(n_559),
.Y(n_661)
);

OAI211xp5_ASAP7_75t_L g662 ( 
.A1(n_616),
.A2(n_585),
.B(n_554),
.C(n_559),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_612),
.Y(n_663)
);

AND2x4_ASAP7_75t_L g664 ( 
.A(n_591),
.B(n_543),
.Y(n_664)
);

INVx2_ASAP7_75t_SL g665 ( 
.A(n_636),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_635),
.B(n_618),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_616),
.B(n_563),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_619),
.B(n_563),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_591),
.Y(n_669)
);

OR2x2_ASAP7_75t_L g670 ( 
.A(n_619),
.B(n_629),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_654),
.B(n_628),
.Y(n_671)
);

OR2x2_ASAP7_75t_L g672 ( 
.A(n_642),
.B(n_625),
.Y(n_672)
);

NOR2x1_ASAP7_75t_SL g673 ( 
.A(n_662),
.B(n_617),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_658),
.B(n_610),
.Y(n_674)
);

AND2x2_ASAP7_75t_L g675 ( 
.A(n_653),
.B(n_648),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_637),
.Y(n_676)
);

BUFx2_ASAP7_75t_L g677 ( 
.A(n_646),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_638),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_655),
.B(n_614),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_637),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_641),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_641),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_653),
.B(n_648),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_661),
.B(n_625),
.Y(n_684)
);

HB1xp67_ASAP7_75t_L g685 ( 
.A(n_656),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_645),
.Y(n_686)
);

OAI22xp5_ASAP7_75t_L g687 ( 
.A1(n_647),
.A2(n_626),
.B1(n_595),
.B2(n_611),
.Y(n_687)
);

BUFx2_ASAP7_75t_L g688 ( 
.A(n_659),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_650),
.B(n_626),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_655),
.B(n_666),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_645),
.Y(n_691)
);

NAND3xp33_ASAP7_75t_L g692 ( 
.A(n_643),
.B(n_606),
.C(n_633),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_650),
.B(n_627),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_649),
.Y(n_694)
);

HB1xp67_ASAP7_75t_L g695 ( 
.A(n_660),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_666),
.B(n_604),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_652),
.B(n_627),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_678),
.Y(n_698)
);

HB1xp67_ASAP7_75t_L g699 ( 
.A(n_685),
.Y(n_699)
);

OR2x2_ASAP7_75t_L g700 ( 
.A(n_677),
.B(n_642),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_682),
.Y(n_701)
);

NAND2x1p5_ASAP7_75t_L g702 ( 
.A(n_688),
.B(n_664),
.Y(n_702)
);

NAND2xp33_ASAP7_75t_L g703 ( 
.A(n_692),
.B(n_592),
.Y(n_703)
);

OR2x2_ASAP7_75t_L g704 ( 
.A(n_677),
.B(n_670),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_682),
.Y(n_705)
);

OR2x2_ASAP7_75t_L g706 ( 
.A(n_695),
.B(n_670),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_675),
.B(n_652),
.Y(n_707)
);

HB1xp67_ASAP7_75t_L g708 ( 
.A(n_688),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_675),
.B(n_668),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_676),
.Y(n_710)
);

OR2x2_ASAP7_75t_L g711 ( 
.A(n_683),
.B(n_649),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_678),
.Y(n_712)
);

AND2x2_ASAP7_75t_L g713 ( 
.A(n_683),
.B(n_668),
.Y(n_713)
);

OR2x2_ASAP7_75t_L g714 ( 
.A(n_672),
.B(n_663),
.Y(n_714)
);

BUFx3_ASAP7_75t_L g715 ( 
.A(n_689),
.Y(n_715)
);

AOI22xp5_ASAP7_75t_L g716 ( 
.A1(n_703),
.A2(n_687),
.B1(n_667),
.B2(n_689),
.Y(n_716)
);

HB1xp67_ASAP7_75t_L g717 ( 
.A(n_708),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_701),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_705),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_710),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_699),
.B(n_686),
.Y(n_721)
);

OR2x2_ASAP7_75t_L g722 ( 
.A(n_704),
.B(n_672),
.Y(n_722)
);

AOI22xp5_ASAP7_75t_L g723 ( 
.A1(n_703),
.A2(n_671),
.B1(n_663),
.B2(n_684),
.Y(n_723)
);

HB1xp67_ASAP7_75t_L g724 ( 
.A(n_708),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_699),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_698),
.Y(n_726)
);

INVx1_ASAP7_75t_SL g727 ( 
.A(n_722),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_718),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_719),
.Y(n_729)
);

INVxp67_ASAP7_75t_L g730 ( 
.A(n_721),
.Y(n_730)
);

NOR3xp33_ASAP7_75t_L g731 ( 
.A(n_716),
.B(n_679),
.C(n_651),
.Y(n_731)
);

OAI321xp33_ASAP7_75t_L g732 ( 
.A1(n_730),
.A2(n_723),
.A3(n_714),
.B1(n_702),
.B2(n_725),
.C(n_721),
.Y(n_732)
);

AND2x2_ASAP7_75t_L g733 ( 
.A(n_727),
.B(n_715),
.Y(n_733)
);

NAND2x1_ASAP7_75t_L g734 ( 
.A(n_728),
.B(n_726),
.Y(n_734)
);

AOI211xp5_ASAP7_75t_L g735 ( 
.A1(n_731),
.A2(n_729),
.B(n_706),
.C(n_696),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_733),
.B(n_615),
.Y(n_736)
);

NOR3x1_ASAP7_75t_L g737 ( 
.A(n_734),
.B(n_674),
.C(n_644),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_735),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_732),
.B(n_715),
.Y(n_739)
);

XNOR2x1_ASAP7_75t_SL g740 ( 
.A(n_738),
.B(n_609),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_739),
.B(n_720),
.Y(n_741)
);

AOI211xp5_ASAP7_75t_L g742 ( 
.A1(n_740),
.A2(n_736),
.B(n_737),
.C(n_644),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_741),
.B(n_724),
.Y(n_743)
);

O2A1O1Ixp33_ASAP7_75t_L g744 ( 
.A1(n_741),
.A2(n_717),
.B(n_669),
.C(n_702),
.Y(n_744)
);

AND3x4_ASAP7_75t_L g745 ( 
.A(n_742),
.B(n_639),
.C(n_669),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_743),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_744),
.Y(n_747)
);

INVx2_ASAP7_75t_SL g748 ( 
.A(n_743),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_743),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_743),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_743),
.Y(n_751)
);

AOI221xp5_ASAP7_75t_L g752 ( 
.A1(n_747),
.A2(n_694),
.B1(n_680),
.B2(n_691),
.C(n_681),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_748),
.Y(n_753)
);

OR2x2_ASAP7_75t_L g754 ( 
.A(n_746),
.B(n_700),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_749),
.Y(n_755)
);

AND3x4_ASAP7_75t_L g756 ( 
.A(n_750),
.B(n_639),
.C(n_664),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_751),
.B(n_713),
.Y(n_757)
);

NOR3xp33_ASAP7_75t_L g758 ( 
.A(n_753),
.B(n_751),
.C(n_745),
.Y(n_758)
);

HB1xp67_ASAP7_75t_L g759 ( 
.A(n_755),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_757),
.Y(n_760)
);

NAND2xp33_ASAP7_75t_L g761 ( 
.A(n_754),
.B(n_534),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_759),
.Y(n_762)
);

AOI22xp5_ASAP7_75t_L g763 ( 
.A1(n_758),
.A2(n_756),
.B1(n_752),
.B2(n_639),
.Y(n_763)
);

INVxp67_ASAP7_75t_L g764 ( 
.A(n_760),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_761),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_759),
.Y(n_766)
);

AOI22xp33_ASAP7_75t_L g767 ( 
.A1(n_762),
.A2(n_630),
.B1(n_665),
.B2(n_697),
.Y(n_767)
);

AOI22xp5_ASAP7_75t_L g768 ( 
.A1(n_766),
.A2(n_665),
.B1(n_657),
.B2(n_712),
.Y(n_768)
);

AOI22xp33_ASAP7_75t_L g769 ( 
.A1(n_765),
.A2(n_693),
.B1(n_697),
.B2(n_684),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_764),
.B(n_698),
.Y(n_770)
);

AOI22xp5_ASAP7_75t_L g771 ( 
.A1(n_763),
.A2(n_712),
.B1(n_693),
.B2(n_690),
.Y(n_771)
);

AOI22xp5_ASAP7_75t_L g772 ( 
.A1(n_771),
.A2(n_590),
.B1(n_709),
.B2(n_707),
.Y(n_772)
);

NAND2xp33_ASAP7_75t_R g773 ( 
.A(n_770),
.B(n_543),
.Y(n_773)
);

CKINVDCx20_ASAP7_75t_R g774 ( 
.A(n_768),
.Y(n_774)
);

AOI22xp5_ASAP7_75t_L g775 ( 
.A1(n_774),
.A2(n_767),
.B1(n_769),
.B2(n_563),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_772),
.Y(n_776)
);

OAI22xp5_ASAP7_75t_L g777 ( 
.A1(n_773),
.A2(n_711),
.B1(n_659),
.B2(n_563),
.Y(n_777)
);

AOI21xp5_ASAP7_75t_L g778 ( 
.A1(n_776),
.A2(n_775),
.B(n_777),
.Y(n_778)
);

AOI222xp33_ASAP7_75t_L g779 ( 
.A1(n_778),
.A2(n_673),
.B1(n_664),
.B2(n_638),
.C1(n_640),
.C2(n_554),
.Y(n_779)
);

OR2x6_ASAP7_75t_L g780 ( 
.A(n_779),
.B(n_513),
.Y(n_780)
);

AOI211xp5_ASAP7_75t_L g781 ( 
.A1(n_780),
.A2(n_547),
.B(n_664),
.C(n_640),
.Y(n_781)
);


endmodule