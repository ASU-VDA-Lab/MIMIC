module real_jpeg_21675_n_17 (n_8, n_0, n_2, n_10, n_9, n_12, n_345, n_6, n_346, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_17);

input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_345;
input n_6;
input n_346;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_0),
.A2(n_70),
.B1(n_71),
.B2(n_130),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_0),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_0),
.A2(n_52),
.B1(n_54),
.B2(n_130),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_0),
.A2(n_32),
.B1(n_33),
.B2(n_130),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_0),
.A2(n_24),
.B1(n_26),
.B2(n_130),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_1),
.A2(n_24),
.B1(n_26),
.B2(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_1),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_1),
.A2(n_32),
.B1(n_33),
.B2(n_63),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_1),
.A2(n_63),
.B1(n_70),
.B2(n_71),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g258 ( 
.A1(n_1),
.A2(n_52),
.B1(n_54),
.B2(n_63),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_2),
.A2(n_24),
.B1(n_26),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_2),
.A2(n_32),
.B1(n_33),
.B2(n_35),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_2),
.A2(n_35),
.B1(n_52),
.B2(n_54),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_2),
.A2(n_35),
.B1(n_70),
.B2(n_71),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_3),
.A2(n_52),
.B1(n_54),
.B2(n_125),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_3),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_3),
.A2(n_70),
.B1(n_71),
.B2(n_125),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_3),
.A2(n_32),
.B1(n_33),
.B2(n_125),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_3),
.A2(n_24),
.B1(n_26),
.B2(n_125),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_4),
.A2(n_23),
.B1(n_24),
.B2(n_26),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_4),
.A2(n_23),
.B1(n_32),
.B2(n_33),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_4),
.A2(n_23),
.B1(n_70),
.B2(n_71),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_4),
.A2(n_23),
.B1(n_52),
.B2(n_54),
.Y(n_290)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_6),
.A2(n_24),
.B1(n_26),
.B2(n_94),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_6),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_6),
.A2(n_70),
.B1(n_71),
.B2(n_94),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_L g221 ( 
.A1(n_6),
.A2(n_52),
.B1(n_54),
.B2(n_94),
.Y(n_221)
);

OAI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_6),
.A2(n_32),
.B1(n_33),
.B2(n_94),
.Y(n_264)
);

A2O1A1O1Ixp25_ASAP7_75t_L g109 ( 
.A1(n_7),
.A2(n_54),
.B(n_66),
.C(n_110),
.D(n_111),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_7),
.B(n_54),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_7),
.B(n_51),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_7),
.Y(n_149)
);

OAI21xp33_ASAP7_75t_L g155 ( 
.A1(n_7),
.A2(n_131),
.B(n_133),
.Y(n_155)
);

A2O1A1O1Ixp25_ASAP7_75t_L g169 ( 
.A1(n_7),
.A2(n_32),
.B(n_48),
.C(n_170),
.D(n_171),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_7),
.B(n_32),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_7),
.B(n_36),
.Y(n_193)
);

AOI21xp33_ASAP7_75t_L g209 ( 
.A1(n_7),
.A2(n_33),
.B(n_210),
.Y(n_209)
);

OAI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_7),
.A2(n_24),
.B1(n_26),
.B2(n_149),
.Y(n_227)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_8),
.Y(n_132)
);

INVx8_ASAP7_75t_L g151 ( 
.A(n_8),
.Y(n_151)
);

BUFx10_ASAP7_75t_L g70 ( 
.A(n_9),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_10),
.A2(n_24),
.B1(n_26),
.B2(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_10),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_10),
.A2(n_61),
.B1(n_70),
.B2(n_71),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_10),
.A2(n_52),
.B1(n_54),
.B2(n_61),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_10),
.A2(n_32),
.B1(n_33),
.B2(n_61),
.Y(n_283)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_12),
.A2(n_52),
.B1(n_54),
.B2(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_12),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_12),
.A2(n_70),
.B1(n_71),
.B2(n_113),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_12),
.A2(n_32),
.B1(n_33),
.B2(n_113),
.Y(n_172)
);

OAI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_12),
.A2(n_24),
.B1(n_26),
.B2(n_113),
.Y(n_230)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_14),
.A2(n_29),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_15),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_40),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_38),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_37),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_21),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_21),
.B(n_39),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_21),
.B(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_21),
.B(n_42),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_27),
.B1(n_34),
.B2(n_36),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_22),
.A2(n_27),
.B1(n_36),
.B2(n_76),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_24),
.Y(n_26)
);

A2O1A1Ixp33_ASAP7_75t_L g28 ( 
.A1(n_24),
.A2(n_29),
.B(n_30),
.C(n_31),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_29),
.Y(n_30)
);

A2O1A1Ixp33_ASAP7_75t_L g208 ( 
.A1(n_24),
.A2(n_29),
.B(n_149),
.C(n_209),
.Y(n_208)
);

BUFx2_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_SL g37 ( 
.A1(n_27),
.A2(n_34),
.B(n_36),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_27),
.A2(n_227),
.B(n_228),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_27),
.B(n_230),
.Y(n_239)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_28),
.A2(n_31),
.B1(n_60),
.B2(n_62),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_28),
.A2(n_31),
.B1(n_60),
.B2(n_93),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_28),
.A2(n_31),
.B1(n_238),
.B2(n_267),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_28),
.A2(n_229),
.B(n_267),
.Y(n_285)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_29),
.Y(n_210)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

OAI21xp33_ASAP7_75t_L g237 ( 
.A1(n_31),
.A2(n_238),
.B(n_239),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_31),
.A2(n_93),
.B(n_239),
.Y(n_309)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

O2A1O1Ixp33_ASAP7_75t_SL g48 ( 
.A1(n_33),
.A2(n_49),
.B(n_50),
.C(n_51),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_49),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_36),
.B(n_230),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_37),
.Y(n_39)
);

OAI21x1_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_80),
.B(n_343),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_75),
.C(n_77),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_43),
.A2(n_44),
.B1(n_83),
.B2(n_85),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_58),
.C(n_64),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_45),
.A2(n_46),
.B1(n_64),
.B2(n_91),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_47),
.A2(n_55),
.B1(n_56),
.B2(n_57),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_47),
.A2(n_55),
.B1(n_56),
.B2(n_98),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_47),
.A2(n_56),
.B1(n_189),
.B2(n_224),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_47),
.A2(n_224),
.B(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_48),
.A2(n_51),
.B(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_48),
.B(n_191),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_48),
.A2(n_51),
.B1(n_264),
.B2(n_283),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_48),
.A2(n_51),
.B1(n_99),
.B2(n_283),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_49),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_51)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_49),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_50),
.Y(n_178)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_52),
.Y(n_54)
);

O2A1O1Ixp33_ASAP7_75t_L g66 ( 
.A1(n_52),
.A2(n_67),
.B(n_68),
.C(n_69),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_67),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_52),
.B(n_53),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_54),
.A2(n_170),
.B1(n_177),
.B2(n_178),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_56),
.B(n_172),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_56),
.A2(n_189),
.B(n_190),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_56),
.A2(n_190),
.B(n_263),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_57),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_58),
.A2(n_59),
.B1(n_89),
.B2(n_90),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_62),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_64),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_64),
.A2(n_91),
.B1(n_96),
.B2(n_97),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_SL g64 ( 
.A1(n_65),
.A2(n_73),
.B(n_74),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_65),
.A2(n_73),
.B1(n_124),
.B2(n_168),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_65),
.A2(n_168),
.B(n_200),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_65),
.A2(n_73),
.B1(n_221),
.B2(n_249),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_65),
.A2(n_73),
.B1(n_249),
.B2(n_258),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_65),
.A2(n_73),
.B1(n_258),
.B2(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_66),
.B(n_127),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_66),
.A2(n_69),
.B1(n_299),
.B2(n_300),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_67),
.A2(n_70),
.B1(n_71),
.B2(n_72),
.Y(n_69)
);

CKINVDCx9p33_ASAP7_75t_R g72 ( 
.A(n_67),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_67),
.B(n_71),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_68),
.A2(n_70),
.B1(n_116),
.B2(n_117),
.Y(n_115)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_69),
.Y(n_73)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_70),
.Y(n_71)
);

NAND2x1_ASAP7_75t_SL g131 ( 
.A(n_70),
.B(n_132),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_71),
.B(n_157),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_73),
.B(n_112),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_73),
.A2(n_124),
.B(n_126),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_73),
.B(n_149),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_73),
.A2(n_126),
.B(n_221),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_74),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_75),
.A2(n_77),
.B1(n_78),
.B2(n_84),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_75),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_100),
.B(n_342),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_86),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_82),
.B(n_86),
.Y(n_342)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_83),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_92),
.C(n_95),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_87),
.A2(n_88),
.B1(n_92),
.B2(n_328),
.Y(n_334)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_91),
.B(n_92),
.C(n_96),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_92),
.A2(n_328),
.B1(n_329),
.B2(n_330),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_92),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_95),
.B(n_334),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

OAI321xp33_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_325),
.A3(n_335),
.B1(n_340),
.B2(n_341),
.C(n_345),
.Y(n_100)
);

AOI321xp33_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_275),
.A3(n_313),
.B1(n_319),
.B2(n_324),
.C(n_346),
.Y(n_101)
);

NOR3xp33_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_232),
.C(n_271),
.Y(n_102)
);

AOI21x1_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_202),
.B(n_231),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_105),
.A2(n_183),
.B(n_201),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_162),
.B(n_182),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_107),
.A2(n_137),
.B(n_161),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_118),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_108),
.B(n_118),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_109),
.B(n_114),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_109),
.A2(n_114),
.B1(n_115),
.B2(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_109),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_110),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_R g200 ( 
.A(n_111),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_112),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_128),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_121),
.B1(n_122),
.B2(n_123),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_120),
.B(n_123),
.C(n_128),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_129),
.A2(n_131),
.B(n_133),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_129),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_131),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_131),
.B(n_135),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_131),
.A2(n_132),
.B1(n_213),
.B2(n_214),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_131),
.A2(n_158),
.B1(n_214),
.B2(n_247),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_131),
.A2(n_151),
.B1(n_247),
.B2(n_256),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_131),
.A2(n_132),
.B(n_256),
.Y(n_288)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_132),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_136),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_136),
.A2(n_140),
.B1(n_142),
.B2(n_143),
.Y(n_139)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_136),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_136),
.A2(n_153),
.B(n_180),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_136),
.A2(n_142),
.B1(n_180),
.B2(n_195),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_146),
.B(n_160),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_144),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_139),
.B(n_144),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_141),
.A2(n_151),
.B(n_152),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_147),
.A2(n_154),
.B(n_159),
.Y(n_146)
);

NOR2x1_ASAP7_75t_R g147 ( 
.A(n_148),
.B(n_150),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_148),
.B(n_150),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_149),
.B(n_158),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_155),
.B(n_156),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_163),
.B(n_164),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_165),
.A2(n_166),
.B1(n_175),
.B2(n_181),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_169),
.B1(n_173),
.B2(n_174),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_167),
.Y(n_174)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_169),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_169),
.B(n_174),
.C(n_181),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_171),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_172),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_175),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_179),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_176),
.B(n_179),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_184),
.B(n_185),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_197),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_186),
.B(n_198),
.C(n_199),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_187),
.A2(n_188),
.B1(n_192),
.B2(n_196),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_187),
.B(n_193),
.C(n_194),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_192),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_194),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_195),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_203),
.B(n_204),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_218),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_215),
.B1(n_216),
.B2(n_217),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_206),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_206),
.B(n_217),
.C(n_218),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_208),
.B1(n_211),
.B2(n_212),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_207),
.B(n_212),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_208),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_212),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_215),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_226),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_220),
.A2(n_222),
.B1(n_223),
.B2(n_225),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_220),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_222),
.B(n_225),
.C(n_226),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_223),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

AOI21xp33_ASAP7_75t_L g320 ( 
.A1(n_233),
.A2(n_321),
.B(n_322),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_251),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_234),
.B(n_251),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_245),
.C(n_250),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_235),
.B(n_274),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_244),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_240),
.B1(n_241),
.B2(n_243),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_237),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_240),
.B(n_243),
.C(n_244),
.Y(n_269)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_245),
.B(n_250),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_248),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_246),
.B(n_248),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_252),
.A2(n_253),
.B1(n_269),
.B2(n_270),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_259),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_254),
.B(n_259),
.C(n_270),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_257),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_255),
.B(n_257),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_260),
.B(n_265),
.C(n_268),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_262),
.A2(n_265),
.B1(n_266),
.B2(n_268),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_262),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_264),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_266),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_269),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_272),
.B(n_273),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_293),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_276),
.B(n_293),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_286),
.C(n_292),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_277),
.A2(n_278),
.B1(n_286),
.B2(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_279),
.B(n_282),
.C(n_284),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_282),
.B1(n_284),
.B2(n_285),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_282),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_286),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_288),
.B1(n_289),
.B2(n_291),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_287),
.A2(n_288),
.B1(n_308),
.B2(n_309),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_287),
.A2(n_305),
.B(n_309),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_288),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_288),
.B(n_289),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_289),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_290),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_292),
.B(n_317),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_294),
.A2(n_295),
.B1(n_311),
.B2(n_312),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_296),
.A2(n_297),
.B1(n_303),
.B2(n_304),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_296),
.B(n_304),
.C(n_312),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_297),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_298),
.A2(n_301),
.B(n_302),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_298),
.B(n_301),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_302),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_302),
.A2(n_327),
.B1(n_331),
.B2(n_339),
.Y(n_338)
);

CKINVDCx16_ASAP7_75t_R g303 ( 
.A(n_304),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_305),
.A2(n_306),
.B1(n_307),
.B2(n_310),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_307),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_309),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_311),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_314),
.A2(n_320),
.B(n_323),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_315),
.B(n_316),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_333),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_326),
.B(n_333),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_331),
.C(n_332),
.Y(n_326)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_327),
.Y(n_339)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_332),
.B(n_338),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_337),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_336),
.B(n_337),
.Y(n_340)
);


endmodule