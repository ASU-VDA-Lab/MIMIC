module fake_netlist_5_1692_n_288 (n_29, n_16, n_43, n_0, n_12, n_9, n_36, n_25, n_18, n_27, n_42, n_22, n_1, n_8, n_10, n_24, n_28, n_21, n_40, n_34, n_38, n_4, n_32, n_35, n_41, n_11, n_17, n_19, n_7, n_37, n_15, n_26, n_30, n_20, n_5, n_33, n_14, n_2, n_31, n_23, n_13, n_3, n_6, n_39, n_288);

input n_29;
input n_16;
input n_43;
input n_0;
input n_12;
input n_9;
input n_36;
input n_25;
input n_18;
input n_27;
input n_42;
input n_22;
input n_1;
input n_8;
input n_10;
input n_24;
input n_28;
input n_21;
input n_40;
input n_34;
input n_38;
input n_4;
input n_32;
input n_35;
input n_41;
input n_11;
input n_17;
input n_19;
input n_7;
input n_37;
input n_15;
input n_26;
input n_30;
input n_20;
input n_5;
input n_33;
input n_14;
input n_2;
input n_31;
input n_23;
input n_13;
input n_3;
input n_6;
input n_39;

output n_288;

wire n_137;
wire n_210;
wire n_168;
wire n_260;
wire n_191;
wire n_164;
wire n_286;
wire n_91;
wire n_208;
wire n_122;
wire n_82;
wire n_194;
wire n_282;
wire n_142;
wire n_176;
wire n_214;
wire n_140;
wire n_248;
wire n_124;
wire n_86;
wire n_146;
wire n_136;
wire n_268;
wire n_182;
wire n_143;
wire n_83;
wire n_132;
wire n_61;
wire n_237;
wire n_90;
wire n_241;
wire n_127;
wire n_75;
wire n_101;
wire n_180;
wire n_184;
wire n_226;
wire n_235;
wire n_65;
wire n_78;
wire n_74;
wire n_144;
wire n_281;
wire n_207;
wire n_240;
wire n_114;
wire n_57;
wire n_96;
wire n_189;
wire n_220;
wire n_165;
wire n_111;
wire n_231;
wire n_108;
wire n_229;
wire n_257;
wire n_213;
wire n_129;
wire n_66;
wire n_98;
wire n_177;
wire n_60;
wire n_155;
wire n_152;
wire n_197;
wire n_107;
wire n_69;
wire n_58;
wire n_236;
wire n_116;
wire n_195;
wire n_227;
wire n_45;
wire n_117;
wire n_249;
wire n_271;
wire n_284;
wire n_46;
wire n_233;
wire n_94;
wire n_203;
wire n_245;
wire n_274;
wire n_205;
wire n_123;
wire n_113;
wire n_139;
wire n_105;
wire n_280;
wire n_246;
wire n_80;
wire n_179;
wire n_125;
wire n_269;
wire n_167;
wire n_128;
wire n_73;
wire n_234;
wire n_277;
wire n_92;
wire n_267;
wire n_149;
wire n_120;
wire n_285;
wire n_232;
wire n_135;
wire n_156;
wire n_126;
wire n_254;
wire n_225;
wire n_84;
wire n_202;
wire n_130;
wire n_266;
wire n_272;
wire n_219;
wire n_258;
wire n_157;
wire n_265;
wire n_79;
wire n_193;
wire n_131;
wire n_151;
wire n_47;
wire n_173;
wire n_192;
wire n_251;
wire n_244;
wire n_53;
wire n_160;
wire n_198;
wire n_223;
wire n_247;
wire n_188;
wire n_190;
wire n_201;
wire n_158;
wire n_263;
wire n_44;
wire n_224;
wire n_154;
wire n_100;
wire n_62;
wire n_138;
wire n_148;
wire n_71;
wire n_228;
wire n_264;
wire n_283;
wire n_109;
wire n_112;
wire n_212;
wire n_85;
wire n_159;
wire n_163;
wire n_276;
wire n_95;
wire n_119;
wire n_183;
wire n_185;
wire n_243;
wire n_239;
wire n_275;
wire n_175;
wire n_252;
wire n_169;
wire n_59;
wire n_262;
wire n_255;
wire n_133;
wire n_238;
wire n_215;
wire n_55;
wire n_196;
wire n_99;
wire n_211;
wire n_218;
wire n_181;
wire n_49;
wire n_54;
wire n_178;
wire n_147;
wire n_221;
wire n_67;
wire n_121;
wire n_242;
wire n_76;
wire n_200;
wire n_87;
wire n_150;
wire n_170;
wire n_162;
wire n_64;
wire n_102;
wire n_77;
wire n_106;
wire n_209;
wire n_161;
wire n_259;
wire n_273;
wire n_287;
wire n_270;
wire n_222;
wire n_230;
wire n_81;
wire n_118;
wire n_89;
wire n_279;
wire n_70;
wire n_115;
wire n_68;
wire n_93;
wire n_261;
wire n_253;
wire n_72;
wire n_186;
wire n_174;
wire n_199;
wire n_134;
wire n_187;
wire n_104;
wire n_172;
wire n_103;
wire n_56;
wire n_51;
wire n_63;
wire n_97;
wire n_166;
wire n_141;
wire n_206;
wire n_217;
wire n_171;
wire n_153;
wire n_145;
wire n_256;
wire n_48;
wire n_204;
wire n_50;
wire n_250;
wire n_52;
wire n_278;
wire n_88;
wire n_110;
wire n_216;

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_13),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_19),
.Y(n_45)
);

CKINVDCx5p33_ASAP7_75t_R g46 ( 
.A(n_23),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

INVxp33_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVxp67_ASAP7_75t_SL g54 ( 
.A(n_39),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_8),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

CKINVDCx14_ASAP7_75t_R g59 ( 
.A(n_1),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_15),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_10),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_14),
.Y(n_65)
);

INVxp67_ASAP7_75t_SL g66 ( 
.A(n_6),
.Y(n_66)
);

BUFx2_ASAP7_75t_SL g67 ( 
.A(n_35),
.Y(n_67)
);

CKINVDCx5p33_ASAP7_75t_R g68 ( 
.A(n_24),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_0),
.Y(n_69)
);

CKINVDCx5p33_ASAP7_75t_R g70 ( 
.A(n_30),
.Y(n_70)
);

CKINVDCx5p33_ASAP7_75t_R g71 ( 
.A(n_11),
.Y(n_71)
);

BUFx2_ASAP7_75t_SL g72 ( 
.A(n_16),
.Y(n_72)
);

INVxp33_ASAP7_75t_SL g73 ( 
.A(n_38),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_18),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_29),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_44),
.B(n_45),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

BUFx8_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_51),
.B(n_0),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_51),
.B(n_1),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_59),
.B(n_2),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_46),
.B(n_2),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_57),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_58),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_46),
.B(n_3),
.Y(n_97)
);

AND2x4_ASAP7_75t_L g98 ( 
.A(n_60),
.B(n_3),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_62),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_63),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_64),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_76),
.B(n_68),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_83),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_79),
.B(n_73),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g106 ( 
.A(n_87),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

INVx2_ASAP7_75t_SL g108 ( 
.A(n_76),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_78),
.B(n_71),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_70),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_79),
.B(n_73),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_91),
.B(n_54),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_91),
.B(n_70),
.Y(n_113)
);

NOR3xp33_ASAP7_75t_L g114 ( 
.A(n_84),
.B(n_74),
.C(n_61),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_93),
.B(n_72),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_90),
.B(n_74),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_67),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_61),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_102),
.Y(n_119)
);

BUFx5_ASAP7_75t_L g120 ( 
.A(n_101),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_85),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_102),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_77),
.Y(n_123)
);

A2O1A1Ixp33_ASAP7_75t_L g124 ( 
.A1(n_85),
.A2(n_4),
.B(n_5),
.C(n_7),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_80),
.Y(n_125)
);

BUFx2_ASAP7_75t_L g126 ( 
.A(n_108),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_109),
.B(n_98),
.Y(n_127)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_104),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_103),
.B(n_98),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_125),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_107),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_123),
.Y(n_132)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_113),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_119),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_120),
.B(n_88),
.Y(n_135)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_122),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_115),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_105),
.B(n_84),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_106),
.Y(n_139)
);

AND2x4_ASAP7_75t_L g140 ( 
.A(n_124),
.B(n_80),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_120),
.B(n_106),
.Y(n_141)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_106),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_120),
.B(n_100),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_110),
.B(n_97),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_117),
.Y(n_145)
);

INVx1_ASAP7_75t_SL g146 ( 
.A(n_126),
.Y(n_146)
);

OA21x2_ASAP7_75t_L g147 ( 
.A1(n_135),
.A2(n_112),
.B(n_82),
.Y(n_147)
);

OR2x6_ASAP7_75t_L g148 ( 
.A(n_138),
.B(n_111),
.Y(n_148)
);

AND2x4_ASAP7_75t_L g149 ( 
.A(n_140),
.B(n_114),
.Y(n_149)
);

INVx2_ASAP7_75t_SL g150 ( 
.A(n_144),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_130),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_129),
.A2(n_116),
.B(n_118),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_138),
.A2(n_121),
.B1(n_82),
.B2(n_96),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_131),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_137),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_130),
.Y(n_156)
);

NAND2x1_ASAP7_75t_L g157 ( 
.A(n_142),
.B(n_99),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_131),
.Y(n_158)
);

BUFx12f_ASAP7_75t_L g159 ( 
.A(n_137),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_134),
.Y(n_160)
);

NOR2xp67_ASAP7_75t_SL g161 ( 
.A(n_133),
.B(n_94),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_133),
.B(n_86),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_137),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_127),
.B(n_106),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_134),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_137),
.B(n_120),
.Y(n_166)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_151),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_151),
.Y(n_168)
);

OAI21x1_ASAP7_75t_L g169 ( 
.A1(n_166),
.A2(n_141),
.B(n_143),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_159),
.Y(n_170)
);

HB1xp67_ASAP7_75t_L g171 ( 
.A(n_146),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_148),
.A2(n_81),
.B1(n_133),
.B2(n_145),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_156),
.Y(n_173)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_156),
.Y(n_174)
);

OR2x2_ASAP7_75t_L g175 ( 
.A(n_150),
.B(n_145),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_160),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_160),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_154),
.Y(n_178)
);

O2A1O1Ixp33_ASAP7_75t_L g179 ( 
.A1(n_150),
.A2(n_140),
.B(n_136),
.C(n_132),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_163),
.A2(n_145),
.B1(n_140),
.B2(n_139),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_159),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_158),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_165),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_155),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_168),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_175),
.B(n_149),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_168),
.Y(n_187)
);

BUFx2_ASAP7_75t_L g188 ( 
.A(n_171),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_173),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_176),
.Y(n_190)
);

INVxp67_ASAP7_75t_SL g191 ( 
.A(n_175),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_178),
.B(n_149),
.Y(n_192)
);

OR2x2_ASAP7_75t_L g193 ( 
.A(n_184),
.B(n_149),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_177),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g195 ( 
.A(n_170),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_183),
.A2(n_148),
.B1(n_152),
.B2(n_182),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_177),
.Y(n_197)
);

BUFx2_ASAP7_75t_L g198 ( 
.A(n_170),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_167),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_178),
.B(n_148),
.Y(n_200)
);

OR2x2_ASAP7_75t_L g201 ( 
.A(n_181),
.B(n_148),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_182),
.Y(n_202)
);

OAI21x1_ASAP7_75t_L g203 ( 
.A1(n_196),
.A2(n_169),
.B(n_179),
.Y(n_203)
);

NOR4xp75_ASAP7_75t_L g204 ( 
.A(n_200),
.B(n_180),
.C(n_172),
.D(n_81),
.Y(n_204)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_188),
.Y(n_205)
);

OR2x2_ASAP7_75t_L g206 ( 
.A(n_191),
.B(n_186),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_192),
.A2(n_153),
.B1(n_183),
.B2(n_164),
.Y(n_207)
);

INVx2_ASAP7_75t_SL g208 ( 
.A(n_193),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_202),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_189),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_190),
.Y(n_211)
);

AOI211xp5_ASAP7_75t_L g212 ( 
.A1(n_201),
.A2(n_162),
.B(n_136),
.C(n_153),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_185),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_186),
.B(n_192),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_185),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_200),
.B(n_174),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_187),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_194),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_198),
.Y(n_219)
);

BUFx2_ASAP7_75t_L g220 ( 
.A(n_195),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_210),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_208),
.B(n_193),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g223 ( 
.A(n_220),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_211),
.Y(n_224)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_205),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_208),
.B(n_196),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_209),
.Y(n_227)
);

NAND2x1p5_ASAP7_75t_L g228 ( 
.A(n_206),
.B(n_199),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_219),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_214),
.B(n_199),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_216),
.B(n_197),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_213),
.Y(n_232)
);

AOI211xp5_ASAP7_75t_SL g233 ( 
.A1(n_212),
.A2(n_174),
.B(n_167),
.C(n_187),
.Y(n_233)
);

INVxp33_ASAP7_75t_L g234 ( 
.A(n_216),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_218),
.B(n_217),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_232),
.Y(n_236)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_228),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_234),
.B(n_217),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_222),
.B(n_215),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_225),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_226),
.B(n_207),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_235),
.B(n_213),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_230),
.B(n_223),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_227),
.B(n_215),
.Y(n_244)
);

NAND4xp75_ASAP7_75t_L g245 ( 
.A(n_231),
.B(n_204),
.C(n_147),
.D(n_17),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_229),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_230),
.B(n_207),
.Y(n_247)
);

OR2x4_ASAP7_75t_L g248 ( 
.A(n_231),
.B(n_161),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_221),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_229),
.B(n_128),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_224),
.Y(n_251)
);

AND2x4_ASAP7_75t_L g252 ( 
.A(n_237),
.B(n_203),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_240),
.B(n_128),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_246),
.B(n_9),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_243),
.B(n_233),
.Y(n_255)
);

NAND2x1p5_ASAP7_75t_L g256 ( 
.A(n_237),
.B(n_203),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_238),
.B(n_147),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_250),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_247),
.B(n_174),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_249),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_249),
.Y(n_261)
);

OAI31xp33_ASAP7_75t_SL g262 ( 
.A1(n_254),
.A2(n_241),
.A3(n_251),
.B(n_245),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_260),
.Y(n_263)
);

OAI211xp5_ASAP7_75t_L g264 ( 
.A1(n_258),
.A2(n_241),
.B(n_246),
.C(n_239),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_261),
.Y(n_265)
);

NAND4xp25_ASAP7_75t_L g266 ( 
.A(n_253),
.B(n_242),
.C(n_244),
.D(n_237),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_255),
.B(n_248),
.Y(n_267)
);

AND2x4_ASAP7_75t_L g268 ( 
.A(n_263),
.B(n_252),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_265),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_267),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_266),
.Y(n_271)
);

OA211x2_ASAP7_75t_L g272 ( 
.A1(n_270),
.A2(n_262),
.B(n_259),
.C(n_257),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_269),
.Y(n_273)
);

NAND4xp75_ASAP7_75t_L g274 ( 
.A(n_271),
.B(n_244),
.C(n_242),
.D(n_264),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_274),
.B(n_268),
.Y(n_275)
);

AOI211xp5_ASAP7_75t_SL g276 ( 
.A1(n_272),
.A2(n_268),
.B(n_252),
.C(n_236),
.Y(n_276)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_273),
.Y(n_277)
);

NOR2x1p5_ASAP7_75t_L g278 ( 
.A(n_277),
.B(n_167),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_275),
.B(n_256),
.Y(n_279)
);

NOR2x1p5_ASAP7_75t_L g280 ( 
.A(n_276),
.B(n_157),
.Y(n_280)
);

BUFx2_ASAP7_75t_L g281 ( 
.A(n_278),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_279),
.B(n_26),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_280),
.B(n_27),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_283),
.A2(n_169),
.B(n_36),
.Y(n_284)
);

OAI21xp33_ASAP7_75t_L g285 ( 
.A1(n_282),
.A2(n_40),
.B(n_43),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_281),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_286),
.Y(n_287)
);

OAI22x1_ASAP7_75t_L g288 ( 
.A1(n_287),
.A2(n_284),
.B1(n_285),
.B2(n_142),
.Y(n_288)
);


endmodule