module fake_jpeg_26664_n_102 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_102);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_102;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_8),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_0),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

INVx11_ASAP7_75t_SL g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_20),
.B(n_13),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_23),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_20),
.B(n_13),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

OR2x2_ASAP7_75t_L g26 ( 
.A(n_20),
.B(n_11),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_29),
.Y(n_35)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_27),
.B(n_28),
.Y(n_39)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_27),
.A2(n_15),
.B1(n_21),
.B2(n_17),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_31),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_26),
.A2(n_21),
.B1(n_14),
.B2(n_17),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_22),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_33),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_27),
.A2(n_19),
.B1(n_16),
.B2(n_12),
.Y(n_33)
);

XOR2xp5_ASAP7_75t_L g37 ( 
.A(n_23),
.B(n_14),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_19),
.C(n_16),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_31),
.C(n_26),
.Y(n_53)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

A2O1A1O1Ixp25_ASAP7_75t_L g43 ( 
.A1(n_37),
.A2(n_26),
.B(n_25),
.C(n_24),
.D(n_29),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_44),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_33),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_34),
.B(n_12),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_46),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_34),
.B(n_7),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_9),
.Y(n_48)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_48),
.B(n_49),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_32),
.B(n_9),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_35),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_51),
.B(n_52),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_35),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_55),
.Y(n_63)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_30),
.Y(n_56)
);

XOR2xp5_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_39),
.Y(n_70)
);

BUFx24_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_59),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_SL g60 ( 
.A1(n_41),
.A2(n_39),
.B(n_25),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_54),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_65),
.Y(n_71)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_64),
.B(n_67),
.Y(n_75)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_70),
.B(n_53),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_68),
.A2(n_56),
.B1(n_57),
.B2(n_52),
.Y(n_73)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

OA21x2_ASAP7_75t_SL g74 ( 
.A1(n_70),
.A2(n_59),
.B(n_60),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_74),
.A2(n_77),
.B(n_50),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_76),
.B(n_62),
.C(n_25),
.Y(n_84)
);

AOI322xp5_ASAP7_75t_SL g77 ( 
.A1(n_69),
.A2(n_50),
.A3(n_58),
.B1(n_59),
.B2(n_6),
.C1(n_4),
.C2(n_5),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_50),
.Y(n_79)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_79),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_81),
.B(n_82),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_76),
.B(n_74),
.C(n_79),
.Y(n_82)
);

A2O1A1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_75),
.A2(n_62),
.B(n_59),
.C(n_64),
.Y(n_83)
);

OAI221xp5_ASAP7_75t_L g90 ( 
.A1(n_83),
.A2(n_71),
.B1(n_78),
.B2(n_11),
.C(n_29),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_84),
.B(n_78),
.Y(n_91)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_80),
.Y(n_87)
);

NOR2xp67_ASAP7_75t_SL g95 ( 
.A(n_87),
.B(n_0),
.Y(n_95)
);

OAI21x1_ASAP7_75t_L g88 ( 
.A1(n_83),
.A2(n_72),
.B(n_75),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_88),
.A2(n_90),
.B1(n_28),
.B2(n_36),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_91),
.B(n_86),
.C(n_85),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_92),
.B(n_93),
.Y(n_98)
);

MAJx2_ASAP7_75t_L g94 ( 
.A(n_89),
.B(n_82),
.C(n_24),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_94),
.B(n_87),
.C(n_38),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_95),
.B(n_0),
.Y(n_97)
);

AOI322xp5_ASAP7_75t_L g99 ( 
.A1(n_96),
.A2(n_97),
.A3(n_28),
.B1(n_2),
.B2(n_3),
.C1(n_4),
.C2(n_5),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_99),
.B(n_100),
.C(n_36),
.Y(n_101)
);

AOI322xp5_ASAP7_75t_L g100 ( 
.A1(n_98),
.A2(n_29),
.A3(n_36),
.B1(n_4),
.B2(n_5),
.C1(n_1),
.C2(n_2),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_1),
.Y(n_102)
);


endmodule