module fake_jpeg_15837_n_56 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_56);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_56;

wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_47;
wire n_22;
wire n_51;
wire n_40;
wire n_19;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_36;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_8),
.B(n_12),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_7),
.B(n_9),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_15),
.B(n_16),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_18),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_23),
.Y(n_28)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_26),
.B(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_SL g35 ( 
.A1(n_31),
.A2(n_26),
.B(n_24),
.Y(n_35)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_L g45 ( 
.A1(n_35),
.A2(n_25),
.B(n_39),
.Y(n_45)
);

OA21x2_ASAP7_75t_L g39 ( 
.A1(n_27),
.A2(n_22),
.B(n_1),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_39),
.A2(n_22),
.B1(n_1),
.B2(n_2),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_44),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_31),
.Y(n_41)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_43),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_33),
.B(n_38),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_21),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g49 ( 
.A(n_45),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_47),
.A2(n_0),
.B(n_3),
.Y(n_52)
);

A2O1A1Ixp33_ASAP7_75t_SL g51 ( 
.A1(n_46),
.A2(n_36),
.B(n_3),
.C(n_4),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_SL g53 ( 
.A1(n_51),
.A2(n_52),
.B(n_46),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_53),
.A2(n_49),
.B1(n_48),
.B2(n_50),
.Y(n_54)
);

A2O1A1Ixp33_ASAP7_75t_L g55 ( 
.A1(n_54),
.A2(n_4),
.B(n_6),
.C(n_10),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_55),
.B(n_11),
.C(n_14),
.Y(n_56)
);


endmodule