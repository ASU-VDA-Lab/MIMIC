module fake_jpeg_6829_n_104 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_104);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_104;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_6),
.Y(n_11)
);

INVxp67_ASAP7_75t_L g12 ( 
.A(n_9),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_10),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_13),
.B(n_1),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_24),
.B(n_25),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_17),
.B(n_2),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_22),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_27),
.A2(n_19),
.B1(n_17),
.B2(n_13),
.Y(n_38)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_29),
.B(n_30),
.Y(n_46)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_30),
.A2(n_22),
.B1(n_23),
.B2(n_14),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_34),
.A2(n_38),
.B1(n_43),
.B2(n_45),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_25),
.B(n_19),
.Y(n_37)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_30),
.A2(n_11),
.B1(n_15),
.B2(n_14),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_29),
.A2(n_28),
.B1(n_27),
.B2(n_15),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_29),
.A2(n_11),
.B1(n_12),
.B2(n_18),
.Y(n_45)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_46),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_54),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_26),
.C(n_24),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_61),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_46),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_50),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_25),
.Y(n_51)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_32),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_53),
.Y(n_62)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_32),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_26),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_56),
.B(n_59),
.Y(n_67)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_58),
.Y(n_65)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_26),
.Y(n_59)
);

MAJx2_ASAP7_75t_L g61 ( 
.A(n_35),
.B(n_12),
.C(n_21),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_40),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_68),
.B(n_72),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g70 ( 
.A(n_49),
.B(n_35),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_61),
.C(n_21),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_55),
.A2(n_44),
.B1(n_33),
.B2(n_31),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_71),
.A2(n_57),
.B1(n_60),
.B2(n_50),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_36),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_73),
.A2(n_78),
.B1(n_80),
.B2(n_63),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_69),
.B(n_48),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_74),
.B(n_77),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_71),
.A2(n_55),
.B1(n_60),
.B2(n_47),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_72),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_65),
.A2(n_47),
.B1(n_44),
.B2(n_52),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_79),
.B(n_81),
.C(n_67),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_66),
.A2(n_33),
.B1(n_31),
.B2(n_40),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_64),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_78),
.A2(n_62),
.B(n_66),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_83),
.B(n_84),
.Y(n_92)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_85),
.Y(n_90)
);

AOI21x1_ASAP7_75t_SL g87 ( 
.A1(n_73),
.A2(n_70),
.B(n_21),
.Y(n_87)
);

A2O1A1O1Ixp25_ASAP7_75t_L g89 ( 
.A1(n_87),
.A2(n_80),
.B(n_75),
.C(n_77),
.D(n_76),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_82),
.B(n_79),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_8),
.Y(n_95)
);

OAI21x1_ASAP7_75t_SL g93 ( 
.A1(n_89),
.A2(n_82),
.B(n_7),
.Y(n_93)
);

AO221x1_ASAP7_75t_L g91 ( 
.A1(n_86),
.A2(n_40),
.B1(n_3),
.B2(n_5),
.C(n_2),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_91),
.B(n_3),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_93),
.B(n_89),
.C(n_7),
.Y(n_99)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_94),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_95),
.B(n_96),
.C(n_88),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_90),
.B(n_5),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_97),
.B(n_99),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_98),
.A2(n_92),
.B(n_95),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_101),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_102),
.A2(n_100),
.B(n_8),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_5),
.Y(n_104)
);


endmodule