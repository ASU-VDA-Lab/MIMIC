module fake_netlist_1_12303_n_12 (n_1, n_2, n_0, n_12);
input n_1;
input n_2;
input n_0;
output n_12;
wire n_11;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_8;
wire n_10;
wire n_7;
INVx3_ASAP7_75t_L g3 ( .A(n_0), .Y(n_3) );
INVx1_ASAP7_75t_L g4 ( .A(n_0), .Y(n_4) );
OAI21x1_ASAP7_75t_L g5 ( .A1(n_3), .A2(n_0), .B(n_1), .Y(n_5) );
AOI22xp33_ASAP7_75t_SL g6 ( .A1(n_4), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_6) );
NOR2x1p5_ASAP7_75t_L g7 ( .A(n_6), .B(n_4), .Y(n_7) );
INVxp67_ASAP7_75t_SL g8 ( .A(n_5), .Y(n_8) );
INVx2_ASAP7_75t_L g9 ( .A(n_8), .Y(n_9) );
AOI22xp5_ASAP7_75t_L g10 ( .A1(n_9), .A2(n_7), .B1(n_4), .B2(n_3), .Y(n_10) );
NOR4xp25_ASAP7_75t_SL g11 ( .A(n_10), .B(n_7), .C(n_5), .D(n_1), .Y(n_11) );
OAI22xp5_ASAP7_75t_L g12 ( .A1(n_11), .A2(n_2), .B1(n_3), .B2(n_9), .Y(n_12) );
endmodule