module real_jpeg_4930_n_7 (n_5, n_4, n_0, n_1, n_51, n_2, n_48, n_6, n_50, n_53, n_3, n_49, n_52, n_7);

input n_5;
input n_4;
input n_0;
input n_1;
input n_51;
input n_2;
input n_48;
input n_6;
input n_50;
input n_53;
input n_3;
input n_49;
input n_52;

output n_7;

wire n_17;
wire n_8;
wire n_43;
wire n_37;
wire n_21;
wire n_33;
wire n_35;
wire n_38;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_44;
wire n_28;
wire n_46;
wire n_23;
wire n_11;
wire n_14;
wire n_45;
wire n_25;
wire n_42;
wire n_22;
wire n_18;
wire n_40;
wire n_39;
wire n_36;
wire n_41;
wire n_26;
wire n_27;
wire n_20;
wire n_19;
wire n_32;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

INVx5_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

OR2x2_ASAP7_75t_L g36 ( 
.A(n_0),
.B(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g10 ( 
.A(n_1),
.B(n_11),
.Y(n_10)
);

AND2x2_ASAP7_75t_L g16 ( 
.A(n_1),
.B(n_11),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_2),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_3),
.B(n_33),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g18 ( 
.A(n_4),
.B(n_19),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_4),
.B(n_19),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_5),
.B(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_5),
.B(n_41),
.Y(n_43)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

XOR2xp5_ASAP7_75t_L g7 ( 
.A(n_8),
.B(n_17),
.Y(n_7)
);

NAND2xp5_ASAP7_75t_SL g8 ( 
.A(n_9),
.B(n_15),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_10),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_13),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_13),
.B(n_34),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_13),
.B(n_42),
.Y(n_41)
);

INVx11_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

CKINVDCx14_ASAP7_75t_R g15 ( 
.A(n_16),
.Y(n_15)
);

OAI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_23),
.B(n_45),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_21),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

AO21x1_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_30),
.B(n_44),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_29),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_26),
.B(n_29),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_28),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_SL g30 ( 
.A1(n_31),
.A2(n_40),
.B(n_43),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_35),
.B(n_39),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_36),
.B(n_38),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_36),
.B(n_38),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_48),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_49),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_50),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_51),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_52),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_53),
.Y(n_42)
);


endmodule