module fake_jpeg_13598_n_181 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_181);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_181;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_9),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_23),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_7),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_46),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

BUFx10_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_12),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_0),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_49),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_39),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_31),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_15),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_29),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_10),
.Y(n_71)
);

CKINVDCx5p33_ASAP7_75t_R g72 ( 
.A(n_3),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_8),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_11),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_26),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_18),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_36),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_16),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_56),
.B(n_0),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_81),
.B(n_82),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_1),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_78),
.Y(n_83)
);

INVx2_ASAP7_75t_SL g100 ( 
.A(n_83),
.Y(n_100)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_78),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_57),
.B(n_1),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_2),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_L g87 ( 
.A1(n_57),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_87),
.A2(n_58),
.B1(n_60),
.B2(n_74),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

CKINVDCx9p33_ASAP7_75t_R g89 ( 
.A(n_72),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_89),
.Y(n_104)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_90),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_84),
.B(n_75),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_98),
.Y(n_107)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_88),
.Y(n_92)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_92),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_93),
.A2(n_77),
.B1(n_80),
.B2(n_71),
.Y(n_118)
);

BUFx10_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_94),
.Y(n_108)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_96),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_82),
.B(n_75),
.Y(n_98)
);

AND2x4_ASAP7_75t_L g99 ( 
.A(n_90),
.B(n_60),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_99),
.B(n_4),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_101),
.B(n_35),
.Y(n_124)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_102),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_98),
.B(n_69),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_105),
.B(n_124),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_91),
.A2(n_79),
.B1(n_63),
.B2(n_55),
.Y(n_109)
);

OA21x2_ASAP7_75t_L g130 ( 
.A1(n_109),
.A2(n_5),
.B(n_6),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_94),
.A2(n_76),
.B1(n_64),
.B2(n_62),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_111),
.Y(n_139)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_112),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_103),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_113),
.B(n_121),
.Y(n_137)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_104),
.Y(n_114)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_114),
.Y(n_131)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_100),
.Y(n_115)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_115),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_99),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_116),
.B(n_117),
.Y(n_125)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_97),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_118),
.A2(n_119),
.B1(n_66),
.B2(n_61),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_93),
.A2(n_69),
.B1(n_73),
.B2(n_70),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_103),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_122),
.B(n_5),
.Y(n_138)
);

INVx11_ASAP7_75t_L g123 ( 
.A(n_94),
.Y(n_123)
);

INVxp33_ASAP7_75t_L g134 ( 
.A(n_123),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_120),
.B(n_68),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_127),
.B(n_128),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_107),
.B(n_67),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_110),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_133),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_106),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_135),
.B(n_138),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_116),
.B(n_6),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_140),
.B(n_142),
.Y(n_157)
);

OAI32xp33_ASAP7_75t_L g141 ( 
.A1(n_111),
.A2(n_7),
.A3(n_13),
.B1(n_14),
.B2(n_20),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_141),
.B(n_143),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_108),
.B(n_114),
.Y(n_142)
);

A2O1A1Ixp33_ASAP7_75t_L g143 ( 
.A1(n_107),
.A2(n_52),
.B(n_22),
.C(n_25),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_137),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_145),
.B(n_147),
.Y(n_166)
);

INVx13_ASAP7_75t_L g146 ( 
.A(n_136),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_146),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_126),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_125),
.A2(n_21),
.B1(n_28),
.B2(n_30),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_148),
.A2(n_40),
.B1(n_42),
.B2(n_43),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_139),
.A2(n_129),
.B(n_134),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_149),
.A2(n_155),
.B(n_158),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_131),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_150),
.B(n_151),
.Y(n_164)
);

AND2x6_ASAP7_75t_L g151 ( 
.A(n_143),
.B(n_130),
.Y(n_151)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_134),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_139),
.B(n_32),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_156),
.B(n_47),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_137),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_144),
.A2(n_33),
.B(n_34),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_159),
.B(n_162),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_163),
.B(n_153),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_152),
.A2(n_48),
.B1(n_50),
.B2(n_51),
.Y(n_165)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_165),
.Y(n_167)
);

FAx1_ASAP7_75t_SL g168 ( 
.A(n_161),
.B(n_157),
.CI(n_151),
.CON(n_168),
.SN(n_168)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_168),
.B(n_169),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_170),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_172),
.B(n_173),
.Y(n_174)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_167),
.Y(n_173)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_174),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_175),
.B(n_154),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_176),
.B(n_166),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_160),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_178),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_179),
.A2(n_171),
.B(n_164),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_180),
.B(n_168),
.Y(n_181)
);


endmodule