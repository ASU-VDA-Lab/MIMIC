module real_jpeg_17876_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_0),
.A2(n_4),
.B1(n_20),
.B2(n_22),
.Y(n_19)
);

INVx2_ASAP7_75t_SL g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_1),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_1),
.Y(n_121)
);

BUFx5_ASAP7_75t_L g153 ( 
.A(n_1),
.Y(n_153)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_1),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_2),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_3),
.Y(n_38)
);

AND2x4_ASAP7_75t_SL g60 ( 
.A(n_3),
.B(n_61),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_3),
.B(n_71),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_3),
.B(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_3),
.B(n_144),
.Y(n_143)
);

AND2x2_ASAP7_75t_SL g170 ( 
.A(n_3),
.B(n_171),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_3),
.B(n_201),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_3),
.B(n_151),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_5),
.B(n_147),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_5),
.A2(n_11),
.B1(n_156),
.B2(n_159),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_5),
.B(n_61),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_5),
.Y(n_196)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_6),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_6),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_6),
.Y(n_87)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_6),
.Y(n_255)
);

BUFx5_ASAP7_75t_L g287 ( 
.A(n_6),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_7),
.B(n_31),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_7),
.B(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_7),
.B(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_7),
.B(n_133),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_7),
.B(n_263),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_7),
.B(n_268),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_7),
.B(n_284),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_8),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_8),
.B(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_8),
.B(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_8),
.B(n_135),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_8),
.B(n_204),
.Y(n_203)
);

BUFx4f_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_9),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g149 ( 
.A(n_9),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_10),
.B(n_123),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_10),
.B(n_151),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_11),
.B(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_11),
.B(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_11),
.B(n_112),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_11),
.B(n_190),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_11),
.B(n_230),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_11),
.B(n_253),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_11),
.B(n_259),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_11),
.B(n_294),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_12),
.B(n_42),
.Y(n_41)
);

AND2x2_ASAP7_75t_SL g53 ( 
.A(n_12),
.B(n_54),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_12),
.B(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_12),
.B(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_13),
.B(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_13),
.B(n_207),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_13),
.B(n_171),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_13),
.B(n_249),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_13),
.B(n_304),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_13),
.B(n_308),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_13),
.B(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_14),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_15),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_15),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_15),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_16),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_16),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_17),
.B(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_18),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g116 ( 
.A(n_18),
.Y(n_116)
);

BUFx5_ASAP7_75t_L g144 ( 
.A(n_18),
.Y(n_144)
);

BUFx12f_ASAP7_75t_SL g20 ( 
.A(n_21),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_214),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_179),
.B(n_212),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_25),
.B(n_180),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_106),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_67),
.C(n_90),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_SL g181 ( 
.A(n_27),
.B(n_182),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_47),
.C(n_55),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

XNOR2x2_ASAP7_75t_L g235 ( 
.A(n_29),
.B(n_236),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_36),
.Y(n_29)
);

MAJx2_ASAP7_75t_L g164 ( 
.A(n_30),
.B(n_41),
.C(n_46),
.Y(n_164)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_34),
.Y(n_251)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_41),
.B1(n_45),
.B2(n_46),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_37),
.Y(n_46)
);

OR2x2_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_39),
.Y(n_37)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_39),
.Y(n_133)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_40),
.Y(n_208)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_44),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_47),
.B(n_56),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_53),
.Y(n_47)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_48),
.B(n_53),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_50),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_51),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_52),
.Y(n_319)
);

BUFx12f_ASAP7_75t_L g204 ( 
.A(n_54),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_60),
.C(n_62),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_57),
.A2(n_60),
.B1(n_224),
.B2(n_225),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_57),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_60),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_60),
.A2(n_225),
.B1(n_302),
.B2(n_303),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_60),
.B(n_298),
.C(n_302),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_62),
.B(n_223),
.Y(n_222)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_65),
.Y(n_304)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_68),
.B(n_90),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_80),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_73),
.C(n_77),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_70),
.B(n_73),
.C(n_77),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_70),
.A2(n_77),
.B1(n_186),
.B2(n_187),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_70),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_70),
.B(n_247),
.Y(n_246)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_73),
.B(n_185),
.Y(n_184)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_77),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_86),
.B1(n_88),
.B2(n_89),
.Y(n_80)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_81),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_81),
.B(n_88),
.C(n_176),
.Y(n_175)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_84),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_85),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_86),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_95),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_96),
.C(n_104),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_100),
.B1(n_104),
.B2(n_105),
.Y(n_95)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_96),
.Y(n_105)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_101),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_101),
.A2(n_104),
.B1(n_228),
.B2(n_278),
.Y(n_277)
);

BUFx5_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_103),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_104),
.B(n_228),
.C(n_229),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_107),
.A2(n_138),
.B1(n_177),
.B2(n_178),
.Y(n_106)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_107),
.Y(n_177)
);

XOR2x2_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_126),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_110),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_117),
.Y(n_110)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_122),
.Y(n_117)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVxp67_ASAP7_75t_SL g126 ( 
.A(n_127),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_131),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_134),
.Y(n_131)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_138),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_165),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_154),
.C(n_164),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_140),
.B(n_210),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_145),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_143),
.B(n_146),
.C(n_150),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_150),
.Y(n_145)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_149),
.Y(n_269)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_154),
.A2(n_155),
.B1(n_164),
.B2(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_155),
.A2(n_189),
.B(n_195),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx6_ASAP7_75t_L g197 ( 
.A(n_157),
.Y(n_197)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_158),
.Y(n_265)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_164),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_175),
.Y(n_165)
);

XNOR2x1_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_170),
.B1(n_173),
.B2(n_174),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_169),
.A2(n_170),
.B1(n_205),
.B2(n_206),
.Y(n_335)
);

INVx2_ASAP7_75t_SL g169 ( 
.A(n_170),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_170),
.B(n_199),
.C(n_205),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_183),
.C(n_209),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_181),
.B(n_238),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_183),
.B(n_209),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_188),
.C(n_198),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_184),
.B(n_188),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_186),
.B(n_248),
.C(n_252),
.Y(n_275)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_198),
.B(n_219),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g334 ( 
.A(n_199),
.B(n_335),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_203),
.Y(n_199)
);

XNOR2x1_ASAP7_75t_SL g282 ( 
.A(n_200),
.B(n_203),
.Y(n_282)
);

INVxp67_ASAP7_75t_SL g292 ( 
.A(n_200),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_SL g312 ( 
.A1(n_200),
.A2(n_292),
.B1(n_293),
.B2(n_313),
.Y(n_312)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_239),
.B(n_349),
.Y(n_214)
);

INVxp33_ASAP7_75t_SL g215 ( 
.A(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_237),
.Y(n_216)
);

NOR2xp67_ASAP7_75t_SL g351 ( 
.A(n_217),
.B(n_237),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_220),
.C(n_235),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_218),
.B(n_347),
.Y(n_346)
);

HB1xp67_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_221),
.B(n_235),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_226),
.C(n_233),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_222),
.B(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_227),
.B(n_234),
.Y(n_340)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_228),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_SL g276 ( 
.A(n_229),
.B(n_277),
.Y(n_276)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx5_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_242),
.A2(n_344),
.B(n_348),
.Y(n_241)
);

AOI21x1_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_329),
.B(n_343),
.Y(n_242)
);

OAI21x1_ASAP7_75t_SL g243 ( 
.A1(n_244),
.A2(n_288),
.B(n_328),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_273),
.Y(n_244)
);

OR2x2_ASAP7_75t_L g328 ( 
.A(n_245),
.B(n_273),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_256),
.C(n_266),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_246),
.B(n_324),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_252),
.Y(n_247)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_256),
.A2(n_257),
.B1(n_266),
.B2(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_262),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_258),
.B(n_262),
.Y(n_299)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_265),
.Y(n_296)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_266),
.Y(n_325)
);

AO22x1_ASAP7_75t_SL g266 ( 
.A1(n_267),
.A2(n_270),
.B1(n_271),
.B2(n_272),
.Y(n_266)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_267),
.Y(n_271)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g272 ( 
.A(n_270),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_270),
.B(n_271),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_272),
.B(n_315),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_279),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_275),
.B(n_279),
.C(n_342),
.Y(n_341)
);

HB1xp67_ASAP7_75t_L g342 ( 
.A(n_276),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_281),
.Y(n_279)
);

MAJx2_ASAP7_75t_L g337 ( 
.A(n_280),
.B(n_282),
.C(n_283),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

BUFx2_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_287),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_289),
.A2(n_322),
.B(n_327),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_290),
.A2(n_305),
.B(n_321),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_297),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_291),
.B(n_297),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_293),
.Y(n_313)
);

BUFx2_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_298),
.A2(n_299),
.B1(n_300),
.B2(n_301),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_306),
.A2(n_314),
.B(n_320),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_312),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_307),
.B(n_312),
.Y(n_320)
);

INVx1_ASAP7_75t_SL g308 ( 
.A(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx2_ASAP7_75t_SL g317 ( 
.A(n_318),
.Y(n_317)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_323),
.B(n_326),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_323),
.B(n_326),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_341),
.Y(n_329)
);

NOR2x1_ASAP7_75t_L g343 ( 
.A(n_330),
.B(n_341),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_331),
.A2(n_332),
.B1(n_338),
.B2(n_339),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_333),
.A2(n_334),
.B1(n_336),
.B2(n_337),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_333),
.B(n_337),
.C(n_338),
.Y(n_345)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

NOR2xp67_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_346),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_345),
.B(n_346),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

HB1xp67_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);


endmodule