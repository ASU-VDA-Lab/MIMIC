module fake_jpeg_5441_n_203 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_203);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_203;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx2_ASAP7_75t_SL g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_34),
.Y(n_44)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_37),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_20),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_38),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_20),
.B(n_17),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_30),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_20),
.Y(n_43)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_40),
.A2(n_30),
.B1(n_19),
.B2(n_27),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_46),
.A2(n_19),
.B1(n_15),
.B2(n_26),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_36),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_47),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_20),
.Y(n_48)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_51),
.B(n_31),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_32),
.B(n_22),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_52),
.B(n_31),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_39),
.A2(n_19),
.B1(n_30),
.B2(n_24),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_53),
.A2(n_21),
.B1(n_29),
.B2(n_25),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_57),
.Y(n_63)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_59),
.B(n_60),
.Y(n_79)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_38),
.B(n_15),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_61),
.B(n_24),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_62),
.B(n_77),
.Y(n_94)
);

BUFx4f_ASAP7_75t_SL g64 ( 
.A(n_50),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_64),
.B(n_66),
.Y(n_86)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_67),
.Y(n_100)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_68),
.B(n_78),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_47),
.A2(n_18),
.B1(n_29),
.B2(n_21),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_69),
.A2(n_80),
.B1(n_22),
.B2(n_23),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_71),
.B(n_73),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_18),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_72),
.B(n_74),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_53),
.B(n_25),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_58),
.A2(n_26),
.B1(n_23),
.B2(n_17),
.Y(n_80)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_82),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_90),
.Y(n_106)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_85),
.B(n_87),
.Y(n_122)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_81),
.B(n_52),
.Y(n_89)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_89),
.Y(n_111)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_70),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_91),
.B(n_99),
.Y(n_112)
);

NAND2xp67_ASAP7_75t_SL g92 ( 
.A(n_77),
.B(n_62),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_72),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_43),
.Y(n_93)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_93),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_51),
.Y(n_96)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_70),
.B(n_42),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_97),
.B(n_62),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_75),
.A2(n_58),
.B1(n_54),
.B2(n_59),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_98),
.A2(n_102),
.B1(n_66),
.B2(n_68),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_64),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_101),
.B(n_42),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_77),
.A2(n_58),
.B1(n_54),
.B2(n_56),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_76),
.B(n_45),
.Y(n_103)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_103),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_105),
.A2(n_100),
.B1(n_101),
.B2(n_54),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_107),
.B(n_118),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_95),
.B(n_75),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_108),
.B(n_109),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_91),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_110),
.Y(n_129)
);

OAI21xp33_ASAP7_75t_L g136 ( 
.A1(n_115),
.A2(n_116),
.B(n_85),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_88),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_83),
.B(n_63),
.Y(n_119)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_119),
.Y(n_125)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_120),
.B(n_55),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_83),
.B(n_99),
.Y(n_121)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_121),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_73),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_123),
.A2(n_124),
.B(n_71),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_97),
.B(n_87),
.C(n_104),
.Y(n_124)
);

AOI322xp5_ASAP7_75t_L g126 ( 
.A1(n_115),
.A2(n_123),
.A3(n_108),
.B1(n_95),
.B2(n_122),
.C1(n_94),
.C2(n_92),
.Y(n_126)
);

BUFx24_ASAP7_75t_SL g151 ( 
.A(n_126),
.Y(n_151)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_128),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_120),
.A2(n_100),
.B(n_94),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_130),
.A2(n_132),
.B(n_137),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_112),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_131),
.B(n_138),
.Y(n_145)
);

AND2x4_ASAP7_75t_L g132 ( 
.A(n_123),
.B(n_95),
.Y(n_132)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_134),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_110),
.B(n_99),
.Y(n_135)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_135),
.Y(n_152)
);

OA21x2_ASAP7_75t_SL g150 ( 
.A1(n_136),
.A2(n_115),
.B(n_118),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_114),
.B(n_90),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_124),
.A2(n_60),
.B1(n_55),
.B2(n_84),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_140),
.A2(n_105),
.B1(n_113),
.B2(n_111),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_106),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_141),
.B(n_142),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_122),
.B(n_84),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_137),
.B(n_109),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_144),
.B(n_155),
.C(n_146),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_132),
.B(n_139),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_148),
.A2(n_153),
.B1(n_125),
.B2(n_133),
.Y(n_164)
);

NOR3xp33_ASAP7_75t_SL g158 ( 
.A(n_150),
.B(n_132),
.C(n_130),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_129),
.B(n_142),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_154),
.B(n_133),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_139),
.B(n_113),
.C(n_111),
.Y(n_155)
);

MAJx2_ASAP7_75t_L g156 ( 
.A(n_132),
.B(n_107),
.C(n_117),
.Y(n_156)
);

MAJx2_ASAP7_75t_L g168 ( 
.A(n_156),
.B(n_114),
.C(n_3),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_140),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_157),
.B(n_141),
.Y(n_163)
);

NOR3xp33_ASAP7_75t_L g179 ( 
.A(n_158),
.B(n_167),
.C(n_6),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_143),
.A2(n_129),
.B1(n_131),
.B2(n_132),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_159),
.A2(n_65),
.B1(n_7),
.B2(n_8),
.Y(n_178)
);

OAI322xp33_ASAP7_75t_L g160 ( 
.A1(n_148),
.A2(n_151),
.A3(n_156),
.B1(n_144),
.B2(n_146),
.C1(n_155),
.C2(n_149),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_160),
.B(n_161),
.C(n_162),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_148),
.B(n_128),
.C(n_127),
.Y(n_162)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_163),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_164),
.A2(n_168),
.B(n_169),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_165),
.B(n_6),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_153),
.B(n_125),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_166),
.B(n_170),
.Y(n_172)
);

NOR2x1_ASAP7_75t_L g167 ( 
.A(n_157),
.B(n_117),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_152),
.B(n_0),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_145),
.B(n_65),
.C(n_9),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_167),
.A2(n_147),
.B1(n_10),
.B2(n_11),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_173),
.B(n_12),
.Y(n_185)
);

AOI31xp67_ASAP7_75t_L g175 ( 
.A1(n_168),
.A2(n_3),
.A3(n_4),
.B(n_5),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_175),
.B(n_179),
.Y(n_181)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_162),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_177),
.B(n_178),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_180),
.B(n_170),
.C(n_166),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_174),
.B(n_161),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_183),
.B(n_188),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_184),
.B(n_176),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_185),
.B(n_7),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_179),
.B(n_158),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_186),
.A2(n_177),
.B(n_14),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_172),
.B(n_10),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_187),
.B(n_182),
.C(n_181),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_171),
.B(n_12),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_190),
.B(n_192),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_191),
.Y(n_197)
);

AOI31xp67_ASAP7_75t_SL g192 ( 
.A1(n_186),
.A2(n_6),
.A3(n_7),
.B(n_8),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_193),
.B(n_194),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_189),
.B(n_182),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_195),
.A2(n_194),
.B(n_181),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_199),
.B(n_197),
.C(n_8),
.Y(n_202)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_196),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_200),
.B(n_198),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_201),
.B(n_202),
.Y(n_203)
);


endmodule