module real_aes_1893_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_801, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_801;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_766;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_791;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_796;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_769;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_785;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_797;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_L g214 ( .A(n_0), .B(n_136), .Y(n_214) );
CKINVDCx20_ASAP7_75t_R g774 ( .A(n_1), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_2), .B(n_797), .Y(n_796) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_3), .B(n_142), .Y(n_155) );
INVx1_ASAP7_75t_L g129 ( .A(n_4), .Y(n_129) );
NAND2xp33_ASAP7_75t_SL g206 ( .A(n_5), .B(n_140), .Y(n_206) );
INVx1_ASAP7_75t_L g187 ( .A(n_6), .Y(n_187) );
NAND2xp5_ASAP7_75t_SL g533 ( .A(n_7), .B(n_160), .Y(n_533) );
INVx1_ASAP7_75t_L g513 ( .A(n_8), .Y(n_513) );
CKINVDCx16_ASAP7_75t_R g797 ( .A(n_9), .Y(n_797) );
AND2x2_ASAP7_75t_L g153 ( .A(n_10), .B(n_146), .Y(n_153) );
CKINVDCx5p33_ASAP7_75t_R g480 ( .A(n_11), .Y(n_480) );
INVx2_ASAP7_75t_L g147 ( .A(n_12), .Y(n_147) );
AOI22xp33_ASAP7_75t_L g100 ( .A1(n_13), .A2(n_101), .B1(n_791), .B2(n_798), .Y(n_100) );
AOI22xp5_ASAP7_75t_L g108 ( .A1(n_14), .A2(n_109), .B1(n_110), .B2(n_765), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g765 ( .A(n_14), .Y(n_765) );
CKINVDCx16_ASAP7_75t_R g112 ( .A(n_15), .Y(n_112) );
NOR2xp33_ASAP7_75t_L g709 ( .A(n_15), .B(n_28), .Y(n_709) );
INVx1_ASAP7_75t_L g541 ( .A(n_16), .Y(n_541) );
OAI22xp5_ASAP7_75t_SL g784 ( .A1(n_17), .A2(n_28), .B1(n_763), .B2(n_785), .Y(n_784) );
CKINVDCx20_ASAP7_75t_R g785 ( .A(n_17), .Y(n_785) );
AOI221x1_ASAP7_75t_L g200 ( .A1(n_18), .A2(n_124), .B1(n_201), .B2(n_203), .C(n_205), .Y(n_200) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_19), .B(n_142), .Y(n_175) );
INVx1_ASAP7_75t_L g106 ( .A(n_20), .Y(n_106) );
INVx1_ASAP7_75t_L g539 ( .A(n_21), .Y(n_539) );
INVx1_ASAP7_75t_SL g462 ( .A(n_22), .Y(n_462) );
NAND2xp5_ASAP7_75t_SL g529 ( .A(n_23), .B(n_143), .Y(n_529) );
AOI21xp5_ASAP7_75t_L g156 ( .A1(n_24), .A2(n_124), .B(n_157), .Y(n_156) );
AOI221xp5_ASAP7_75t_SL g167 ( .A1(n_25), .A2(n_41), .B1(n_124), .B2(n_142), .C(n_168), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_26), .B(n_136), .Y(n_158) );
AOI33xp33_ASAP7_75t_L g499 ( .A1(n_27), .A2(n_52), .A3(n_190), .B1(n_196), .B2(n_500), .B3(n_501), .Y(n_499) );
INVx1_ASAP7_75t_L g763 ( .A(n_28), .Y(n_763) );
INVx1_ASAP7_75t_L g473 ( .A(n_29), .Y(n_473) );
OR2x2_ASAP7_75t_L g148 ( .A(n_30), .B(n_89), .Y(n_148) );
OA21x2_ASAP7_75t_L g181 ( .A1(n_30), .A2(n_89), .B(n_147), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_31), .B(n_132), .Y(n_179) );
INVxp67_ASAP7_75t_L g199 ( .A(n_32), .Y(n_199) );
AND2x2_ASAP7_75t_L g230 ( .A(n_33), .B(n_145), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_34), .B(n_188), .Y(n_459) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_35), .A2(n_124), .B(n_213), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_36), .B(n_132), .Y(n_169) );
AND2x2_ASAP7_75t_L g125 ( .A(n_37), .B(n_126), .Y(n_125) );
AND2x2_ASAP7_75t_L g140 ( .A(n_37), .B(n_129), .Y(n_140) );
INVx1_ASAP7_75t_L g195 ( .A(n_37), .Y(n_195) );
OR2x6_ASAP7_75t_L g104 ( .A(n_38), .B(n_105), .Y(n_104) );
NOR3xp33_ASAP7_75t_L g795 ( .A(n_38), .B(n_112), .C(n_796), .Y(n_795) );
CKINVDCx20_ASAP7_75t_R g475 ( .A(n_39), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_40), .B(n_188), .Y(n_487) );
AOI22xp5_ASAP7_75t_L g522 ( .A1(n_42), .A2(n_160), .B1(n_204), .B2(n_523), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_43), .B(n_531), .Y(n_530) );
AOI22xp5_ASAP7_75t_L g266 ( .A1(n_44), .A2(n_81), .B1(n_124), .B2(n_193), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_45), .B(n_143), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_46), .B(n_136), .Y(n_228) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_47), .B(n_180), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_48), .B(n_143), .Y(n_514) );
CKINVDCx5p33_ASAP7_75t_R g526 ( .A(n_49), .Y(n_526) );
AND2x2_ASAP7_75t_L g217 ( .A(n_50), .B(n_145), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_51), .B(n_145), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_53), .B(n_143), .Y(n_491) );
INVx1_ASAP7_75t_L g128 ( .A(n_54), .Y(n_128) );
INVx1_ASAP7_75t_L g138 ( .A(n_54), .Y(n_138) );
AND2x2_ASAP7_75t_L g492 ( .A(n_55), .B(n_145), .Y(n_492) );
AOI221xp5_ASAP7_75t_L g511 ( .A1(n_56), .A2(n_74), .B1(n_188), .B2(n_193), .C(n_512), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_57), .B(n_188), .Y(n_456) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_58), .B(n_142), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_59), .B(n_204), .Y(n_482) );
AOI21xp5_ASAP7_75t_SL g451 ( .A1(n_60), .A2(n_193), .B(n_452), .Y(n_451) );
AND2x2_ASAP7_75t_L g149 ( .A(n_61), .B(n_145), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_62), .B(n_132), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_63), .B(n_136), .Y(n_135) );
AND2x2_ASAP7_75t_SL g182 ( .A(n_64), .B(n_146), .Y(n_182) );
INVx1_ASAP7_75t_L g536 ( .A(n_65), .Y(n_536) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_66), .A2(n_124), .B(n_226), .Y(n_225) );
INVx1_ASAP7_75t_L g490 ( .A(n_67), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_68), .B(n_132), .Y(n_159) );
AND2x2_ASAP7_75t_SL g267 ( .A(n_69), .B(n_180), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_70), .B(n_767), .Y(n_766) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_71), .A2(n_193), .B(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g126 ( .A(n_72), .Y(n_126) );
INVx1_ASAP7_75t_L g134 ( .A(n_72), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_73), .B(n_188), .Y(n_502) );
AND2x2_ASAP7_75t_L g464 ( .A(n_75), .B(n_203), .Y(n_464) );
INVx1_ASAP7_75t_L g537 ( .A(n_76), .Y(n_537) );
AOI21xp5_ASAP7_75t_L g460 ( .A1(n_77), .A2(n_193), .B(n_461), .Y(n_460) );
A2O1A1Ixp33_ASAP7_75t_L g527 ( .A1(n_78), .A2(n_193), .B(n_263), .C(n_528), .Y(n_527) );
NAND2xp5_ASAP7_75t_SL g141 ( .A(n_79), .B(n_142), .Y(n_141) );
AOI22xp5_ASAP7_75t_L g265 ( .A1(n_80), .A2(n_84), .B1(n_142), .B2(n_188), .Y(n_265) );
INVx1_ASAP7_75t_L g107 ( .A(n_82), .Y(n_107) );
AND2x2_ASAP7_75t_SL g449 ( .A(n_83), .B(n_203), .Y(n_449) );
AOI22xp5_ASAP7_75t_L g496 ( .A1(n_85), .A2(n_193), .B1(n_497), .B2(n_498), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_86), .B(n_136), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_87), .B(n_136), .Y(n_170) );
AOI21xp5_ASAP7_75t_L g123 ( .A1(n_88), .A2(n_124), .B(n_130), .Y(n_123) );
INVx1_ASAP7_75t_L g453 ( .A(n_90), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_91), .B(n_132), .Y(n_131) );
AND2x2_ASAP7_75t_L g503 ( .A(n_92), .B(n_203), .Y(n_503) );
A2O1A1Ixp33_ASAP7_75t_L g470 ( .A1(n_93), .A2(n_471), .B(n_472), .C(n_474), .Y(n_470) );
INVxp67_ASAP7_75t_L g202 ( .A(n_94), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_95), .B(n_142), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_96), .B(n_132), .Y(n_227) );
AOI21xp5_ASAP7_75t_L g176 ( .A1(n_97), .A2(n_124), .B(n_177), .Y(n_176) );
BUFx2_ASAP7_75t_L g778 ( .A(n_98), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_99), .B(n_143), .Y(n_455) );
OA21x2_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_769), .B(n_779), .Y(n_101) );
OAI21x1_ASAP7_75t_L g102 ( .A1(n_103), .A2(n_108), .B(n_766), .Y(n_102) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_103), .B(n_112), .Y(n_773) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_104), .Y(n_103) );
OR2x2_ASAP7_75t_L g768 ( .A(n_104), .B(n_112), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_106), .B(n_107), .Y(n_105) );
NOR2xp33_ASAP7_75t_L g794 ( .A(n_106), .B(n_107), .Y(n_794) );
INVx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
OAI21x1_ASAP7_75t_L g110 ( .A1(n_111), .A2(n_113), .B(n_439), .Y(n_110) );
HB1xp67_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
CKINVDCx16_ASAP7_75t_R g764 ( .A(n_112), .Y(n_764) );
AND2x4_ASAP7_75t_L g113 ( .A(n_114), .B(n_378), .Y(n_113) );
NOR3xp33_ASAP7_75t_L g114 ( .A(n_115), .B(n_271), .C(n_322), .Y(n_114) );
OAI211xp5_ASAP7_75t_SL g115 ( .A1(n_116), .A2(n_161), .B(n_218), .C(n_249), .Y(n_115) );
INVxp67_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
NOR2xp33_ASAP7_75t_L g117 ( .A(n_118), .B(n_150), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
HB1xp67_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_120), .B(n_223), .Y(n_386) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
AND2x2_ASAP7_75t_L g231 ( .A(n_121), .B(n_152), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_121), .B(n_238), .Y(n_237) );
OR2x2_ASAP7_75t_L g248 ( .A(n_121), .B(n_238), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_121), .B(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g285 ( .A(n_121), .B(n_261), .Y(n_285) );
INVx2_ASAP7_75t_L g311 ( .A(n_121), .Y(n_311) );
AND2x4_ASAP7_75t_L g320 ( .A(n_121), .B(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g425 ( .A(n_121), .B(n_292), .Y(n_425) );
AO21x2_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_144), .B(n_149), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g122 ( .A(n_123), .B(n_141), .Y(n_122) );
AND2x6_ASAP7_75t_L g124 ( .A(n_125), .B(n_127), .Y(n_124) );
BUFx3_ASAP7_75t_L g192 ( .A(n_125), .Y(n_192) );
AND2x6_ASAP7_75t_L g136 ( .A(n_126), .B(n_137), .Y(n_136) );
INVx2_ASAP7_75t_L g197 ( .A(n_126), .Y(n_197) );
AND2x4_ASAP7_75t_L g193 ( .A(n_127), .B(n_194), .Y(n_193) );
AND2x2_ASAP7_75t_L g127 ( .A(n_128), .B(n_129), .Y(n_127) );
AND2x4_ASAP7_75t_L g132 ( .A(n_128), .B(n_133), .Y(n_132) );
INVx2_ASAP7_75t_L g190 ( .A(n_128), .Y(n_190) );
HB1xp67_ASAP7_75t_L g191 ( .A(n_129), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_135), .B(n_139), .Y(n_130) );
INVxp67_ASAP7_75t_L g542 ( .A(n_132), .Y(n_542) );
AND2x4_ASAP7_75t_L g143 ( .A(n_133), .B(n_137), .Y(n_143) );
INVx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVxp67_ASAP7_75t_L g540 ( .A(n_136), .Y(n_540) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
AOI21xp5_ASAP7_75t_L g157 ( .A1(n_139), .A2(n_158), .B(n_159), .Y(n_157) );
AOI21xp5_ASAP7_75t_L g168 ( .A1(n_139), .A2(n_169), .B(n_170), .Y(n_168) );
AOI21xp5_ASAP7_75t_L g177 ( .A1(n_139), .A2(n_178), .B(n_179), .Y(n_177) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_139), .A2(n_214), .B(n_215), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_139), .A2(n_227), .B(n_228), .Y(n_226) );
O2A1O1Ixp33_ASAP7_75t_L g452 ( .A1(n_139), .A2(n_453), .B(n_454), .C(n_455), .Y(n_452) );
O2A1O1Ixp33_ASAP7_75t_SL g461 ( .A1(n_139), .A2(n_454), .B(n_462), .C(n_463), .Y(n_461) );
O2A1O1Ixp33_ASAP7_75t_L g489 ( .A1(n_139), .A2(n_454), .B(n_490), .C(n_491), .Y(n_489) );
INVx1_ASAP7_75t_L g497 ( .A(n_139), .Y(n_497) );
O2A1O1Ixp33_ASAP7_75t_SL g512 ( .A1(n_139), .A2(n_454), .B(n_513), .C(n_514), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_139), .A2(n_529), .B(n_530), .Y(n_528) );
NOR2xp33_ASAP7_75t_L g543 ( .A(n_139), .B(n_160), .Y(n_543) );
INVx5_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
AND2x4_ASAP7_75t_L g142 ( .A(n_140), .B(n_143), .Y(n_142) );
HB1xp67_ASAP7_75t_L g474 ( .A(n_140), .Y(n_474) );
INVx1_ASAP7_75t_L g207 ( .A(n_143), .Y(n_207) );
AO21x2_ASAP7_75t_L g223 ( .A1(n_144), .A2(n_224), .B(n_230), .Y(n_223) );
AO21x2_ASAP7_75t_L g238 ( .A1(n_144), .A2(n_224), .B(n_230), .Y(n_238) );
AO21x2_ASAP7_75t_L g457 ( .A1(n_144), .A2(n_458), .B(n_464), .Y(n_457) );
CKINVDCx5p33_ASAP7_75t_R g144 ( .A(n_145), .Y(n_144) );
OA21x2_ASAP7_75t_L g166 ( .A1(n_145), .A2(n_167), .B(n_171), .Y(n_166) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
AND2x2_ASAP7_75t_SL g146 ( .A(n_147), .B(n_148), .Y(n_146) );
AND2x4_ASAP7_75t_L g160 ( .A(n_147), .B(n_148), .Y(n_160) );
AND2x2_ASAP7_75t_L g309 ( .A(n_150), .B(n_310), .Y(n_309) );
OAI32xp33_ASAP7_75t_L g392 ( .A1(n_150), .A2(n_314), .A3(n_318), .B1(n_325), .B2(n_393), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_150), .B(n_425), .Y(n_424) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
AND2x2_ASAP7_75t_L g246 ( .A(n_151), .B(n_247), .Y(n_246) );
NAND3xp33_ASAP7_75t_L g319 ( .A(n_151), .B(n_241), .C(n_320), .Y(n_319) );
OR2x2_ASAP7_75t_L g345 ( .A(n_151), .B(n_248), .Y(n_345) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
HB1xp67_ASAP7_75t_L g235 ( .A(n_152), .Y(n_235) );
INVx5_ASAP7_75t_L g270 ( .A(n_152), .Y(n_270) );
AND2x4_ASAP7_75t_L g326 ( .A(n_152), .B(n_238), .Y(n_326) );
OR2x2_ASAP7_75t_L g341 ( .A(n_152), .B(n_261), .Y(n_341) );
OR2x2_ASAP7_75t_L g367 ( .A(n_152), .B(n_223), .Y(n_367) );
AND2x2_ASAP7_75t_L g375 ( .A(n_152), .B(n_321), .Y(n_375) );
AND2x4_ASAP7_75t_SL g400 ( .A(n_152), .B(n_320), .Y(n_400) );
OR2x6_ASAP7_75t_L g152 ( .A(n_153), .B(n_154), .Y(n_152) );
AOI21xp5_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_156), .B(n_160), .Y(n_154) );
NOR2xp33_ASAP7_75t_L g186 ( .A(n_160), .B(n_187), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g198 ( .A(n_160), .B(n_199), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g201 ( .A(n_160), .B(n_202), .Y(n_201) );
NOR3xp33_ASAP7_75t_L g205 ( .A(n_160), .B(n_206), .C(n_207), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g450 ( .A1(n_160), .A2(n_451), .B(n_456), .Y(n_450) );
INVx1_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_162), .B(n_320), .Y(n_396) );
AND2x2_ASAP7_75t_L g162 ( .A(n_163), .B(n_172), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_163), .B(n_295), .Y(n_294) );
INVx1_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
OR2x6_ASAP7_75t_SL g220 ( .A(n_164), .B(n_221), .Y(n_220) );
INVxp67_ASAP7_75t_SL g164 ( .A(n_165), .Y(n_164) );
INVx1_ASAP7_75t_L g245 ( .A(n_165), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_165), .B(n_280), .Y(n_298) );
HB1xp67_ASAP7_75t_L g436 ( .A(n_165), .Y(n_436) );
INVx1_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx2_ASAP7_75t_L g253 ( .A(n_166), .Y(n_253) );
AND2x2_ASAP7_75t_L g278 ( .A(n_166), .B(n_209), .Y(n_278) );
INVx2_ASAP7_75t_L g306 ( .A(n_166), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_166), .B(n_173), .Y(n_347) );
BUFx3_ASAP7_75t_L g371 ( .A(n_166), .Y(n_371) );
OR2x2_ASAP7_75t_L g383 ( .A(n_166), .B(n_173), .Y(n_383) );
HB1xp67_ASAP7_75t_L g391 ( .A(n_166), .Y(n_391) );
AOI22xp5_ASAP7_75t_L g413 ( .A1(n_172), .A2(n_414), .B1(n_417), .B2(n_418), .Y(n_413) );
AND2x2_ASAP7_75t_L g172 ( .A(n_173), .B(n_183), .Y(n_172) );
INVx1_ASAP7_75t_L g241 ( .A(n_173), .Y(n_241) );
OR2x2_ASAP7_75t_L g252 ( .A(n_173), .B(n_253), .Y(n_252) );
INVx2_ASAP7_75t_L g259 ( .A(n_173), .Y(n_259) );
AND2x4_ASAP7_75t_SL g276 ( .A(n_173), .B(n_184), .Y(n_276) );
AND2x4_ASAP7_75t_L g281 ( .A(n_173), .B(n_282), .Y(n_281) );
INVx2_ASAP7_75t_L g290 ( .A(n_173), .Y(n_290) );
OR2x2_ASAP7_75t_L g296 ( .A(n_173), .B(n_184), .Y(n_296) );
OR2x2_ASAP7_75t_L g297 ( .A(n_173), .B(n_298), .Y(n_297) );
HB1xp67_ASAP7_75t_L g408 ( .A(n_173), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_173), .B(n_278), .Y(n_412) );
OR2x2_ASAP7_75t_L g428 ( .A(n_173), .B(n_331), .Y(n_428) );
OR2x6_ASAP7_75t_L g173 ( .A(n_174), .B(n_182), .Y(n_173) );
AOI21xp5_ASAP7_75t_L g174 ( .A1(n_175), .A2(n_176), .B(n_180), .Y(n_174) );
INVx2_ASAP7_75t_SL g263 ( .A(n_180), .Y(n_263) );
OA21x2_ASAP7_75t_L g510 ( .A1(n_180), .A2(n_511), .B(n_515), .Y(n_510) );
BUFx4f_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx3_ASAP7_75t_L g204 ( .A(n_181), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_183), .B(n_241), .Y(n_240) );
INVx1_ASAP7_75t_L g254 ( .A(n_183), .Y(n_254) );
AND2x2_ASAP7_75t_SL g361 ( .A(n_183), .B(n_245), .Y(n_361) );
AND2x4_ASAP7_75t_L g183 ( .A(n_184), .B(n_208), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_184), .B(n_209), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_184), .B(n_243), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_184), .B(n_253), .Y(n_257) );
INVx3_ASAP7_75t_L g282 ( .A(n_184), .Y(n_282) );
INVx1_ASAP7_75t_L g315 ( .A(n_184), .Y(n_315) );
AND2x2_ASAP7_75t_L g395 ( .A(n_184), .B(n_259), .Y(n_395) );
AND2x4_ASAP7_75t_L g184 ( .A(n_185), .B(n_200), .Y(n_184) );
AOI22xp5_ASAP7_75t_L g185 ( .A1(n_186), .A2(n_188), .B1(n_193), .B2(n_198), .Y(n_185) );
INVx1_ASAP7_75t_L g483 ( .A(n_188), .Y(n_483) );
AND2x4_ASAP7_75t_L g188 ( .A(n_189), .B(n_192), .Y(n_188) );
INVx1_ASAP7_75t_L g524 ( .A(n_189), .Y(n_524) );
AND2x2_ASAP7_75t_L g189 ( .A(n_190), .B(n_191), .Y(n_189) );
OR2x6_ASAP7_75t_L g454 ( .A(n_190), .B(n_197), .Y(n_454) );
INVxp33_ASAP7_75t_L g500 ( .A(n_190), .Y(n_500) );
INVx1_ASAP7_75t_L g525 ( .A(n_192), .Y(n_525) );
INVxp67_ASAP7_75t_L g481 ( .A(n_193), .Y(n_481) );
NOR2x1p5_ASAP7_75t_L g194 ( .A(n_195), .B(n_196), .Y(n_194) );
INVx1_ASAP7_75t_L g501 ( .A(n_196), .Y(n_501) );
INVx3_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
OAI22xp5_ASAP7_75t_L g469 ( .A1(n_203), .A2(n_470), .B1(n_475), .B2(n_476), .Y(n_469) );
INVx3_ASAP7_75t_L g476 ( .A(n_203), .Y(n_476) );
INVx4_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
AOI21x1_ASAP7_75t_L g210 ( .A1(n_204), .A2(n_211), .B(n_217), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_204), .B(n_479), .Y(n_478) );
NOR2xp33_ASAP7_75t_L g472 ( .A(n_207), .B(n_473), .Y(n_472) );
OAI22xp5_ASAP7_75t_L g535 ( .A1(n_207), .A2(n_454), .B1(n_536), .B2(n_537), .Y(n_535) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_209), .B(n_259), .Y(n_258) );
INVx1_ASAP7_75t_L g280 ( .A(n_209), .Y(n_280) );
AND2x2_ASAP7_75t_L g305 ( .A(n_209), .B(n_306), .Y(n_305) );
OR2x2_ASAP7_75t_L g331 ( .A(n_209), .B(n_253), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_209), .B(n_282), .Y(n_348) );
INVx1_ASAP7_75t_L g354 ( .A(n_209), .Y(n_354) );
INVx3_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_212), .B(n_216), .Y(n_211) );
AOI222xp33_ASAP7_75t_SL g218 ( .A1(n_219), .A2(n_222), .B1(n_232), .B2(n_239), .C1(n_242), .C2(n_246), .Y(n_218) );
CKINVDCx16_ASAP7_75t_R g219 ( .A(n_220), .Y(n_219) );
AND2x2_ASAP7_75t_L g222 ( .A(n_223), .B(n_231), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g343 ( .A(n_223), .B(n_292), .Y(n_343) );
AND2x4_ASAP7_75t_L g359 ( .A(n_223), .B(n_270), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_225), .B(n_229), .Y(n_224) );
INVx2_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_234), .B(n_236), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
AND2x2_ASAP7_75t_L g284 ( .A(n_235), .B(n_285), .Y(n_284) );
AOI222xp33_ASAP7_75t_L g249 ( .A1(n_236), .A2(n_250), .B1(n_255), .B2(n_260), .C1(n_268), .C2(n_801), .Y(n_249) );
INVx1_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
OR2x2_ASAP7_75t_L g388 ( .A(n_237), .B(n_292), .Y(n_388) );
OR2x2_ASAP7_75t_L g431 ( .A(n_237), .B(n_337), .Y(n_431) );
AND2x2_ASAP7_75t_L g260 ( .A(n_238), .B(n_261), .Y(n_260) );
INVx2_ASAP7_75t_L g321 ( .A(n_238), .Y(n_321) );
HB1xp67_ASAP7_75t_L g336 ( .A(n_238), .Y(n_336) );
O2A1O1Ixp33_ASAP7_75t_L g349 ( .A1(n_239), .A2(n_350), .B(n_355), .C(n_356), .Y(n_349) );
INVx1_ASAP7_75t_SL g239 ( .A(n_240), .Y(n_239) );
INVx1_ASAP7_75t_L g377 ( .A(n_241), .Y(n_377) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
HB1xp67_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
INVx2_ASAP7_75t_L g307 ( .A(n_246), .Y(n_307) );
AND2x2_ASAP7_75t_L g291 ( .A(n_247), .B(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g300 ( .A(n_247), .B(n_301), .Y(n_300) );
INVx2_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
OAI31xp33_ASAP7_75t_L g342 ( .A1(n_250), .A2(n_268), .A3(n_343), .B(n_344), .Y(n_342) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
A2O1A1Ixp33_ASAP7_75t_L g344 ( .A1(n_251), .A2(n_301), .B(n_345), .C(n_346), .Y(n_344) );
OR2x2_ASAP7_75t_L g251 ( .A(n_252), .B(n_254), .Y(n_251) );
OR2x2_ASAP7_75t_L g333 ( .A(n_252), .B(n_282), .Y(n_333) );
INVx2_ASAP7_75t_SL g255 ( .A(n_256), .Y(n_255) );
OR2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_258), .Y(n_256) );
BUFx2_ASAP7_75t_L g301 ( .A(n_261), .Y(n_301) );
AND2x2_ASAP7_75t_L g310 ( .A(n_261), .B(n_311), .Y(n_310) );
INVx2_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
BUFx6f_ASAP7_75t_L g292 ( .A(n_262), .Y(n_292) );
AOI21x1_ASAP7_75t_L g262 ( .A1(n_263), .A2(n_264), .B(n_267), .Y(n_262) );
AO21x2_ASAP7_75t_L g494 ( .A1(n_263), .A2(n_495), .B(n_503), .Y(n_494) );
AO21x2_ASAP7_75t_L g554 ( .A1(n_263), .A2(n_495), .B(n_503), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_270), .B(n_327), .Y(n_419) );
OAI211xp5_ASAP7_75t_L g271 ( .A1(n_272), .A2(n_283), .B(n_286), .C(n_308), .Y(n_271) );
INVxp33_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
NAND2xp5_ASAP7_75t_SL g273 ( .A(n_274), .B(n_279), .Y(n_273) );
OR2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_277), .Y(n_274) );
INVx1_ASAP7_75t_SL g275 ( .A(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g312 ( .A(n_276), .B(n_305), .Y(n_312) );
OR2x2_ASAP7_75t_L g288 ( .A(n_277), .B(n_289), .Y(n_288) );
OR2x2_ASAP7_75t_L g318 ( .A(n_277), .B(n_292), .Y(n_318) );
INVx2_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g394 ( .A(n_278), .B(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g417 ( .A(n_279), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_281), .B(n_330), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_281), .B(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g429 ( .A(n_281), .B(n_305), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_281), .B(n_435), .Y(n_434) );
AND2x2_ASAP7_75t_L g372 ( .A(n_282), .B(n_354), .Y(n_372) );
INVx1_ASAP7_75t_SL g283 ( .A(n_284), .Y(n_283) );
AOI322xp5_ASAP7_75t_L g426 ( .A1(n_285), .A2(n_305), .A3(n_359), .B1(n_384), .B2(n_427), .C1(n_429), .C2(n_430), .Y(n_426) );
AOI211xp5_ASAP7_75t_SL g286 ( .A1(n_287), .A2(n_291), .B(n_293), .C(n_302), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_289), .B(n_317), .Y(n_339) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g304 ( .A(n_290), .B(n_305), .Y(n_304) );
NOR2x1p5_ASAP7_75t_L g370 ( .A(n_290), .B(n_371), .Y(n_370) );
HB1xp67_ASAP7_75t_L g403 ( .A(n_290), .Y(n_403) );
O2A1O1Ixp33_ASAP7_75t_L g308 ( .A1(n_291), .A2(n_309), .B(n_312), .C(n_313), .Y(n_308) );
AND2x4_ASAP7_75t_L g327 ( .A(n_292), .B(n_311), .Y(n_327) );
INVx2_ASAP7_75t_L g337 ( .A(n_292), .Y(n_337) );
NAND2xp5_ASAP7_75t_SL g357 ( .A(n_292), .B(n_326), .Y(n_357) );
AND2x2_ASAP7_75t_L g399 ( .A(n_292), .B(n_400), .Y(n_399) );
NOR2xp33_ASAP7_75t_L g437 ( .A(n_292), .B(n_416), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_292), .B(n_320), .Y(n_438) );
AOI21xp33_ASAP7_75t_L g293 ( .A1(n_294), .A2(n_297), .B(n_299), .Y(n_293) );
AND2x2_ASAP7_75t_L g389 ( .A(n_295), .B(n_390), .Y(n_389) );
INVx1_ASAP7_75t_SL g295 ( .A(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g317 ( .A(n_298), .Y(n_317) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
NOR2xp33_ASAP7_75t_L g302 ( .A(n_303), .B(n_307), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_310), .B(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g404 ( .A(n_310), .Y(n_404) );
O2A1O1Ixp33_ASAP7_75t_SL g313 ( .A1(n_314), .A2(n_316), .B(n_318), .C(n_319), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
HB1xp67_ASAP7_75t_L g401 ( .A(n_317), .Y(n_401) );
INVx3_ASAP7_75t_SL g416 ( .A(n_320), .Y(n_416) );
NAND5xp2_ASAP7_75t_L g322 ( .A(n_323), .B(n_342), .C(n_349), .D(n_362), .E(n_373), .Y(n_322) );
AOI222xp33_ASAP7_75t_L g323 ( .A1(n_324), .A2(n_328), .B1(n_332), .B2(n_334), .C1(n_338), .C2(n_340), .Y(n_323) );
NOR2xp33_ASAP7_75t_L g324 ( .A(n_325), .B(n_327), .Y(n_324) );
AOI22xp5_ASAP7_75t_L g405 ( .A1(n_325), .A2(n_406), .B1(n_410), .B2(n_411), .Y(n_405) );
INVx2_ASAP7_75t_SL g325 ( .A(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g355 ( .A(n_326), .B(n_327), .Y(n_355) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_SL g332 ( .A(n_333), .Y(n_332) );
NOR2xp33_ASAP7_75t_L g334 ( .A(n_335), .B(n_337), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
NAND2xp5_ASAP7_75t_SL g422 ( .A(n_336), .B(n_423), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_337), .B(n_359), .Y(n_358) );
AND2x2_ASAP7_75t_L g374 ( .A(n_337), .B(n_375), .Y(n_374) );
OR2x2_ASAP7_75t_L g385 ( .A(n_337), .B(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_SL g340 ( .A(n_341), .Y(n_340) );
OR2x2_ASAP7_75t_L g415 ( .A(n_341), .B(n_416), .Y(n_415) );
OR2x2_ASAP7_75t_L g346 ( .A(n_347), .B(n_348), .Y(n_346) );
INVx1_ASAP7_75t_L g363 ( .A(n_348), .Y(n_363) );
INVxp67_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVxp67_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
AOI21xp33_ASAP7_75t_L g356 ( .A1(n_357), .A2(n_358), .B(n_360), .Y(n_356) );
AOI22xp33_ASAP7_75t_L g362 ( .A1(n_359), .A2(n_363), .B1(n_364), .B2(n_368), .Y(n_362) );
HB1xp67_ASAP7_75t_L g410 ( .A(n_359), .Y(n_410) );
INVx2_ASAP7_75t_SL g360 ( .A(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g376 ( .A(n_361), .B(n_377), .Y(n_376) );
AND2x2_ASAP7_75t_L g381 ( .A(n_363), .B(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_SL g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_370), .B(n_372), .Y(n_369) );
INVx1_ASAP7_75t_SL g409 ( .A(n_372), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_374), .B(n_376), .Y(n_373) );
NOR3xp33_ASAP7_75t_L g378 ( .A(n_379), .B(n_397), .C(n_420), .Y(n_378) );
NAND2xp5_ASAP7_75t_SL g379 ( .A(n_380), .B(n_396), .Y(n_379) );
AOI221xp5_ASAP7_75t_L g380 ( .A1(n_381), .A2(n_384), .B1(n_387), .B2(n_389), .C(n_392), .Y(n_380) );
INVx1_ASAP7_75t_SL g382 ( .A(n_383), .Y(n_382) );
OR2x2_ASAP7_75t_L g421 ( .A(n_383), .B(n_409), .Y(n_421) );
INVx1_ASAP7_75t_SL g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_SL g387 ( .A(n_388), .Y(n_387) );
HB1xp67_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_SL g393 ( .A(n_394), .Y(n_393) );
OAI321xp33_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_401), .A3(n_402), .B1(n_404), .B2(n_405), .C(n_413), .Y(n_397) );
INVx1_ASAP7_75t_SL g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_SL g406 ( .A(n_407), .Y(n_406) );
OR2x2_ASAP7_75t_L g407 ( .A(n_408), .B(n_409), .Y(n_407) );
AOI22xp33_ASAP7_75t_L g432 ( .A1(n_411), .A2(n_433), .B1(n_437), .B2(n_438), .Y(n_432) );
INVx1_ASAP7_75t_SL g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
OAI211xp5_ASAP7_75t_SL g420 ( .A1(n_421), .A2(n_422), .B(n_426), .C(n_432), .Y(n_420) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_SL g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVxp67_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
NOR2x1_ASAP7_75t_L g439 ( .A(n_440), .B(n_760), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_441), .B(n_710), .Y(n_440) );
OAI21xp5_ASAP7_75t_L g441 ( .A1(n_442), .A2(n_650), .B(n_709), .Y(n_441) );
NOR3xp33_ASAP7_75t_L g760 ( .A(n_442), .B(n_711), .C(n_761), .Y(n_760) );
INVx1_ASAP7_75t_L g788 ( .A(n_442), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_443), .B(n_614), .Y(n_442) );
NOR3xp33_ASAP7_75t_L g443 ( .A(n_444), .B(n_555), .C(n_584), .Y(n_443) );
NAND2xp5_ASAP7_75t_SL g444 ( .A(n_445), .B(n_544), .Y(n_444) );
AOI22xp5_ASAP7_75t_L g445 ( .A1(n_446), .A2(n_465), .B1(n_504), .B2(n_516), .Y(n_445) );
NAND2x1_ASAP7_75t_L g746 ( .A(n_446), .B(n_545), .Y(n_746) );
INVx2_ASAP7_75t_SL g446 ( .A(n_447), .Y(n_446) );
OR2x2_ASAP7_75t_L g447 ( .A(n_448), .B(n_457), .Y(n_447) );
INVx2_ASAP7_75t_L g518 ( .A(n_448), .Y(n_518) );
INVx4_ASAP7_75t_L g560 ( .A(n_448), .Y(n_560) );
BUFx6f_ASAP7_75t_L g580 ( .A(n_448), .Y(n_580) );
AND2x4_ASAP7_75t_L g591 ( .A(n_448), .B(n_559), .Y(n_591) );
AND2x2_ASAP7_75t_L g597 ( .A(n_448), .B(n_521), .Y(n_597) );
NOR2x1_ASAP7_75t_SL g670 ( .A(n_448), .B(n_532), .Y(n_670) );
OR2x6_ASAP7_75t_L g448 ( .A(n_449), .B(n_450), .Y(n_448) );
INVxp67_ASAP7_75t_L g471 ( .A(n_454), .Y(n_471) );
INVx2_ASAP7_75t_L g531 ( .A(n_454), .Y(n_531) );
INVx2_ASAP7_75t_L g563 ( .A(n_457), .Y(n_563) );
HB1xp67_ASAP7_75t_L g577 ( .A(n_457), .Y(n_577) );
INVx1_ASAP7_75t_L g588 ( .A(n_457), .Y(n_588) );
HB1xp67_ASAP7_75t_L g600 ( .A(n_457), .Y(n_600) );
AND2x2_ASAP7_75t_L g632 ( .A(n_457), .B(n_532), .Y(n_632) );
INVx1_ASAP7_75t_L g658 ( .A(n_457), .Y(n_658) );
AND2x2_ASAP7_75t_L g720 ( .A(n_457), .B(n_548), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_459), .B(n_460), .Y(n_458) );
AND2x2_ASAP7_75t_L g465 ( .A(n_466), .B(n_484), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
AND2x2_ASAP7_75t_L g613 ( .A(n_467), .B(n_552), .Y(n_613) );
INVx2_ASAP7_75t_L g655 ( .A(n_467), .Y(n_655) );
AND2x2_ASAP7_75t_L g757 ( .A(n_467), .B(n_484), .Y(n_757) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_468), .B(n_507), .Y(n_551) );
INVx2_ASAP7_75t_L g572 ( .A(n_468), .Y(n_572) );
AND2x4_ASAP7_75t_L g594 ( .A(n_468), .B(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g629 ( .A(n_468), .Y(n_629) );
AND2x2_ASAP7_75t_L g753 ( .A(n_468), .B(n_510), .Y(n_753) );
OR2x2_ASAP7_75t_L g468 ( .A(n_469), .B(n_477), .Y(n_468) );
AO21x2_ASAP7_75t_L g485 ( .A1(n_476), .A2(n_486), .B(n_492), .Y(n_485) );
AO21x2_ASAP7_75t_L g507 ( .A1(n_476), .A2(n_486), .B(n_492), .Y(n_507) );
OAI22xp5_ASAP7_75t_L g477 ( .A1(n_478), .A2(n_481), .B1(n_482), .B2(n_483), .Y(n_477) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx1_ASAP7_75t_L g727 ( .A(n_484), .Y(n_727) );
AND2x2_ASAP7_75t_L g484 ( .A(n_485), .B(n_493), .Y(n_484) );
NOR2xp67_ASAP7_75t_L g602 ( .A(n_485), .B(n_572), .Y(n_602) );
AND2x2_ASAP7_75t_L g607 ( .A(n_485), .B(n_572), .Y(n_607) );
INVx2_ASAP7_75t_L g620 ( .A(n_485), .Y(n_620) );
NOR2x1_ASAP7_75t_L g685 ( .A(n_485), .B(n_686), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_487), .B(n_488), .Y(n_486) );
AND2x4_ASAP7_75t_L g593 ( .A(n_493), .B(n_506), .Y(n_593) );
AND2x2_ASAP7_75t_L g608 ( .A(n_493), .B(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g663 ( .A(n_493), .Y(n_663) );
INVx2_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_494), .B(n_510), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_494), .B(n_507), .Y(n_661) );
NAND2xp5_ASAP7_75t_SL g495 ( .A(n_496), .B(n_502), .Y(n_495) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVxp33_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
NAND2x1p5_ASAP7_75t_L g505 ( .A(n_506), .B(n_508), .Y(n_505) );
INVx3_ASAP7_75t_L g569 ( .A(n_506), .Y(n_569) );
INVx3_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
HB1xp67_ASAP7_75t_L g567 ( .A(n_507), .Y(n_567) );
AND2x2_ASAP7_75t_L g681 ( .A(n_507), .B(n_682), .Y(n_681) );
INVx3_ASAP7_75t_L g624 ( .A(n_508), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_508), .B(n_663), .Y(n_704) );
BUFx3_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
AND2x2_ASAP7_75t_L g571 ( .A(n_509), .B(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
AND2x4_ASAP7_75t_L g552 ( .A(n_510), .B(n_553), .Y(n_552) );
INVx2_ASAP7_75t_L g595 ( .A(n_510), .Y(n_595) );
INVxp67_ASAP7_75t_L g609 ( .A(n_510), .Y(n_609) );
HB1xp67_ASAP7_75t_L g682 ( .A(n_510), .Y(n_682) );
INVx1_ASAP7_75t_L g686 ( .A(n_510), .Y(n_686) );
INVx1_ASAP7_75t_L g664 ( .A(n_516), .Y(n_664) );
NOR2x1_ASAP7_75t_L g516 ( .A(n_517), .B(n_519), .Y(n_516) );
NOR2x1_ASAP7_75t_L g641 ( .A(n_517), .B(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
AND2x2_ASAP7_75t_L g706 ( .A(n_518), .B(n_547), .Y(n_706) );
OR2x2_ASAP7_75t_L g758 ( .A(n_519), .B(n_759), .Y(n_758) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
AND2x2_ASAP7_75t_L g657 ( .A(n_520), .B(n_658), .Y(n_657) );
AND2x2_ASAP7_75t_L g693 ( .A(n_520), .B(n_580), .Y(n_693) );
AND2x2_ASAP7_75t_L g520 ( .A(n_521), .B(n_532), .Y(n_520) );
AND2x4_ASAP7_75t_L g547 ( .A(n_521), .B(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g559 ( .A(n_521), .Y(n_559) );
INVx2_ASAP7_75t_L g576 ( .A(n_521), .Y(n_576) );
HB1xp67_ASAP7_75t_L g702 ( .A(n_521), .Y(n_702) );
AND2x2_ASAP7_75t_L g521 ( .A(n_522), .B(n_527), .Y(n_521) );
NOR3xp33_ASAP7_75t_L g523 ( .A(n_524), .B(n_525), .C(n_526), .Y(n_523) );
INVx3_ASAP7_75t_L g548 ( .A(n_532), .Y(n_548) );
INVx2_ASAP7_75t_L g642 ( .A(n_532), .Y(n_642) );
AND2x4_ASAP7_75t_L g532 ( .A(n_533), .B(n_534), .Y(n_532) );
OAI21xp5_ASAP7_75t_L g534 ( .A1(n_535), .A2(n_538), .B(n_543), .Y(n_534) );
OAI22xp5_ASAP7_75t_L g538 ( .A1(n_539), .A2(n_540), .B1(n_541), .B2(n_542), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_545), .B(n_549), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
NOR2xp33_ASAP7_75t_L g639 ( .A(n_546), .B(n_622), .Y(n_639) );
NOR2x1_ASAP7_75t_L g731 ( .A(n_546), .B(n_560), .Y(n_731) );
INVx4_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_547), .B(n_622), .Y(n_708) );
AND2x2_ASAP7_75t_L g575 ( .A(n_548), .B(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g589 ( .A(n_548), .Y(n_589) );
AOI22xp5_ASAP7_75t_SL g637 ( .A1(n_549), .A2(n_638), .B1(n_639), .B2(n_640), .Y(n_637) );
AND2x2_ASAP7_75t_L g549 ( .A(n_550), .B(n_552), .Y(n_549) );
NAND2x1p5_ASAP7_75t_L g634 ( .A(n_550), .B(n_608), .Y(n_634) );
INVx2_ASAP7_75t_SL g550 ( .A(n_551), .Y(n_550) );
OR2x2_ASAP7_75t_L g742 ( .A(n_551), .B(n_583), .Y(n_742) );
AND2x2_ASAP7_75t_L g565 ( .A(n_552), .B(n_566), .Y(n_565) );
AND2x4_ASAP7_75t_L g601 ( .A(n_552), .B(n_602), .Y(n_601) );
AND2x2_ASAP7_75t_L g744 ( .A(n_552), .B(n_655), .Y(n_744) );
INVx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
AND2x4_ASAP7_75t_L g619 ( .A(n_554), .B(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g645 ( .A(n_554), .Y(n_645) );
AND2x2_ASAP7_75t_L g680 ( .A(n_554), .B(n_572), .Y(n_680) );
OAI221xp5_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_564), .B1(n_568), .B2(n_573), .C(n_578), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_561), .Y(n_557) );
INVx1_ASAP7_75t_L g636 ( .A(n_558), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_558), .B(n_632), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_558), .B(n_720), .Y(n_719) );
AND2x4_ASAP7_75t_L g558 ( .A(n_559), .B(n_560), .Y(n_558) );
NOR2xp67_ASAP7_75t_SL g604 ( .A(n_560), .B(n_605), .Y(n_604) );
HB1xp67_ASAP7_75t_L g617 ( .A(n_560), .Y(n_617) );
AND2x4_ASAP7_75t_SL g701 ( .A(n_560), .B(n_702), .Y(n_701) );
OR2x2_ASAP7_75t_L g748 ( .A(n_560), .B(n_749), .Y(n_748) );
HB1xp67_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx3_ASAP7_75t_L g622 ( .A(n_562), .Y(n_622) );
INVx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
HB1xp67_ASAP7_75t_L g759 ( .A(n_563), .Y(n_759) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
AOI221x1_ASAP7_75t_L g712 ( .A1(n_565), .A2(n_713), .B1(n_715), .B2(n_716), .C(n_718), .Y(n_712) );
AND2x2_ASAP7_75t_L g638 ( .A(n_566), .B(n_594), .Y(n_638) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
OR2x2_ASAP7_75t_L g568 ( .A(n_569), .B(n_570), .Y(n_568) );
AND2x2_ASAP7_75t_L g581 ( .A(n_569), .B(n_582), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_569), .B(n_571), .Y(n_755) );
INVx2_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx2_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_575), .B(n_577), .Y(n_574) );
AND2x2_ASAP7_75t_SL g579 ( .A(n_575), .B(n_580), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_575), .B(n_588), .Y(n_605) );
INVx2_ASAP7_75t_L g612 ( .A(n_575), .Y(n_612) );
INVx1_ASAP7_75t_L g674 ( .A(n_576), .Y(n_674) );
BUFx2_ASAP7_75t_L g694 ( .A(n_577), .Y(n_694) );
NAND2xp33_ASAP7_75t_SL g578 ( .A(n_579), .B(n_581), .Y(n_578) );
OR2x6_ASAP7_75t_L g611 ( .A(n_580), .B(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g740 ( .A(n_580), .B(n_632), .Y(n_740) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_585), .B(n_603), .Y(n_584) );
AOI22xp5_ASAP7_75t_L g585 ( .A1(n_586), .A2(n_592), .B1(n_596), .B2(n_601), .Y(n_585) );
NOR2xp33_ASAP7_75t_L g586 ( .A(n_587), .B(n_590), .Y(n_586) );
AND2x2_ASAP7_75t_SL g649 ( .A(n_587), .B(n_591), .Y(n_649) );
AND2x4_ASAP7_75t_L g715 ( .A(n_587), .B(n_673), .Y(n_715) );
AND2x4_ASAP7_75t_SL g587 ( .A(n_588), .B(n_589), .Y(n_587) );
HB1xp67_ASAP7_75t_L g730 ( .A(n_588), .Y(n_730) );
INVx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g630 ( .A(n_591), .B(n_631), .Y(n_630) );
HB1xp67_ASAP7_75t_L g683 ( .A(n_591), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_591), .B(n_622), .Y(n_714) );
AND2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
AND2x2_ASAP7_75t_L g735 ( .A(n_593), .B(n_654), .Y(n_735) );
INVx3_ASAP7_75t_L g646 ( .A(n_594), .Y(n_646) );
AND2x2_ASAP7_75t_L g667 ( .A(n_594), .B(n_619), .Y(n_667) );
NAND2x1_ASAP7_75t_SL g738 ( .A(n_594), .B(n_645), .Y(n_738) );
AND2x2_ASAP7_75t_L g596 ( .A(n_597), .B(n_598), .Y(n_596) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
AOI22xp5_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_606), .B1(n_610), .B2(n_613), .Y(n_603) );
BUFx2_ASAP7_75t_L g659 ( .A(n_605), .Y(n_659) );
AOI22xp33_ASAP7_75t_L g705 ( .A1(n_606), .A2(n_697), .B1(n_706), .B2(n_707), .Y(n_705) );
AND2x2_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .Y(n_606) );
NAND2x1p5_ASAP7_75t_L g662 ( .A(n_607), .B(n_663), .Y(n_662) );
AND2x2_ASAP7_75t_L g627 ( .A(n_608), .B(n_628), .Y(n_627) );
INVx2_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
NAND3xp33_ASAP7_75t_L g691 ( .A(n_612), .B(n_692), .C(n_694), .Y(n_691) );
INVx1_ASAP7_75t_L g647 ( .A(n_613), .Y(n_647) );
AOI211x1_ASAP7_75t_L g614 ( .A1(n_615), .A2(n_623), .B(n_625), .C(n_643), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_617), .B(n_618), .Y(n_616) );
NAND2xp5_ASAP7_75t_SL g725 ( .A(n_618), .B(n_706), .Y(n_725) );
AND2x2_ASAP7_75t_L g618 ( .A(n_619), .B(n_621), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_619), .B(n_654), .Y(n_653) );
AND2x2_ASAP7_75t_L g697 ( .A(n_619), .B(n_655), .Y(n_697) );
AND2x2_ASAP7_75t_L g752 ( .A(n_619), .B(n_753), .Y(n_752) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g675 ( .A(n_622), .Y(n_675) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
OR2x2_ASAP7_75t_L g717 ( .A(n_624), .B(n_662), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_626), .B(n_637), .Y(n_625) );
AOI22xp5_ASAP7_75t_SL g626 ( .A1(n_627), .A2(n_630), .B1(n_633), .B2(n_635), .Y(n_626) );
BUFx2_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
AND2x2_ASAP7_75t_L g690 ( .A(n_629), .B(n_685), .Y(n_690) );
INVx1_ASAP7_75t_SL g732 ( .A(n_629), .Y(n_732) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
AND2x2_ASAP7_75t_SL g700 ( .A(n_632), .B(n_701), .Y(n_700) );
INVx3_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVxp67_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
HB1xp67_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
AND2x2_ASAP7_75t_L g736 ( .A(n_641), .B(n_658), .Y(n_736) );
AOI21xp5_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_647), .B(n_648), .Y(n_643) );
OR2x2_ASAP7_75t_L g644 ( .A(n_645), .B(n_646), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_645), .B(n_690), .Y(n_689) );
OR2x2_ASAP7_75t_L g660 ( .A(n_646), .B(n_661), .Y(n_660) );
INVx1_ASAP7_75t_SL g648 ( .A(n_649), .Y(n_648) );
INVxp67_ASAP7_75t_SL g790 ( .A(n_650), .Y(n_790) );
NAND3x1_ASAP7_75t_L g650 ( .A(n_651), .B(n_687), .C(n_695), .Y(n_650) );
NAND4xp25_ASAP7_75t_L g761 ( .A(n_651), .B(n_687), .C(n_695), .D(n_762), .Y(n_761) );
NOR2x1_ASAP7_75t_L g651 ( .A(n_652), .B(n_665), .Y(n_651) );
OAI222xp33_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_656), .B1(n_659), .B2(n_660), .C1(n_662), .C2(n_664), .Y(n_652) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
OAI21xp5_ASAP7_75t_SL g739 ( .A1(n_657), .A2(n_740), .B(n_741), .Y(n_739) );
NAND2xp5_ASAP7_75t_SL g722 ( .A(n_658), .B(n_673), .Y(n_722) );
OAI22xp5_ASAP7_75t_L g718 ( .A1(n_661), .A2(n_719), .B1(n_721), .B2(n_722), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_666), .B(n_676), .Y(n_665) );
NAND2xp5_ASAP7_75t_SL g666 ( .A(n_667), .B(n_668), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_669), .B(n_671), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_669), .B(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_672), .B(n_675), .Y(n_671) );
INVx2_ASAP7_75t_SL g672 ( .A(n_673), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_673), .B(n_675), .Y(n_678) );
INVx2_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
AOI22xp5_ASAP7_75t_L g676 ( .A1(n_677), .A2(n_679), .B1(n_683), .B2(n_684), .Y(n_676) );
AND2x4_ASAP7_75t_L g679 ( .A(n_680), .B(n_681), .Y(n_679) );
AND2x2_ASAP7_75t_L g684 ( .A(n_680), .B(n_685), .Y(n_684) );
NAND2xp5_ASAP7_75t_SL g687 ( .A(n_688), .B(n_691), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g721 ( .A(n_690), .Y(n_721) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
AND2x2_ASAP7_75t_L g695 ( .A(n_696), .B(n_705), .Y(n_695) );
AOI22xp5_ASAP7_75t_SL g696 ( .A1(n_697), .A2(n_698), .B1(n_700), .B2(n_703), .Y(n_696) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVxp67_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
NAND2xp33_ASAP7_75t_L g710 ( .A(n_709), .B(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g789 ( .A(n_711), .Y(n_789) );
NAND3x1_ASAP7_75t_L g711 ( .A(n_712), .B(n_723), .C(n_743), .Y(n_711) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
AOI22xp5_ASAP7_75t_L g734 ( .A1(n_715), .A2(n_735), .B1(n_736), .B2(n_737), .Y(n_734) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_SL g749 ( .A(n_720), .Y(n_749) );
NOR2x1_ASAP7_75t_L g723 ( .A(n_724), .B(n_733), .Y(n_723) );
AOI21xp5_ASAP7_75t_SL g724 ( .A1(n_725), .A2(n_726), .B(n_732), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_727), .B(n_728), .Y(n_726) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_730), .B(n_731), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_734), .B(n_739), .Y(n_733) );
INVx2_ASAP7_75t_SL g737 ( .A(n_738), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_738), .B(n_751), .Y(n_750) );
INVx1_ASAP7_75t_SL g741 ( .A(n_742), .Y(n_741) );
AOI221xp5_ASAP7_75t_L g743 ( .A1(n_744), .A2(n_745), .B1(n_747), .B2(n_750), .C(n_754), .Y(n_743) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVxp67_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx2_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
AOI21xp5_ASAP7_75t_L g754 ( .A1(n_755), .A2(n_756), .B(n_758), .Y(n_754) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
NOR2xp33_ASAP7_75t_L g762 ( .A(n_763), .B(n_764), .Y(n_762) );
INVx3_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
NAND2xp5_ASAP7_75t_SL g769 ( .A(n_770), .B(n_775), .Y(n_769) );
INVxp67_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
AOI21xp33_ASAP7_75t_SL g781 ( .A1(n_771), .A2(n_772), .B(n_782), .Y(n_781) );
NOR2xp33_ASAP7_75t_SL g771 ( .A(n_772), .B(n_774), .Y(n_771) );
BUFx2_ASAP7_75t_R g772 ( .A(n_773), .Y(n_772) );
CKINVDCx11_ASAP7_75t_R g775 ( .A(n_776), .Y(n_775) );
BUFx3_ASAP7_75t_L g780 ( .A(n_776), .Y(n_780) );
CKINVDCx20_ASAP7_75t_R g776 ( .A(n_777), .Y(n_776) );
HB1xp67_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_780), .B(n_781), .Y(n_779) );
OAI22xp5_ASAP7_75t_L g782 ( .A1(n_783), .A2(n_784), .B1(n_786), .B2(n_787), .Y(n_782) );
INVx1_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
INVx1_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
AND3x2_ASAP7_75t_L g787 ( .A(n_788), .B(n_789), .C(n_790), .Y(n_787) );
CKINVDCx5p33_ASAP7_75t_R g791 ( .A(n_792), .Y(n_791) );
INVx2_ASAP7_75t_L g799 ( .A(n_792), .Y(n_799) );
INVx3_ASAP7_75t_SL g792 ( .A(n_793), .Y(n_792) );
AND2x2_ASAP7_75t_SL g793 ( .A(n_794), .B(n_795), .Y(n_793) );
INVx1_ASAP7_75t_SL g798 ( .A(n_799), .Y(n_798) );
endmodule