module fake_jpeg_13925_n_557 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_557);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_557;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_18),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx24_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

BUFx16f_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

CKINVDCx14_ASAP7_75t_R g42 ( 
.A(n_2),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_8),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_R g51 ( 
.A(n_14),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

INVx11_ASAP7_75t_SL g53 ( 
.A(n_7),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_2),
.B(n_12),
.Y(n_54)
);

CKINVDCx14_ASAP7_75t_R g55 ( 
.A(n_3),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_5),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_15),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_58),
.Y(n_134)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_59),
.Y(n_131)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_60),
.Y(n_139)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g180 ( 
.A(n_61),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_62),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g133 ( 
.A(n_63),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_64),
.Y(n_165)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_65),
.Y(n_138)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_66),
.Y(n_161)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_29),
.Y(n_67)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_67),
.Y(n_136)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_68),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_26),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_69),
.Y(n_175)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_33),
.Y(n_70)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_70),
.Y(n_140)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_24),
.Y(n_71)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_71),
.Y(n_149)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_30),
.Y(n_72)
);

INVx5_ASAP7_75t_SL g177 ( 
.A(n_72),
.Y(n_177)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_24),
.Y(n_73)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_73),
.Y(n_151)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_30),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g186 ( 
.A(n_74),
.Y(n_186)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_33),
.Y(n_75)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_75),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_26),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_76),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_28),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_77),
.Y(n_189)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_24),
.Y(n_78)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_78),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_33),
.Y(n_79)
);

INVx5_ASAP7_75t_L g194 ( 
.A(n_79),
.Y(n_194)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_21),
.Y(n_80)
);

INVx5_ASAP7_75t_L g195 ( 
.A(n_80),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_28),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_81),
.Y(n_207)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_33),
.Y(n_82)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_82),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_28),
.Y(n_83)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_83),
.Y(n_150)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_21),
.Y(n_84)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_84),
.Y(n_163)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_21),
.Y(n_85)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_85),
.Y(n_199)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_23),
.Y(n_86)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_86),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_22),
.Y(n_87)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_87),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_28),
.Y(n_88)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_88),
.Y(n_166)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_20),
.Y(n_89)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_89),
.Y(n_190)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_23),
.Y(n_90)
);

INVx6_ASAP7_75t_L g188 ( 
.A(n_90),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_38),
.Y(n_91)
);

INVx6_ASAP7_75t_L g210 ( 
.A(n_91),
.Y(n_210)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_20),
.Y(n_92)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_92),
.Y(n_200)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

INVx8_ASAP7_75t_L g141 ( 
.A(n_93),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_38),
.Y(n_94)
);

INVx8_ASAP7_75t_L g143 ( 
.A(n_94),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_53),
.Y(n_95)
);

INVx13_ASAP7_75t_L g147 ( 
.A(n_95),
.Y(n_147)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_27),
.Y(n_96)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_96),
.Y(n_201)
);

BUFx5_ASAP7_75t_L g97 ( 
.A(n_22),
.Y(n_97)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_97),
.Y(n_206)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_25),
.Y(n_98)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_98),
.Y(n_197)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_41),
.Y(n_99)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_99),
.Y(n_204)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_41),
.Y(n_100)
);

HB1xp67_ASAP7_75t_L g142 ( 
.A(n_100),
.Y(n_142)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_27),
.Y(n_101)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_101),
.Y(n_203)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_25),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g144 ( 
.A(n_102),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_54),
.B(n_0),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_103),
.B(n_118),
.Y(n_129)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_31),
.Y(n_104)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_104),
.Y(n_205)
);

INVx3_ASAP7_75t_SL g105 ( 
.A(n_25),
.Y(n_105)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_105),
.Y(n_137)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_31),
.Y(n_106)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_106),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_38),
.Y(n_107)
);

INVx8_ASAP7_75t_L g202 ( 
.A(n_107),
.Y(n_202)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_38),
.Y(n_108)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_108),
.Y(n_155)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_37),
.B(n_18),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_109),
.B(n_116),
.Y(n_130)
);

INVxp67_ASAP7_75t_SL g110 ( 
.A(n_41),
.Y(n_110)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_110),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_22),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_111),
.B(n_115),
.Y(n_162)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_37),
.Y(n_112)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_112),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_40),
.Y(n_113)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_113),
.Y(n_185)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_35),
.Y(n_114)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_114),
.Y(n_193)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_39),
.Y(n_115)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_40),
.Y(n_116)
);

INVx3_ASAP7_75t_SL g117 ( 
.A(n_40),
.Y(n_117)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_117),
.Y(n_192)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_40),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_39),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_119),
.B(n_120),
.Y(n_153)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_43),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_43),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_121),
.B(n_122),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_47),
.Y(n_122)
);

BUFx24_ASAP7_75t_L g123 ( 
.A(n_42),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_123),
.B(n_51),
.Y(n_172)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_45),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_124),
.B(n_125),
.Y(n_174)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_47),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_61),
.A2(n_35),
.B1(n_44),
.B2(n_47),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_126),
.A2(n_128),
.B1(n_145),
.B2(n_146),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_123),
.A2(n_23),
.B1(n_50),
.B2(n_55),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_127),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_66),
.A2(n_35),
.B1(n_44),
.B2(n_56),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_103),
.A2(n_54),
.B1(n_50),
.B2(n_19),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_132),
.A2(n_135),
.B1(n_196),
.B2(n_94),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_109),
.A2(n_50),
.B1(n_19),
.B2(n_44),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_110),
.A2(n_47),
.B1(n_56),
.B2(n_45),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_60),
.A2(n_56),
.B1(n_46),
.B2(n_49),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_58),
.A2(n_56),
.B1(n_46),
.B2(n_49),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_156),
.A2(n_158),
.B1(n_159),
.B2(n_211),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_80),
.A2(n_52),
.B1(n_48),
.B2(n_57),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_114),
.A2(n_52),
.B1(n_48),
.B2(n_57),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_95),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_168),
.B(n_178),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_105),
.A2(n_55),
.B1(n_51),
.B2(n_42),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_171),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_172),
.B(n_130),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_85),
.B(n_34),
.Y(n_178)
);

OA22x2_ASAP7_75t_L g179 ( 
.A1(n_62),
.A2(n_34),
.B1(n_32),
.B2(n_41),
.Y(n_179)
);

OAI32xp33_ASAP7_75t_L g264 ( 
.A1(n_179),
.A2(n_13),
.A3(n_15),
.B1(n_16),
.B2(n_180),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_117),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_181),
.B(n_182),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_118),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_125),
.B(n_32),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_184),
.B(n_191),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_64),
.B(n_18),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_187),
.B(n_208),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_69),
.B(n_17),
.Y(n_191)
);

OAI22xp33_ASAP7_75t_L g196 ( 
.A1(n_76),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_77),
.B(n_3),
.C(n_5),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_198),
.B(n_179),
.C(n_145),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_81),
.B(n_5),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_83),
.B(n_5),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_209),
.B(n_10),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_88),
.A2(n_122),
.B1(n_113),
.B2(n_107),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_134),
.Y(n_212)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_212),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_214),
.B(n_223),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_142),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_215),
.B(n_230),
.Y(n_290)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_154),
.Y(n_216)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_216),
.Y(n_284)
);

BUFx10_ASAP7_75t_L g217 ( 
.A(n_192),
.Y(n_217)
);

BUFx24_ASAP7_75t_L g325 ( 
.A(n_217),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_129),
.A2(n_91),
.B1(n_7),
.B2(n_8),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_218),
.A2(n_250),
.B1(n_264),
.B2(n_269),
.Y(n_309)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_155),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g292 ( 
.A(n_219),
.Y(n_292)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_176),
.Y(n_220)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_220),
.Y(n_291)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_137),
.Y(n_221)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_221),
.Y(n_293)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_170),
.Y(n_222)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_222),
.Y(n_289)
);

AND2x2_ASAP7_75t_SL g223 ( 
.A(n_153),
.B(n_6),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_149),
.Y(n_224)
);

INVx3_ASAP7_75t_L g315 ( 
.A(n_224),
.Y(n_315)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_195),
.Y(n_225)
);

INVx4_ASAP7_75t_L g314 ( 
.A(n_225),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_196),
.A2(n_6),
.B1(n_9),
.B2(n_10),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_227),
.A2(n_228),
.B1(n_252),
.B2(n_258),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_174),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_228)
);

BUFx2_ASAP7_75t_L g229 ( 
.A(n_164),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_229),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_142),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_231),
.B(n_235),
.Y(n_299)
);

BUFx2_ASAP7_75t_L g232 ( 
.A(n_164),
.Y(n_232)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_232),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_160),
.B(n_9),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_233),
.B(n_240),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_144),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_162),
.B(n_16),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_236),
.B(n_238),
.Y(n_310)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_141),
.Y(n_237)
);

INVx4_ASAP7_75t_L g331 ( 
.A(n_237),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_177),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_144),
.Y(n_241)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_241),
.Y(n_305)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_190),
.Y(n_242)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_242),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_204),
.B(n_11),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_243),
.B(n_248),
.Y(n_319)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_200),
.Y(n_244)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_244),
.Y(n_317)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_201),
.Y(n_245)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_245),
.Y(n_332)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_151),
.Y(n_246)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_246),
.Y(n_334)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_203),
.Y(n_247)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_247),
.Y(n_335)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_185),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_136),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_249),
.B(n_254),
.Y(n_327)
);

OAI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_158),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_197),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_251),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_173),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_252)
);

INVx8_ASAP7_75t_L g253 ( 
.A(n_157),
.Y(n_253)
);

INVx6_ASAP7_75t_L g287 ( 
.A(n_253),
.Y(n_287)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_167),
.Y(n_254)
);

INVx4_ASAP7_75t_L g255 ( 
.A(n_133),
.Y(n_255)
);

BUFx4f_ASAP7_75t_L g318 ( 
.A(n_255),
.Y(n_318)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_141),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g294 ( 
.A1(n_256),
.A2(n_257),
.B1(n_262),
.B2(n_263),
.Y(n_294)
);

INVx5_ASAP7_75t_L g257 ( 
.A(n_163),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_162),
.A2(n_205),
.B1(n_179),
.B2(n_188),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_147),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_260),
.Y(n_312)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_148),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_261),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_157),
.Y(n_262)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_199),
.Y(n_263)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_169),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_265),
.A2(n_266),
.B1(n_268),
.B2(n_272),
.Y(n_302)
);

BUFx2_ASAP7_75t_L g266 ( 
.A(n_161),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_267),
.B(n_165),
.C(n_175),
.Y(n_313)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_140),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_211),
.A2(n_159),
.B1(n_126),
.B2(n_128),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_152),
.B(n_15),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_271),
.B(n_281),
.Y(n_295)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_188),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_131),
.B(n_138),
.Y(n_273)
);

NOR2x1_ASAP7_75t_L g333 ( 
.A(n_273),
.B(n_282),
.Y(n_333)
);

CKINVDCx6p67_ASAP7_75t_R g274 ( 
.A(n_147),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g303 ( 
.A1(n_274),
.A2(n_275),
.B1(n_276),
.B2(n_277),
.Y(n_303)
);

INVx5_ASAP7_75t_L g275 ( 
.A(n_163),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_206),
.A2(n_180),
.B1(n_194),
.B2(n_193),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_210),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_210),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_SL g326 ( 
.A1(n_278),
.A2(n_279),
.B1(n_183),
.B2(n_189),
.Y(n_326)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_150),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_177),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_156),
.Y(n_282)
);

A2O1A1Ixp33_ASAP7_75t_L g288 ( 
.A1(n_230),
.A2(n_146),
.B(n_186),
.C(n_139),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_288),
.B(n_297),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_223),
.B(n_213),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_270),
.A2(n_186),
.B(n_133),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_298),
.A2(n_275),
.B(n_257),
.Y(n_346)
);

AOI22xp33_ASAP7_75t_L g301 ( 
.A1(n_234),
.A2(n_202),
.B1(n_143),
.B2(n_150),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_301),
.A2(n_322),
.B1(n_330),
.B2(n_336),
.Y(n_369)
);

O2A1O1Ixp33_ASAP7_75t_SL g304 ( 
.A1(n_270),
.A2(n_143),
.B(n_202),
.C(n_206),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_304),
.B(n_274),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_223),
.B(n_267),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_306),
.B(n_313),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_226),
.B(n_166),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_307),
.B(n_311),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_228),
.B(n_236),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_252),
.B(n_166),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_320),
.B(n_328),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_280),
.A2(n_165),
.B1(n_175),
.B2(n_183),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_326),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_264),
.B(n_189),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_214),
.B(n_207),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_329),
.B(n_253),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_258),
.A2(n_259),
.B1(n_283),
.B2(n_227),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_L g336 ( 
.A1(n_217),
.A2(n_133),
.B1(n_207),
.B2(n_259),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_272),
.A2(n_276),
.B1(n_239),
.B2(n_261),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_337),
.A2(n_238),
.B1(n_232),
.B2(n_229),
.Y(n_340)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_293),
.Y(n_338)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_338),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_328),
.A2(n_217),
.B1(n_266),
.B2(n_225),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g382 ( 
.A1(n_339),
.A2(n_340),
.B(n_346),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_343),
.B(n_352),
.Y(n_386)
);

BUFx24_ASAP7_75t_L g344 ( 
.A(n_325),
.Y(n_344)
);

BUFx3_ASAP7_75t_L g408 ( 
.A(n_344),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_292),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_345),
.B(n_363),
.Y(n_383)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_293),
.Y(n_347)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_347),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_306),
.B(n_221),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_348),
.B(n_360),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_SL g349 ( 
.A1(n_333),
.A2(n_274),
.B(n_219),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g379 ( 
.A1(n_349),
.A2(n_354),
.B(n_303),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_309),
.A2(n_329),
.B1(n_330),
.B2(n_300),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_350),
.A2(n_353),
.B1(n_355),
.B2(n_357),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_297),
.B(n_249),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_309),
.A2(n_248),
.B1(n_262),
.B2(n_265),
.Y(n_353)
);

OAI22xp33_ASAP7_75t_SL g355 ( 
.A1(n_333),
.A2(n_237),
.B1(n_256),
.B2(n_263),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_SL g356 ( 
.A(n_300),
.B(n_212),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_356),
.B(n_289),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_300),
.A2(n_255),
.B1(n_313),
.B2(n_320),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_307),
.B(n_312),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_358),
.B(n_365),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_311),
.A2(n_298),
.B1(n_323),
.B2(n_304),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_359),
.A2(n_357),
.B1(n_369),
.B2(n_342),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_290),
.B(n_310),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_299),
.B(n_322),
.Y(n_361)
);

CKINVDCx14_ASAP7_75t_R g393 ( 
.A(n_361),
.Y(n_393)
);

CKINVDCx16_ASAP7_75t_R g363 ( 
.A(n_325),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_323),
.A2(n_337),
.B1(n_304),
.B2(n_288),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_364),
.A2(n_367),
.B1(n_368),
.B2(n_296),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_295),
.B(n_319),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_295),
.B(n_308),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_366),
.B(n_370),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_284),
.A2(n_291),
.B1(n_335),
.B2(n_317),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_284),
.A2(n_291),
.B1(n_335),
.B2(n_317),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_327),
.B(n_332),
.Y(n_370)
);

INVx1_ASAP7_75t_SL g371 ( 
.A(n_325),
.Y(n_371)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_371),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_285),
.B(n_305),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_372),
.B(n_375),
.Y(n_409)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_316),
.Y(n_373)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_373),
.Y(n_395)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_316),
.Y(n_374)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_374),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_305),
.B(n_332),
.Y(n_375)
);

AOI22xp33_ASAP7_75t_L g376 ( 
.A1(n_324),
.A2(n_314),
.B1(n_331),
.B2(n_334),
.Y(n_376)
);

AOI22xp33_ASAP7_75t_SL g391 ( 
.A1(n_376),
.A2(n_296),
.B1(n_287),
.B2(n_321),
.Y(n_391)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_334),
.Y(n_378)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_378),
.Y(n_405)
);

AOI21xp5_ASAP7_75t_L g439 ( 
.A1(n_379),
.A2(n_397),
.B(n_401),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_L g380 ( 
.A1(n_341),
.A2(n_302),
.B(n_294),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_L g413 ( 
.A1(n_380),
.A2(n_406),
.B(n_410),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_385),
.A2(n_407),
.B1(n_361),
.B2(n_356),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_364),
.A2(n_287),
.B1(n_331),
.B2(n_314),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_387),
.B(n_389),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_L g389 ( 
.A1(n_362),
.A2(n_339),
.B1(n_354),
.B2(n_341),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_367),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_390),
.B(n_370),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g437 ( 
.A(n_391),
.Y(n_437)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_349),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_392),
.B(n_360),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_396),
.B(n_410),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_SL g397 ( 
.A1(n_346),
.A2(n_286),
.B(n_318),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_362),
.A2(n_289),
.B1(n_315),
.B2(n_286),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_398),
.B(n_403),
.Y(n_422)
);

AOI22xp33_ASAP7_75t_SL g401 ( 
.A1(n_377),
.A2(n_321),
.B1(n_315),
.B2(n_318),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_351),
.A2(n_318),
.B1(n_350),
.B2(n_358),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_404),
.A2(n_366),
.B1(n_374),
.B2(n_373),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_359),
.A2(n_361),
.B1(n_369),
.B2(n_353),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_L g407 ( 
.A1(n_351),
.A2(n_343),
.B1(n_340),
.B2(n_365),
.Y(n_407)
);

AND2x2_ASAP7_75t_SL g410 ( 
.A(n_342),
.B(n_348),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_412),
.A2(n_384),
.B1(n_380),
.B2(n_386),
.Y(n_443)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_414),
.Y(n_449)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_395),
.Y(n_415)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_415),
.Y(n_457)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_395),
.Y(n_416)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_416),
.Y(n_464)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_402),
.Y(n_417)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_417),
.Y(n_467)
);

OAI21xp5_ASAP7_75t_L g419 ( 
.A1(n_379),
.A2(n_372),
.B(n_375),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_L g446 ( 
.A1(n_419),
.A2(n_397),
.B(n_382),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_409),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_420),
.B(n_428),
.Y(n_455)
);

INVxp67_ASAP7_75t_L g463 ( 
.A(n_421),
.Y(n_463)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_402),
.Y(n_423)
);

INVx1_ASAP7_75t_SL g460 ( 
.A(n_423),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_400),
.B(n_352),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_SL g442 ( 
.A(n_424),
.B(n_388),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_410),
.B(n_399),
.C(n_396),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_425),
.B(n_427),
.C(n_432),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_SL g451 ( 
.A(n_426),
.B(n_386),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_399),
.B(n_356),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_409),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_429),
.A2(n_430),
.B1(n_433),
.B2(n_411),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_406),
.A2(n_368),
.B1(n_338),
.B2(n_347),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_405),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_431),
.B(n_434),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_410),
.B(n_378),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_406),
.A2(n_404),
.B1(n_384),
.B2(n_390),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_383),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_388),
.B(n_345),
.Y(n_435)
);

NAND3xp33_ASAP7_75t_L g447 ( 
.A(n_435),
.B(n_440),
.C(n_424),
.Y(n_447)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_405),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_436),
.B(n_441),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_396),
.B(n_371),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_438),
.B(n_407),
.C(n_403),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_400),
.B(n_363),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_381),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_442),
.B(n_447),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_443),
.B(n_451),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_445),
.B(n_448),
.C(n_459),
.Y(n_474)
);

OAI21xp5_ASAP7_75t_L g481 ( 
.A1(n_446),
.A2(n_439),
.B(n_401),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_425),
.B(n_389),
.C(n_385),
.Y(n_448)
);

OR2x2_ASAP7_75t_L g450 ( 
.A(n_430),
.B(n_382),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_450),
.Y(n_476)
);

INVxp67_ASAP7_75t_SL g452 ( 
.A(n_419),
.Y(n_452)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_452),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_420),
.B(n_383),
.Y(n_453)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_453),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_422),
.Y(n_454)
);

AOI22xp33_ASAP7_75t_L g485 ( 
.A1(n_454),
.A2(n_415),
.B1(n_423),
.B2(n_417),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_428),
.B(n_398),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_456),
.B(n_458),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_434),
.B(n_394),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_426),
.B(n_387),
.C(n_393),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_SL g461 ( 
.A(n_429),
.B(n_394),
.Y(n_461)
);

CKINVDCx16_ASAP7_75t_R g487 ( 
.A(n_461),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_432),
.B(n_393),
.C(n_381),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_462),
.B(n_427),
.C(n_441),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_L g470 ( 
.A1(n_468),
.A2(n_418),
.B1(n_412),
.B2(n_422),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_443),
.A2(n_433),
.B1(n_418),
.B2(n_413),
.Y(n_469)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_469),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_470),
.A2(n_486),
.B1(n_490),
.B2(n_460),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_454),
.A2(n_413),
.B1(n_437),
.B2(n_439),
.Y(n_472)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_472),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_444),
.B(n_438),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_473),
.B(n_480),
.Y(n_493)
);

HB1xp67_ASAP7_75t_L g475 ( 
.A(n_449),
.Y(n_475)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_475),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_466),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_479),
.B(n_484),
.Y(n_492)
);

OR2x6_ASAP7_75t_SL g494 ( 
.A(n_481),
.B(n_459),
.Y(n_494)
);

OAI21xp5_ASAP7_75t_L g484 ( 
.A1(n_446),
.A2(n_411),
.B(n_436),
.Y(n_484)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_485),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_461),
.A2(n_416),
.B1(n_431),
.B2(n_408),
.Y(n_486)
);

AOI21xp5_ASAP7_75t_L g488 ( 
.A1(n_450),
.A2(n_391),
.B(n_371),
.Y(n_488)
);

INVxp67_ASAP7_75t_SL g505 ( 
.A(n_488),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_444),
.B(n_344),
.C(n_408),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_489),
.B(n_448),
.C(n_462),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_455),
.A2(n_344),
.B1(n_408),
.B2(n_445),
.Y(n_490)
);

AOI21xp5_ASAP7_75t_L g513 ( 
.A1(n_494),
.A2(n_472),
.B(n_481),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_SL g495 ( 
.A(n_471),
.B(n_451),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g519 ( 
.A(n_495),
.B(n_497),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_SL g507 ( 
.A1(n_499),
.A2(n_469),
.B1(n_468),
.B2(n_450),
.Y(n_507)
);

CKINVDCx14_ASAP7_75t_R g500 ( 
.A(n_478),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_500),
.B(n_449),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_SL g501 ( 
.A(n_471),
.B(n_455),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_501),
.B(n_502),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_482),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_482),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_503),
.B(n_458),
.Y(n_512)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_473),
.B(n_453),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_504),
.B(n_480),
.C(n_474),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_507),
.A2(n_498),
.B1(n_496),
.B2(n_476),
.Y(n_523)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_496),
.A2(n_487),
.B1(n_470),
.B2(n_483),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_SL g530 ( 
.A1(n_508),
.A2(n_477),
.B1(n_476),
.B2(n_494),
.Y(n_530)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_491),
.Y(n_509)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_509),
.Y(n_528)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_492),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_510),
.B(n_512),
.Y(n_529)
);

AOI21x1_ASAP7_75t_L g525 ( 
.A1(n_513),
.A2(n_488),
.B(n_498),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_SL g521 ( 
.A1(n_514),
.A2(n_465),
.B1(n_477),
.B2(n_506),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_515),
.B(n_493),
.Y(n_520)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_492),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_L g524 ( 
.A1(n_516),
.A2(n_518),
.B1(n_505),
.B2(n_506),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_493),
.B(n_474),
.C(n_489),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_517),
.B(n_497),
.C(n_504),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_L g518 ( 
.A1(n_499),
.A2(n_487),
.B1(n_483),
.B2(n_479),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_520),
.B(n_522),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_521),
.B(n_524),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_L g534 ( 
.A1(n_523),
.A2(n_510),
.B1(n_516),
.B2(n_513),
.Y(n_534)
);

OAI21xp5_ASAP7_75t_L g539 ( 
.A1(n_525),
.A2(n_456),
.B(n_501),
.Y(n_539)
);

XNOR2xp5_ASAP7_75t_L g526 ( 
.A(n_515),
.B(n_517),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_526),
.B(n_527),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_L g527 ( 
.A(n_508),
.B(n_490),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_530),
.B(n_465),
.Y(n_537)
);

AOI21xp5_ASAP7_75t_SL g532 ( 
.A1(n_529),
.A2(n_514),
.B(n_511),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_532),
.B(n_442),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_534),
.B(n_537),
.Y(n_546)
);

AOI21xp5_ASAP7_75t_L g535 ( 
.A1(n_526),
.A2(n_519),
.B(n_494),
.Y(n_535)
);

AOI21xp5_ASAP7_75t_L g540 ( 
.A1(n_535),
.A2(n_536),
.B(n_539),
.Y(n_540)
);

OAI21xp5_ASAP7_75t_L g536 ( 
.A1(n_522),
.A2(n_507),
.B(n_484),
.Y(n_536)
);

INVx1_ASAP7_75t_SL g541 ( 
.A(n_531),
.Y(n_541)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_541),
.Y(n_548)
);

AOI22xp5_ASAP7_75t_SL g542 ( 
.A1(n_533),
.A2(n_463),
.B1(n_527),
.B2(n_528),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_542),
.B(n_486),
.C(n_495),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_SL g543 ( 
.A(n_538),
.B(n_520),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_543),
.B(n_523),
.Y(n_547)
);

NOR2xp67_ASAP7_75t_SL g549 ( 
.A(n_544),
.B(n_545),
.Y(n_549)
);

NOR2xp67_ASAP7_75t_SL g545 ( 
.A(n_533),
.B(n_519),
.Y(n_545)
);

INVxp67_ASAP7_75t_SL g551 ( 
.A(n_547),
.Y(n_551)
);

AOI211x1_ASAP7_75t_L g552 ( 
.A1(n_550),
.A2(n_540),
.B(n_549),
.C(n_546),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_552),
.B(n_548),
.C(n_466),
.Y(n_553)
);

OAI21xp5_ASAP7_75t_SL g554 ( 
.A1(n_553),
.A2(n_551),
.B(n_460),
.Y(n_554)
);

A2O1A1O1Ixp25_ASAP7_75t_L g555 ( 
.A1(n_554),
.A2(n_467),
.B(n_457),
.C(n_464),
.D(n_344),
.Y(n_555)
);

AOI21xp5_ASAP7_75t_SL g556 ( 
.A1(n_555),
.A2(n_457),
.B(n_464),
.Y(n_556)
);

OAI21xp33_ASAP7_75t_L g557 ( 
.A1(n_556),
.A2(n_467),
.B(n_460),
.Y(n_557)
);


endmodule