module real_aes_2678_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_793, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_793;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_635;
wire n_503;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_666;
wire n_551;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_746;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_769;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_617;
wire n_552;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_288;
wire n_147;
wire n_756;
wire n_150;
wire n_404;
wire n_598;
wire n_728;
wire n_713;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_789;
wire n_268;
wire n_544;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_753;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_SL g178 ( .A(n_0), .B(n_136), .Y(n_178) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_1), .A2(n_149), .B(n_228), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g787 ( .A(n_2), .B(n_788), .Y(n_787) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_3), .B(n_136), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_4), .B(n_158), .Y(n_477) );
NAND2xp5_ASAP7_75t_SL g157 ( .A(n_5), .B(n_158), .Y(n_157) );
INVx1_ASAP7_75t_L g143 ( .A(n_6), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_7), .B(n_158), .Y(n_236) );
CKINVDCx16_ASAP7_75t_R g788 ( .A(n_8), .Y(n_788) );
CKINVDCx20_ASAP7_75t_R g790 ( .A(n_9), .Y(n_790) );
NAND2xp33_ASAP7_75t_L g221 ( .A(n_10), .B(n_156), .Y(n_221) );
AND2x2_ASAP7_75t_L g479 ( .A(n_11), .B(n_215), .Y(n_479) );
AND2x2_ASAP7_75t_L g489 ( .A(n_12), .B(n_180), .Y(n_489) );
INVx2_ASAP7_75t_L g147 ( .A(n_13), .Y(n_147) );
AOI221x1_ASAP7_75t_L g165 ( .A1(n_14), .A2(n_25), .B1(n_136), .B2(n_149), .C(n_166), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_15), .B(n_158), .Y(n_539) );
CKINVDCx16_ASAP7_75t_R g116 ( .A(n_16), .Y(n_116) );
AND3x1_ASAP7_75t_L g785 ( .A(n_16), .B(n_37), .C(n_786), .Y(n_785) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_17), .B(n_136), .Y(n_217) );
AO21x2_ASAP7_75t_L g214 ( .A1(n_18), .A2(n_215), .B(n_216), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_19), .B(n_163), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_20), .B(n_158), .Y(n_209) );
AO21x1_ASAP7_75t_L g135 ( .A1(n_21), .A2(n_136), .B(n_144), .Y(n_135) );
NAND2xp5_ASAP7_75t_SL g544 ( .A(n_22), .B(n_136), .Y(n_544) );
INVx1_ASAP7_75t_L g120 ( .A(n_23), .Y(n_120) );
AOI22xp33_ASAP7_75t_L g493 ( .A1(n_24), .A2(n_91), .B1(n_136), .B2(n_494), .Y(n_493) );
NAND2x1_ASAP7_75t_L g176 ( .A(n_26), .B(n_158), .Y(n_176) );
NAND2x1_ASAP7_75t_L g235 ( .A(n_27), .B(n_156), .Y(n_235) );
OR2x2_ASAP7_75t_L g146 ( .A(n_28), .B(n_88), .Y(n_146) );
OA21x2_ASAP7_75t_L g182 ( .A1(n_28), .A2(n_88), .B(n_147), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_29), .B(n_156), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_30), .B(n_158), .Y(n_220) );
AO21x2_ASAP7_75t_L g534 ( .A1(n_31), .A2(n_180), .B(n_535), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_32), .B(n_156), .Y(n_155) );
AOI21xp5_ASAP7_75t_L g474 ( .A1(n_33), .A2(n_149), .B(n_475), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_34), .B(n_158), .Y(n_558) );
AOI21xp5_ASAP7_75t_L g188 ( .A1(n_35), .A2(n_149), .B(n_189), .Y(n_188) );
AND2x2_ASAP7_75t_L g142 ( .A(n_36), .B(n_143), .Y(n_142) );
AND2x2_ASAP7_75t_L g150 ( .A(n_36), .B(n_151), .Y(n_150) );
INVx1_ASAP7_75t_L g502 ( .A(n_36), .Y(n_502) );
OR2x6_ASAP7_75t_L g118 ( .A(n_37), .B(n_119), .Y(n_118) );
NAND2xp5_ASAP7_75t_SL g192 ( .A(n_38), .B(n_136), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_39), .B(n_136), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_40), .B(n_158), .Y(n_531) );
CKINVDCx20_ASAP7_75t_R g213 ( .A(n_41), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_42), .B(n_156), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_43), .B(n_136), .Y(n_465) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_44), .Y(n_122) );
AOI22xp5_ASAP7_75t_SL g750 ( .A1(n_45), .A2(n_66), .B1(n_751), .B2(n_752), .Y(n_750) );
CKINVDCx20_ASAP7_75t_R g751 ( .A(n_45), .Y(n_751) );
AOI22xp5_ASAP7_75t_L g771 ( .A1(n_46), .A2(n_86), .B1(n_772), .B2(n_773), .Y(n_771) );
CKINVDCx20_ASAP7_75t_R g773 ( .A(n_46), .Y(n_773) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_47), .A2(n_149), .B(n_485), .Y(n_484) );
AOI21xp5_ASAP7_75t_L g233 ( .A1(n_48), .A2(n_149), .B(n_234), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_49), .B(n_156), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_50), .B(n_156), .Y(n_177) );
NAND2xp5_ASAP7_75t_SL g536 ( .A(n_51), .B(n_136), .Y(n_536) );
XNOR2xp5_ASAP7_75t_L g749 ( .A(n_52), .B(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g139 ( .A(n_53), .Y(n_139) );
INVx1_ASAP7_75t_L g153 ( .A(n_53), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_54), .B(n_158), .Y(n_487) );
AND2x2_ASAP7_75t_L g526 ( .A(n_55), .B(n_163), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_56), .B(n_156), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_57), .B(n_158), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_58), .B(n_156), .Y(n_557) );
AOI21xp5_ASAP7_75t_L g174 ( .A1(n_59), .A2(n_149), .B(n_175), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g488 ( .A(n_60), .B(n_136), .Y(n_488) );
NAND2xp5_ASAP7_75t_SL g528 ( .A(n_61), .B(n_136), .Y(n_528) );
AOI21xp5_ASAP7_75t_L g555 ( .A1(n_62), .A2(n_149), .B(n_556), .Y(n_555) );
AO21x1_ASAP7_75t_L g148 ( .A1(n_63), .A2(n_149), .B(n_154), .Y(n_148) );
AND2x2_ASAP7_75t_L g550 ( .A(n_64), .B(n_164), .Y(n_550) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_65), .B(n_136), .Y(n_226) );
CKINVDCx20_ASAP7_75t_R g752 ( .A(n_66), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_67), .B(n_156), .Y(n_532) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_68), .B(n_136), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_69), .B(n_156), .Y(n_540) );
AOI22xp5_ASAP7_75t_L g499 ( .A1(n_70), .A2(n_95), .B1(n_149), .B2(n_500), .Y(n_499) );
AND2x2_ASAP7_75t_L g193 ( .A(n_71), .B(n_164), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_72), .B(n_158), .Y(n_547) );
INVx1_ASAP7_75t_L g141 ( .A(n_73), .Y(n_141) );
INVx1_ASAP7_75t_L g151 ( .A(n_73), .Y(n_151) );
AND2x2_ASAP7_75t_L g239 ( .A(n_74), .B(n_180), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_75), .B(n_156), .Y(n_476) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_76), .A2(n_149), .B(n_530), .Y(n_529) );
AOI21xp5_ASAP7_75t_L g466 ( .A1(n_77), .A2(n_149), .B(n_467), .Y(n_466) );
AOI21xp5_ASAP7_75t_L g537 ( .A1(n_78), .A2(n_149), .B(n_538), .Y(n_537) );
AND2x2_ASAP7_75t_L g560 ( .A(n_79), .B(n_164), .Y(n_560) );
CKINVDCx20_ASAP7_75t_R g760 ( .A(n_80), .Y(n_760) );
NAND2xp5_ASAP7_75t_SL g491 ( .A(n_81), .B(n_163), .Y(n_491) );
INVx1_ASAP7_75t_L g121 ( .A(n_82), .Y(n_121) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_83), .B(n_136), .Y(n_211) );
AND2x2_ASAP7_75t_L g224 ( .A(n_84), .B(n_180), .Y(n_224) );
AND2x2_ASAP7_75t_L g470 ( .A(n_85), .B(n_215), .Y(n_470) );
CKINVDCx20_ASAP7_75t_R g772 ( .A(n_86), .Y(n_772) );
AND2x2_ASAP7_75t_L g144 ( .A(n_87), .B(n_145), .Y(n_144) );
AND2x2_ASAP7_75t_L g183 ( .A(n_89), .B(n_180), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_90), .B(n_156), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_92), .B(n_158), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_93), .B(n_156), .Y(n_167) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_94), .A2(n_149), .B(n_208), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g545 ( .A1(n_96), .A2(n_149), .B(n_546), .Y(n_545) );
OAI22xp5_ASAP7_75t_SL g769 ( .A1(n_97), .A2(n_770), .B1(n_771), .B2(n_774), .Y(n_769) );
CKINVDCx20_ASAP7_75t_R g774 ( .A(n_97), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_98), .B(n_158), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_99), .B(n_158), .Y(n_229) );
BUFx2_ASAP7_75t_L g549 ( .A(n_100), .Y(n_549) );
BUFx2_ASAP7_75t_L g108 ( .A(n_101), .Y(n_108) );
BUFx2_ASAP7_75t_SL g765 ( .A(n_101), .Y(n_765) );
AOI21xp5_ASAP7_75t_L g218 ( .A1(n_102), .A2(n_149), .B(n_219), .Y(n_218) );
AOI21xp33_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_779), .B(n_789), .Y(n_103) );
OA21x2_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_123), .B(n_763), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_106), .B(n_109), .Y(n_105) );
HB1xp67_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
HB1xp67_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVxp67_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
AOI21xp5_ASAP7_75t_L g766 ( .A1(n_110), .A2(n_767), .B(n_776), .Y(n_766) );
NOR2xp33_ASAP7_75t_SL g110 ( .A(n_111), .B(n_122), .Y(n_110) );
INVx1_ASAP7_75t_SL g111 ( .A(n_112), .Y(n_111) );
BUFx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g113 ( .A(n_114), .Y(n_113) );
BUFx3_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
BUFx2_ASAP7_75t_R g778 ( .A(n_115), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_116), .B(n_117), .Y(n_115) );
OR2x6_ASAP7_75t_SL g452 ( .A(n_116), .B(n_117), .Y(n_452) );
AND2x6_ASAP7_75t_SL g748 ( .A(n_116), .B(n_118), .Y(n_748) );
OR2x2_ASAP7_75t_L g762 ( .A(n_116), .B(n_118), .Y(n_762) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_L g784 ( .A(n_119), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g119 ( .A(n_120), .B(n_121), .Y(n_119) );
OAI21xp5_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_749), .B(n_753), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
OAI22xp5_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_452), .B1(n_453), .B2(n_747), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
OAI22x1_ASAP7_75t_L g754 ( .A1(n_127), .A2(n_452), .B1(n_755), .B2(n_756), .Y(n_754) );
AND2x4_ASAP7_75t_L g127 ( .A(n_128), .B(n_351), .Y(n_127) );
NOR3xp33_ASAP7_75t_L g128 ( .A(n_129), .B(n_288), .C(n_311), .Y(n_128) );
NAND3xp33_ASAP7_75t_SL g129 ( .A(n_130), .B(n_240), .C(n_257), .Y(n_129) );
OAI31xp33_ASAP7_75t_SL g130 ( .A1(n_131), .A2(n_170), .A3(n_194), .B(n_201), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_131), .B(n_315), .Y(n_314) );
INVx1_ASAP7_75t_SL g131 ( .A(n_132), .Y(n_131) );
OR2x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_162), .Y(n_132) );
AND2x4_ASAP7_75t_L g243 ( .A(n_133), .B(n_162), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_133), .B(n_185), .Y(n_272) );
AND2x4_ASAP7_75t_L g274 ( .A(n_133), .B(n_268), .Y(n_274) );
AND2x2_ASAP7_75t_L g405 ( .A(n_133), .B(n_198), .Y(n_405) );
INVx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx2_ASAP7_75t_L g250 ( .A(n_134), .Y(n_250) );
OAI21x1_ASAP7_75t_SL g134 ( .A1(n_135), .A2(n_148), .B(n_160), .Y(n_134) );
AND2x4_ASAP7_75t_L g136 ( .A(n_137), .B(n_142), .Y(n_136) );
AND2x4_ASAP7_75t_L g137 ( .A(n_138), .B(n_140), .Y(n_137) );
AND2x6_ASAP7_75t_L g156 ( .A(n_138), .B(n_151), .Y(n_156) );
INVx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
AND2x4_ASAP7_75t_L g158 ( .A(n_140), .B(n_153), .Y(n_158) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx5_ASAP7_75t_L g159 ( .A(n_142), .Y(n_159) );
AND2x2_ASAP7_75t_L g152 ( .A(n_143), .B(n_153), .Y(n_152) );
HB1xp67_ASAP7_75t_L g497 ( .A(n_143), .Y(n_497) );
INVx1_ASAP7_75t_L g161 ( .A(n_144), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_145), .B(n_161), .Y(n_160) );
INVx1_ASAP7_75t_SL g205 ( .A(n_145), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_145), .A2(n_217), .B(n_218), .Y(n_216) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_145), .A2(n_528), .B(n_529), .Y(n_527) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_145), .A2(n_536), .B(n_537), .Y(n_535) );
AND2x4_ASAP7_75t_L g145 ( .A(n_146), .B(n_147), .Y(n_145) );
AND2x2_ASAP7_75t_SL g164 ( .A(n_146), .B(n_147), .Y(n_164) );
AND2x6_ASAP7_75t_L g149 ( .A(n_150), .B(n_152), .Y(n_149) );
BUFx3_ASAP7_75t_L g498 ( .A(n_150), .Y(n_498) );
INVx2_ASAP7_75t_L g504 ( .A(n_151), .Y(n_504) );
AND2x4_ASAP7_75t_L g500 ( .A(n_152), .B(n_501), .Y(n_500) );
INVx2_ASAP7_75t_L g496 ( .A(n_153), .Y(n_496) );
AOI21xp5_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_157), .B(n_159), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_156), .B(n_549), .Y(n_548) );
AOI21xp5_ASAP7_75t_L g166 ( .A1(n_159), .A2(n_167), .B(n_168), .Y(n_166) );
AOI21xp5_ASAP7_75t_L g175 ( .A1(n_159), .A2(n_176), .B(n_177), .Y(n_175) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_159), .A2(n_190), .B(n_191), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_159), .A2(n_209), .B(n_210), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_159), .A2(n_220), .B(n_221), .Y(n_219) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_159), .A2(n_229), .B(n_230), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_159), .A2(n_235), .B(n_236), .Y(n_234) );
AOI21xp5_ASAP7_75t_L g467 ( .A1(n_159), .A2(n_468), .B(n_469), .Y(n_467) );
AOI21xp5_ASAP7_75t_L g475 ( .A1(n_159), .A2(n_476), .B(n_477), .Y(n_475) );
AOI21xp5_ASAP7_75t_L g485 ( .A1(n_159), .A2(n_486), .B(n_487), .Y(n_485) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_159), .A2(n_531), .B(n_532), .Y(n_530) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_159), .A2(n_539), .B(n_540), .Y(n_538) );
AOI21xp5_ASAP7_75t_L g546 ( .A1(n_159), .A2(n_547), .B(n_548), .Y(n_546) );
AOI21xp5_ASAP7_75t_L g556 ( .A1(n_159), .A2(n_557), .B(n_558), .Y(n_556) );
AND2x2_ASAP7_75t_L g184 ( .A(n_162), .B(n_185), .Y(n_184) );
AND2x2_ASAP7_75t_SL g341 ( .A(n_162), .B(n_249), .Y(n_341) );
AND2x2_ASAP7_75t_L g347 ( .A(n_162), .B(n_186), .Y(n_347) );
AND2x2_ASAP7_75t_L g436 ( .A(n_162), .B(n_437), .Y(n_436) );
OA21x2_ASAP7_75t_L g162 ( .A1(n_163), .A2(n_165), .B(n_169), .Y(n_162) );
OA21x2_ASAP7_75t_L g196 ( .A1(n_163), .A2(n_165), .B(n_169), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_163), .A2(n_226), .B(n_227), .Y(n_225) );
CKINVDCx5p33_ASAP7_75t_R g238 ( .A(n_163), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g464 ( .A1(n_163), .A2(n_465), .B(n_466), .Y(n_464) );
AO21x2_ASAP7_75t_L g492 ( .A1(n_163), .A2(n_493), .B(n_499), .Y(n_492) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx1_ASAP7_75t_SL g418 ( .A(n_170), .Y(n_418) );
AND2x2_ASAP7_75t_L g170 ( .A(n_171), .B(n_184), .Y(n_170) );
BUFx2_ASAP7_75t_L g247 ( .A(n_171), .Y(n_247) );
AND2x2_ASAP7_75t_L g281 ( .A(n_171), .B(n_185), .Y(n_281) );
AND2x2_ASAP7_75t_L g330 ( .A(n_171), .B(n_186), .Y(n_330) );
INVx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
AND2x2_ASAP7_75t_L g287 ( .A(n_172), .B(n_186), .Y(n_287) );
INVxp67_ASAP7_75t_L g299 ( .A(n_172), .Y(n_299) );
BUFx3_ASAP7_75t_L g344 ( .A(n_172), .Y(n_344) );
AO21x2_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_179), .B(n_183), .Y(n_172) );
AO21x2_ASAP7_75t_L g198 ( .A1(n_173), .A2(n_179), .B(n_183), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_174), .B(n_178), .Y(n_173) );
AO21x2_ASAP7_75t_L g186 ( .A1(n_179), .A2(n_187), .B(n_193), .Y(n_186) );
AO21x2_ASAP7_75t_L g200 ( .A1(n_179), .A2(n_187), .B(n_193), .Y(n_200) );
AO21x2_ASAP7_75t_L g553 ( .A1(n_179), .A2(n_554), .B(n_560), .Y(n_553) );
AO21x1_ASAP7_75t_SL g577 ( .A1(n_179), .A2(n_554), .B(n_560), .Y(n_577) );
INVx3_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx4_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
AO21x2_ASAP7_75t_L g482 ( .A1(n_181), .A2(n_483), .B(n_489), .Y(n_482) );
INVx3_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
BUFx4f_ASAP7_75t_L g215 ( .A(n_182), .Y(n_215) );
OAI31xp33_ASAP7_75t_L g240 ( .A1(n_184), .A2(n_241), .A3(n_246), .B(n_251), .Y(n_240) );
AND2x2_ASAP7_75t_L g248 ( .A(n_185), .B(n_249), .Y(n_248) );
INVx2_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
AND2x2_ASAP7_75t_L g267 ( .A(n_186), .B(n_268), .Y(n_267) );
NAND2xp5_ASAP7_75t_SL g187 ( .A(n_188), .B(n_192), .Y(n_187) );
AOI322xp5_ASAP7_75t_L g441 ( .A1(n_194), .A2(n_316), .A3(n_345), .B1(n_350), .B2(n_442), .C1(n_445), .C2(n_446), .Y(n_441) );
AND2x2_ASAP7_75t_L g194 ( .A(n_195), .B(n_197), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_195), .B(n_287), .Y(n_292) );
NAND2x1_ASAP7_75t_L g329 ( .A(n_195), .B(n_330), .Y(n_329) );
AND2x4_ASAP7_75t_L g373 ( .A(n_195), .B(n_277), .Y(n_373) );
INVx1_ASAP7_75t_SL g387 ( .A(n_195), .Y(n_387) );
INVx2_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
INVx2_ASAP7_75t_L g268 ( .A(n_196), .Y(n_268) );
HB1xp67_ASAP7_75t_L g411 ( .A(n_196), .Y(n_411) );
AND2x2_ASAP7_75t_L g340 ( .A(n_197), .B(n_341), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_197), .B(n_387), .Y(n_386) );
AND2x4_ASAP7_75t_SL g197 ( .A(n_198), .B(n_199), .Y(n_197) );
BUFx2_ASAP7_75t_L g245 ( .A(n_198), .Y(n_245) );
INVx1_ASAP7_75t_L g437 ( .A(n_198), .Y(n_437) );
OR2x2_ASAP7_75t_L g304 ( .A(n_199), .B(n_249), .Y(n_304) );
NAND2xp5_ASAP7_75t_SL g338 ( .A(n_199), .B(n_274), .Y(n_338) );
INVx2_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
AND2x4_ASAP7_75t_L g277 ( .A(n_200), .B(n_249), .Y(n_277) );
AND2x2_ASAP7_75t_L g201 ( .A(n_202), .B(n_222), .Y(n_201) );
INVxp67_ASAP7_75t_SL g202 ( .A(n_203), .Y(n_202) );
INVx1_ASAP7_75t_L g333 ( .A(n_203), .Y(n_333) );
OR2x2_ASAP7_75t_L g360 ( .A(n_203), .B(n_361), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_204), .B(n_214), .Y(n_203) );
NOR2x1_ASAP7_75t_SL g254 ( .A(n_204), .B(n_223), .Y(n_254) );
AND2x2_ASAP7_75t_L g261 ( .A(n_204), .B(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g433 ( .A(n_204), .B(n_295), .Y(n_433) );
AO21x2_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_206), .B(n_212), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g212 ( .A(n_205), .B(n_213), .Y(n_212) );
AO21x2_ASAP7_75t_L g310 ( .A1(n_205), .A2(n_206), .B(n_212), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_207), .B(n_211), .Y(n_206) );
OR2x2_ASAP7_75t_L g255 ( .A(n_214), .B(n_256), .Y(n_255) );
BUFx3_ASAP7_75t_L g264 ( .A(n_214), .Y(n_264) );
INVx2_ASAP7_75t_L g295 ( .A(n_214), .Y(n_295) );
INVx1_ASAP7_75t_L g336 ( .A(n_214), .Y(n_336) );
AND2x2_ASAP7_75t_L g367 ( .A(n_214), .B(n_223), .Y(n_367) );
AND2x2_ASAP7_75t_L g398 ( .A(n_214), .B(n_325), .Y(n_398) );
AOI21xp5_ASAP7_75t_L g543 ( .A1(n_215), .A2(n_544), .B(n_545), .Y(n_543) );
AND2x2_ASAP7_75t_L g294 ( .A(n_222), .B(n_295), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_222), .B(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_SL g397 ( .A(n_222), .B(n_398), .Y(n_397) );
AND2x2_ASAP7_75t_L g402 ( .A(n_222), .B(n_264), .Y(n_402) );
AND2x2_ASAP7_75t_L g222 ( .A(n_223), .B(n_231), .Y(n_222) );
INVx5_ASAP7_75t_L g262 ( .A(n_223), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_223), .B(n_256), .Y(n_334) );
BUFx2_ASAP7_75t_L g394 ( .A(n_223), .Y(n_394) );
OR2x6_ASAP7_75t_L g223 ( .A(n_224), .B(n_225), .Y(n_223) );
INVx4_ASAP7_75t_L g256 ( .A(n_231), .Y(n_256) );
AND2x2_ASAP7_75t_L g379 ( .A(n_231), .B(n_262), .Y(n_379) );
AO21x2_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_238), .B(n_239), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_233), .B(n_237), .Y(n_232) );
AOI21x1_ASAP7_75t_L g472 ( .A1(n_238), .A2(n_473), .B(n_479), .Y(n_472) );
INVx1_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
OAI221xp5_ASAP7_75t_L g368 ( .A1(n_242), .A2(n_369), .B1(n_372), .B2(n_374), .C(n_375), .Y(n_368) );
NAND2xp5_ASAP7_75t_SL g242 ( .A(n_243), .B(n_244), .Y(n_242) );
AND2x2_ASAP7_75t_L g390 ( .A(n_243), .B(n_281), .Y(n_390) );
INVx1_ASAP7_75t_SL g416 ( .A(n_243), .Y(n_416) );
AND2x2_ASAP7_75t_L g401 ( .A(n_244), .B(n_373), .Y(n_401) );
INVx2_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g346 ( .A(n_245), .B(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g246 ( .A(n_247), .B(n_248), .Y(n_246) );
AND2x2_ASAP7_75t_L g270 ( .A(n_247), .B(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g276 ( .A(n_247), .B(n_277), .Y(n_276) );
INVx1_ASAP7_75t_L g300 ( .A(n_248), .Y(n_300) );
AND2x2_ASAP7_75t_L g358 ( .A(n_248), .B(n_286), .Y(n_358) );
INVx2_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
BUFx2_ASAP7_75t_L g283 ( .A(n_250), .Y(n_283) );
INVx1_ASAP7_75t_SL g251 ( .A(n_252), .Y(n_251) );
OR2x2_ASAP7_75t_L g252 ( .A(n_253), .B(n_255), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
INVx2_ASAP7_75t_L g279 ( .A(n_255), .Y(n_279) );
OR2x2_ASAP7_75t_L g447 ( .A(n_255), .B(n_448), .Y(n_447) );
INVx2_ASAP7_75t_L g263 ( .A(n_256), .Y(n_263) );
AND2x4_ASAP7_75t_L g319 ( .A(n_256), .B(n_320), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_256), .B(n_324), .Y(n_323) );
NAND2x1p5_ASAP7_75t_L g361 ( .A(n_256), .B(n_262), .Y(n_361) );
AND2x2_ASAP7_75t_L g421 ( .A(n_256), .B(n_324), .Y(n_421) );
AOI22xp33_ASAP7_75t_L g257 ( .A1(n_258), .A2(n_265), .B1(n_278), .B2(n_280), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_258), .B(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
INVx2_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
AND3x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_263), .C(n_264), .Y(n_260) );
AND2x4_ASAP7_75t_L g278 ( .A(n_261), .B(n_279), .Y(n_278) );
INVx4_ASAP7_75t_L g318 ( .A(n_262), .Y(n_318) );
AND2x2_ASAP7_75t_SL g451 ( .A(n_262), .B(n_319), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_263), .B(n_427), .Y(n_426) );
INVx2_ASAP7_75t_L g363 ( .A(n_264), .Y(n_363) );
AOI322xp5_ASAP7_75t_L g428 ( .A1(n_264), .A2(n_393), .A3(n_429), .B1(n_431), .B2(n_434), .C1(n_438), .C2(n_439), .Y(n_428) );
NAND4xp25_ASAP7_75t_SL g265 ( .A(n_266), .B(n_269), .C(n_273), .D(n_275), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_SL g395 ( .A(n_267), .B(n_283), .Y(n_395) );
BUFx2_ASAP7_75t_L g286 ( .A(n_268), .Y(n_286) );
INVx1_ASAP7_75t_SL g269 ( .A(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g410 ( .A(n_271), .B(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
OR2x2_ASAP7_75t_L g424 ( .A(n_272), .B(n_299), .Y(n_424) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g290 ( .A(n_274), .B(n_291), .Y(n_290) );
OAI211xp5_ASAP7_75t_L g342 ( .A1(n_274), .A2(n_343), .B(n_345), .C(n_348), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_274), .B(n_281), .Y(n_400) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
AOI22xp5_ASAP7_75t_L g357 ( .A1(n_276), .A2(n_358), .B1(n_359), .B2(n_362), .Y(n_357) );
AOI22xp5_ASAP7_75t_L g312 ( .A1(n_277), .A2(n_313), .B1(n_317), .B2(n_321), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_277), .B(n_366), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_277), .B(n_414), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_277), .B(n_436), .Y(n_435) );
INVx2_ASAP7_75t_L g444 ( .A(n_277), .Y(n_444) );
INVx1_ASAP7_75t_L g383 ( .A(n_278), .Y(n_383) );
OAI21xp33_ASAP7_75t_SL g280 ( .A1(n_281), .A2(n_282), .B(n_284), .Y(n_280) );
INVx1_ASAP7_75t_L g291 ( .A(n_281), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_281), .B(n_286), .Y(n_440) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g376 ( .A(n_283), .B(n_287), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_285), .B(n_287), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_285), .B(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
OR2x2_ASAP7_75t_L g443 ( .A(n_286), .B(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g417 ( .A(n_287), .Y(n_417) );
A2O1A1Ixp33_ASAP7_75t_L g288 ( .A1(n_289), .A2(n_292), .B(n_293), .C(n_296), .Y(n_288) );
INVxp67_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
OAI22xp33_ASAP7_75t_SL g403 ( .A1(n_291), .A2(n_322), .B1(n_369), .B2(n_404), .Y(n_403) );
INVx1_ASAP7_75t_SL g293 ( .A(n_294), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_295), .B(n_318), .Y(n_326) );
OR2x2_ASAP7_75t_L g355 ( .A(n_295), .B(n_356), .Y(n_355) );
OAI21xp5_ASAP7_75t_SL g296 ( .A1(n_297), .A2(n_301), .B(n_305), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
OR2x2_ASAP7_75t_L g298 ( .A(n_299), .B(n_300), .Y(n_298) );
INVx1_ASAP7_75t_L g316 ( .A(n_299), .Y(n_316) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
OAI211xp5_ASAP7_75t_SL g354 ( .A1(n_302), .A2(n_355), .B(n_357), .C(n_365), .Y(n_354) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
NOR2xp67_ASAP7_75t_SL g388 ( .A(n_307), .B(n_334), .Y(n_388) );
INVx1_ASAP7_75t_L g391 ( .A(n_307), .Y(n_391) );
INVx2_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_309), .B(n_318), .Y(n_448) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g320 ( .A(n_310), .Y(n_320) );
INVx2_ASAP7_75t_L g325 ( .A(n_310), .Y(n_325) );
NAND4xp25_ASAP7_75t_L g311 ( .A(n_312), .B(n_327), .C(n_339), .D(n_342), .Y(n_311) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
OAI22xp33_ASAP7_75t_L g446 ( .A1(n_315), .A2(n_447), .B1(n_449), .B2(n_450), .Y(n_446) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
AND2x4_ASAP7_75t_L g414 ( .A(n_318), .B(n_344), .Y(n_414) );
AND2x2_ASAP7_75t_L g335 ( .A(n_319), .B(n_336), .Y(n_335) );
INVx2_ASAP7_75t_L g356 ( .A(n_319), .Y(n_356) );
AND2x2_ASAP7_75t_L g366 ( .A(n_319), .B(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
OR2x2_ASAP7_75t_L g322 ( .A(n_323), .B(n_326), .Y(n_322) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_325), .Y(n_380) );
INVx1_ASAP7_75t_L g370 ( .A(n_326), .Y(n_370) );
AOI32xp33_ASAP7_75t_L g327 ( .A1(n_328), .A2(n_331), .A3(n_334), .B1(n_335), .B2(n_337), .Y(n_327) );
OAI21xp33_ASAP7_75t_L g375 ( .A1(n_328), .A2(n_376), .B(n_377), .Y(n_375) );
INVx2_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
AOI221xp5_ASAP7_75t_L g407 ( .A1(n_331), .A2(n_408), .B1(n_410), .B2(n_412), .C(n_415), .Y(n_407) );
INVx1_ASAP7_75t_SL g331 ( .A(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g392 ( .A(n_333), .B(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g350 ( .A(n_334), .Y(n_350) );
AOI22xp5_ASAP7_75t_L g422 ( .A1(n_335), .A2(n_373), .B1(n_423), .B2(n_425), .Y(n_422) );
INVx1_ASAP7_75t_L g349 ( .A(n_336), .Y(n_349) );
AND2x2_ASAP7_75t_L g427 ( .A(n_336), .B(n_380), .Y(n_427) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
NAND2xp5_ASAP7_75t_SL g430 ( .A(n_343), .B(n_395), .Y(n_430) );
INVx1_ASAP7_75t_L g449 ( .A(n_343), .Y(n_449) );
INVx1_ASAP7_75t_SL g343 ( .A(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g348 ( .A(n_349), .B(n_350), .Y(n_348) );
NOR2xp67_ASAP7_75t_L g351 ( .A(n_352), .B(n_406), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_353), .B(n_396), .Y(n_352) );
NOR3xp33_ASAP7_75t_SL g353 ( .A(n_354), .B(n_368), .C(n_381), .Y(n_353) );
INVx1_ASAP7_75t_L g371 ( .A(n_356), .Y(n_371) );
INVx1_ASAP7_75t_SL g382 ( .A(n_358), .Y(n_382) );
INVx2_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx2_ASAP7_75t_L g364 ( .A(n_361), .Y(n_364) );
INVx2_ASAP7_75t_L g374 ( .A(n_362), .Y(n_374) );
AND2x2_ASAP7_75t_L g362 ( .A(n_363), .B(n_364), .Y(n_362) );
AND2x4_ASAP7_75t_L g420 ( .A(n_363), .B(n_421), .Y(n_420) );
AND2x4_ASAP7_75t_L g438 ( .A(n_367), .B(n_421), .Y(n_438) );
NAND2xp5_ASAP7_75t_SL g369 ( .A(n_370), .B(n_371), .Y(n_369) );
INVx1_ASAP7_75t_SL g372 ( .A(n_373), .Y(n_372) );
NOR2xp33_ASAP7_75t_L g377 ( .A(n_378), .B(n_380), .Y(n_377) );
AOI32xp33_ASAP7_75t_L g389 ( .A1(n_378), .A2(n_390), .A3(n_391), .B1(n_392), .B2(n_395), .Y(n_389) );
NOR2xp33_ASAP7_75t_SL g408 ( .A(n_378), .B(n_409), .Y(n_408) );
INVx2_ASAP7_75t_SL g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g409 ( .A(n_380), .Y(n_409) );
OAI211xp5_ASAP7_75t_SL g381 ( .A1(n_382), .A2(n_383), .B(n_384), .C(n_389), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_385), .B(n_388), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
AND2x2_ASAP7_75t_L g445 ( .A(n_393), .B(n_433), .Y(n_445) );
INVx2_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_394), .B(n_433), .Y(n_432) );
AOI221xp5_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_399), .B1(n_401), .B2(n_402), .C(n_403), .Y(n_396) );
INVx1_ASAP7_75t_SL g399 ( .A(n_400), .Y(n_399) );
CKINVDCx16_ASAP7_75t_R g404 ( .A(n_405), .Y(n_404) );
NAND4xp25_ASAP7_75t_L g406 ( .A(n_407), .B(n_422), .C(n_428), .D(n_441), .Y(n_406) );
INVxp33_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
O2A1O1Ixp33_ASAP7_75t_L g415 ( .A1(n_416), .A2(n_417), .B(n_418), .C(n_419), .Y(n_415) );
INVx2_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_SL g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_SL g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx3_ASAP7_75t_SL g450 ( .A(n_451), .Y(n_450) );
AOI22x1_ASAP7_75t_SL g768 ( .A1(n_453), .A2(n_454), .B1(n_769), .B2(n_775), .Y(n_768) );
INVx3_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
BUFx2_ASAP7_75t_L g755 ( .A(n_454), .Y(n_755) );
AND2x4_ASAP7_75t_L g454 ( .A(n_455), .B(n_660), .Y(n_454) );
NOR4xp75_ASAP7_75t_L g455 ( .A(n_456), .B(n_583), .C(n_608), .D(n_635), .Y(n_455) );
OAI21xp5_ASAP7_75t_L g456 ( .A1(n_457), .A2(n_521), .B(n_561), .Y(n_456) );
NOR4xp25_ASAP7_75t_L g457 ( .A(n_458), .B(n_505), .C(n_512), .D(n_516), .Y(n_457) );
INVx1_ASAP7_75t_SL g458 ( .A(n_459), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_460), .B(n_480), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_462), .B(n_471), .Y(n_461) );
NAND2x1p5_ASAP7_75t_L g623 ( .A(n_462), .B(n_624), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_462), .B(n_509), .Y(n_654) );
AND2x2_ASAP7_75t_L g679 ( .A(n_462), .B(n_680), .Y(n_679) );
AND2x2_ASAP7_75t_L g704 ( .A(n_462), .B(n_490), .Y(n_704) );
AND2x2_ASAP7_75t_L g745 ( .A(n_462), .B(n_514), .Y(n_745) );
INVx4_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
AND2x4_ASAP7_75t_SL g518 ( .A(n_463), .B(n_511), .Y(n_518) );
AND2x2_ASAP7_75t_L g520 ( .A(n_463), .B(n_482), .Y(n_520) );
NOR2x1_ASAP7_75t_L g569 ( .A(n_463), .B(n_570), .Y(n_569) );
INVx1_ASAP7_75t_L g580 ( .A(n_463), .Y(n_580) );
AND2x2_ASAP7_75t_L g586 ( .A(n_463), .B(n_514), .Y(n_586) );
BUFx2_ASAP7_75t_L g599 ( .A(n_463), .Y(n_599) );
AND2x4_ASAP7_75t_L g630 ( .A(n_463), .B(n_631), .Y(n_630) );
AND2x2_ASAP7_75t_L g677 ( .A(n_463), .B(n_678), .Y(n_677) );
OR2x6_ASAP7_75t_L g463 ( .A(n_464), .B(n_470), .Y(n_463) );
INVx1_ASAP7_75t_L g671 ( .A(n_471), .Y(n_671) );
HB1xp67_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx3_ASAP7_75t_L g511 ( .A(n_472), .Y(n_511) );
AND2x2_ASAP7_75t_L g514 ( .A(n_472), .B(n_482), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_474), .B(n_478), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_480), .B(n_689), .Y(n_742) );
INVx2_ASAP7_75t_SL g480 ( .A(n_481), .Y(n_480) );
OR2x2_ASAP7_75t_L g579 ( .A(n_481), .B(n_580), .Y(n_579) );
OR2x2_ASAP7_75t_L g481 ( .A(n_482), .B(n_490), .Y(n_481) );
INVx2_ASAP7_75t_L g510 ( .A(n_482), .Y(n_510) );
INVx2_ASAP7_75t_L g570 ( .A(n_482), .Y(n_570) );
AND2x2_ASAP7_75t_L g680 ( .A(n_482), .B(n_511), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_484), .B(n_488), .Y(n_483) );
INVx2_ASAP7_75t_L g568 ( .A(n_490), .Y(n_568) );
BUFx3_ASAP7_75t_L g585 ( .A(n_490), .Y(n_585) );
AND2x2_ASAP7_75t_L g612 ( .A(n_490), .B(n_613), .Y(n_612) );
AND2x4_ASAP7_75t_L g490 ( .A(n_491), .B(n_492), .Y(n_490) );
AND2x4_ASAP7_75t_L g507 ( .A(n_491), .B(n_492), .Y(n_507) );
AND2x4_ASAP7_75t_L g494 ( .A(n_495), .B(n_498), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_496), .B(n_497), .Y(n_495) );
NOR2x1p5_ASAP7_75t_L g501 ( .A(n_502), .B(n_503), .Y(n_501) );
INVx3_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
NOR2x1_ASAP7_75t_L g505 ( .A(n_506), .B(n_508), .Y(n_505) );
INVx2_ASAP7_75t_L g515 ( .A(n_506), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_506), .B(n_671), .Y(n_670) );
OR2x2_ASAP7_75t_L g683 ( .A(n_506), .B(n_623), .Y(n_683) );
AND2x2_ASAP7_75t_L g707 ( .A(n_506), .B(n_518), .Y(n_707) );
INVx3_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
AND2x2_ASAP7_75t_L g603 ( .A(n_507), .B(n_510), .Y(n_603) );
AND2x2_ASAP7_75t_L g685 ( .A(n_507), .B(n_678), .Y(n_685) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx1_ASAP7_75t_SL g728 ( .A(n_509), .Y(n_728) );
AND2x2_ASAP7_75t_L g509 ( .A(n_510), .B(n_511), .Y(n_509) );
INVx1_ASAP7_75t_L g613 ( .A(n_510), .Y(n_613) );
HB1xp67_ASAP7_75t_L g617 ( .A(n_511), .Y(n_617) );
INVx2_ASAP7_75t_L g625 ( .A(n_511), .Y(n_625) );
INVx1_ASAP7_75t_L g631 ( .A(n_511), .Y(n_631) );
AOI222xp33_ASAP7_75t_SL g561 ( .A1(n_512), .A2(n_562), .B1(n_566), .B2(n_571), .C1(n_578), .C2(n_581), .Y(n_561) );
INVx1_ASAP7_75t_SL g512 ( .A(n_513), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_514), .B(n_515), .Y(n_513) );
INVx1_ASAP7_75t_L g638 ( .A(n_514), .Y(n_638) );
BUFx2_ASAP7_75t_L g667 ( .A(n_514), .Y(n_667) );
OAI211xp5_ASAP7_75t_L g661 ( .A1(n_515), .A2(n_662), .B(n_666), .C(n_674), .Y(n_661) );
OR2x2_ASAP7_75t_L g732 ( .A(n_515), .B(n_733), .Y(n_732) );
AND2x2_ASAP7_75t_L g740 ( .A(n_515), .B(n_645), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_517), .B(n_519), .Y(n_516) );
INVx2_ASAP7_75t_SL g517 ( .A(n_518), .Y(n_517) );
AND2x2_ASAP7_75t_SL g697 ( .A(n_518), .B(n_698), .Y(n_697) );
AND2x2_ASAP7_75t_L g715 ( .A(n_518), .B(n_603), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_518), .B(n_695), .Y(n_722) );
OR2x2_ASAP7_75t_L g723 ( .A(n_519), .B(n_585), .Y(n_723) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
AND2x2_ASAP7_75t_L g645 ( .A(n_520), .B(n_617), .Y(n_645) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_523), .B(n_541), .Y(n_522) );
INVx1_ASAP7_75t_L g739 ( .A(n_523), .Y(n_739) );
NOR2xp67_ASAP7_75t_L g523 ( .A(n_524), .B(n_533), .Y(n_523) );
AND2x2_ASAP7_75t_L g582 ( .A(n_524), .B(n_542), .Y(n_582) );
INVx1_ASAP7_75t_L g659 ( .A(n_524), .Y(n_659) );
OR2x2_ASAP7_75t_L g718 ( .A(n_524), .B(n_542), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_524), .B(n_590), .Y(n_724) );
INVx4_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx2_ASAP7_75t_L g565 ( .A(n_525), .Y(n_565) );
OR2x2_ASAP7_75t_L g597 ( .A(n_525), .B(n_552), .Y(n_597) );
AND2x2_ASAP7_75t_L g606 ( .A(n_525), .B(n_534), .Y(n_606) );
NAND2x1_ASAP7_75t_L g634 ( .A(n_525), .B(n_542), .Y(n_634) );
AND2x2_ASAP7_75t_L g681 ( .A(n_525), .B(n_576), .Y(n_681) );
OR2x6_ASAP7_75t_L g525 ( .A(n_526), .B(n_527), .Y(n_525) );
HB1xp67_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx1_ASAP7_75t_L g564 ( .A(n_534), .Y(n_564) );
INVx1_ASAP7_75t_L g574 ( .A(n_534), .Y(n_574) );
AND2x2_ASAP7_75t_L g590 ( .A(n_534), .B(n_577), .Y(n_590) );
INVx2_ASAP7_75t_L g595 ( .A(n_534), .Y(n_595) );
OR2x2_ASAP7_75t_L g691 ( .A(n_534), .B(n_542), .Y(n_691) );
AND2x2_ASAP7_75t_L g541 ( .A(n_542), .B(n_551), .Y(n_541) );
NOR2x1_ASAP7_75t_SL g576 ( .A(n_542), .B(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g594 ( .A(n_542), .B(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g607 ( .A(n_542), .B(n_552), .Y(n_607) );
BUFx2_ASAP7_75t_L g626 ( .A(n_542), .Y(n_626) );
INVx2_ASAP7_75t_SL g653 ( .A(n_542), .Y(n_653) );
OR2x6_ASAP7_75t_L g542 ( .A(n_543), .B(n_550), .Y(n_542) );
INVx2_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g563 ( .A(n_552), .B(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g709 ( .A(n_552), .B(n_651), .Y(n_709) );
INVx3_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_555), .B(n_559), .Y(n_554) );
AOI211xp5_ASAP7_75t_L g725 ( .A1(n_562), .A2(n_586), .B(n_726), .C(n_730), .Y(n_725) );
AND2x2_ASAP7_75t_L g562 ( .A(n_563), .B(n_565), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_563), .B(n_641), .Y(n_676) );
BUFx2_ASAP7_75t_L g640 ( .A(n_564), .Y(n_640) );
OR2x2_ASAP7_75t_L g588 ( .A(n_565), .B(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_L g673 ( .A(n_565), .B(n_607), .Y(n_673) );
AND2x2_ASAP7_75t_L g694 ( .A(n_565), .B(n_650), .Y(n_694) );
INVx2_ASAP7_75t_L g701 ( .A(n_565), .Y(n_701) );
OAI21xp5_ASAP7_75t_SL g706 ( .A1(n_566), .A2(n_707), .B(n_708), .Y(n_706) );
AND2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_569), .Y(n_566) );
AND2x2_ASAP7_75t_L g648 ( .A(n_567), .B(n_630), .Y(n_648) );
OR2x2_ASAP7_75t_L g727 ( .A(n_567), .B(n_728), .Y(n_727) );
INVx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_568), .B(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_570), .Y(n_601) );
AND2x2_ASAP7_75t_L g678 ( .A(n_570), .B(n_625), .Y(n_678) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
OR2x2_ASAP7_75t_L g572 ( .A(n_573), .B(n_575), .Y(n_572) );
AND2x2_ASAP7_75t_L g663 ( .A(n_573), .B(n_664), .Y(n_663) );
AND2x4_ASAP7_75t_SL g672 ( .A(n_573), .B(n_673), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_573), .B(n_582), .Y(n_705) );
INVx3_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g581 ( .A(n_574), .B(n_582), .Y(n_581) );
OR2x2_ASAP7_75t_L g700 ( .A(n_575), .B(n_701), .Y(n_700) );
INVx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g650 ( .A(n_576), .B(n_651), .Y(n_650) );
AND2x2_ASAP7_75t_L g620 ( .A(n_577), .B(n_595), .Y(n_620) );
OAI31xp33_ASAP7_75t_L g627 ( .A1(n_578), .A2(n_628), .A3(n_630), .B(n_632), .Y(n_627) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
NAND2xp5_ASAP7_75t_SL g629 ( .A(n_580), .B(n_603), .Y(n_629) );
AO21x1_ASAP7_75t_L g583 ( .A1(n_584), .A2(n_587), .B(n_591), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_585), .B(n_586), .Y(n_584) );
OR2x2_ASAP7_75t_L g639 ( .A(n_585), .B(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g744 ( .A(n_585), .Y(n_744) );
INVx2_ASAP7_75t_SL g729 ( .A(n_586), .Y(n_729) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
OR2x2_ASAP7_75t_L g633 ( .A(n_589), .B(n_634), .Y(n_633) );
OR2x2_ASAP7_75t_L g717 ( .A(n_589), .B(n_718), .Y(n_717) );
INVx2_ASAP7_75t_SL g589 ( .A(n_590), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_590), .B(n_653), .Y(n_734) );
OAI22xp5_ASAP7_75t_L g591 ( .A1(n_592), .A2(n_598), .B1(n_602), .B2(n_604), .Y(n_591) );
AOI21xp33_ASAP7_75t_L g710 ( .A1(n_592), .A2(n_711), .B(n_712), .Y(n_710) );
INVx3_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
AND2x4_ASAP7_75t_L g593 ( .A(n_594), .B(n_596), .Y(n_593) );
INVx1_ASAP7_75t_L g651 ( .A(n_595), .Y(n_651) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
OR2x2_ASAP7_75t_L g665 ( .A(n_597), .B(n_626), .Y(n_665) );
OR2x2_ASAP7_75t_L g690 ( .A(n_597), .B(n_691), .Y(n_690) );
OR2x2_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_599), .B(n_603), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_599), .B(n_612), .Y(n_611) );
INVx2_ASAP7_75t_L g689 ( .A(n_599), .Y(n_689) );
INVx2_ASAP7_75t_L g618 ( .A(n_600), .Y(n_618) );
INVx1_ASAP7_75t_L g698 ( .A(n_601), .Y(n_698) );
AND2x2_ASAP7_75t_L g621 ( .A(n_603), .B(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g695 ( .A(n_603), .Y(n_695) );
INVx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_606), .B(n_607), .Y(n_605) );
NAND2xp5_ASAP7_75t_SL g608 ( .A(n_609), .B(n_627), .Y(n_608) );
OAI321xp33_ASAP7_75t_L g609 ( .A1(n_610), .A2(n_614), .A3(n_619), .B1(n_620), .B2(n_621), .C(n_626), .Y(n_609) );
AOI322xp5_ASAP7_75t_L g735 ( .A1(n_610), .A2(n_641), .A3(n_736), .B1(n_738), .B2(n_740), .C1(n_741), .C2(n_746), .Y(n_735) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
BUFx2_ASAP7_75t_L g688 ( .A(n_613), .Y(n_688) );
AND2x2_ASAP7_75t_L g614 ( .A(n_615), .B(n_618), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_615), .B(n_695), .Y(n_712) );
INVx2_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx2_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g720 ( .A(n_618), .Y(n_720) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
NAND2xp33_ASAP7_75t_SL g652 ( .A(n_620), .B(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
OAI21xp33_ASAP7_75t_SL g719 ( .A1(n_623), .A2(n_629), .B(n_720), .Y(n_719) );
INVx1_ASAP7_75t_SL g624 ( .A(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx2_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx3_ASAP7_75t_L g641 ( .A(n_634), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_636), .B(n_655), .Y(n_635) );
AOI221xp5_ASAP7_75t_L g636 ( .A1(n_637), .A2(n_641), .B1(n_642), .B2(n_643), .C(n_646), .Y(n_636) );
NOR2xp33_ASAP7_75t_L g637 ( .A(n_638), .B(n_639), .Y(n_637) );
HB1xp67_ASAP7_75t_L g657 ( .A(n_638), .Y(n_657) );
AND2x2_ASAP7_75t_L g642 ( .A(n_640), .B(n_641), .Y(n_642) );
INVx2_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
OAI22xp33_ASAP7_75t_SL g646 ( .A1(n_647), .A2(n_649), .B1(n_652), .B2(n_654), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
AND2x2_ASAP7_75t_L g658 ( .A(n_650), .B(n_659), .Y(n_658) );
OAI21xp33_ASAP7_75t_L g741 ( .A1(n_653), .A2(n_742), .B(n_743), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_656), .B(n_658), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
NOR3xp33_ASAP7_75t_SL g660 ( .A(n_661), .B(n_692), .C(n_713), .Y(n_660) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_SL g664 ( .A(n_665), .Y(n_664) );
OAI22xp5_ASAP7_75t_L g726 ( .A1(n_665), .A2(n_700), .B1(n_727), .B2(n_729), .Y(n_726) );
OAI21xp33_ASAP7_75t_SL g666 ( .A1(n_667), .A2(n_668), .B(n_672), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_667), .B(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
HB1xp67_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
AOI221xp5_ASAP7_75t_L g714 ( .A1(n_673), .A2(n_715), .B1(n_716), .B2(n_719), .C(n_721), .Y(n_714) );
AOI221xp5_ASAP7_75t_L g674 ( .A1(n_675), .A2(n_677), .B1(n_679), .B2(n_681), .C(n_682), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g711 ( .A(n_677), .Y(n_711) );
INVx1_ASAP7_75t_L g733 ( .A(n_678), .Y(n_733) );
INVx1_ASAP7_75t_SL g731 ( .A(n_679), .Y(n_731) );
AOI31xp33_ASAP7_75t_L g682 ( .A1(n_683), .A2(n_684), .A3(n_686), .B(n_690), .Y(n_682) );
OAI221xp5_ASAP7_75t_L g692 ( .A1(n_683), .A2(n_693), .B1(n_695), .B2(n_696), .C(n_793), .Y(n_692) );
INVx2_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_687), .B(n_689), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
AOI211xp5_ASAP7_75t_L g696 ( .A1(n_697), .A2(n_699), .B(n_702), .C(n_710), .Y(n_696) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
AND2x2_ASAP7_75t_L g708 ( .A(n_701), .B(n_709), .Y(n_708) );
OAI21xp5_ASAP7_75t_SL g702 ( .A1(n_703), .A2(n_705), .B(n_706), .Y(n_702) );
INVx1_ASAP7_75t_L g737 ( .A(n_709), .Y(n_737) );
BUFx2_ASAP7_75t_SL g746 ( .A(n_709), .Y(n_746) );
NAND3xp33_ASAP7_75t_SL g713 ( .A(n_714), .B(n_725), .C(n_735), .Y(n_713) );
INVx2_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
AOI21xp33_ASAP7_75t_L g721 ( .A1(n_722), .A2(n_723), .B(n_724), .Y(n_721) );
AOI21xp33_ASAP7_75t_L g730 ( .A1(n_731), .A2(n_732), .B(n_734), .Y(n_730) );
HB1xp67_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVxp67_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_744), .B(n_745), .Y(n_743) );
CKINVDCx11_ASAP7_75t_R g747 ( .A(n_748), .Y(n_747) );
CKINVDCx5p33_ASAP7_75t_R g758 ( .A(n_748), .Y(n_758) );
AOI21xp5_ASAP7_75t_L g753 ( .A1(n_749), .A2(n_754), .B(n_759), .Y(n_753) );
CKINVDCx6p67_ASAP7_75t_R g756 ( .A(n_757), .Y(n_756) );
INVx3_ASAP7_75t_SL g757 ( .A(n_758), .Y(n_757) );
NOR2xp33_ASAP7_75t_L g759 ( .A(n_760), .B(n_761), .Y(n_759) );
BUFx2_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_764), .B(n_766), .Y(n_763) );
INVx1_ASAP7_75t_SL g764 ( .A(n_765), .Y(n_764) );
INVx1_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
INVx1_ASAP7_75t_L g775 ( .A(n_769), .Y(n_775) );
INVx1_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
INVx1_ASAP7_75t_SL g776 ( .A(n_777), .Y(n_776) );
INVx1_ASAP7_75t_SL g777 ( .A(n_778), .Y(n_777) );
INVx1_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
INVx1_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
INVx1_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
INVx1_ASAP7_75t_SL g791 ( .A(n_782), .Y(n_791) );
CKINVDCx5p33_ASAP7_75t_R g782 ( .A(n_783), .Y(n_782) );
AND2x2_ASAP7_75t_SL g783 ( .A(n_784), .B(n_785), .Y(n_783) );
INVx2_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
NOR2xp33_ASAP7_75t_L g789 ( .A(n_790), .B(n_791), .Y(n_789) );
endmodule