module fake_jpeg_1958_n_111 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_111);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_111;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx5_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_6),
.B(n_18),
.Y(n_30)
);

CKINVDCx14_ASAP7_75t_R g31 ( 
.A(n_23),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_17),
.Y(n_32)
);

CKINVDCx14_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_28),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_33),
.Y(n_52)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_39),
.Y(n_42)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

CKINVDCx9p33_ASAP7_75t_R g54 ( 
.A(n_44),
.Y(n_54)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_45),
.B(n_32),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_41),
.A2(n_37),
.B1(n_33),
.B2(n_31),
.Y(n_46)
);

AO22x1_ASAP7_75t_SL g55 ( 
.A1(n_46),
.A2(n_43),
.B1(n_37),
.B2(n_42),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_47),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_40),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_50),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_45),
.B(n_31),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_52),
.B(n_30),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_55),
.A2(n_63),
.B1(n_46),
.B2(n_53),
.Y(n_65)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

NAND3xp33_ASAP7_75t_L g74 ( 
.A(n_57),
.B(n_64),
.C(n_58),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_47),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_60),
.B(n_61),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_15),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_49),
.A2(n_42),
.B1(n_44),
.B2(n_35),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_47),
.B(n_0),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_62),
.B(n_53),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_67),
.B(n_72),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_59),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_68),
.B(n_73),
.Y(n_76)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_51),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_74),
.B(n_0),
.Y(n_84)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_75),
.Y(n_79)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

CKINVDCx10_ASAP7_75t_R g81 ( 
.A(n_75),
.Y(n_81)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

FAx1_ASAP7_75t_SL g83 ( 
.A(n_74),
.B(n_58),
.CI(n_51),
.CON(n_83),
.SN(n_83)
);

OAI321xp33_ASAP7_75t_L g87 ( 
.A1(n_83),
.A2(n_26),
.A3(n_25),
.B1(n_24),
.B2(n_22),
.C(n_20),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_84),
.B(n_19),
.Y(n_88)
);

OAI32xp33_ASAP7_75t_L g85 ( 
.A1(n_66),
.A2(n_29),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_85),
.B(n_86),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_71),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_87),
.A2(n_93),
.B1(n_95),
.B2(n_96),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_78),
.B(n_1),
.Y(n_90)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_90),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_82),
.B(n_71),
.C(n_16),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_91),
.B(n_81),
.C(n_77),
.Y(n_98)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_77),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_76),
.A2(n_5),
.B(n_8),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_98),
.B(n_99),
.C(n_91),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_89),
.B(n_83),
.C(n_85),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_102),
.B(n_103),
.Y(n_104)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_100),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_104),
.B(n_101),
.Y(n_105)
);

AOI322xp5_ASAP7_75t_L g106 ( 
.A1(n_105),
.A2(n_96),
.A3(n_94),
.B1(n_92),
.B2(n_97),
.C1(n_83),
.C2(n_12),
.Y(n_106)
);

NOR2x1p5_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_94),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_12),
.C(n_9),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_8),
.C(n_9),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_10),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_110),
.B(n_11),
.Y(n_111)
);


endmodule