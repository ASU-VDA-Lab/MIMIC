module real_jpeg_1848_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_202;
wire n_128;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx2_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_2),
.A2(n_39),
.B1(n_40),
.B2(n_42),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_2),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_2),
.A2(n_39),
.B1(n_60),
.B2(n_61),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_2),
.A2(n_23),
.B1(n_24),
.B2(n_39),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_2),
.A2(n_39),
.B1(n_72),
.B2(n_75),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_2),
.B(n_61),
.C(n_69),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_2),
.B(n_67),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_2),
.B(n_40),
.C(n_55),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_2),
.B(n_24),
.C(n_46),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_2),
.B(n_53),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_2),
.B(n_31),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_2),
.B(n_50),
.Y(n_239)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_3),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_4),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_5),
.A2(n_72),
.B1(n_74),
.B2(n_75),
.Y(n_71)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_5),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_5),
.A2(n_60),
.B1(n_61),
.B2(n_74),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_5),
.A2(n_40),
.B1(n_42),
.B2(n_74),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_5),
.A2(n_23),
.B1(n_24),
.B2(n_74),
.Y(n_217)
);

BUFx16f_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_7),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g22 ( 
.A1(n_8),
.A2(n_23),
.B1(n_24),
.B2(n_28),
.Y(n_22)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_8),
.A2(n_28),
.B1(n_40),
.B2(n_42),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_8),
.A2(n_28),
.B1(n_60),
.B2(n_61),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_8),
.A2(n_28),
.B1(n_72),
.B2(n_75),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_9),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_10),
.A2(n_23),
.B1(n_24),
.B2(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_10),
.A2(n_35),
.B1(n_40),
.B2(n_42),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_10),
.A2(n_35),
.B1(n_72),
.B2(n_75),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_10),
.A2(n_35),
.B1(n_60),
.B2(n_61),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_SL g12 ( 
.A(n_13),
.B(n_264),
.C(n_320),
.Y(n_12)
);

OA21x2_ASAP7_75t_SL g13 ( 
.A1(n_14),
.A2(n_319),
.B(n_324),
.Y(n_13)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_311),
.B(n_318),
.Y(n_14)
);

OAI21xp5_ASAP7_75t_SL g15 ( 
.A1(n_16),
.A2(n_273),
.B(n_308),
.Y(n_15)
);

A2O1A1O1Ixp25_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_135),
.B(n_253),
.C(n_254),
.D(n_272),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_113),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_18),
.B(n_113),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_80),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_19),
.B(n_81),
.C(n_107),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_52),
.C(n_64),
.Y(n_19)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_20),
.B(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_36),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_21),
.B(n_36),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_29),
.B(n_32),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_22),
.A2(n_30),
.B(n_88),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_23),
.A2(n_24),
.B1(n_45),
.B2(n_46),
.Y(n_48)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_24),
.B(n_235),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_29),
.B(n_34),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_29),
.A2(n_30),
.B(n_87),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_29),
.B(n_87),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_29),
.B(n_217),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_30),
.B(n_34),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_30),
.B(n_217),
.Y(n_231)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_31),
.B(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_32),
.B(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_33),
.B(n_216),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_37),
.B(n_49),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_37),
.B(n_202),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_43),
.Y(n_37)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_38),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_38),
.B(n_50),
.Y(n_188)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_40),
.A2(n_42),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_40),
.A2(n_42),
.B1(n_55),
.B2(n_56),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_40),
.B(n_211),
.Y(n_210)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_43),
.B(n_51),
.Y(n_92)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_43),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_43),
.B(n_190),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_48),
.Y(n_43)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_48),
.Y(n_50)
);

OAI21x1_ASAP7_75t_SL g110 ( 
.A1(n_49),
.A2(n_91),
.B(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_49),
.B(n_189),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_50),
.B(n_51),
.Y(n_49)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_50),
.B(n_190),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_52),
.A2(n_64),
.B1(n_65),
.B2(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_52),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_52),
.A2(n_117),
.B1(n_315),
.B2(n_316),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_52),
.B(n_315),
.C(n_317),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_57),
.B(n_63),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_53),
.B(n_63),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_53),
.B(n_128),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_53),
.A2(n_154),
.B(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_54),
.B(n_59),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_54),
.B(n_103),
.Y(n_102)
);

INVx3_ASAP7_75t_SL g56 ( 
.A(n_55),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_55),
.A2(n_56),
.B1(n_60),
.B2(n_61),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_57),
.B(n_63),
.Y(n_105)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_58),
.B(n_127),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_58),
.B(n_103),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_58),
.A2(n_287),
.B(n_288),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_60),
.A2(n_61),
.B1(n_68),
.B2(n_69),
.Y(n_67)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_61),
.B(n_185),
.Y(n_184)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_76),
.Y(n_65)
);

CKINVDCx14_ASAP7_75t_R g147 ( 
.A(n_66),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_71),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_67),
.B(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_67),
.B(n_79),
.Y(n_121)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_67),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_68),
.A2(n_69),
.B1(n_72),
.B2(n_75),
.Y(n_78)
);

INVx6_ASAP7_75t_SL g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_71),
.B(n_77),
.Y(n_99)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_72),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_72),
.B(n_132),
.Y(n_131)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_76),
.A2(n_265),
.B(n_301),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_76),
.B(n_96),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_77),
.B(n_79),
.Y(n_76)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_77),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_81),
.A2(n_82),
.B1(n_106),
.B2(n_107),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_93),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_83),
.B(n_94),
.C(n_101),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_89),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_84),
.B(n_89),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_88),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_85),
.B(n_215),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_88),
.B(n_230),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_91),
.B(n_92),
.Y(n_89)
);

AOI21x1_ASAP7_75t_SL g151 ( 
.A1(n_90),
.A2(n_111),
.B(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_92),
.B(n_202),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_92),
.B(n_188),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_94),
.A2(n_95),
.B1(n_100),
.B2(n_101),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_99),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_98),
.B(n_149),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_98),
.A2(n_149),
.B(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_99),
.B(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_104),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_102),
.B(n_126),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_102),
.Y(n_288)
);

INVxp33_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_105),
.B(n_156),
.Y(n_203)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_109),
.B1(n_110),
.B2(n_112),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_108),
.A2(n_109),
.B1(n_183),
.B2(n_184),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_108),
.A2(n_109),
.B1(n_263),
.B2(n_264),
.Y(n_262)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_109),
.B(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_109),
.B(n_110),
.Y(n_261)
);

AOI21xp33_ASAP7_75t_L g277 ( 
.A1(n_109),
.A2(n_261),
.B(n_263),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_110),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_118),
.C(n_134),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_114),
.A2(n_115),
.B1(n_134),
.B2(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_139),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_122),
.C(n_129),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_119),
.A2(n_120),
.B1(n_122),
.B2(n_123),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_121),
.B(n_283),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_121),
.A2(n_149),
.B(n_301),
.Y(n_315)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_125),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g306 ( 
.A(n_124),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_129),
.B(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_133),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_130),
.A2(n_131),
.B1(n_133),
.B2(n_167),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_133),
.Y(n_167)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_134),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_157),
.B(n_250),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_137),
.A2(n_251),
.B(n_252),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_138),
.B(n_141),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_138),
.B(n_141),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_144),
.C(n_145),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_142),
.B(n_160),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_144),
.B(n_145),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_150),
.C(n_153),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_146),
.B(n_164),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_148),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_148),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_150),
.A2(n_151),
.B1(n_153),
.B2(n_165),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_150),
.A2(n_151),
.B1(n_286),
.B2(n_289),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_150),
.A2(n_151),
.B1(n_304),
.B2(n_305),
.Y(n_303)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_151),
.B(n_281),
.C(n_286),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_151),
.B(n_305),
.C(n_307),
.Y(n_317)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_153),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_154),
.B(n_155),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_154),
.B(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_175),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_159),
.B(n_161),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_159),
.B(n_161),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_166),
.C(n_168),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_162),
.A2(n_163),
.B1(n_192),
.B2(n_193),
.Y(n_191)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_166),
.B(n_168),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.C(n_171),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_169),
.B(n_180),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_170),
.A2(n_171),
.B1(n_172),
.B2(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_170),
.Y(n_181)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_174),
.B(n_231),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_194),
.B(n_249),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_191),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_177),
.B(n_191),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_182),
.C(n_186),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_178),
.A2(n_179),
.B1(n_197),
.B2(n_199),
.Y(n_196)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_182),
.A2(n_186),
.B1(n_187),
.B2(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_182),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_189),
.Y(n_187)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

AOI21x1_ASAP7_75t_SL g194 ( 
.A1(n_195),
.A2(n_205),
.B(n_248),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_196),
.B(n_200),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_196),
.B(n_200),
.Y(n_248)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_197),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_203),
.C(n_204),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_201),
.B(n_203),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_204),
.B(n_246),
.Y(n_245)
);

OAI21x1_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_243),
.B(n_247),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_225),
.B(n_242),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_213),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_208),
.B(n_213),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_212),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_209),
.A2(n_210),
.B1(n_212),
.B2(n_228),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_212),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_218),
.B1(n_219),
.B2(n_224),
.Y(n_213)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_214),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_220),
.A2(n_221),
.B1(n_222),
.B2(n_223),
.Y(n_219)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_220),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_221),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_221),
.B(n_222),
.C(n_224),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_226),
.A2(n_232),
.B(n_241),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_227),
.B(n_229),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_227),
.B(n_229),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_237),
.B(n_240),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_236),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_238),
.B(n_239),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_244),
.B(n_245),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_255),
.B(n_256),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_257),
.B(n_259),
.C(n_267),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_259),
.A2(n_260),
.B1(n_266),
.B2(n_267),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_268),
.A2(n_269),
.B(n_271),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_268),
.B(n_269),
.Y(n_271)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_270),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_271),
.A2(n_279),
.B1(n_280),
.B2(n_290),
.Y(n_278)
);

CKINVDCx14_ASAP7_75t_R g290 ( 
.A(n_271),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_271),
.B(n_277),
.C(n_279),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_291),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_275),
.B(n_276),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_282),
.B1(n_284),
.B2(n_285),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_281),
.A2(n_282),
.B1(n_298),
.B2(n_299),
.Y(n_297)
);

CKINVDCx14_ASAP7_75t_R g281 ( 
.A(n_282),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_282),
.B(n_294),
.C(n_298),
.Y(n_312)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_286),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_291),
.A2(n_309),
.B(n_310),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_292),
.B(n_293),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_294),
.A2(n_295),
.B1(n_296),
.B2(n_297),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_300),
.A2(n_302),
.B1(n_303),
.B2(n_307),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_300),
.Y(n_307)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_312),
.B(n_313),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_312),
.B(n_313),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_317),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_315),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_322),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_321),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_321),
.B(n_323),
.Y(n_325)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_323),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);


endmodule