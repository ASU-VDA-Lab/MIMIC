module real_aes_17276_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_800;
wire n_778;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_852;
wire n_766;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_549;
wire n_376;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_528;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_872;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_656;
wire n_532;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_102;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_867;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_546;
wire n_151;
wire n_639;
wire n_587;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
AND2x4_ASAP7_75t_L g111 ( .A(n_0), .B(n_112), .Y(n_111) );
AOI22xp5_ASAP7_75t_L g264 ( .A1(n_1), .A2(n_4), .B1(n_265), .B2(n_266), .Y(n_264) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_2), .A2(n_44), .B1(n_136), .B2(n_165), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g251 ( .A1(n_3), .A2(n_25), .B1(n_165), .B2(n_246), .Y(n_251) );
AOI22xp5_ASAP7_75t_L g607 ( .A1(n_5), .A2(n_16), .B1(n_525), .B2(n_608), .Y(n_607) );
AOI22xp5_ASAP7_75t_L g121 ( .A1(n_6), .A2(n_31), .B1(n_122), .B2(n_123), .Y(n_121) );
INVx1_ASAP7_75t_L g123 ( .A(n_6), .Y(n_123) );
AOI22xp33_ASAP7_75t_L g201 ( .A1(n_7), .A2(n_62), .B1(n_173), .B2(n_202), .Y(n_201) );
AOI22xp5_ASAP7_75t_L g135 ( .A1(n_8), .A2(n_17), .B1(n_136), .B2(n_138), .Y(n_135) );
INVx1_ASAP7_75t_L g112 ( .A(n_9), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g245 ( .A(n_10), .Y(n_245) );
CKINVDCx5p33_ASAP7_75t_R g578 ( .A(n_11), .Y(n_578) );
AOI22xp5_ASAP7_75t_L g545 ( .A1(n_12), .A2(n_19), .B1(n_546), .B2(n_547), .Y(n_545) );
BUFx2_ASAP7_75t_L g115 ( .A(n_13), .Y(n_115) );
OR2x2_ASAP7_75t_L g846 ( .A(n_13), .B(n_39), .Y(n_846) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_14), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g610 ( .A(n_15), .Y(n_610) );
AOI21xp5_ASAP7_75t_L g860 ( .A1(n_18), .A2(n_861), .B(n_868), .Y(n_860) );
AOI22xp5_ASAP7_75t_L g524 ( .A1(n_20), .A2(n_99), .B1(n_266), .B2(n_525), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_21), .A2(n_40), .B1(n_208), .B2(n_582), .Y(n_606) );
NAND2xp5_ASAP7_75t_SL g579 ( .A(n_22), .B(n_207), .Y(n_579) );
OAI21x1_ASAP7_75t_L g148 ( .A1(n_23), .A2(n_59), .B(n_149), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g255 ( .A(n_24), .Y(n_255) );
CKINVDCx5p33_ASAP7_75t_R g530 ( .A(n_26), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_27), .B(n_141), .Y(n_221) );
INVx4_ASAP7_75t_R g189 ( .A(n_28), .Y(n_189) );
AOI22xp33_ASAP7_75t_L g561 ( .A1(n_29), .A2(n_48), .B1(n_143), .B2(n_263), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_30), .A2(n_55), .B1(n_143), .B2(n_525), .Y(n_535) );
INVx1_ASAP7_75t_L g122 ( .A(n_31), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g594 ( .A(n_32), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_33), .B(n_582), .Y(n_581) );
CKINVDCx5p33_ASAP7_75t_R g571 ( .A(n_34), .Y(n_571) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_35), .B(n_165), .Y(n_228) );
INVx1_ASAP7_75t_L g270 ( .A(n_36), .Y(n_270) );
A2O1A1Ixp33_ASAP7_75t_SL g243 ( .A1(n_37), .A2(n_136), .B(n_140), .C(n_244), .Y(n_243) );
AOI22xp33_ASAP7_75t_L g252 ( .A1(n_38), .A2(n_56), .B1(n_136), .B2(n_143), .Y(n_252) );
HB1xp67_ASAP7_75t_L g117 ( .A(n_39), .Y(n_117) );
AOI22xp5_ASAP7_75t_L g590 ( .A1(n_41), .A2(n_87), .B1(n_136), .B2(n_591), .Y(n_590) );
CKINVDCx5p33_ASAP7_75t_R g241 ( .A(n_42), .Y(n_241) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_43), .A2(n_47), .B1(n_136), .B2(n_138), .Y(n_548) );
OAI22xp5_ASAP7_75t_L g851 ( .A1(n_45), .A2(n_69), .B1(n_852), .B2(n_853), .Y(n_851) );
CKINVDCx5p33_ASAP7_75t_R g853 ( .A(n_45), .Y(n_853) );
AOI22xp33_ASAP7_75t_L g526 ( .A1(n_46), .A2(n_60), .B1(n_525), .B2(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g872 ( .A(n_49), .Y(n_872) );
INVx1_ASAP7_75t_L g225 ( .A(n_50), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_51), .B(n_136), .Y(n_227) );
CKINVDCx5p33_ASAP7_75t_R g163 ( .A(n_52), .Y(n_163) );
INVx2_ASAP7_75t_L g841 ( .A(n_53), .Y(n_841) );
INVx1_ASAP7_75t_L g107 ( .A(n_54), .Y(n_107) );
BUFx3_ASAP7_75t_L g844 ( .A(n_54), .Y(n_844) );
CKINVDCx5p33_ASAP7_75t_R g191 ( .A(n_57), .Y(n_191) );
AOI22xp33_ASAP7_75t_L g142 ( .A1(n_58), .A2(n_88), .B1(n_136), .B2(n_143), .Y(n_142) );
CKINVDCx20_ASAP7_75t_R g870 ( .A(n_61), .Y(n_870) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_63), .A2(n_76), .B1(n_263), .B2(n_527), .Y(n_534) );
CKINVDCx5p33_ASAP7_75t_R g154 ( .A(n_64), .Y(n_154) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_65), .A2(n_79), .B1(n_136), .B2(n_138), .Y(n_569) );
AOI22xp5_ASAP7_75t_L g568 ( .A1(n_66), .A2(n_97), .B1(n_525), .B2(n_547), .Y(n_568) );
INVx1_ASAP7_75t_L g149 ( .A(n_67), .Y(n_149) );
AND2x4_ASAP7_75t_L g151 ( .A(n_68), .B(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g852 ( .A(n_69), .Y(n_852) );
AOI22xp33_ASAP7_75t_L g262 ( .A1(n_70), .A2(n_90), .B1(n_143), .B2(n_263), .Y(n_262) );
AO22x1_ASAP7_75t_L g205 ( .A1(n_71), .A2(n_77), .B1(n_206), .B2(n_208), .Y(n_205) );
INVx1_ASAP7_75t_L g152 ( .A(n_72), .Y(n_152) );
AND2x2_ASAP7_75t_L g247 ( .A(n_73), .B(n_159), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_74), .B(n_173), .Y(n_172) );
CKINVDCx5p33_ASAP7_75t_R g238 ( .A(n_75), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_78), .B(n_165), .Y(n_164) );
INVx2_ASAP7_75t_L g141 ( .A(n_80), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g186 ( .A(n_81), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_82), .B(n_159), .Y(n_218) );
AOI22xp33_ASAP7_75t_L g592 ( .A1(n_83), .A2(n_98), .B1(n_143), .B2(n_173), .Y(n_592) );
CKINVDCx5p33_ASAP7_75t_R g537 ( .A(n_84), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_85), .B(n_147), .Y(n_203) );
CKINVDCx5p33_ASAP7_75t_R g563 ( .A(n_86), .Y(n_563) );
NAND2xp5_ASAP7_75t_SL g585 ( .A(n_89), .B(n_159), .Y(n_585) );
CKINVDCx5p33_ASAP7_75t_R g551 ( .A(n_91), .Y(n_551) );
NAND2xp5_ASAP7_75t_SL g158 ( .A(n_92), .B(n_159), .Y(n_158) );
INVx1_ASAP7_75t_L g110 ( .A(n_93), .Y(n_110) );
NOR2xp33_ASAP7_75t_L g858 ( .A(n_93), .B(n_859), .Y(n_858) );
NAND2xp33_ASAP7_75t_L g583 ( .A(n_94), .B(n_207), .Y(n_583) );
A2O1A1Ixp33_ASAP7_75t_L g183 ( .A1(n_95), .A2(n_145), .B(n_173), .C(n_184), .Y(n_183) );
AND2x2_ASAP7_75t_L g193 ( .A(n_96), .B(n_194), .Y(n_193) );
NAND2xp33_ASAP7_75t_L g170 ( .A(n_100), .B(n_171), .Y(n_170) );
AOI21xp5_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_118), .B(n_871), .Y(n_101) );
NOR2xp33_ASAP7_75t_R g871 ( .A(n_102), .B(n_872), .Y(n_871) );
CKINVDCx10_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
OR2x6_ASAP7_75t_L g103 ( .A(n_104), .B(n_113), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
NOR2x1p5_ASAP7_75t_L g105 ( .A(n_106), .B(n_108), .Y(n_105) );
HB1xp67_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g859 ( .A(n_107), .Y(n_859) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_109), .B(n_111), .Y(n_108) );
BUFx6f_ASAP7_75t_L g835 ( .A(n_109), .Y(n_835) );
BUFx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
INVx2_ASAP7_75t_L g512 ( .A(n_110), .Y(n_512) );
INVx1_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
NOR2xp33_ASAP7_75t_L g114 ( .A(n_115), .B(n_116), .Y(n_114) );
INVxp33_ASAP7_75t_SL g116 ( .A(n_117), .Y(n_116) );
AO21x2_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_837), .B(n_847), .Y(n_118) );
OAI22xp5_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_121), .B1(n_124), .B2(n_836), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx2_ASAP7_75t_L g836 ( .A(n_124), .Y(n_836) );
OAI22x1_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_510), .B1(n_513), .B2(n_834), .Y(n_124) );
AND2x2_ASAP7_75t_L g125 ( .A(n_126), .B(n_419), .Y(n_125) );
NOR3xp33_ASAP7_75t_L g126 ( .A(n_127), .B(n_335), .C(n_366), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_128), .B(n_301), .Y(n_127) );
AOI211x1_ASAP7_75t_SL g128 ( .A1(n_129), .A2(n_213), .B(n_256), .C(n_287), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_131), .B(n_177), .Y(n_130) );
AND2x2_ASAP7_75t_L g442 ( .A(n_131), .B(n_317), .Y(n_442) );
AND2x2_ASAP7_75t_L g131 ( .A(n_132), .B(n_156), .Y(n_131) );
INVx1_ASAP7_75t_L g327 ( .A(n_132), .Y(n_327) );
OR2x2_ASAP7_75t_L g448 ( .A(n_132), .B(n_299), .Y(n_448) );
INVx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
AND2x2_ASAP7_75t_L g284 ( .A(n_133), .B(n_157), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_133), .B(n_299), .Y(n_298) );
INVx2_ASAP7_75t_L g316 ( .A(n_133), .Y(n_316) );
OR2x2_ASAP7_75t_L g347 ( .A(n_133), .B(n_178), .Y(n_347) );
AND2x2_ASAP7_75t_L g361 ( .A(n_133), .B(n_178), .Y(n_361) );
AND2x2_ASAP7_75t_L g398 ( .A(n_133), .B(n_354), .Y(n_398) );
AO31x2_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_146), .A3(n_150), .B(n_153), .Y(n_133) );
OAI22x1_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_139), .B1(n_142), .B2(n_144), .Y(n_134) );
INVx4_ASAP7_75t_L g138 ( .A(n_136), .Y(n_138) );
INVx1_ASAP7_75t_L g527 ( .A(n_136), .Y(n_527) );
INVx1_ASAP7_75t_L g547 ( .A(n_136), .Y(n_547) );
INVx3_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_137), .Y(n_143) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_137), .Y(n_165) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_137), .Y(n_171) );
INVx1_ASAP7_75t_L g173 ( .A(n_137), .Y(n_173) );
INVx1_ASAP7_75t_L g185 ( .A(n_137), .Y(n_185) );
INVx1_ASAP7_75t_L g190 ( .A(n_137), .Y(n_190) );
BUFx6f_ASAP7_75t_L g207 ( .A(n_137), .Y(n_207) );
INVx1_ASAP7_75t_L g209 ( .A(n_137), .Y(n_209) );
INVx1_ASAP7_75t_L g240 ( .A(n_137), .Y(n_240) );
INVx2_ASAP7_75t_L g246 ( .A(n_137), .Y(n_246) );
O2A1O1Ixp33_ASAP7_75t_L g162 ( .A1(n_138), .A2(n_163), .B(n_164), .C(n_166), .Y(n_162) );
O2A1O1Ixp5_ASAP7_75t_L g577 ( .A1(n_138), .A2(n_140), .B(n_578), .C(n_579), .Y(n_577) );
OAI22xp5_ASAP7_75t_L g250 ( .A1(n_139), .A2(n_199), .B1(n_251), .B2(n_252), .Y(n_250) );
OAI22xp5_ASAP7_75t_L g261 ( .A1(n_139), .A2(n_144), .B1(n_262), .B2(n_264), .Y(n_261) );
OAI22xp5_ASAP7_75t_L g523 ( .A1(n_139), .A2(n_524), .B1(n_526), .B2(n_528), .Y(n_523) );
OAI22xp5_ASAP7_75t_L g533 ( .A1(n_139), .A2(n_528), .B1(n_534), .B2(n_535), .Y(n_533) );
OAI22xp5_ASAP7_75t_L g544 ( .A1(n_139), .A2(n_545), .B1(n_548), .B2(n_549), .Y(n_544) );
OAI22xp5_ASAP7_75t_L g559 ( .A1(n_139), .A2(n_528), .B1(n_560), .B2(n_561), .Y(n_559) );
OAI22xp5_ASAP7_75t_L g567 ( .A1(n_139), .A2(n_549), .B1(n_568), .B2(n_569), .Y(n_567) );
AOI21xp5_ASAP7_75t_L g580 ( .A1(n_139), .A2(n_581), .B(n_583), .Y(n_580) );
OAI22xp5_ASAP7_75t_L g589 ( .A1(n_139), .A2(n_144), .B1(n_590), .B2(n_592), .Y(n_589) );
OAI22xp5_ASAP7_75t_L g605 ( .A1(n_139), .A2(n_528), .B1(n_606), .B2(n_607), .Y(n_605) );
INVx6_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
AOI21xp5_ASAP7_75t_L g169 ( .A1(n_140), .A2(n_170), .B(n_172), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_140), .B(n_205), .Y(n_204) );
A2O1A1Ixp33_ASAP7_75t_L g300 ( .A1(n_140), .A2(n_198), .B(n_205), .C(n_211), .Y(n_300) );
BUFx8_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx1_ASAP7_75t_L g145 ( .A(n_141), .Y(n_145) );
INVx2_ASAP7_75t_L g168 ( .A(n_141), .Y(n_168) );
INVx1_ASAP7_75t_L g224 ( .A(n_141), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_143), .B(n_223), .Y(n_222) );
INVx2_ASAP7_75t_L g265 ( .A(n_143), .Y(n_265) );
NAND2xp5_ASAP7_75t_SL g187 ( .A(n_144), .B(n_188), .Y(n_187) );
INVx1_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx1_ASAP7_75t_SL g549 ( .A(n_145), .Y(n_549) );
NOR2xp33_ASAP7_75t_L g529 ( .A(n_146), .B(n_530), .Y(n_529) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_146), .B(n_537), .Y(n_536) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx2_ASAP7_75t_L g155 ( .A(n_147), .Y(n_155) );
INVx2_ASAP7_75t_L g181 ( .A(n_147), .Y(n_181) );
OAI21xp33_ASAP7_75t_L g211 ( .A1(n_147), .A2(n_203), .B(n_212), .Y(n_211) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_148), .Y(n_160) );
INVx2_ASAP7_75t_L g192 ( .A(n_150), .Y(n_192) );
AO31x2_ASAP7_75t_L g543 ( .A1(n_150), .A2(n_234), .A3(n_544), .B(n_550), .Y(n_543) );
AO31x2_ASAP7_75t_L g558 ( .A1(n_150), .A2(n_253), .A3(n_559), .B(n_562), .Y(n_558) );
AO31x2_ASAP7_75t_L g604 ( .A1(n_150), .A2(n_588), .A3(n_605), .B(n_609), .Y(n_604) );
BUFx10_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
BUFx10_ASAP7_75t_L g176 ( .A(n_151), .Y(n_176) );
INVx1_ASAP7_75t_L g212 ( .A(n_151), .Y(n_212) );
INVx1_ASAP7_75t_L g268 ( .A(n_151), .Y(n_268) );
NOR2xp33_ASAP7_75t_L g153 ( .A(n_154), .B(n_155), .Y(n_153) );
INVx2_ASAP7_75t_L g194 ( .A(n_155), .Y(n_194) );
BUFx2_ASAP7_75t_L g234 ( .A(n_155), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g254 ( .A(n_155), .B(n_255), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g269 ( .A(n_155), .B(n_270), .Y(n_269) );
BUFx2_ASAP7_75t_L g278 ( .A(n_156), .Y(n_278) );
AND2x2_ASAP7_75t_L g329 ( .A(n_156), .B(n_195), .Y(n_329) );
AND2x2_ASAP7_75t_L g472 ( .A(n_156), .B(n_178), .Y(n_472) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
BUFx3_ASAP7_75t_L g296 ( .A(n_157), .Y(n_296) );
AND2x2_ASAP7_75t_L g315 ( .A(n_157), .B(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g352 ( .A(n_157), .Y(n_352) );
AND2x2_ASAP7_75t_L g376 ( .A(n_157), .B(n_178), .Y(n_376) );
NAND2x1p5_ASAP7_75t_L g157 ( .A(n_158), .B(n_161), .Y(n_157) );
NOR2x1_ASAP7_75t_L g174 ( .A(n_159), .B(n_175), .Y(n_174) );
INVx2_ASAP7_75t_L g253 ( .A(n_159), .Y(n_253) );
INVx4_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
AND2x2_ASAP7_75t_L g229 ( .A(n_160), .B(n_176), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g562 ( .A(n_160), .B(n_563), .Y(n_562) );
NOR2xp33_ASAP7_75t_L g570 ( .A(n_160), .B(n_571), .Y(n_570) );
INVx2_ASAP7_75t_SL g575 ( .A(n_160), .Y(n_575) );
BUFx3_ASAP7_75t_L g588 ( .A(n_160), .Y(n_588) );
NOR2xp33_ASAP7_75t_L g609 ( .A(n_160), .B(n_610), .Y(n_609) );
OAI21x1_ASAP7_75t_L g161 ( .A1(n_162), .A2(n_169), .B(n_174), .Y(n_161) );
NOR2xp33_ASAP7_75t_L g237 ( .A(n_165), .B(n_238), .Y(n_237) );
INVx2_ASAP7_75t_SL g166 ( .A(n_167), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
BUFx3_ASAP7_75t_L g200 ( .A(n_168), .Y(n_200) );
OAI22xp33_ASAP7_75t_L g188 ( .A1(n_171), .A2(n_189), .B1(n_190), .B2(n_191), .Y(n_188) );
INVx2_ASAP7_75t_L g263 ( .A(n_171), .Y(n_263) );
INVx1_ASAP7_75t_L g582 ( .A(n_171), .Y(n_582) );
INVx1_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
AO31x2_ASAP7_75t_L g249 ( .A1(n_176), .A2(n_250), .A3(n_253), .B(n_254), .Y(n_249) );
HB1xp67_ASAP7_75t_L g276 ( .A(n_177), .Y(n_276) );
AND2x2_ASAP7_75t_L g337 ( .A(n_177), .B(n_326), .Y(n_337) );
INVx2_ASAP7_75t_L g469 ( .A(n_177), .Y(n_469) );
AND2x2_ASAP7_75t_L g177 ( .A(n_178), .B(n_195), .Y(n_177) );
INVx1_ASAP7_75t_L g274 ( .A(n_178), .Y(n_274) );
AND2x4_ASAP7_75t_L g286 ( .A(n_178), .B(n_196), .Y(n_286) );
INVx2_ASAP7_75t_L g354 ( .A(n_178), .Y(n_354) );
AO21x2_ASAP7_75t_L g178 ( .A1(n_179), .A2(n_182), .B(n_193), .Y(n_178) );
AO31x2_ASAP7_75t_L g521 ( .A1(n_179), .A2(n_522), .A3(n_523), .B(n_529), .Y(n_521) );
AO31x2_ASAP7_75t_L g532 ( .A1(n_179), .A2(n_267), .A3(n_533), .B(n_536), .Y(n_532) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
NOR2xp33_ASAP7_75t_SL g550 ( .A(n_181), .B(n_551), .Y(n_550) );
NOR2xp33_ASAP7_75t_L g593 ( .A(n_181), .B(n_594), .Y(n_593) );
AOI21xp5_ASAP7_75t_L g182 ( .A1(n_183), .A2(n_187), .B(n_192), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g184 ( .A(n_185), .B(n_186), .Y(n_184) );
INVx2_ASAP7_75t_L g202 ( .A(n_185), .Y(n_202) );
INVx1_ASAP7_75t_L g608 ( .A(n_190), .Y(n_608) );
INVx1_ASAP7_75t_L g522 ( .A(n_192), .Y(n_522) );
AND2x2_ASAP7_75t_L g353 ( .A(n_195), .B(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g360 ( .A(n_195), .Y(n_360) );
INVx2_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
AND2x2_ASAP7_75t_L g438 ( .A(n_196), .B(n_354), .Y(n_438) );
AOI21x1_ASAP7_75t_L g196 ( .A1(n_197), .A2(n_204), .B(n_210), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
OAI21x1_ASAP7_75t_L g198 ( .A1(n_199), .A2(n_201), .B(n_203), .Y(n_198) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_199), .A2(n_227), .B(n_228), .Y(n_226) );
INVx2_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
INVx2_ASAP7_75t_L g528 ( .A(n_200), .Y(n_528) );
INVx1_ASAP7_75t_L g546 ( .A(n_202), .Y(n_546) );
INVxp67_ASAP7_75t_SL g206 ( .A(n_207), .Y(n_206) );
INVx3_ASAP7_75t_L g525 ( .A(n_207), .Y(n_525) );
OAI21xp33_ASAP7_75t_SL g220 ( .A1(n_208), .A2(n_221), .B(n_222), .Y(n_220) );
INVx1_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx1_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_212), .A2(n_236), .B(n_243), .Y(n_235) );
INVx1_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_215), .B(n_230), .Y(n_214) );
OR2x2_ASAP7_75t_L g343 ( .A(n_215), .B(n_231), .Y(n_343) );
AND2x2_ASAP7_75t_L g481 ( .A(n_215), .B(n_425), .Y(n_481) );
INVx2_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
AND2x4_ASAP7_75t_L g258 ( .A(n_216), .B(n_259), .Y(n_258) );
OR2x2_ASAP7_75t_L g363 ( .A(n_216), .B(n_364), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_216), .B(n_305), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_216), .B(n_281), .Y(n_418) );
INVx3_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx1_ASAP7_75t_L g275 ( .A(n_217), .Y(n_275) );
AND2x2_ASAP7_75t_L g291 ( .A(n_217), .B(n_292), .Y(n_291) );
NAND2x1p5_ASAP7_75t_SL g304 ( .A(n_217), .B(n_305), .Y(n_304) );
OR2x2_ASAP7_75t_L g312 ( .A(n_217), .B(n_313), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_217), .B(n_281), .Y(n_383) );
AND2x2_ASAP7_75t_L g431 ( .A(n_217), .B(n_260), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_217), .B(n_259), .Y(n_474) );
BUFx2_ASAP7_75t_L g493 ( .A(n_217), .Y(n_493) );
AND2x4_ASAP7_75t_L g217 ( .A(n_218), .B(n_219), .Y(n_217) );
OAI21xp5_ASAP7_75t_L g219 ( .A1(n_220), .A2(n_226), .B(n_229), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_224), .B(n_225), .Y(n_223) );
BUFx4f_ASAP7_75t_L g242 ( .A(n_224), .Y(n_242) );
INVx1_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
OR2x2_ASAP7_75t_L g277 ( .A(n_231), .B(n_278), .Y(n_277) );
INVx2_ASAP7_75t_L g390 ( .A(n_231), .Y(n_390) );
OR2x2_ASAP7_75t_L g231 ( .A(n_232), .B(n_248), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g293 ( .A(n_232), .B(n_260), .Y(n_293) );
INVx2_ASAP7_75t_L g305 ( .A(n_232), .Y(n_305) );
AND2x2_ASAP7_75t_L g341 ( .A(n_232), .B(n_249), .Y(n_341) );
INVx2_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
INVx1_ASAP7_75t_L g281 ( .A(n_233), .Y(n_281) );
AOI21x1_ASAP7_75t_L g233 ( .A1(n_234), .A2(n_235), .B(n_247), .Y(n_233) );
AO31x2_ASAP7_75t_L g260 ( .A1(n_234), .A2(n_261), .A3(n_267), .B(n_269), .Y(n_260) );
AO31x2_ASAP7_75t_L g566 ( .A1(n_234), .A2(n_522), .A3(n_567), .B(n_570), .Y(n_566) );
OAI21xp5_ASAP7_75t_L g236 ( .A1(n_237), .A2(n_239), .B(n_242), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_240), .B(n_241), .Y(n_239) );
INVx2_ASAP7_75t_L g266 ( .A(n_240), .Y(n_266) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_245), .B(n_246), .Y(n_244) );
INVx2_ASAP7_75t_SL g591 ( .A(n_246), .Y(n_591) );
INVx1_ASAP7_75t_L g365 ( .A(n_248), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_248), .B(n_260), .Y(n_382) );
INVx2_ASAP7_75t_SL g248 ( .A(n_249), .Y(n_248) );
BUFx2_ASAP7_75t_L g292 ( .A(n_249), .Y(n_292) );
OR2x2_ASAP7_75t_L g324 ( .A(n_249), .B(n_260), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_249), .B(n_260), .Y(n_402) );
OAI22xp5_ASAP7_75t_L g256 ( .A1(n_257), .A2(n_277), .B1(n_279), .B2(n_283), .Y(n_256) );
AOI22xp5_ASAP7_75t_L g257 ( .A1(n_258), .A2(n_271), .B1(n_275), .B2(n_276), .Y(n_257) );
INVx2_ASAP7_75t_L g282 ( .A(n_258), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_258), .B(n_341), .Y(n_355) );
AND2x2_ASAP7_75t_L g389 ( .A(n_258), .B(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
INVx1_ASAP7_75t_L g307 ( .A(n_260), .Y(n_307) );
INVx1_ASAP7_75t_L g313 ( .A(n_260), .Y(n_313) );
AO31x2_ASAP7_75t_L g587 ( .A1(n_267), .A2(n_588), .A3(n_589), .B(n_593), .Y(n_587) );
INVx2_ASAP7_75t_SL g267 ( .A(n_268), .Y(n_267) );
INVx2_ASAP7_75t_SL g584 ( .A(n_268), .Y(n_584) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
OR2x2_ASAP7_75t_L g447 ( .A(n_273), .B(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
INVx1_ASAP7_75t_L g328 ( .A(n_274), .Y(n_328) );
AND3x1_ASAP7_75t_L g432 ( .A(n_274), .B(n_295), .C(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g388 ( .A(n_275), .Y(n_388) );
AND2x4_ASAP7_75t_L g424 ( .A(n_275), .B(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g462 ( .A(n_278), .Y(n_462) );
INVx1_ASAP7_75t_L g466 ( .A(n_279), .Y(n_466) );
OR2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_282), .Y(n_279) );
OR2x2_ASAP7_75t_L g439 ( .A(n_280), .B(n_440), .Y(n_439) );
INVxp67_ASAP7_75t_SL g487 ( .A(n_280), .Y(n_487) );
INVxp67_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
OR2x2_ASAP7_75t_L g387 ( .A(n_281), .B(n_365), .Y(n_387) );
AND2x2_ASAP7_75t_L g429 ( .A(n_281), .B(n_296), .Y(n_429) );
HB1xp67_ASAP7_75t_L g433 ( .A(n_281), .Y(n_433) );
NAND2xp5_ASAP7_75t_SL g283 ( .A(n_284), .B(n_285), .Y(n_283) );
O2A1O1Ixp33_ASAP7_75t_L g348 ( .A1(n_284), .A2(n_285), .B(n_349), .C(n_355), .Y(n_348) );
NAND2x1_ASAP7_75t_L g392 ( .A(n_284), .B(n_393), .Y(n_392) );
NOR2xp33_ASAP7_75t_L g488 ( .A(n_284), .B(n_442), .Y(n_488) );
INVx3_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_286), .B(n_315), .Y(n_334) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
NAND2xp5_ASAP7_75t_SL g288 ( .A(n_289), .B(n_294), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_291), .B(n_293), .Y(n_290) );
INVx2_ASAP7_75t_L g310 ( .A(n_292), .Y(n_310) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_293), .Y(n_371) );
NOR2xp33_ASAP7_75t_L g435 ( .A(n_294), .B(n_436), .Y(n_435) );
AND2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_297), .Y(n_294) );
AND2x2_ASAP7_75t_L g344 ( .A(n_295), .B(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_295), .B(n_361), .Y(n_408) );
NAND2x1p5_ASAP7_75t_L g414 ( .A(n_295), .B(n_415), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_295), .B(n_353), .Y(n_509) );
INVx3_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
BUFx2_ASAP7_75t_L g492 ( .A(n_296), .Y(n_492) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx2_ASAP7_75t_L g318 ( .A(n_299), .Y(n_318) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
AOI21xp5_ASAP7_75t_L g301 ( .A1(n_302), .A2(n_314), .B(n_319), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_303), .B(n_308), .Y(n_302) );
OR2x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_306), .Y(n_303) );
OAI33xp33_ASAP7_75t_L g368 ( .A1(n_304), .A2(n_309), .A3(n_369), .B1(n_370), .B2(n_372), .B3(n_373), .Y(n_368) );
OR2x2_ASAP7_75t_L g500 ( .A(n_304), .B(n_324), .Y(n_500) );
INVx2_ASAP7_75t_L g502 ( .A(n_304), .Y(n_502) );
INVx1_ASAP7_75t_L g323 ( .A(n_305), .Y(n_323) );
OR2x2_ASAP7_75t_L g364 ( .A(n_305), .B(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_309), .B(n_311), .Y(n_308) );
INVx1_ASAP7_75t_L g372 ( .A(n_309), .Y(n_372) );
NOR3xp33_ASAP7_75t_L g490 ( .A(n_309), .B(n_491), .C(n_493), .Y(n_490) );
INVx2_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
NOR2xp33_ASAP7_75t_L g449 ( .A(n_310), .B(n_450), .Y(n_449) );
NOR2xp33_ASAP7_75t_L g478 ( .A(n_310), .B(n_474), .Y(n_478) );
AND2x4_ASAP7_75t_L g507 ( .A(n_310), .B(n_508), .Y(n_507) );
INVxp67_ASAP7_75t_SL g311 ( .A(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g333 ( .A(n_312), .Y(n_333) );
OR2x2_ASAP7_75t_L g339 ( .A(n_312), .B(n_340), .Y(n_339) );
OR2x2_ASAP7_75t_L g452 ( .A(n_312), .B(n_387), .Y(n_452) );
INVx1_ASAP7_75t_L g508 ( .A(n_312), .Y(n_508) );
AND2x4_ASAP7_75t_SL g314 ( .A(n_315), .B(n_317), .Y(n_314) );
INVx1_ASAP7_75t_L g331 ( .A(n_315), .Y(n_331) );
INVx1_ASAP7_75t_L g374 ( .A(n_316), .Y(n_374) );
AND2x2_ASAP7_75t_L g415 ( .A(n_316), .B(n_318), .Y(n_415) );
INVx1_ASAP7_75t_L g455 ( .A(n_317), .Y(n_455) );
INVx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
OR2x2_ASAP7_75t_L g346 ( .A(n_318), .B(n_347), .Y(n_346) );
OAI22xp33_ASAP7_75t_L g319 ( .A1(n_320), .A2(n_325), .B1(n_332), .B2(n_334), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx2_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
OR2x2_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
INVx2_ASAP7_75t_L g411 ( .A(n_324), .Y(n_411) );
INVx2_ASAP7_75t_L g425 ( .A(n_324), .Y(n_425) );
AOI211xp5_ASAP7_75t_L g325 ( .A1(n_326), .A2(n_328), .B(n_329), .C(n_330), .Y(n_325) );
INVx1_ASAP7_75t_L g369 ( .A(n_326), .Y(n_369) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_327), .B(n_352), .Y(n_454) );
OR2x2_ASAP7_75t_L g470 ( .A(n_327), .B(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g483 ( .A(n_327), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_329), .B(n_397), .Y(n_458) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
NAND2xp5_ASAP7_75t_SL g335 ( .A(n_336), .B(n_356), .Y(n_335) );
AOI221xp5_ASAP7_75t_L g336 ( .A1(n_337), .A2(n_338), .B1(n_342), .B2(n_344), .C(n_348), .Y(n_336) );
INVx2_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
OAI32xp33_ASAP7_75t_L g505 ( .A1(n_339), .A2(n_436), .A3(n_454), .B1(n_506), .B2(n_509), .Y(n_505) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g475 ( .A(n_341), .Y(n_475) );
INVx2_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
OAI21xp5_ASAP7_75t_L g356 ( .A1(n_344), .A2(n_357), .B(n_362), .Y(n_356) );
NAND2x1_ASAP7_75t_L g504 ( .A(n_345), .B(n_492), .Y(n_504) );
INVx2_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx2_ASAP7_75t_L g379 ( .A(n_347), .Y(n_379) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_351), .B(n_353), .Y(n_350) );
AND2x2_ASAP7_75t_L g498 ( .A(n_351), .B(n_379), .Y(n_498) );
INVx2_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g446 ( .A(n_352), .Y(n_446) );
INVx2_ASAP7_75t_L g399 ( .A(n_353), .Y(n_399) );
INVx2_ASAP7_75t_SL g357 ( .A(n_358), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_359), .B(n_361), .Y(n_358) );
AND2x2_ASAP7_75t_L g375 ( .A(n_359), .B(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx2_ASAP7_75t_L g394 ( .A(n_360), .Y(n_394) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
NAND4xp25_ASAP7_75t_L g366 ( .A(n_367), .B(n_384), .C(n_395), .D(n_406), .Y(n_366) );
AOI22xp5_ASAP7_75t_L g367 ( .A1(n_368), .A2(n_375), .B1(n_377), .B2(n_380), .Y(n_367) );
OAI22xp5_ASAP7_75t_L g496 ( .A1(n_369), .A2(n_497), .B1(n_499), .B2(n_500), .Y(n_496) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
AND2x2_ASAP7_75t_L g479 ( .A(n_374), .B(n_438), .Y(n_479) );
AND2x2_ASAP7_75t_L g482 ( .A(n_376), .B(n_483), .Y(n_482) );
AOI22xp5_ASAP7_75t_L g395 ( .A1(n_377), .A2(n_396), .B1(n_400), .B2(n_403), .Y(n_395) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx2_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
OR2x2_ASAP7_75t_L g381 ( .A(n_382), .B(n_383), .Y(n_381) );
OR2x2_ASAP7_75t_L g417 ( .A(n_382), .B(n_418), .Y(n_417) );
OR2x2_ASAP7_75t_L g401 ( .A(n_383), .B(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g412 ( .A(n_383), .Y(n_412) );
OAI21xp5_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_389), .B(n_391), .Y(n_384) );
O2A1O1Ixp33_ASAP7_75t_L g489 ( .A1(n_385), .A2(n_490), .B(n_494), .C(n_496), .Y(n_489) );
AND2x2_ASAP7_75t_L g385 ( .A(n_386), .B(n_388), .Y(n_385) );
INVxp67_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g464 ( .A(n_387), .Y(n_464) );
AND2x4_ASAP7_75t_L g457 ( .A(n_390), .B(n_431), .Y(n_457) );
INVx2_ASAP7_75t_SL g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_397), .B(n_399), .Y(n_396) );
OAI21xp33_ASAP7_75t_L g422 ( .A1(n_397), .A2(n_423), .B(n_426), .Y(n_422) );
INVx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
AND2x2_ASAP7_75t_L g428 ( .A(n_398), .B(n_429), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_398), .B(n_462), .Y(n_461) );
INVx2_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
OR2x2_ASAP7_75t_L g404 ( .A(n_402), .B(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
OAI22xp5_ASAP7_75t_L g434 ( .A1(n_404), .A2(n_435), .B1(n_439), .B2(n_441), .Y(n_434) );
AOI22xp33_ASAP7_75t_L g406 ( .A1(n_407), .A2(n_409), .B1(n_413), .B2(n_416), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_411), .B(n_412), .Y(n_410) );
HB1xp67_ASAP7_75t_L g427 ( .A(n_411), .Y(n_427) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
NOR2xp33_ASAP7_75t_L g419 ( .A(n_420), .B(n_484), .Y(n_419) );
NAND4xp25_ASAP7_75t_L g420 ( .A(n_421), .B(n_443), .C(n_459), .D(n_476), .Y(n_420) );
NOR2xp33_ASAP7_75t_L g421 ( .A(n_422), .B(n_434), .Y(n_421) );
INVx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
AND2x2_ASAP7_75t_L g486 ( .A(n_424), .B(n_487), .Y(n_486) );
AOI22xp5_ASAP7_75t_L g426 ( .A1(n_427), .A2(n_428), .B1(n_430), .B2(n_432), .Y(n_426) );
INVxp67_ASAP7_75t_L g450 ( .A(n_430), .Y(n_450) );
BUFx2_ASAP7_75t_SL g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g440 ( .A(n_431), .Y(n_440) );
AND2x2_ASAP7_75t_L g463 ( .A(n_431), .B(n_464), .Y(n_463) );
INVx3_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
AOI21xp5_ASAP7_75t_L g443 ( .A1(n_444), .A2(n_449), .B(n_451), .Y(n_443) );
NOR2x1_ASAP7_75t_L g444 ( .A(n_445), .B(n_447), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
OR2x6_ASAP7_75t_L g468 ( .A(n_446), .B(n_469), .Y(n_468) );
INVx3_ASAP7_75t_L g465 ( .A(n_447), .Y(n_465) );
OAI32xp33_ASAP7_75t_L g451 ( .A1(n_452), .A2(n_453), .A3(n_455), .B1(n_456), .B2(n_458), .Y(n_451) );
INVx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
AOI221xp5_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_463), .B1(n_465), .B2(n_466), .C(n_467), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
AOI21xp5_ASAP7_75t_L g467 ( .A1(n_468), .A2(n_470), .B(n_473), .Y(n_467) );
INVx2_ASAP7_75t_SL g471 ( .A(n_472), .Y(n_471) );
OR2x2_ASAP7_75t_L g473 ( .A(n_474), .B(n_475), .Y(n_473) );
NOR2x1_ASAP7_75t_L g476 ( .A(n_477), .B(n_480), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_478), .B(n_479), .Y(n_477) );
INVx1_ASAP7_75t_L g499 ( .A(n_478), .Y(n_499) );
INVx1_ASAP7_75t_L g495 ( .A(n_479), .Y(n_495) );
AND2x2_ASAP7_75t_L g480 ( .A(n_481), .B(n_482), .Y(n_480) );
OAI211xp5_ASAP7_75t_SL g484 ( .A1(n_485), .A2(n_488), .B(n_489), .C(n_501), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVxp67_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx1_ASAP7_75t_SL g497 ( .A(n_498), .Y(n_497) );
AOI21xp33_ASAP7_75t_L g501 ( .A1(n_502), .A2(n_503), .B(n_505), .Y(n_501) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
CKINVDCx5p33_ASAP7_75t_R g510 ( .A(n_511), .Y(n_510) );
BUFx8_ASAP7_75t_SL g511 ( .A(n_512), .Y(n_511) );
AND2x2_ASAP7_75t_L g866 ( .A(n_512), .B(n_867), .Y(n_866) );
XNOR2x1_ASAP7_75t_L g850 ( .A(n_513), .B(n_851), .Y(n_850) );
AND3x4_ASAP7_75t_L g513 ( .A(n_514), .B(n_696), .C(n_750), .Y(n_513) );
NOR2x1_ASAP7_75t_L g514 ( .A(n_515), .B(n_656), .Y(n_514) );
NAND3xp33_ASAP7_75t_L g515 ( .A(n_516), .B(n_595), .C(n_638), .Y(n_515) );
OAI21xp33_ASAP7_75t_L g516 ( .A1(n_517), .A2(n_538), .B(n_553), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
HB1xp67_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
OR2x2_ASAP7_75t_L g688 ( .A(n_519), .B(n_599), .Y(n_688) );
INVx2_ASAP7_75t_L g714 ( .A(n_519), .Y(n_714) );
OR2x2_ASAP7_75t_L g519 ( .A(n_520), .B(n_531), .Y(n_519) );
INVx1_ASAP7_75t_L g613 ( .A(n_520), .Y(n_613) );
INVx2_ASAP7_75t_L g728 ( .A(n_520), .Y(n_728) );
INVx2_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx2_ASAP7_75t_L g541 ( .A(n_521), .Y(n_541) );
AND2x4_ASAP7_75t_L g671 ( .A(n_521), .B(n_633), .Y(n_671) );
INVx1_ASAP7_75t_L g724 ( .A(n_531), .Y(n_724) );
INVx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g552 ( .A(n_532), .Y(n_552) );
AND2x4_ASAP7_75t_L g602 ( .A(n_532), .B(n_603), .Y(n_602) );
HB1xp67_ASAP7_75t_L g630 ( .A(n_532), .Y(n_630) );
INVx2_ASAP7_75t_L g633 ( .A(n_532), .Y(n_633) );
OR2x2_ASAP7_75t_L g647 ( .A(n_532), .B(n_604), .Y(n_647) );
AND2x2_ASAP7_75t_L g749 ( .A(n_532), .B(n_543), .Y(n_749) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g804 ( .A(n_539), .B(n_805), .Y(n_804) );
OR2x2_ASAP7_75t_L g539 ( .A(n_540), .B(n_542), .Y(n_539) );
OR2x2_ASAP7_75t_L g631 ( .A(n_540), .B(n_632), .Y(n_631) );
NAND2xp5_ASAP7_75t_SL g695 ( .A(n_540), .B(n_650), .Y(n_695) );
AND2x2_ASAP7_75t_L g760 ( .A(n_540), .B(n_736), .Y(n_760) );
INVx4_ASAP7_75t_L g794 ( .A(n_540), .Y(n_794) );
INVx3_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g629 ( .A(n_541), .B(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g667 ( .A(n_541), .B(n_601), .Y(n_667) );
AND2x2_ASAP7_75t_L g777 ( .A(n_541), .B(n_604), .Y(n_777) );
AND2x2_ASAP7_75t_L g811 ( .A(n_541), .B(n_633), .Y(n_811) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_543), .B(n_552), .Y(n_542) );
INVx4_ASAP7_75t_SL g601 ( .A(n_543), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_543), .B(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g712 ( .A(n_543), .B(n_604), .Y(n_712) );
BUFx2_ASAP7_75t_L g730 ( .A(n_543), .Y(n_730) );
AOI222xp33_ASAP7_75t_L g638 ( .A1(n_552), .A2(n_639), .B1(n_644), .B2(n_645), .C1(n_648), .C2(n_652), .Y(n_638) );
INVx1_ASAP7_75t_L g769 ( .A(n_552), .Y(n_769) );
AND2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_564), .Y(n_553) );
AND2x2_ASAP7_75t_L g806 ( .A(n_554), .B(n_618), .Y(n_806) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g827 ( .A(n_555), .B(n_828), .Y(n_827) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
AND2x4_ASAP7_75t_L g636 ( .A(n_556), .B(n_637), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_556), .B(n_619), .Y(n_775) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_557), .B(n_623), .Y(n_665) );
AND2x2_ASAP7_75t_L g693 ( .A(n_557), .B(n_573), .Y(n_693) );
INVx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
AND2x2_ASAP7_75t_L g622 ( .A(n_558), .B(n_623), .Y(n_622) );
OR2x2_ASAP7_75t_L g655 ( .A(n_558), .B(n_587), .Y(n_655) );
INVx1_ASAP7_75t_L g683 ( .A(n_558), .Y(n_683) );
HB1xp67_ASAP7_75t_L g789 ( .A(n_558), .Y(n_789) );
AOI222xp33_ASAP7_75t_L g738 ( .A1(n_564), .A2(n_681), .B1(n_739), .B2(n_740), .C1(n_742), .C2(n_744), .Y(n_738) );
AND2x4_ASAP7_75t_L g564 ( .A(n_565), .B(n_572), .Y(n_564) );
INVx1_ASAP7_75t_L g673 ( .A(n_565), .Y(n_673) );
BUFx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx3_ASAP7_75t_L g619 ( .A(n_566), .Y(n_619) );
AND2x2_ASAP7_75t_L g624 ( .A(n_566), .B(n_587), .Y(n_624) );
AND2x2_ASAP7_75t_L g684 ( .A(n_566), .B(n_586), .Y(n_684) );
AND2x2_ASAP7_75t_L g672 ( .A(n_572), .B(n_673), .Y(n_672) );
AND2x4_ASAP7_75t_L g767 ( .A(n_572), .B(n_683), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_572), .B(n_774), .Y(n_773) );
AND3x1_ASAP7_75t_L g832 ( .A(n_572), .B(n_602), .C(n_833), .Y(n_832) );
AND2x4_ASAP7_75t_L g572 ( .A(n_573), .B(n_586), .Y(n_572) );
AND2x2_ASAP7_75t_L g653 ( .A(n_573), .B(n_619), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g802 ( .A(n_573), .B(n_755), .Y(n_802) );
INVx2_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
BUFx2_ASAP7_75t_L g616 ( .A(n_574), .Y(n_616) );
OAI21x1_ASAP7_75t_L g574 ( .A1(n_575), .A2(n_576), .B(n_585), .Y(n_574) );
OAI21x1_ASAP7_75t_L g623 ( .A1(n_575), .A2(n_576), .B(n_585), .Y(n_623) );
OAI21x1_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_580), .B(n_584), .Y(n_576) );
INVx2_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
AND2x4_ASAP7_75t_L g618 ( .A(n_587), .B(n_619), .Y(n_618) );
OR2x2_ASAP7_75t_L g651 ( .A(n_587), .B(n_637), .Y(n_651) );
INVx1_ASAP7_75t_L g661 ( .A(n_587), .Y(n_661) );
BUFx2_ASAP7_75t_L g755 ( .A(n_587), .Y(n_755) );
AOI21xp5_ASAP7_75t_L g595 ( .A1(n_596), .A2(n_614), .B(n_620), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
NAND2x1_ASAP7_75t_L g597 ( .A(n_598), .B(n_611), .Y(n_597) );
AOI221xp5_ASAP7_75t_SL g678 ( .A1(n_598), .A2(n_679), .B1(n_685), .B2(n_689), .C(n_694), .Y(n_678) );
AND2x4_ASAP7_75t_L g598 ( .A(n_599), .B(n_602), .Y(n_598) );
INVx2_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_600), .B(n_613), .Y(n_799) );
INVx2_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_601), .B(n_633), .Y(n_632) );
AND2x4_ASAP7_75t_L g641 ( .A(n_601), .B(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g677 ( .A(n_601), .Y(n_677) );
INVx1_ASAP7_75t_L g687 ( .A(n_601), .Y(n_687) );
AND2x2_ASAP7_75t_L g706 ( .A(n_601), .B(n_707), .Y(n_706) );
OR2x2_ASAP7_75t_L g718 ( .A(n_601), .B(n_719), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g831 ( .A(n_601), .B(n_724), .Y(n_831) );
INVx2_ASAP7_75t_L g666 ( .A(n_602), .Y(n_666) );
AND2x2_ASAP7_75t_L g676 ( .A(n_602), .B(n_677), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_602), .B(n_687), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g819 ( .A(n_602), .B(n_820), .Y(n_819) );
INVx2_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g627 ( .A(n_604), .Y(n_627) );
HB1xp67_ASAP7_75t_L g670 ( .A(n_604), .Y(n_670) );
INVx1_ASAP7_75t_L g707 ( .A(n_604), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_604), .B(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
OR2x2_ASAP7_75t_L g646 ( .A(n_612), .B(n_647), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_612), .B(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
HB1xp67_ASAP7_75t_L g705 ( .A(n_613), .Y(n_705) );
NOR2xp33_ASAP7_75t_R g614 ( .A(n_615), .B(n_617), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
NOR3xp33_ASAP7_75t_L g694 ( .A(n_616), .B(n_686), .C(n_695), .Y(n_694) );
AND2x2_ASAP7_75t_L g717 ( .A(n_616), .B(n_624), .Y(n_717) );
AND2x2_ASAP7_75t_L g746 ( .A(n_616), .B(n_716), .Y(n_746) );
OR2x2_ASAP7_75t_L g813 ( .A(n_616), .B(n_814), .Y(n_813) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
AND2x4_ASAP7_75t_L g739 ( .A(n_618), .B(n_622), .Y(n_739) );
INVx2_ASAP7_75t_SL g823 ( .A(n_618), .Y(n_823) );
INVx2_ASAP7_75t_L g650 ( .A(n_619), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_619), .B(n_664), .Y(n_663) );
INVx3_ASAP7_75t_L g692 ( .A(n_619), .Y(n_692) );
HB1xp67_ASAP7_75t_L g765 ( .A(n_619), .Y(n_765) );
OAI32xp33_ASAP7_75t_L g620 ( .A1(n_621), .A2(n_625), .A3(n_628), .B1(n_631), .B2(n_634), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_622), .B(n_624), .Y(n_621) );
AND2x2_ASAP7_75t_L g644 ( .A(n_622), .B(n_624), .Y(n_644) );
AND2x2_ASAP7_75t_L g702 ( .A(n_622), .B(n_684), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_622), .B(n_684), .Y(n_710) );
INVx1_ASAP7_75t_L g637 ( .A(n_623), .Y(n_637) );
AND2x4_ASAP7_75t_SL g635 ( .A(n_624), .B(n_636), .Y(n_635) );
INVx1_ASAP7_75t_SL g779 ( .A(n_624), .Y(n_779) );
INVx2_ASAP7_75t_L g814 ( .A(n_624), .Y(n_814) );
AND2x2_ASAP7_75t_L g826 ( .A(n_624), .B(n_693), .Y(n_826) );
NOR3xp33_ASAP7_75t_L g756 ( .A(n_625), .B(n_747), .C(n_757), .Y(n_756) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g642 ( .A(n_627), .Y(n_642) );
AOI321xp33_ASAP7_75t_L g825 ( .A1(n_628), .A2(n_687), .A3(n_826), .B1(n_827), .B2(n_829), .C(n_832), .Y(n_825) );
INVx2_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g643 ( .A(n_630), .Y(n_643) );
OAI22xp5_ASAP7_75t_L g829 ( .A1(n_632), .A2(n_651), .B1(n_830), .B2(n_831), .Y(n_829) );
INVx3_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_L g732 ( .A(n_636), .B(n_691), .Y(n_732) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
NAND2xp5_ASAP7_75t_SL g640 ( .A(n_641), .B(n_643), .Y(n_640) );
INVx1_ASAP7_75t_L g766 ( .A(n_641), .Y(n_766) );
NAND2x1_ASAP7_75t_L g793 ( .A(n_641), .B(n_794), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g810 ( .A(n_641), .B(n_811), .Y(n_810) );
AND2x2_ASAP7_75t_L g791 ( .A(n_643), .B(n_777), .Y(n_791) );
INVx2_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx2_ASAP7_75t_L g731 ( .A(n_647), .Y(n_731) );
OR2x2_ASAP7_75t_L g798 ( .A(n_647), .B(n_799), .Y(n_798) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
OR2x2_ASAP7_75t_L g649 ( .A(n_650), .B(n_651), .Y(n_649) );
NOR2xp33_ASAP7_75t_L g675 ( .A(n_650), .B(n_651), .Y(n_675) );
NOR2x1p5_ASAP7_75t_L g716 ( .A(n_650), .B(n_655), .Y(n_716) );
INVx1_ASAP7_75t_L g786 ( .A(n_650), .Y(n_786) );
NOR2x1_ASAP7_75t_L g787 ( .A(n_651), .B(n_788), .Y(n_787) );
AND2x2_ASAP7_75t_L g652 ( .A(n_653), .B(n_654), .Y(n_652) );
INVxp67_ASAP7_75t_SL g830 ( .A(n_653), .Y(n_830) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
NAND3xp33_ASAP7_75t_L g656 ( .A(n_657), .B(n_668), .C(n_678), .Y(n_656) );
NAND3xp33_ASAP7_75t_L g657 ( .A(n_658), .B(n_666), .C(n_667), .Y(n_657) );
AND2x4_ASAP7_75t_L g658 ( .A(n_659), .B(n_662), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
BUFx2_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g808 ( .A(n_662), .Y(n_808) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVxp67_ASAP7_75t_SL g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g700 ( .A(n_665), .Y(n_700) );
INVx1_ASAP7_75t_L g736 ( .A(n_665), .Y(n_736) );
NAND2xp33_ASAP7_75t_L g740 ( .A(n_666), .B(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g744 ( .A(n_666), .Y(n_744) );
INVx1_ASAP7_75t_L g770 ( .A(n_667), .Y(n_770) );
AOI21xp5_ASAP7_75t_L g668 ( .A1(n_669), .A2(n_672), .B(n_674), .Y(n_668) );
AND2x4_ASAP7_75t_L g669 ( .A(n_670), .B(n_671), .Y(n_669) );
INVx3_ASAP7_75t_L g719 ( .A(n_671), .Y(n_719) );
AND2x2_ASAP7_75t_L g674 ( .A(n_675), .B(n_676), .Y(n_674) );
INVxp67_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
AND2x2_ASAP7_75t_L g681 ( .A(n_682), .B(n_684), .Y(n_681) );
INVx2_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
AND2x2_ASAP7_75t_L g796 ( .A(n_683), .B(n_786), .Y(n_796) );
AND2x2_ASAP7_75t_L g699 ( .A(n_684), .B(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g764 ( .A(n_684), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_686), .B(n_688), .Y(n_685) );
OR2x2_ASAP7_75t_L g722 ( .A(n_687), .B(n_723), .Y(n_722) );
INVx2_ASAP7_75t_L g701 ( .A(n_688), .Y(n_701) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_691), .B(n_693), .Y(n_690) );
INVx2_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
AND2x4_ASAP7_75t_L g735 ( .A(n_692), .B(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g824 ( .A(n_693), .Y(n_824) );
NOR2xp67_ASAP7_75t_L g696 ( .A(n_697), .B(n_733), .Y(n_696) );
NAND3xp33_ASAP7_75t_SL g697 ( .A(n_698), .B(n_708), .C(n_720), .Y(n_697) );
AOI22xp33_ASAP7_75t_L g698 ( .A1(n_699), .A2(n_701), .B1(n_702), .B2(n_703), .Y(n_698) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_705), .B(n_706), .Y(n_704) );
INVx1_ASAP7_75t_L g741 ( .A(n_706), .Y(n_741) );
AND2x2_ASAP7_75t_L g816 ( .A(n_706), .B(n_727), .Y(n_816) );
INVx1_ASAP7_75t_L g763 ( .A(n_707), .Y(n_763) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
OAI32xp33_ASAP7_75t_L g709 ( .A1(n_710), .A2(n_711), .A3(n_713), .B1(n_715), .B2(n_718), .Y(n_709) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx2_ASAP7_75t_L g743 ( .A(n_712), .Y(n_743) );
NAND2x1_ASAP7_75t_L g781 ( .A(n_712), .B(n_782), .Y(n_781) );
HB1xp67_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
AND2x2_ASAP7_75t_L g742 ( .A(n_714), .B(n_743), .Y(n_742) );
NOR2x1_ASAP7_75t_L g715 ( .A(n_716), .B(n_717), .Y(n_715) );
OAI211xp5_ASAP7_75t_SL g768 ( .A1(n_719), .A2(n_762), .B(n_769), .C(n_770), .Y(n_768) );
INVx2_ASAP7_75t_L g782 ( .A(n_719), .Y(n_782) );
OAI21xp5_ASAP7_75t_L g720 ( .A1(n_721), .A2(n_725), .B(n_732), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
HB1xp67_ASAP7_75t_L g737 ( .A(n_726), .Y(n_737) );
NAND2x1_ASAP7_75t_L g726 ( .A(n_727), .B(n_729), .Y(n_726) );
INVx2_ASAP7_75t_L g820 ( .A(n_727), .Y(n_820) );
INVx3_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
AND2x2_ASAP7_75t_L g828 ( .A(n_728), .B(n_763), .Y(n_828) );
AND2x2_ASAP7_75t_L g833 ( .A(n_728), .B(n_789), .Y(n_833) );
AND2x4_ASAP7_75t_L g729 ( .A(n_730), .B(n_731), .Y(n_729) );
INVx1_ASAP7_75t_L g758 ( .A(n_731), .Y(n_758) );
OAI211xp5_ASAP7_75t_L g733 ( .A1(n_734), .A2(n_737), .B(n_738), .C(n_745), .Y(n_733) );
INVxp67_ASAP7_75t_SL g734 ( .A(n_735), .Y(n_734) );
NAND2x1p5_ASAP7_75t_L g752 ( .A(n_735), .B(n_753), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_746), .B(n_747), .Y(n_745) );
INVx2_ASAP7_75t_SL g747 ( .A(n_748), .Y(n_747) );
NOR3xp33_ASAP7_75t_L g750 ( .A(n_751), .B(n_783), .C(n_812), .Y(n_750) );
OAI211xp5_ASAP7_75t_L g751 ( .A1(n_752), .A2(n_756), .B(n_759), .C(n_771), .Y(n_751) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
AOI22xp5_ASAP7_75t_L g795 ( .A1(n_757), .A2(n_796), .B1(n_797), .B2(n_800), .Y(n_795) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
AOI22xp5_ASAP7_75t_L g759 ( .A1(n_760), .A2(n_761), .B1(n_767), .B2(n_768), .Y(n_759) );
OAI22xp33_ASAP7_75t_L g761 ( .A1(n_762), .A2(n_764), .B1(n_765), .B2(n_766), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g805 ( .A(n_762), .B(n_794), .Y(n_805) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
AND2x2_ASAP7_75t_L g776 ( .A(n_769), .B(n_777), .Y(n_776) );
AOI22xp5_ASAP7_75t_L g771 ( .A1(n_772), .A2(n_776), .B1(n_778), .B2(n_780), .Y(n_771) );
INVx1_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
INVx1_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
OR2x2_ASAP7_75t_L g801 ( .A(n_775), .B(n_802), .Y(n_801) );
INVx2_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
INVx1_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
OAI211xp5_ASAP7_75t_SL g783 ( .A1(n_784), .A2(n_790), .B(n_795), .C(n_803), .Y(n_783) );
INVx2_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
AND2x2_ASAP7_75t_L g785 ( .A(n_786), .B(n_787), .Y(n_785) );
INVx1_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
NOR2xp33_ASAP7_75t_L g790 ( .A(n_791), .B(n_792), .Y(n_790) );
INVx2_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
INVx1_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
INVx2_ASAP7_75t_SL g800 ( .A(n_801), .Y(n_800) );
AOI22xp5_ASAP7_75t_L g803 ( .A1(n_804), .A2(n_806), .B1(n_807), .B2(n_809), .Y(n_803) );
INVx1_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
INVx1_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
OAI211xp5_ASAP7_75t_SL g812 ( .A1(n_813), .A2(n_815), .B(n_817), .C(n_825), .Y(n_812) );
INVxp67_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
NAND2xp5_ASAP7_75t_L g817 ( .A(n_818), .B(n_821), .Y(n_817) );
INVx1_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
INVx1_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
OR2x2_ASAP7_75t_L g822 ( .A(n_823), .B(n_824), .Y(n_822) );
INVx4_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
INVx1_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
INVx4_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
AND2x6_ASAP7_75t_SL g839 ( .A(n_840), .B(n_842), .Y(n_839) );
BUFx3_ASAP7_75t_L g848 ( .A(n_840), .Y(n_848) );
INVx1_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
NOR2xp33_ASAP7_75t_L g864 ( .A(n_841), .B(n_865), .Y(n_864) );
NAND2xp5_ASAP7_75t_L g842 ( .A(n_843), .B(n_845), .Y(n_842) );
INVx1_ASAP7_75t_L g843 ( .A(n_844), .Y(n_843) );
NOR2x1_ASAP7_75t_L g867 ( .A(n_844), .B(n_846), .Y(n_867) );
AND2x6_ASAP7_75t_SL g857 ( .A(n_845), .B(n_858), .Y(n_857) );
INVx1_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
OAI21xp5_ASAP7_75t_L g847 ( .A1(n_848), .A2(n_849), .B(n_860), .Y(n_847) );
NAND2xp5_ASAP7_75t_L g849 ( .A(n_850), .B(n_854), .Y(n_849) );
INVx3_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
INVx3_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
CKINVDCx8_ASAP7_75t_R g856 ( .A(n_857), .Y(n_856) );
CKINVDCx5p33_ASAP7_75t_R g869 ( .A(n_857), .Y(n_869) );
INVx3_ASAP7_75t_L g861 ( .A(n_862), .Y(n_861) );
INVx6_ASAP7_75t_L g862 ( .A(n_863), .Y(n_862) );
BUFx10_ASAP7_75t_L g863 ( .A(n_864), .Y(n_863) );
INVx1_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
NOR2xp33_ASAP7_75t_L g868 ( .A(n_869), .B(n_870), .Y(n_868) );
endmodule