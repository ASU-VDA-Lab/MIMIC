module fake_netlist_1_7169_n_717 (n_44, n_81, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_717);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_717;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_560;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_415;
wire n_235;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_363;
wire n_409;
wire n_315;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_498;
wire n_349;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_494;
wire n_223;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g82 ( .A(n_12), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_21), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_78), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_25), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_61), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_69), .Y(n_87) );
INVxp67_ASAP7_75t_L g88 ( .A(n_8), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_41), .Y(n_89) );
CKINVDCx20_ASAP7_75t_R g90 ( .A(n_19), .Y(n_90) );
CKINVDCx5p33_ASAP7_75t_R g91 ( .A(n_11), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_70), .Y(n_92) );
CKINVDCx14_ASAP7_75t_R g93 ( .A(n_31), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_21), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_46), .Y(n_95) );
INVxp33_ASAP7_75t_SL g96 ( .A(n_6), .Y(n_96) );
CKINVDCx5p33_ASAP7_75t_R g97 ( .A(n_77), .Y(n_97) );
CKINVDCx5p33_ASAP7_75t_R g98 ( .A(n_8), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_81), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_15), .Y(n_100) );
INVxp33_ASAP7_75t_SL g101 ( .A(n_22), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_74), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_51), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_11), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_45), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_66), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_19), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_24), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_35), .Y(n_109) );
INVxp67_ASAP7_75t_SL g110 ( .A(n_43), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_73), .Y(n_111) );
INVxp33_ASAP7_75t_SL g112 ( .A(n_16), .Y(n_112) );
NOR2xp33_ASAP7_75t_L g113 ( .A(n_63), .B(n_57), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_14), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_20), .Y(n_115) );
BUFx6f_ASAP7_75t_L g116 ( .A(n_13), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_56), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_18), .Y(n_118) );
HB1xp67_ASAP7_75t_L g119 ( .A(n_29), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_55), .Y(n_120) );
INVxp67_ASAP7_75t_SL g121 ( .A(n_4), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_28), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_27), .Y(n_123) );
BUFx3_ASAP7_75t_L g124 ( .A(n_12), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_17), .Y(n_125) );
INVxp67_ASAP7_75t_L g126 ( .A(n_10), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_44), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_59), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_52), .Y(n_129) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_60), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_39), .Y(n_131) );
AND2x2_ASAP7_75t_L g132 ( .A(n_119), .B(n_0), .Y(n_132) );
INVx1_ASAP7_75t_SL g133 ( .A(n_91), .Y(n_133) );
AND2x2_ASAP7_75t_L g134 ( .A(n_93), .B(n_0), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_130), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_130), .Y(n_136) );
AND2x2_ASAP7_75t_L g137 ( .A(n_124), .B(n_1), .Y(n_137) );
INVxp67_ASAP7_75t_L g138 ( .A(n_124), .Y(n_138) );
AND2x2_ASAP7_75t_L g139 ( .A(n_82), .B(n_1), .Y(n_139) );
NAND2xp5_ASAP7_75t_SL g140 ( .A(n_130), .B(n_2), .Y(n_140) );
INVx6_ASAP7_75t_L g141 ( .A(n_130), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_89), .Y(n_142) );
BUFx2_ASAP7_75t_L g143 ( .A(n_91), .Y(n_143) );
INVx3_ASAP7_75t_L g144 ( .A(n_116), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_130), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_82), .B(n_2), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_131), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_89), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_92), .Y(n_149) );
NAND2x1_ASAP7_75t_L g150 ( .A(n_83), .B(n_3), .Y(n_150) );
AND2x2_ASAP7_75t_L g151 ( .A(n_83), .B(n_3), .Y(n_151) );
INVx3_ASAP7_75t_L g152 ( .A(n_116), .Y(n_152) );
CKINVDCx8_ASAP7_75t_R g153 ( .A(n_97), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_131), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_92), .Y(n_155) );
INVx1_ASAP7_75t_SL g156 ( .A(n_98), .Y(n_156) );
AND2x4_ASAP7_75t_L g157 ( .A(n_94), .B(n_4), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_94), .B(n_5), .Y(n_158) );
HB1xp67_ASAP7_75t_L g159 ( .A(n_98), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_95), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_107), .B(n_5), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_95), .Y(n_162) );
INVx5_ASAP7_75t_L g163 ( .A(n_116), .Y(n_163) );
INVx1_ASAP7_75t_SL g164 ( .A(n_125), .Y(n_164) );
CKINVDCx5p33_ASAP7_75t_R g165 ( .A(n_97), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_99), .Y(n_166) );
AND2x6_ASAP7_75t_L g167 ( .A(n_99), .B(n_40), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_127), .Y(n_168) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_116), .Y(n_169) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_116), .Y(n_170) );
AND2x4_ASAP7_75t_L g171 ( .A(n_107), .B(n_6), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_127), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_84), .Y(n_173) );
BUFx8_ASAP7_75t_L g174 ( .A(n_85), .Y(n_174) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_86), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_87), .Y(n_176) );
INVx3_ASAP7_75t_L g177 ( .A(n_157), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_175), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_163), .Y(n_179) );
BUFx2_ASAP7_75t_L g180 ( .A(n_143), .Y(n_180) );
INVx1_ASAP7_75t_SL g181 ( .A(n_143), .Y(n_181) );
BUFx6f_ASAP7_75t_L g182 ( .A(n_169), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_163), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_163), .Y(n_184) );
INVx1_ASAP7_75t_SL g185 ( .A(n_133), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_175), .Y(n_186) );
AND2x4_ASAP7_75t_L g187 ( .A(n_157), .B(n_100), .Y(n_187) );
INVx1_ASAP7_75t_SL g188 ( .A(n_133), .Y(n_188) );
INVx3_ASAP7_75t_L g189 ( .A(n_157), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_175), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g191 ( .A(n_165), .B(n_101), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_175), .Y(n_192) );
BUFx3_ASAP7_75t_L g193 ( .A(n_167), .Y(n_193) );
BUFx6f_ASAP7_75t_L g194 ( .A(n_169), .Y(n_194) );
INVx3_ASAP7_75t_L g195 ( .A(n_157), .Y(n_195) );
AND2x2_ASAP7_75t_L g196 ( .A(n_138), .B(n_125), .Y(n_196) );
BUFx6f_ASAP7_75t_L g197 ( .A(n_169), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_169), .Y(n_198) );
BUFx3_ASAP7_75t_L g199 ( .A(n_167), .Y(n_199) );
INVx2_ASAP7_75t_L g200 ( .A(n_169), .Y(n_200) );
INVx3_ASAP7_75t_L g201 ( .A(n_171), .Y(n_201) );
AND2x6_ASAP7_75t_L g202 ( .A(n_171), .B(n_102), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_175), .Y(n_203) );
AND2x4_ASAP7_75t_L g204 ( .A(n_171), .B(n_114), .Y(n_204) );
AOI22xp5_ASAP7_75t_L g205 ( .A1(n_171), .A2(n_112), .B1(n_96), .B2(n_121), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_169), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_175), .Y(n_207) );
A2O1A1Ixp33_ASAP7_75t_L g208 ( .A1(n_142), .A2(n_111), .B(n_109), .C(n_105), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_155), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_163), .Y(n_210) );
INVx1_ASAP7_75t_SL g211 ( .A(n_156), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g212 ( .A(n_138), .B(n_120), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_170), .Y(n_213) );
CKINVDCx16_ASAP7_75t_R g214 ( .A(n_159), .Y(n_214) );
BUFx6f_ASAP7_75t_L g215 ( .A(n_170), .Y(n_215) );
NOR2xp33_ASAP7_75t_SL g216 ( .A(n_153), .B(n_129), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_170), .Y(n_217) );
BUFx2_ASAP7_75t_L g218 ( .A(n_134), .Y(n_218) );
BUFx6f_ASAP7_75t_L g219 ( .A(n_170), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g220 ( .A(n_173), .B(n_122), .Y(n_220) );
AND2x2_ASAP7_75t_L g221 ( .A(n_156), .B(n_164), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_155), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_163), .Y(n_223) );
INVx4_ASAP7_75t_L g224 ( .A(n_167), .Y(n_224) );
AND2x6_ASAP7_75t_L g225 ( .A(n_137), .B(n_123), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_163), .Y(n_226) );
INVx4_ASAP7_75t_L g227 ( .A(n_167), .Y(n_227) );
NOR2xp33_ASAP7_75t_SL g228 ( .A(n_153), .B(n_129), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_155), .Y(n_229) );
BUFx10_ASAP7_75t_L g230 ( .A(n_167), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_162), .Y(n_231) );
INVx3_ASAP7_75t_L g232 ( .A(n_147), .Y(n_232) );
AO22x1_ASAP7_75t_L g233 ( .A1(n_167), .A2(n_110), .B1(n_117), .B2(n_118), .Y(n_233) );
INVx2_ASAP7_75t_L g234 ( .A(n_170), .Y(n_234) );
BUFx6f_ASAP7_75t_L g235 ( .A(n_170), .Y(n_235) );
INVxp67_ASAP7_75t_SL g236 ( .A(n_134), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_163), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_173), .B(n_128), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_162), .Y(n_239) );
OR2x2_ASAP7_75t_L g240 ( .A(n_164), .B(n_88), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_176), .B(n_108), .Y(n_241) );
BUFx3_ASAP7_75t_L g242 ( .A(n_167), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_162), .Y(n_243) );
NAND2xp5_ASAP7_75t_SL g244 ( .A(n_224), .B(n_174), .Y(n_244) );
INVx2_ASAP7_75t_L g245 ( .A(n_209), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_241), .B(n_132), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_209), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_222), .Y(n_248) );
BUFx2_ASAP7_75t_L g249 ( .A(n_181), .Y(n_249) );
NOR2xp33_ASAP7_75t_R g250 ( .A(n_214), .B(n_153), .Y(n_250) );
NAND2xp5_ASAP7_75t_SL g251 ( .A(n_224), .B(n_174), .Y(n_251) );
INVx2_ASAP7_75t_L g252 ( .A(n_222), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_229), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_229), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_238), .B(n_132), .Y(n_255) );
OR2x6_ASAP7_75t_L g256 ( .A(n_180), .B(n_150), .Y(n_256) );
CKINVDCx5p33_ASAP7_75t_R g257 ( .A(n_214), .Y(n_257) );
INVxp67_ASAP7_75t_SL g258 ( .A(n_180), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_196), .B(n_174), .Y(n_259) );
CKINVDCx5p33_ASAP7_75t_R g260 ( .A(n_185), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_231), .Y(n_261) );
BUFx6f_ASAP7_75t_L g262 ( .A(n_230), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_231), .Y(n_263) );
INVx1_ASAP7_75t_SL g264 ( .A(n_188), .Y(n_264) );
INVx3_ASAP7_75t_L g265 ( .A(n_232), .Y(n_265) );
AOI22xp33_ASAP7_75t_L g266 ( .A1(n_202), .A2(n_142), .B1(n_148), .B2(n_160), .Y(n_266) );
AND2x4_ASAP7_75t_L g267 ( .A(n_236), .B(n_139), .Y(n_267) );
INVx4_ASAP7_75t_L g268 ( .A(n_202), .Y(n_268) );
AO22x1_ASAP7_75t_L g269 ( .A1(n_211), .A2(n_174), .B1(n_167), .B2(n_103), .Y(n_269) );
INVx2_ASAP7_75t_L g270 ( .A(n_239), .Y(n_270) );
INVx1_ASAP7_75t_SL g271 ( .A(n_221), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_196), .B(n_148), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_239), .Y(n_273) );
INVx2_ASAP7_75t_L g274 ( .A(n_243), .Y(n_274) );
AOI22xp33_ASAP7_75t_L g275 ( .A1(n_202), .A2(n_168), .B1(n_160), .B2(n_149), .Y(n_275) );
OR2x2_ASAP7_75t_L g276 ( .A(n_240), .B(n_146), .Y(n_276) );
OR2x2_ASAP7_75t_L g277 ( .A(n_240), .B(n_146), .Y(n_277) );
NOR2xp33_ASAP7_75t_L g278 ( .A(n_187), .B(n_176), .Y(n_278) );
HB1xp67_ASAP7_75t_L g279 ( .A(n_221), .Y(n_279) );
A2O1A1Ixp33_ASAP7_75t_L g280 ( .A1(n_177), .A2(n_189), .B(n_195), .C(n_201), .Y(n_280) );
AND2x6_ASAP7_75t_L g281 ( .A(n_193), .B(n_137), .Y(n_281) );
INVx5_ASAP7_75t_L g282 ( .A(n_202), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_218), .B(n_149), .Y(n_283) );
AND2x4_ASAP7_75t_L g284 ( .A(n_187), .B(n_139), .Y(n_284) );
AOI22xp5_ASAP7_75t_L g285 ( .A1(n_205), .A2(n_151), .B1(n_150), .B2(n_168), .Y(n_285) );
AND2x2_ASAP7_75t_L g286 ( .A(n_218), .B(n_151), .Y(n_286) );
INVx4_ASAP7_75t_L g287 ( .A(n_202), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_187), .B(n_172), .Y(n_288) );
BUFx8_ASAP7_75t_L g289 ( .A(n_225), .Y(n_289) );
NOR2xp33_ASAP7_75t_L g290 ( .A(n_187), .B(n_161), .Y(n_290) );
CKINVDCx20_ASAP7_75t_R g291 ( .A(n_205), .Y(n_291) );
INVx3_ASAP7_75t_L g292 ( .A(n_232), .Y(n_292) );
BUFx4f_ASAP7_75t_L g293 ( .A(n_225), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_204), .B(n_172), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_243), .Y(n_295) );
INVx2_ASAP7_75t_SL g296 ( .A(n_204), .Y(n_296) );
AOI22xp33_ASAP7_75t_L g297 ( .A1(n_202), .A2(n_172), .B1(n_166), .B2(n_154), .Y(n_297) );
BUFx2_ASAP7_75t_L g298 ( .A(n_225), .Y(n_298) );
AOI22x1_ASAP7_75t_L g299 ( .A1(n_224), .A2(n_166), .B1(n_147), .B2(n_154), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_232), .Y(n_300) );
NAND2xp5_ASAP7_75t_SL g301 ( .A(n_224), .B(n_166), .Y(n_301) );
INVx2_ASAP7_75t_SL g302 ( .A(n_204), .Y(n_302) );
BUFx12f_ASAP7_75t_L g303 ( .A(n_204), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_212), .B(n_161), .Y(n_304) );
AND2x4_ASAP7_75t_L g305 ( .A(n_202), .B(n_158), .Y(n_305) );
AOI22xp5_ASAP7_75t_L g306 ( .A1(n_225), .A2(n_126), .B1(n_158), .B2(n_140), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_225), .B(n_128), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_225), .B(n_108), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_178), .Y(n_309) );
INVx4_ASAP7_75t_L g310 ( .A(n_225), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_232), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_177), .B(n_106), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_177), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_177), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_178), .Y(n_315) );
CKINVDCx5p33_ASAP7_75t_R g316 ( .A(n_250), .Y(n_316) );
INVx3_ASAP7_75t_L g317 ( .A(n_310), .Y(n_317) );
AND2x2_ASAP7_75t_L g318 ( .A(n_264), .B(n_191), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_276), .B(n_277), .Y(n_319) );
OAI21xp5_ASAP7_75t_L g320 ( .A1(n_280), .A2(n_227), .B(n_189), .Y(n_320) );
BUFx3_ASAP7_75t_L g321 ( .A(n_289), .Y(n_321) );
A2O1A1Ixp33_ASAP7_75t_L g322 ( .A1(n_280), .A2(n_201), .B(n_195), .C(n_189), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_245), .Y(n_323) );
BUFx6f_ASAP7_75t_L g324 ( .A(n_268), .Y(n_324) );
BUFx6f_ASAP7_75t_L g325 ( .A(n_268), .Y(n_325) );
OAI22xp5_ASAP7_75t_L g326 ( .A1(n_271), .A2(n_189), .B1(n_195), .B2(n_201), .Y(n_326) );
O2A1O1Ixp33_ASAP7_75t_L g327 ( .A1(n_279), .A2(n_208), .B(n_201), .C(n_195), .Y(n_327) );
AND2x4_ASAP7_75t_L g328 ( .A(n_310), .B(n_227), .Y(n_328) );
BUFx2_ASAP7_75t_L g329 ( .A(n_249), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_288), .Y(n_330) );
OR2x2_ASAP7_75t_L g331 ( .A(n_260), .B(n_220), .Y(n_331) );
NOR2x1_ASAP7_75t_R g332 ( .A(n_260), .B(n_103), .Y(n_332) );
INVx3_ASAP7_75t_SL g333 ( .A(n_257), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_258), .B(n_216), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_245), .Y(n_335) );
BUFx2_ASAP7_75t_R g336 ( .A(n_257), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_294), .Y(n_337) );
BUFx6f_ASAP7_75t_L g338 ( .A(n_287), .Y(n_338) );
INVxp67_ASAP7_75t_L g339 ( .A(n_296), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_247), .Y(n_340) );
OAI221xp5_ASAP7_75t_L g341 ( .A1(n_285), .A2(n_228), .B1(n_104), .B2(n_115), .C(n_227), .Y(n_341) );
BUFx6f_ASAP7_75t_L g342 ( .A(n_287), .Y(n_342) );
BUFx12f_ASAP7_75t_L g343 ( .A(n_303), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_284), .B(n_233), .Y(n_344) );
AND2x4_ASAP7_75t_L g345 ( .A(n_267), .B(n_227), .Y(n_345) );
HAxp5_ASAP7_75t_L g346 ( .A(n_291), .B(n_90), .CON(n_346), .SN(n_346) );
INVx3_ASAP7_75t_L g347 ( .A(n_289), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_284), .B(n_233), .Y(n_348) );
BUFx6f_ASAP7_75t_L g349 ( .A(n_282), .Y(n_349) );
OR2x2_ASAP7_75t_L g350 ( .A(n_256), .B(n_147), .Y(n_350) );
AOI22xp5_ASAP7_75t_L g351 ( .A1(n_303), .A2(n_193), .B1(n_199), .B2(n_242), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_247), .Y(n_352) );
AOI22xp33_ASAP7_75t_L g353 ( .A1(n_290), .A2(n_242), .B1(n_193), .B2(n_199), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_252), .Y(n_354) );
BUFx6f_ASAP7_75t_L g355 ( .A(n_282), .Y(n_355) );
AOI22xp33_ASAP7_75t_L g356 ( .A1(n_290), .A2(n_242), .B1(n_199), .B2(n_154), .Y(n_356) );
BUFx12f_ASAP7_75t_L g357 ( .A(n_289), .Y(n_357) );
BUFx2_ASAP7_75t_L g358 ( .A(n_250), .Y(n_358) );
BUFx6f_ASAP7_75t_L g359 ( .A(n_282), .Y(n_359) );
AND2x4_ASAP7_75t_L g360 ( .A(n_284), .B(n_106), .Y(n_360) );
AO22x1_ASAP7_75t_L g361 ( .A1(n_281), .A2(n_113), .B1(n_9), .B2(n_10), .Y(n_361) );
A2O1A1Ixp33_ASAP7_75t_L g362 ( .A1(n_278), .A2(n_272), .B(n_304), .C(n_261), .Y(n_362) );
OR2x6_ASAP7_75t_L g363 ( .A(n_298), .B(n_237), .Y(n_363) );
INVx5_ASAP7_75t_L g364 ( .A(n_281), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_252), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_254), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_254), .Y(n_367) );
AOI22xp33_ASAP7_75t_L g368 ( .A1(n_305), .A2(n_230), .B1(n_152), .B2(n_144), .Y(n_368) );
INVx3_ASAP7_75t_L g369 ( .A(n_270), .Y(n_369) );
INVx3_ASAP7_75t_L g370 ( .A(n_270), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_267), .B(n_230), .Y(n_371) );
AOI22xp5_ASAP7_75t_L g372 ( .A1(n_305), .A2(n_230), .B1(n_190), .B2(n_203), .Y(n_372) );
OAI22xp33_ASAP7_75t_L g373 ( .A1(n_329), .A2(n_291), .B1(n_293), .B2(n_256), .Y(n_373) );
OAI22xp5_ASAP7_75t_L g374 ( .A1(n_362), .A2(n_266), .B1(n_275), .B2(n_293), .Y(n_374) );
O2A1O1Ixp33_ASAP7_75t_L g375 ( .A1(n_362), .A2(n_283), .B(n_255), .C(n_246), .Y(n_375) );
AND2x4_ASAP7_75t_L g376 ( .A(n_347), .B(n_282), .Y(n_376) );
AOI21xp33_ASAP7_75t_L g377 ( .A1(n_327), .A2(n_259), .B(n_299), .Y(n_377) );
AND2x4_ASAP7_75t_L g378 ( .A(n_347), .B(n_302), .Y(n_378) );
AOI22xp33_ASAP7_75t_L g379 ( .A1(n_319), .A2(n_305), .B1(n_256), .B2(n_267), .Y(n_379) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_343), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_323), .Y(n_381) );
AOI21xp5_ASAP7_75t_L g382 ( .A1(n_322), .A2(n_301), .B(n_244), .Y(n_382) );
INVx3_ASAP7_75t_L g383 ( .A(n_324), .Y(n_383) );
OAI21xp33_ASAP7_75t_SL g384 ( .A1(n_340), .A2(n_275), .B(n_266), .Y(n_384) );
BUFx2_ASAP7_75t_L g385 ( .A(n_343), .Y(n_385) );
INVxp67_ASAP7_75t_L g386 ( .A(n_332), .Y(n_386) );
OAI22xp33_ASAP7_75t_L g387 ( .A1(n_333), .A2(n_306), .B1(n_312), .B2(n_307), .Y(n_387) );
BUFx3_ASAP7_75t_L g388 ( .A(n_324), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_323), .Y(n_389) );
AOI22xp33_ASAP7_75t_SL g390 ( .A1(n_360), .A2(n_286), .B1(n_281), .B2(n_278), .Y(n_390) );
NAND3x1_ASAP7_75t_L g391 ( .A(n_334), .B(n_308), .C(n_248), .Y(n_391) );
AOI22xp33_ASAP7_75t_L g392 ( .A1(n_360), .A2(n_281), .B1(n_314), .B2(n_313), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_335), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_335), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_330), .B(n_274), .Y(n_395) );
AOI22xp33_ASAP7_75t_L g396 ( .A1(n_360), .A2(n_281), .B1(n_251), .B2(n_244), .Y(n_396) );
O2A1O1Ixp33_ASAP7_75t_SL g397 ( .A1(n_322), .A2(n_251), .B(n_263), .C(n_273), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_365), .Y(n_398) );
AND2x4_ASAP7_75t_L g399 ( .A(n_321), .B(n_274), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_365), .Y(n_400) );
A2O1A1Ixp33_ASAP7_75t_L g401 ( .A1(n_320), .A2(n_253), .B(n_295), .C(n_297), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_337), .B(n_297), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_352), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_354), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_369), .Y(n_405) );
INVx3_ASAP7_75t_L g406 ( .A(n_324), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_369), .Y(n_407) );
AOI21xp5_ASAP7_75t_L g408 ( .A1(n_397), .A2(n_269), .B(n_367), .Y(n_408) );
AOI22xp33_ASAP7_75t_L g409 ( .A1(n_390), .A2(n_331), .B1(n_341), .B2(n_318), .Y(n_409) );
AOI22xp33_ASAP7_75t_SL g410 ( .A1(n_374), .A2(n_357), .B1(n_358), .B2(n_316), .Y(n_410) );
AOI22xp33_ASAP7_75t_SL g411 ( .A1(n_374), .A2(n_357), .B1(n_316), .B2(n_321), .Y(n_411) );
AOI22xp33_ASAP7_75t_L g412 ( .A1(n_373), .A2(n_333), .B1(n_345), .B2(n_350), .Y(n_412) );
OAI22xp5_ASAP7_75t_SL g413 ( .A1(n_379), .A2(n_346), .B1(n_364), .B2(n_336), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_389), .Y(n_414) );
NOR2x1_ASAP7_75t_L g415 ( .A(n_387), .B(n_366), .Y(n_415) );
OAI22xp5_ASAP7_75t_L g416 ( .A1(n_375), .A2(n_364), .B1(n_370), .B2(n_348), .Y(n_416) );
BUFx3_ASAP7_75t_L g417 ( .A(n_388), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_395), .B(n_370), .Y(n_418) );
AOI21xp5_ASAP7_75t_L g419 ( .A1(n_375), .A2(n_344), .B(n_326), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_395), .B(n_345), .Y(n_420) );
AOI221xp5_ASAP7_75t_L g421 ( .A1(n_384), .A2(n_361), .B1(n_339), .B2(n_346), .C(n_356), .Y(n_421) );
OR2x2_ASAP7_75t_L g422 ( .A(n_403), .B(n_363), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_389), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_381), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_389), .Y(n_425) );
AOI22xp33_ASAP7_75t_L g426 ( .A1(n_399), .A2(n_364), .B1(n_339), .B2(n_363), .Y(n_426) );
NOR2x1_ASAP7_75t_L g427 ( .A(n_381), .B(n_363), .Y(n_427) );
AND2x4_ASAP7_75t_L g428 ( .A(n_403), .B(n_364), .Y(n_428) );
AOI22xp33_ASAP7_75t_L g429 ( .A1(n_399), .A2(n_265), .B1(n_292), .B2(n_317), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_394), .B(n_265), .Y(n_430) );
INVx1_ASAP7_75t_SL g431 ( .A(n_399), .Y(n_431) );
NAND2xp5_ASAP7_75t_SL g432 ( .A(n_399), .B(n_324), .Y(n_432) );
OAI222xp33_ASAP7_75t_L g433 ( .A1(n_396), .A2(n_356), .B1(n_368), .B2(n_292), .C1(n_300), .C2(n_311), .Y(n_433) );
AO31x2_ASAP7_75t_L g434 ( .A1(n_401), .A2(n_135), .A3(n_136), .B(n_145), .Y(n_434) );
AOI22xp33_ASAP7_75t_L g435 ( .A1(n_402), .A2(n_317), .B1(n_371), .B2(n_368), .Y(n_435) );
AOI21xp5_ASAP7_75t_L g436 ( .A1(n_377), .A2(n_301), .B(n_353), .Y(n_436) );
AOI22xp33_ASAP7_75t_L g437 ( .A1(n_402), .A2(n_328), .B1(n_325), .B2(n_342), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_424), .B(n_394), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_424), .B(n_398), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_414), .Y(n_440) );
NAND4xp25_ASAP7_75t_L g441 ( .A(n_409), .B(n_386), .C(n_385), .D(n_392), .Y(n_441) );
INVxp67_ASAP7_75t_L g442 ( .A(n_418), .Y(n_442) );
OAI221xp5_ASAP7_75t_L g443 ( .A1(n_421), .A2(n_384), .B1(n_385), .B2(n_377), .C(n_380), .Y(n_443) );
OAI21xp5_ASAP7_75t_SL g444 ( .A1(n_411), .A2(n_376), .B(n_378), .Y(n_444) );
OAI22xp5_ASAP7_75t_L g445 ( .A1(n_421), .A2(n_404), .B1(n_391), .B2(n_400), .Y(n_445) );
NAND3xp33_ASAP7_75t_L g446 ( .A(n_410), .B(n_382), .C(n_400), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_414), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_418), .B(n_398), .Y(n_448) );
OAI211xp5_ASAP7_75t_SL g449 ( .A1(n_412), .A2(n_144), .B(n_152), .C(n_404), .Y(n_449) );
NAND4xp25_ASAP7_75t_SL g450 ( .A(n_413), .B(n_382), .C(n_393), .D(n_391), .Y(n_450) );
AOI221xp5_ASAP7_75t_L g451 ( .A1(n_413), .A2(n_378), .B1(n_393), .B2(n_407), .C(n_405), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_414), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_423), .B(n_393), .Y(n_453) );
OR2x2_ASAP7_75t_L g454 ( .A(n_431), .B(n_405), .Y(n_454) );
INVx3_ASAP7_75t_L g455 ( .A(n_428), .Y(n_455) );
OAI211xp5_ASAP7_75t_L g456 ( .A1(n_426), .A2(n_144), .B(n_152), .C(n_136), .Y(n_456) );
AOI22xp5_ASAP7_75t_L g457 ( .A1(n_420), .A2(n_378), .B1(n_391), .B2(n_405), .Y(n_457) );
OAI31xp33_ASAP7_75t_L g458 ( .A1(n_433), .A2(n_378), .A3(n_376), .B(n_388), .Y(n_458) );
NOR2x1_ASAP7_75t_L g459 ( .A(n_427), .B(n_388), .Y(n_459) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_415), .A2(n_376), .B1(n_407), .B2(n_383), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_423), .B(n_407), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_420), .B(n_376), .Y(n_462) );
AOI22xp33_ASAP7_75t_L g463 ( .A1(n_415), .A2(n_406), .B1(n_383), .B2(n_325), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_423), .Y(n_464) );
OAI22xp5_ASAP7_75t_L g465 ( .A1(n_422), .A2(n_406), .B1(n_383), .B2(n_353), .Y(n_465) );
AOI222xp33_ASAP7_75t_L g466 ( .A1(n_416), .A2(n_144), .B1(n_152), .B2(n_406), .C1(n_383), .C2(n_145), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_425), .B(n_406), .Y(n_467) );
AOI31xp33_ASAP7_75t_L g468 ( .A1(n_427), .A2(n_7), .A3(n_9), .B(n_13), .Y(n_468) );
AOI22xp33_ASAP7_75t_SL g469 ( .A1(n_428), .A2(n_338), .B1(n_342), .B2(n_325), .Y(n_469) );
OAI332xp33_ASAP7_75t_L g470 ( .A1(n_422), .A2(n_135), .A3(n_136), .B1(n_145), .B2(n_207), .B3(n_203), .C1(n_186), .C2(n_190), .Y(n_470) );
NAND4xp25_ASAP7_75t_L g471 ( .A(n_419), .B(n_135), .C(n_207), .D(n_192), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_425), .Y(n_472) );
NAND3xp33_ASAP7_75t_L g473 ( .A(n_416), .B(n_192), .C(n_186), .Y(n_473) );
AOI211xp5_ASAP7_75t_SL g474 ( .A1(n_428), .A2(n_351), .B(n_328), .C(n_372), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_438), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_440), .Y(n_476) );
OAI22xp5_ASAP7_75t_L g477 ( .A1(n_468), .A2(n_431), .B1(n_437), .B2(n_435), .Y(n_477) );
OR2x2_ASAP7_75t_L g478 ( .A(n_440), .B(n_425), .Y(n_478) );
AND2x2_ASAP7_75t_SL g479 ( .A(n_457), .B(n_428), .Y(n_479) );
AOI22xp5_ASAP7_75t_L g480 ( .A1(n_441), .A2(n_429), .B1(n_430), .B2(n_432), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_447), .Y(n_481) );
AND2x4_ASAP7_75t_L g482 ( .A(n_455), .B(n_417), .Y(n_482) );
BUFx3_ASAP7_75t_L g483 ( .A(n_453), .Y(n_483) );
OR2x2_ASAP7_75t_L g484 ( .A(n_452), .B(n_434), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_448), .B(n_434), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_452), .Y(n_486) );
NAND3xp33_ASAP7_75t_L g487 ( .A(n_443), .B(n_436), .C(n_408), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_464), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_448), .B(n_434), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_464), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_472), .Y(n_491) );
INVx3_ASAP7_75t_L g492 ( .A(n_472), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_438), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_439), .B(n_430), .Y(n_494) );
OAI33xp33_ASAP7_75t_L g495 ( .A1(n_445), .A2(n_7), .A3(n_14), .B1(n_15), .B2(n_16), .B3(n_17), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_439), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_453), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_461), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_461), .B(n_434), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_467), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_467), .Y(n_501) );
OAI22xp33_ASAP7_75t_L g502 ( .A1(n_444), .A2(n_417), .B1(n_325), .B2(n_338), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_442), .B(n_417), .Y(n_503) );
OAI211xp5_ASAP7_75t_SL g504 ( .A1(n_458), .A2(n_217), .B(n_198), .C(n_200), .Y(n_504) );
AOI22xp33_ASAP7_75t_L g505 ( .A1(n_449), .A2(n_141), .B1(n_342), .B2(n_338), .Y(n_505) );
INVx2_ASAP7_75t_L g506 ( .A(n_454), .Y(n_506) );
OAI211xp5_ASAP7_75t_SL g507 ( .A1(n_451), .A2(n_217), .B(n_198), .C(n_200), .Y(n_507) );
OAI33xp33_ASAP7_75t_L g508 ( .A1(n_465), .A2(n_18), .A3(n_20), .B1(n_234), .B2(n_217), .B3(n_213), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_462), .Y(n_509) );
OAI221xp5_ASAP7_75t_L g510 ( .A1(n_446), .A2(n_141), .B1(n_234), .B2(n_213), .C(n_206), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_454), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_455), .B(n_434), .Y(n_512) );
OAI221xp5_ASAP7_75t_SL g513 ( .A1(n_457), .A2(n_434), .B1(n_234), .B2(n_213), .C(n_206), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_455), .B(n_23), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_460), .B(n_26), .Y(n_515) );
BUFx3_ASAP7_75t_L g516 ( .A(n_446), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_459), .B(n_30), .Y(n_517) );
OAI211xp5_ASAP7_75t_SL g518 ( .A1(n_474), .A2(n_466), .B(n_463), .C(n_459), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_469), .B(n_32), .Y(n_519) );
NOR2xp67_ASAP7_75t_L g520 ( .A(n_450), .B(n_33), .Y(n_520) );
OAI321xp33_ASAP7_75t_L g521 ( .A1(n_471), .A2(n_198), .A3(n_200), .B1(n_206), .B2(n_182), .C(n_194), .Y(n_521) );
INVx4_ASAP7_75t_L g522 ( .A(n_470), .Y(n_522) );
OR2x2_ASAP7_75t_L g523 ( .A(n_473), .B(n_34), .Y(n_523) );
AND2x2_ASAP7_75t_SL g524 ( .A(n_456), .B(n_342), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_485), .B(n_141), .Y(n_525) );
NAND3xp33_ASAP7_75t_L g526 ( .A(n_487), .B(n_219), .C(n_194), .Y(n_526) );
INVx1_ASAP7_75t_SL g527 ( .A(n_483), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_485), .B(n_489), .Y(n_528) );
OAI33xp33_ASAP7_75t_L g529 ( .A1(n_477), .A2(n_141), .A3(n_37), .B1(n_38), .B2(n_42), .B3(n_47), .Y(n_529) );
HB1xp67_ASAP7_75t_L g530 ( .A(n_483), .Y(n_530) );
INVxp67_ASAP7_75t_L g531 ( .A(n_478), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_489), .B(n_141), .Y(n_532) );
OR2x6_ASAP7_75t_L g533 ( .A(n_481), .B(n_338), .Y(n_533) );
INVx4_ASAP7_75t_L g534 ( .A(n_524), .Y(n_534) );
INVx2_ASAP7_75t_SL g535 ( .A(n_478), .Y(n_535) );
OR2x2_ASAP7_75t_L g536 ( .A(n_506), .B(n_36), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_475), .B(n_48), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_476), .Y(n_538) );
OR2x2_ASAP7_75t_L g539 ( .A(n_506), .B(n_49), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_476), .Y(n_540) );
HB1xp67_ASAP7_75t_L g541 ( .A(n_481), .Y(n_541) );
NAND3xp33_ASAP7_75t_L g542 ( .A(n_518), .B(n_219), .C(n_194), .Y(n_542) );
NAND2xp5_ASAP7_75t_SL g543 ( .A(n_502), .B(n_524), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_499), .B(n_50), .Y(n_544) );
AOI211xp5_ASAP7_75t_L g545 ( .A1(n_520), .A2(n_235), .B(n_194), .C(n_197), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_499), .B(n_53), .Y(n_546) );
OAI221xp5_ASAP7_75t_L g547 ( .A1(n_522), .A2(n_219), .B1(n_194), .B2(n_197), .C(n_235), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_512), .B(n_54), .Y(n_548) );
OR2x2_ASAP7_75t_L g549 ( .A(n_511), .B(n_58), .Y(n_549) );
NOR2xp67_ASAP7_75t_L g550 ( .A(n_519), .B(n_62), .Y(n_550) );
HB1xp67_ASAP7_75t_L g551 ( .A(n_492), .Y(n_551) );
OAI31xp33_ASAP7_75t_L g552 ( .A1(n_519), .A2(n_328), .A3(n_237), .B(n_67), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_493), .Y(n_553) );
HB1xp67_ASAP7_75t_L g554 ( .A(n_492), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_512), .B(n_64), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_500), .B(n_65), .Y(n_556) );
NAND4xp75_ASAP7_75t_L g557 ( .A(n_479), .B(n_68), .C(n_71), .D(n_72), .Y(n_557) );
NAND3xp33_ASAP7_75t_L g558 ( .A(n_480), .B(n_215), .C(n_235), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_493), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_496), .Y(n_560) );
AOI21xp5_ASAP7_75t_L g561 ( .A1(n_521), .A2(n_359), .B(n_355), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_500), .B(n_75), .Y(n_562) );
HB1xp67_ASAP7_75t_L g563 ( .A(n_492), .Y(n_563) );
NOR3xp33_ASAP7_75t_L g564 ( .A(n_495), .B(n_184), .C(n_226), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_501), .B(n_76), .Y(n_565) );
INVx2_ASAP7_75t_L g566 ( .A(n_486), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_501), .B(n_79), .Y(n_567) );
OR2x2_ASAP7_75t_L g568 ( .A(n_511), .B(n_80), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_509), .B(n_215), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_498), .B(n_197), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_486), .Y(n_571) );
INVx2_ASAP7_75t_L g572 ( .A(n_488), .Y(n_572) );
AOI221xp5_ASAP7_75t_L g573 ( .A1(n_522), .A2(n_197), .B1(n_182), .B2(n_215), .C(n_194), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_498), .B(n_235), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_494), .B(n_497), .Y(n_575) );
INVx1_ASAP7_75t_SL g576 ( .A(n_482), .Y(n_576) );
AOI211xp5_ASAP7_75t_L g577 ( .A1(n_516), .A2(n_235), .B(n_182), .C(n_219), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_497), .B(n_235), .Y(n_578) );
OR2x2_ASAP7_75t_L g579 ( .A(n_488), .B(n_215), .Y(n_579) );
OR2x6_ASAP7_75t_L g580 ( .A(n_516), .B(n_359), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_490), .Y(n_581) );
OAI211xp5_ASAP7_75t_L g582 ( .A1(n_522), .A2(n_359), .B(n_349), .C(n_355), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_490), .B(n_182), .Y(n_583) );
OR2x2_ASAP7_75t_L g584 ( .A(n_535), .B(n_491), .Y(n_584) );
AND2x2_ASAP7_75t_L g585 ( .A(n_527), .B(n_479), .Y(n_585) );
NOR2xp33_ASAP7_75t_L g586 ( .A(n_560), .B(n_508), .Y(n_586) );
AOI211xp5_ASAP7_75t_SL g587 ( .A1(n_582), .A2(n_513), .B(n_523), .C(n_517), .Y(n_587) );
INVxp67_ASAP7_75t_SL g588 ( .A(n_541), .Y(n_588) );
INVx3_ASAP7_75t_L g589 ( .A(n_534), .Y(n_589) );
INVxp67_ASAP7_75t_L g590 ( .A(n_530), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_528), .B(n_503), .Y(n_591) );
NOR2xp33_ASAP7_75t_L g592 ( .A(n_575), .B(n_515), .Y(n_592) );
INVx2_ASAP7_75t_L g593 ( .A(n_566), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_528), .B(n_484), .Y(n_594) );
NAND2xp5_ASAP7_75t_SL g595 ( .A(n_534), .B(n_482), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_538), .Y(n_596) );
OR2x2_ASAP7_75t_L g597 ( .A(n_531), .B(n_484), .Y(n_597) );
INVxp67_ASAP7_75t_L g598 ( .A(n_525), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_553), .B(n_482), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_559), .B(n_517), .Y(n_600) );
OR2x2_ASAP7_75t_L g601 ( .A(n_576), .B(n_523), .Y(n_601) );
INVxp67_ASAP7_75t_L g602 ( .A(n_532), .Y(n_602) );
INVxp67_ASAP7_75t_L g603 ( .A(n_532), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_548), .B(n_514), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_548), .B(n_514), .Y(n_605) );
OAI22xp5_ASAP7_75t_L g606 ( .A1(n_550), .A2(n_505), .B1(n_515), .B2(n_510), .Y(n_606) );
AND2x2_ASAP7_75t_L g607 ( .A(n_555), .B(n_219), .Y(n_607) );
OAI31xp33_ASAP7_75t_L g608 ( .A1(n_543), .A2(n_507), .A3(n_504), .B(n_237), .Y(n_608) );
NAND3xp33_ASAP7_75t_L g609 ( .A(n_542), .B(n_182), .C(n_197), .Y(n_609) );
INVx2_ASAP7_75t_L g610 ( .A(n_572), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_540), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_571), .B(n_215), .Y(n_612) );
OR2x2_ASAP7_75t_L g613 ( .A(n_572), .B(n_197), .Y(n_613) );
NOR2xp33_ASAP7_75t_L g614 ( .A(n_529), .B(n_215), .Y(n_614) );
NAND4xp25_ASAP7_75t_L g615 ( .A(n_552), .B(n_179), .C(n_183), .D(n_210), .Y(n_615) );
NOR2xp67_ASAP7_75t_SL g616 ( .A(n_557), .B(n_359), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_581), .Y(n_617) );
NAND2xp5_ASAP7_75t_SL g618 ( .A(n_534), .B(n_355), .Y(n_618) );
INVxp67_ASAP7_75t_L g619 ( .A(n_551), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_554), .Y(n_620) );
OAI22xp33_ASAP7_75t_L g621 ( .A1(n_536), .A2(n_355), .B1(n_349), .B2(n_179), .Y(n_621) );
AOI21xp5_ASAP7_75t_L g622 ( .A1(n_545), .A2(n_349), .B(n_309), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_563), .Y(n_623) );
NOR2xp33_ASAP7_75t_R g624 ( .A(n_544), .B(n_349), .Y(n_624) );
AND2x4_ASAP7_75t_L g625 ( .A(n_580), .B(n_219), .Y(n_625) );
NAND2xp5_ASAP7_75t_SL g626 ( .A(n_558), .B(n_210), .Y(n_626) );
AND2x2_ASAP7_75t_L g627 ( .A(n_544), .B(n_223), .Y(n_627) );
AND2x2_ASAP7_75t_L g628 ( .A(n_546), .B(n_223), .Y(n_628) );
AND2x2_ASAP7_75t_L g629 ( .A(n_546), .B(n_315), .Y(n_629) );
INVx2_ASAP7_75t_L g630 ( .A(n_593), .Y(n_630) );
INVxp67_ASAP7_75t_SL g631 ( .A(n_588), .Y(n_631) );
NOR2xp33_ASAP7_75t_L g632 ( .A(n_590), .B(n_547), .Y(n_632) );
XOR2x2_ASAP7_75t_L g633 ( .A(n_595), .B(n_557), .Y(n_633) );
AOI22x1_ASAP7_75t_SL g634 ( .A1(n_589), .A2(n_573), .B1(n_577), .B2(n_580), .Y(n_634) );
AND3x1_ASAP7_75t_L g635 ( .A(n_589), .B(n_562), .C(n_556), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_596), .Y(n_636) );
NOR2xp33_ASAP7_75t_L g637 ( .A(n_586), .B(n_537), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_594), .B(n_574), .Y(n_638) );
INVxp67_ASAP7_75t_SL g639 ( .A(n_588), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_611), .Y(n_640) );
INVx2_ASAP7_75t_SL g641 ( .A(n_584), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_586), .B(n_570), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_620), .B(n_570), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_617), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_623), .B(n_578), .Y(n_645) );
OAI211xp5_ASAP7_75t_L g646 ( .A1(n_624), .A2(n_539), .B(n_549), .C(n_536), .Y(n_646) );
NAND3xp33_ASAP7_75t_L g647 ( .A(n_619), .B(n_564), .C(n_526), .Y(n_647) );
AOI221xp5_ASAP7_75t_L g648 ( .A1(n_598), .A2(n_565), .B1(n_567), .B2(n_556), .C(n_569), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_592), .B(n_565), .Y(n_649) );
NAND2xp5_ASAP7_75t_SL g650 ( .A(n_624), .B(n_549), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_592), .B(n_539), .Y(n_651) );
AND2x4_ASAP7_75t_L g652 ( .A(n_589), .B(n_580), .Y(n_652) );
XOR2x2_ASAP7_75t_L g653 ( .A(n_595), .B(n_568), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_597), .Y(n_654) );
A2O1A1Ixp33_ASAP7_75t_L g655 ( .A1(n_587), .A2(n_568), .B(n_561), .C(n_579), .Y(n_655) );
INVx1_ASAP7_75t_SL g656 ( .A(n_607), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_599), .Y(n_657) );
AOI211xp5_ASAP7_75t_L g658 ( .A1(n_618), .A2(n_583), .B(n_533), .C(n_315), .Y(n_658) );
XOR2x2_ASAP7_75t_L g659 ( .A(n_585), .B(n_583), .Y(n_659) );
AO22x1_ASAP7_75t_L g660 ( .A1(n_604), .A2(n_262), .B1(n_533), .B2(n_605), .Y(n_660) );
AND2x2_ASAP7_75t_L g661 ( .A(n_602), .B(n_533), .Y(n_661) );
NAND2xp33_ASAP7_75t_SL g662 ( .A(n_618), .B(n_262), .Y(n_662) );
OA222x2_ASAP7_75t_L g663 ( .A1(n_603), .A2(n_262), .B1(n_601), .B2(n_600), .C1(n_610), .C2(n_616), .Y(n_663) );
AOI21xp33_ASAP7_75t_SL g664 ( .A1(n_606), .A2(n_621), .B(n_608), .Y(n_664) );
INVxp33_ASAP7_75t_SL g665 ( .A(n_627), .Y(n_665) );
OAI22xp5_ASAP7_75t_L g666 ( .A1(n_621), .A2(n_609), .B1(n_626), .B2(n_629), .Y(n_666) );
OAI22xp33_ASAP7_75t_L g667 ( .A1(n_626), .A2(n_628), .B1(n_613), .B2(n_614), .Y(n_667) );
NAND3xp33_ASAP7_75t_L g668 ( .A(n_614), .B(n_612), .C(n_625), .Y(n_668) );
INVx1_ASAP7_75t_SL g669 ( .A(n_625), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_625), .Y(n_670) );
INVx1_ASAP7_75t_SL g671 ( .A(n_622), .Y(n_671) );
NOR3xp33_ASAP7_75t_SL g672 ( .A(n_615), .B(n_586), .C(n_413), .Y(n_672) );
XNOR2xp5_ASAP7_75t_L g673 ( .A(n_591), .B(n_380), .Y(n_673) );
INVx3_ASAP7_75t_L g674 ( .A(n_589), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_596), .Y(n_675) );
OAI211xp5_ASAP7_75t_L g676 ( .A1(n_624), .A2(n_582), .B(n_595), .C(n_587), .Y(n_676) );
OA22x2_ASAP7_75t_L g677 ( .A1(n_595), .A2(n_589), .B1(n_527), .B2(n_590), .Y(n_677) );
AOI22xp5_ASAP7_75t_L g678 ( .A1(n_586), .A2(n_592), .B1(n_413), .B2(n_598), .Y(n_678) );
NAND2xp33_ASAP7_75t_SL g679 ( .A(n_624), .B(n_595), .Y(n_679) );
AOI221xp5_ASAP7_75t_L g680 ( .A1(n_637), .A2(n_664), .B1(n_642), .B2(n_678), .C(n_667), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_641), .B(n_657), .Y(n_681) );
OAI32xp33_ASAP7_75t_L g682 ( .A1(n_679), .A2(n_674), .A3(n_662), .B1(n_665), .B2(n_666), .Y(n_682) );
OAI21xp5_ASAP7_75t_L g683 ( .A1(n_677), .A2(n_655), .B(n_676), .Y(n_683) );
HB1xp67_ASAP7_75t_L g684 ( .A(n_639), .Y(n_684) );
AOI221xp5_ASAP7_75t_L g685 ( .A1(n_637), .A2(n_654), .B1(n_632), .B2(n_675), .C(n_640), .Y(n_685) );
AOI21xp33_ASAP7_75t_L g686 ( .A1(n_632), .A2(n_671), .B(n_677), .Y(n_686) );
NOR2xp33_ASAP7_75t_L g687 ( .A(n_673), .B(n_641), .Y(n_687) );
AOI21xp33_ASAP7_75t_L g688 ( .A1(n_676), .A2(n_668), .B(n_647), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_636), .Y(n_689) );
NAND3xp33_ASAP7_75t_L g690 ( .A(n_672), .B(n_655), .C(n_658), .Y(n_690) );
OAI21xp5_ASAP7_75t_SL g691 ( .A1(n_666), .A2(n_646), .B(n_674), .Y(n_691) );
HB1xp67_ASAP7_75t_L g692 ( .A(n_631), .Y(n_692) );
HB1xp67_ASAP7_75t_L g693 ( .A(n_630), .Y(n_693) );
INVx2_ASAP7_75t_L g694 ( .A(n_693), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_684), .Y(n_695) );
NOR2xp33_ASAP7_75t_SL g696 ( .A(n_682), .B(n_669), .Y(n_696) );
OAI211xp5_ASAP7_75t_L g697 ( .A1(n_683), .A2(n_650), .B(n_670), .C(n_648), .Y(n_697) );
OAI311xp33_ASAP7_75t_L g698 ( .A1(n_680), .A2(n_663), .A3(n_633), .B1(n_649), .C1(n_651), .Y(n_698) );
NAND4xp25_ASAP7_75t_SL g699 ( .A(n_688), .B(n_633), .C(n_656), .D(n_635), .Y(n_699) );
AOI321xp33_ASAP7_75t_L g700 ( .A1(n_685), .A2(n_650), .A3(n_661), .B1(n_652), .B2(n_645), .C(n_643), .Y(n_700) );
AOI22xp5_ASAP7_75t_L g701 ( .A1(n_690), .A2(n_653), .B1(n_659), .B2(n_634), .Y(n_701) );
NAND3xp33_ASAP7_75t_SL g702 ( .A(n_691), .B(n_638), .C(n_660), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_695), .Y(n_703) );
INVx2_ASAP7_75t_L g704 ( .A(n_694), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_697), .Y(n_705) );
INVxp33_ASAP7_75t_L g706 ( .A(n_696), .Y(n_706) );
INVxp33_ASAP7_75t_SL g707 ( .A(n_701), .Y(n_707) );
AOI22xp5_ASAP7_75t_L g708 ( .A1(n_707), .A2(n_699), .B1(n_702), .B2(n_686), .Y(n_708) );
NAND3xp33_ASAP7_75t_L g709 ( .A(n_705), .B(n_700), .C(n_692), .Y(n_709) );
AND2x4_ASAP7_75t_L g710 ( .A(n_703), .B(n_687), .Y(n_710) );
INVx2_ASAP7_75t_L g711 ( .A(n_710), .Y(n_711) );
AND3x1_ASAP7_75t_L g712 ( .A(n_708), .B(n_705), .C(n_703), .Y(n_712) );
OR2x6_ASAP7_75t_L g713 ( .A(n_711), .B(n_709), .Y(n_713) );
INVxp67_ASAP7_75t_SL g714 ( .A(n_712), .Y(n_714) );
OAI21xp5_ASAP7_75t_L g715 ( .A1(n_714), .A2(n_706), .B(n_699), .Y(n_715) );
OAI22xp33_ASAP7_75t_L g716 ( .A1(n_715), .A2(n_713), .B1(n_704), .B2(n_698), .Y(n_716) );
AOI222xp33_ASAP7_75t_L g717 ( .A1(n_716), .A2(n_704), .B1(n_689), .B2(n_681), .C1(n_693), .C2(n_644), .Y(n_717) );
endmodule