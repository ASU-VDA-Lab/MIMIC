module fake_netlist_1_8116_n_13 (n_1, n_2, n_0, n_13);
input n_1;
input n_2;
input n_0;
output n_13;
wire n_11;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_8;
wire n_10;
wire n_7;
OR2x2_ASAP7_75t_L g3 ( .A(n_0), .B(n_2), .Y(n_3) );
INVx1_ASAP7_75t_L g4 ( .A(n_2), .Y(n_4) );
OR2x6_ASAP7_75t_L g5 ( .A(n_3), .B(n_0), .Y(n_5) );
OAI21x1_ASAP7_75t_L g6 ( .A1(n_4), .A2(n_3), .B(n_1), .Y(n_6) );
OR2x2_ASAP7_75t_L g7 ( .A(n_5), .B(n_0), .Y(n_7) );
AND2x2_ASAP7_75t_L g8 ( .A(n_5), .B(n_0), .Y(n_8) );
AOI211x1_ASAP7_75t_L g9 ( .A1(n_8), .A2(n_5), .B(n_6), .C(n_1), .Y(n_9) );
AOI31xp33_ASAP7_75t_L g10 ( .A1(n_9), .A2(n_7), .A3(n_5), .B(n_2), .Y(n_10) );
OAI21xp5_ASAP7_75t_L g11 ( .A1(n_9), .A2(n_6), .B(n_5), .Y(n_11) );
NAND3xp33_ASAP7_75t_SL g12 ( .A(n_11), .B(n_1), .C(n_6), .Y(n_12) );
OA21x2_ASAP7_75t_L g13 ( .A1(n_12), .A2(n_10), .B(n_1), .Y(n_13) );
endmodule