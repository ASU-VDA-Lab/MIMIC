module fake_netlist_6_3982_n_179 (n_16, n_1, n_9, n_8, n_18, n_10, n_21, n_24, n_6, n_15, n_27, n_3, n_14, n_0, n_4, n_22, n_26, n_13, n_11, n_28, n_17, n_23, n_12, n_20, n_7, n_30, n_2, n_5, n_19, n_29, n_31, n_25, n_179);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_6;
input n_15;
input n_27;
input n_3;
input n_14;
input n_0;
input n_4;
input n_22;
input n_26;
input n_13;
input n_11;
input n_28;
input n_17;
input n_23;
input n_12;
input n_20;
input n_7;
input n_30;
input n_2;
input n_5;
input n_19;
input n_29;
input n_31;
input n_25;

output n_179;

wire n_52;
wire n_91;
wire n_119;
wire n_46;
wire n_146;
wire n_163;
wire n_147;
wire n_154;
wire n_88;
wire n_98;
wire n_113;
wire n_39;
wire n_63;
wire n_73;
wire n_148;
wire n_138;
wire n_161;
wire n_68;
wire n_166;
wire n_50;
wire n_158;
wire n_49;
wire n_83;
wire n_167;
wire n_101;
wire n_144;
wire n_174;
wire n_127;
wire n_125;
wire n_153;
wire n_168;
wire n_178;
wire n_77;
wire n_156;
wire n_149;
wire n_152;
wire n_106;
wire n_92;
wire n_145;
wire n_42;
wire n_133;
wire n_96;
wire n_90;
wire n_160;
wire n_131;
wire n_105;
wire n_54;
wire n_132;
wire n_102;
wire n_87;
wire n_32;
wire n_66;
wire n_99;
wire n_130;
wire n_78;
wire n_84;
wire n_85;
wire n_164;
wire n_100;
wire n_129;
wire n_121;
wire n_137;
wire n_142;
wire n_143;
wire n_47;
wire n_62;
wire n_155;
wire n_75;
wire n_109;
wire n_150;
wire n_122;
wire n_45;
wire n_34;
wire n_140;
wire n_70;
wire n_120;
wire n_37;
wire n_67;
wire n_33;
wire n_82;
wire n_38;
wire n_110;
wire n_151;
wire n_61;
wire n_112;
wire n_172;
wire n_81;
wire n_59;
wire n_76;
wire n_36;
wire n_124;
wire n_55;
wire n_126;
wire n_94;
wire n_97;
wire n_108;
wire n_58;
wire n_116;
wire n_64;
wire n_117;
wire n_118;
wire n_175;
wire n_48;
wire n_65;
wire n_40;
wire n_93;
wire n_80;
wire n_141;
wire n_135;
wire n_165;
wire n_139;
wire n_41;
wire n_134;
wire n_177;
wire n_176;
wire n_114;
wire n_86;
wire n_104;
wire n_95;
wire n_107;
wire n_71;
wire n_74;
wire n_123;
wire n_136;
wire n_72;
wire n_89;
wire n_173;
wire n_103;
wire n_111;
wire n_60;
wire n_159;
wire n_157;
wire n_162;
wire n_170;
wire n_35;
wire n_115;
wire n_69;
wire n_128;
wire n_79;
wire n_43;
wire n_171;
wire n_57;
wire n_169;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

INVxp67_ASAP7_75t_SL g32 ( 
.A(n_22),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

CKINVDCx5p33_ASAP7_75t_R g36 ( 
.A(n_25),
.Y(n_36)
);

CKINVDCx5p33_ASAP7_75t_R g37 ( 
.A(n_5),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_31),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_4),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_1),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

CKINVDCx5p33_ASAP7_75t_R g46 ( 
.A(n_23),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_15),
.Y(n_50)
);

CKINVDCx5p33_ASAP7_75t_R g51 ( 
.A(n_7),
.Y(n_51)
);

INVxp67_ASAP7_75t_SL g52 ( 
.A(n_6),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_35),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_35),
.B(n_2),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_4),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_34),
.B(n_5),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_47),
.B(n_6),
.Y(n_65)
);

AND2x6_ASAP7_75t_L g66 ( 
.A(n_33),
.B(n_30),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_7),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_8),
.Y(n_68)
);

AND2x4_ASAP7_75t_SL g69 ( 
.A(n_40),
.B(n_9),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_38),
.B(n_12),
.Y(n_70)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVxp67_ASAP7_75t_SL g73 ( 
.A(n_45),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_49),
.B(n_14),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_53),
.B(n_17),
.Y(n_75)
);

NOR3xp33_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_52),
.C(n_51),
.Y(n_76)
);

NAND2x1p5_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_50),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

NOR2xp67_ASAP7_75t_L g80 ( 
.A(n_61),
.B(n_46),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_64),
.A2(n_37),
.B1(n_51),
.B2(n_42),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_73),
.A2(n_32),
.B(n_46),
.Y(n_82)
);

AOI21x1_ASAP7_75t_L g83 ( 
.A1(n_74),
.A2(n_18),
.B(n_19),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_60),
.A2(n_37),
.B(n_43),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

OA22x2_ASAP7_75t_L g86 ( 
.A1(n_63),
.A2(n_27),
.B1(n_29),
.B2(n_65),
.Y(n_86)
);

A2O1A1Ixp33_ASAP7_75t_L g87 ( 
.A1(n_63),
.A2(n_65),
.B(n_55),
.C(n_56),
.Y(n_87)
);

OAI21x1_ASAP7_75t_L g88 ( 
.A1(n_72),
.A2(n_58),
.B(n_70),
.Y(n_88)
);

NAND2x1p5_ASAP7_75t_L g89 ( 
.A(n_61),
.B(n_71),
.Y(n_89)
);

CKINVDCx5p33_ASAP7_75t_R g90 ( 
.A(n_71),
.Y(n_90)
);

CKINVDCx10_ASAP7_75t_R g91 ( 
.A(n_69),
.Y(n_91)
);

AND2x4_ASAP7_75t_L g92 ( 
.A(n_71),
.B(n_59),
.Y(n_92)
);

BUFx10_ASAP7_75t_L g93 ( 
.A(n_90),
.Y(n_93)
);

AOI21x1_ASAP7_75t_L g94 ( 
.A1(n_78),
.A2(n_58),
.B(n_59),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_92),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_92),
.B(n_75),
.Y(n_96)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

AND2x4_ASAP7_75t_L g98 ( 
.A(n_87),
.B(n_69),
.Y(n_98)
);

AND2x4_ASAP7_75t_L g99 ( 
.A(n_87),
.B(n_66),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

NOR2x1_ASAP7_75t_SL g101 ( 
.A(n_83),
.B(n_62),
.Y(n_101)
);

BUFx2_ASAP7_75t_L g102 ( 
.A(n_89),
.Y(n_102)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_89),
.A2(n_68),
.B1(n_67),
.B2(n_72),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_94),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_94),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_103),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_103),
.Y(n_108)
);

INVx2_ASAP7_75t_SL g109 ( 
.A(n_97),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_102),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_98),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_95),
.B(n_86),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_110),
.B(n_95),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_112),
.A2(n_111),
.B(n_76),
.Y(n_114)
);

AOI221xp5_ASAP7_75t_L g115 ( 
.A1(n_112),
.A2(n_81),
.B1(n_76),
.B2(n_97),
.C(n_84),
.Y(n_115)
);

NAND4xp25_ASAP7_75t_L g116 ( 
.A(n_110),
.B(n_67),
.C(n_56),
.D(n_55),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_109),
.B(n_97),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_110),
.B(n_93),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_109),
.A2(n_97),
.B1(n_99),
.B2(n_66),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_117),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_118),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_113),
.B(n_93),
.Y(n_122)
);

OR2x6_ASAP7_75t_L g123 ( 
.A(n_114),
.B(n_97),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_116),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_123),
.B(n_115),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_123),
.B(n_98),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_122),
.B(n_91),
.Y(n_127)
);

AND2x4_ASAP7_75t_L g128 ( 
.A(n_123),
.B(n_98),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_121),
.B(n_98),
.Y(n_129)
);

INVx1_ASAP7_75t_SL g130 ( 
.A(n_124),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_120),
.B(n_102),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_124),
.Y(n_132)
);

INVx1_ASAP7_75t_SL g133 ( 
.A(n_124),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_121),
.B(n_93),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_124),
.Y(n_135)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_129),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_131),
.B(n_77),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_132),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_131),
.B(n_93),
.Y(n_139)
);

INVx1_ASAP7_75t_SL g140 ( 
.A(n_130),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_125),
.B(n_77),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_129),
.B(n_80),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_138),
.Y(n_143)
);

NAND4xp25_ASAP7_75t_L g144 ( 
.A(n_137),
.B(n_132),
.C(n_130),
.D(n_133),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_136),
.Y(n_145)
);

NAND2x1p5_ASAP7_75t_L g146 ( 
.A(n_140),
.B(n_128),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_136),
.Y(n_147)
);

OAI221xp5_ASAP7_75t_L g148 ( 
.A1(n_139),
.A2(n_127),
.B1(n_134),
.B2(n_125),
.C(n_135),
.Y(n_148)
);

NAND3xp33_ASAP7_75t_L g149 ( 
.A(n_141),
.B(n_104),
.C(n_96),
.Y(n_149)
);

AO21x1_ASAP7_75t_L g150 ( 
.A1(n_139),
.A2(n_128),
.B(n_126),
.Y(n_150)
);

NOR3x1_ASAP7_75t_L g151 ( 
.A(n_142),
.B(n_107),
.C(n_108),
.Y(n_151)
);

NOR3xp33_ASAP7_75t_L g152 ( 
.A(n_142),
.B(n_126),
.C(n_128),
.Y(n_152)
);

INVxp67_ASAP7_75t_SL g153 ( 
.A(n_145),
.Y(n_153)
);

NOR2x1_ASAP7_75t_L g154 ( 
.A(n_144),
.B(n_128),
.Y(n_154)
);

OAI22xp33_ASAP7_75t_L g155 ( 
.A1(n_148),
.A2(n_72),
.B1(n_62),
.B2(n_100),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_143),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_145),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_152),
.A2(n_66),
.B1(n_99),
.B2(n_119),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_147),
.Y(n_159)
);

AND2x4_ASAP7_75t_L g160 ( 
.A(n_151),
.B(n_79),
.Y(n_160)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_146),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_149),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_156),
.Y(n_163)
);

AND2x2_ASAP7_75t_SL g164 ( 
.A(n_162),
.B(n_150),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_159),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_157),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_153),
.Y(n_167)
);

NOR2xp67_ASAP7_75t_L g168 ( 
.A(n_160),
.B(n_100),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_161),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_161),
.B(n_85),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_164),
.A2(n_154),
.B1(n_155),
.B2(n_160),
.Y(n_171)
);

OAI222xp33_ASAP7_75t_L g172 ( 
.A1(n_170),
.A2(n_158),
.B1(n_119),
.B2(n_82),
.C1(n_99),
.C2(n_105),
.Y(n_172)
);

NAND5xp2_ASAP7_75t_L g173 ( 
.A(n_167),
.B(n_108),
.C(n_107),
.D(n_105),
.E(n_66),
.Y(n_173)
);

OAI21xp33_ASAP7_75t_L g174 ( 
.A1(n_170),
.A2(n_169),
.B(n_163),
.Y(n_174)
);

OAI221xp5_ASAP7_75t_L g175 ( 
.A1(n_174),
.A2(n_171),
.B1(n_168),
.B2(n_165),
.C(n_166),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_172),
.B(n_168),
.Y(n_176)
);

AO21x2_ASAP7_75t_L g177 ( 
.A1(n_173),
.A2(n_101),
.B(n_106),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_175),
.A2(n_99),
.B1(n_106),
.B2(n_66),
.Y(n_178)
);

AOI221xp5_ASAP7_75t_L g179 ( 
.A1(n_178),
.A2(n_176),
.B1(n_177),
.B2(n_103),
.C(n_66),
.Y(n_179)
);


endmodule