module fake_netlist_6_4453_n_1851 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1851);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1851;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_1810;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_535;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

BUFx10_ASAP7_75t_L g173 ( 
.A(n_151),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_113),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_33),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_135),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_90),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_95),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_144),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_141),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_150),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_17),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_6),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_58),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_76),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_56),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_54),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_155),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_6),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_1),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_26),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_51),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_101),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_166),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_16),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_108),
.Y(n_196)
);

BUFx10_ASAP7_75t_L g197 ( 
.A(n_83),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_106),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_70),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_5),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_120),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_72),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_37),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_53),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_170),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_51),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_22),
.Y(n_207)
);

BUFx10_ASAP7_75t_L g208 ( 
.A(n_147),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_29),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_114),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_45),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_161),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_87),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_4),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_118),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_154),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_124),
.Y(n_217)
);

BUFx2_ASAP7_75t_SL g218 ( 
.A(n_130),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_19),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_53),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_105),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_115),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_62),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_41),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_3),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_159),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_139),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_21),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_33),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_7),
.Y(n_230)
);

INVx2_ASAP7_75t_SL g231 ( 
.A(n_41),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_44),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_81),
.Y(n_233)
);

BUFx2_ASAP7_75t_L g234 ( 
.A(n_35),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_56),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_30),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_93),
.Y(n_237)
);

BUFx2_ASAP7_75t_L g238 ( 
.A(n_47),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_165),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_143),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_19),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_26),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_140),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_0),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_30),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_132),
.Y(n_246)
);

BUFx8_ASAP7_75t_SL g247 ( 
.A(n_133),
.Y(n_247)
);

INVxp67_ASAP7_75t_SL g248 ( 
.A(n_80),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_152),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_69),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_46),
.Y(n_251)
);

INVx2_ASAP7_75t_SL g252 ( 
.A(n_121),
.Y(n_252)
);

BUFx3_ASAP7_75t_L g253 ( 
.A(n_39),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_164),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_103),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_52),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_47),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_79),
.Y(n_258)
);

BUFx10_ASAP7_75t_L g259 ( 
.A(n_40),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_134),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_45),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_157),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_54),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_60),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_66),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_13),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_21),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_156),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_43),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_11),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_97),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_82),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_171),
.Y(n_273)
);

BUFx10_ASAP7_75t_L g274 ( 
.A(n_49),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_22),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_0),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_160),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_49),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_168),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_127),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_129),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_20),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_142),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_119),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_123),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_38),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_16),
.Y(n_287)
);

INVxp33_ASAP7_75t_L g288 ( 
.A(n_136),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_77),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_7),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_65),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_107),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_125),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_146),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_137),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_86),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_167),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_99),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_61),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_64),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_28),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_98),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_43),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_94),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_2),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_78),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_74),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_131),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_158),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_88),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_12),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_73),
.Y(n_312)
);

INVx2_ASAP7_75t_SL g313 ( 
.A(n_68),
.Y(n_313)
);

INVx2_ASAP7_75t_SL g314 ( 
.A(n_36),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_17),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_91),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_14),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_46),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_112),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_9),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_145),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_24),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_44),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_18),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_28),
.Y(n_325)
);

BUFx3_ASAP7_75t_L g326 ( 
.A(n_39),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_10),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_13),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_149),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_89),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_52),
.Y(n_331)
);

BUFx2_ASAP7_75t_SL g332 ( 
.A(n_169),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_59),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_34),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_117),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_31),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_37),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_34),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_122),
.Y(n_339)
);

INVx1_ASAP7_75t_SL g340 ( 
.A(n_84),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_20),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_104),
.Y(n_342)
);

BUFx3_ASAP7_75t_L g343 ( 
.A(n_63),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_40),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_27),
.Y(n_345)
);

INVxp67_ASAP7_75t_SL g346 ( 
.A(n_194),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_183),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_247),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_183),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_183),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_174),
.Y(n_351)
);

INVxp67_ASAP7_75t_SL g352 ( 
.A(n_194),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_183),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_183),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_303),
.Y(n_355)
);

INVxp67_ASAP7_75t_SL g356 ( 
.A(n_249),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_176),
.Y(n_357)
);

INVxp33_ASAP7_75t_SL g358 ( 
.A(n_234),
.Y(n_358)
);

HB1xp67_ASAP7_75t_L g359 ( 
.A(n_234),
.Y(n_359)
);

INVxp67_ASAP7_75t_SL g360 ( 
.A(n_249),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_303),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_303),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_303),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_181),
.Y(n_364)
);

INVx1_ASAP7_75t_SL g365 ( 
.A(n_238),
.Y(n_365)
);

BUFx3_ASAP7_75t_L g366 ( 
.A(n_343),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_303),
.Y(n_367)
);

INVxp33_ASAP7_75t_SL g368 ( 
.A(n_238),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_178),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_190),
.Y(n_370)
);

INVxp33_ASAP7_75t_SL g371 ( 
.A(n_182),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_285),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_186),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_190),
.Y(n_374)
);

CKINVDCx16_ASAP7_75t_R g375 ( 
.A(n_175),
.Y(n_375)
);

CKINVDCx16_ASAP7_75t_R g376 ( 
.A(n_175),
.Y(n_376)
);

HB1xp67_ASAP7_75t_L g377 ( 
.A(n_203),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_339),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_200),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_180),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_227),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_180),
.Y(n_382)
);

INVxp67_ASAP7_75t_SL g383 ( 
.A(n_343),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_199),
.Y(n_384)
);

CKINVDCx16_ASAP7_75t_R g385 ( 
.A(n_203),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_200),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_215),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_245),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_245),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_201),
.Y(n_390)
);

INVxp67_ASAP7_75t_SL g391 ( 
.A(n_296),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_202),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_263),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_263),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_186),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_184),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_215),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_187),
.Y(n_398)
);

CKINVDCx16_ASAP7_75t_R g399 ( 
.A(n_241),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_187),
.Y(n_400)
);

HB1xp67_ASAP7_75t_L g401 ( 
.A(n_241),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_204),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_204),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_206),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_210),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_206),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_216),
.Y(n_407)
);

BUFx3_ASAP7_75t_L g408 ( 
.A(n_173),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_222),
.Y(n_409)
);

HB1xp67_ASAP7_75t_L g410 ( 
.A(n_275),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_223),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_207),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_207),
.Y(n_413)
);

CKINVDCx16_ASAP7_75t_R g414 ( 
.A(n_275),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_226),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_242),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_242),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_233),
.Y(n_418)
);

INVxp33_ASAP7_75t_SL g419 ( 
.A(n_191),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_251),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_227),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_251),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_237),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_305),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_239),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_305),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_320),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_240),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_320),
.Y(n_429)
);

INVxp67_ASAP7_75t_SL g430 ( 
.A(n_335),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_324),
.Y(n_431)
);

AND2x4_ASAP7_75t_L g432 ( 
.A(n_353),
.B(n_252),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_347),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_421),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_421),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_347),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_358),
.A2(n_286),
.B1(n_232),
.B2(n_317),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_SL g438 ( 
.A(n_365),
.B(n_301),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_421),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_351),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_346),
.B(n_252),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_349),
.Y(n_442)
);

INVx3_ASAP7_75t_L g443 ( 
.A(n_421),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_349),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_352),
.B(n_253),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_356),
.B(n_313),
.Y(n_446)
);

INVx6_ASAP7_75t_L g447 ( 
.A(n_381),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_421),
.Y(n_448)
);

AND2x4_ASAP7_75t_L g449 ( 
.A(n_353),
.B(n_313),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g450 ( 
.A(n_360),
.B(n_253),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_421),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_357),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_369),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_381),
.Y(n_454)
);

INVx3_ASAP7_75t_L g455 ( 
.A(n_381),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_383),
.B(n_326),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_381),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_368),
.B(n_301),
.Y(n_458)
);

AND2x4_ASAP7_75t_L g459 ( 
.A(n_350),
.B(n_354),
.Y(n_459)
);

BUFx2_ASAP7_75t_L g460 ( 
.A(n_380),
.Y(n_460)
);

BUFx3_ASAP7_75t_L g461 ( 
.A(n_381),
.Y(n_461)
);

BUFx2_ASAP7_75t_L g462 ( 
.A(n_382),
.Y(n_462)
);

OAI21x1_ASAP7_75t_L g463 ( 
.A1(n_396),
.A2(n_179),
.B(n_177),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_350),
.Y(n_464)
);

HB1xp67_ASAP7_75t_L g465 ( 
.A(n_377),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_354),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_355),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_387),
.A2(n_282),
.B1(n_236),
.B2(n_344),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_355),
.B(n_250),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_361),
.B(n_362),
.Y(n_470)
);

HB1xp67_ASAP7_75t_L g471 ( 
.A(n_401),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_384),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_396),
.B(n_326),
.Y(n_473)
);

HB1xp67_ASAP7_75t_L g474 ( 
.A(n_410),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_361),
.Y(n_475)
);

AND2x4_ASAP7_75t_L g476 ( 
.A(n_362),
.B(n_177),
.Y(n_476)
);

HB1xp67_ASAP7_75t_L g477 ( 
.A(n_359),
.Y(n_477)
);

NOR2x1_ASAP7_75t_L g478 ( 
.A(n_363),
.B(n_218),
.Y(n_478)
);

HB1xp67_ASAP7_75t_L g479 ( 
.A(n_366),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_SL g480 ( 
.A1(n_375),
.A2(n_331),
.B1(n_325),
.B2(n_324),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_366),
.B(n_184),
.Y(n_481)
);

BUFx3_ASAP7_75t_L g482 ( 
.A(n_363),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_390),
.Y(n_483)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_367),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_392),
.Y(n_485)
);

HB1xp67_ASAP7_75t_L g486 ( 
.A(n_375),
.Y(n_486)
);

INVx3_ASAP7_75t_L g487 ( 
.A(n_367),
.Y(n_487)
);

OAI21x1_ASAP7_75t_L g488 ( 
.A1(n_389),
.A2(n_185),
.B(n_179),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_407),
.Y(n_489)
);

AND2x4_ASAP7_75t_L g490 ( 
.A(n_389),
.B(n_185),
.Y(n_490)
);

BUFx12f_ASAP7_75t_L g491 ( 
.A(n_348),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_395),
.Y(n_492)
);

AND2x6_ASAP7_75t_L g493 ( 
.A(n_408),
.B(n_227),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_395),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_398),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_370),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_370),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_376),
.A2(n_325),
.B1(n_331),
.B2(n_189),
.Y(n_498)
);

INVx3_ASAP7_75t_L g499 ( 
.A(n_374),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_374),
.Y(n_500)
);

AND2x4_ASAP7_75t_L g501 ( 
.A(n_398),
.B(n_188),
.Y(n_501)
);

HB1xp67_ASAP7_75t_L g502 ( 
.A(n_376),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_391),
.B(n_430),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_379),
.B(n_193),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_379),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_400),
.Y(n_506)
);

AND2x4_ASAP7_75t_L g507 ( 
.A(n_400),
.B(n_188),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_402),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_459),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_459),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_459),
.Y(n_511)
);

OR2x2_ASAP7_75t_L g512 ( 
.A(n_477),
.B(n_385),
.Y(n_512)
);

INVx4_ASAP7_75t_L g513 ( 
.A(n_457),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_503),
.B(n_409),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_440),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_452),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_482),
.Y(n_517)
);

BUFx3_ASAP7_75t_L g518 ( 
.A(n_461),
.Y(n_518)
);

INVx3_ASAP7_75t_L g519 ( 
.A(n_434),
.Y(n_519)
);

INVx3_ASAP7_75t_L g520 ( 
.A(n_434),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_457),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_469),
.B(n_411),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_459),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_482),
.Y(n_524)
);

NAND3xp33_ASAP7_75t_L g525 ( 
.A(n_441),
.B(n_446),
.C(n_445),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_482),
.Y(n_526)
);

NOR2x1p5_ASAP7_75t_L g527 ( 
.A(n_453),
.B(n_408),
.Y(n_527)
);

INVx5_ASAP7_75t_L g528 ( 
.A(n_434),
.Y(n_528)
);

BUFx2_ASAP7_75t_L g529 ( 
.A(n_486),
.Y(n_529)
);

AND2x2_ASAP7_75t_SL g530 ( 
.A(n_438),
.B(n_198),
.Y(n_530)
);

INVx2_ASAP7_75t_SL g531 ( 
.A(n_479),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_459),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_433),
.Y(n_533)
);

OR2x2_ASAP7_75t_L g534 ( 
.A(n_477),
.B(n_385),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_457),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_433),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_464),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_436),
.Y(n_538)
);

HB1xp67_ASAP7_75t_L g539 ( 
.A(n_486),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_436),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_464),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_442),
.Y(n_542)
);

INVx2_ASAP7_75t_SL g543 ( 
.A(n_479),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_464),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_503),
.B(n_445),
.Y(n_545)
);

BUFx10_ASAP7_75t_L g546 ( 
.A(n_472),
.Y(n_546)
);

XNOR2xp5_ASAP7_75t_L g547 ( 
.A(n_437),
.B(n_364),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_442),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_464),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_444),
.Y(n_550)
);

INVx2_ASAP7_75t_SL g551 ( 
.A(n_445),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_444),
.Y(n_552)
);

INVx3_ASAP7_75t_L g553 ( 
.A(n_434),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_434),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_466),
.Y(n_555)
);

AOI22xp33_ASAP7_75t_L g556 ( 
.A1(n_450),
.A2(n_231),
.B1(n_314),
.B2(n_332),
.Y(n_556)
);

INVx3_ASAP7_75t_L g557 ( 
.A(n_434),
.Y(n_557)
);

OAI22xp33_ASAP7_75t_L g558 ( 
.A1(n_438),
.A2(n_399),
.B1(n_414),
.B2(n_288),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_450),
.B(n_415),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_466),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_467),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_467),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_475),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_434),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_475),
.Y(n_565)
);

NAND2xp33_ASAP7_75t_R g566 ( 
.A(n_460),
.B(n_371),
.Y(n_566)
);

BUFx3_ASAP7_75t_L g567 ( 
.A(n_461),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_483),
.B(n_418),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_496),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_490),
.Y(n_570)
);

OAI21xp33_ASAP7_75t_SL g571 ( 
.A1(n_458),
.A2(n_314),
.B(n_231),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_450),
.B(n_423),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_485),
.B(n_419),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_496),
.Y(n_574)
);

BUFx6f_ASAP7_75t_L g575 ( 
.A(n_457),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_489),
.B(n_425),
.Y(n_576)
);

OR2x2_ASAP7_75t_L g577 ( 
.A(n_465),
.B(n_399),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_496),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_441),
.B(n_428),
.Y(n_579)
);

INVx4_ASAP7_75t_L g580 ( 
.A(n_457),
.Y(n_580)
);

NAND2xp33_ASAP7_75t_L g581 ( 
.A(n_493),
.B(n_227),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_446),
.B(n_405),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_496),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_490),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_457),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_497),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_456),
.B(n_340),
.Y(n_587)
);

OAI22xp5_ASAP7_75t_L g588 ( 
.A1(n_458),
.A2(n_414),
.B1(n_219),
.B2(n_397),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_490),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_497),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_456),
.B(n_478),
.Y(n_591)
);

NOR2x1p5_ASAP7_75t_L g592 ( 
.A(n_491),
.B(n_192),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_456),
.B(n_254),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_497),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_497),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_478),
.B(n_255),
.Y(n_596)
);

OAI22xp33_ASAP7_75t_SL g597 ( 
.A1(n_468),
.A2(n_271),
.B1(n_243),
.B2(n_329),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_432),
.B(n_258),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_500),
.Y(n_599)
);

INVx2_ASAP7_75t_SL g600 ( 
.A(n_465),
.Y(n_600)
);

AOI21x1_ASAP7_75t_L g601 ( 
.A1(n_463),
.A2(n_196),
.B(n_193),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_500),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_490),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_500),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_500),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_505),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_505),
.Y(n_607)
);

INVx2_ASAP7_75t_SL g608 ( 
.A(n_471),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_505),
.Y(n_609)
);

NAND3xp33_ASAP7_75t_L g610 ( 
.A(n_504),
.B(n_373),
.C(n_205),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_432),
.B(n_260),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_481),
.B(n_386),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_505),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_490),
.Y(n_614)
);

INVx2_ASAP7_75t_SL g615 ( 
.A(n_471),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_484),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_432),
.B(n_262),
.Y(n_617)
);

BUFx10_ASAP7_75t_L g618 ( 
.A(n_502),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_484),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_476),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_476),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_SL g622 ( 
.A(n_480),
.B(n_173),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_484),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_484),
.Y(n_624)
);

INVx1_ASAP7_75t_SL g625 ( 
.A(n_502),
.Y(n_625)
);

BUFx3_ASAP7_75t_L g626 ( 
.A(n_461),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_476),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_484),
.Y(n_628)
);

INVx4_ASAP7_75t_L g629 ( 
.A(n_457),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_491),
.Y(n_630)
);

OAI22xp33_ASAP7_75t_L g631 ( 
.A1(n_468),
.A2(n_266),
.B1(n_345),
.B2(n_269),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_432),
.B(n_264),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_474),
.B(n_372),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_449),
.B(n_272),
.Y(n_634)
);

OAI21xp33_ASAP7_75t_SL g635 ( 
.A1(n_504),
.A2(n_403),
.B(n_402),
.Y(n_635)
);

BUFx6f_ASAP7_75t_L g636 ( 
.A(n_457),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_487),
.Y(n_637)
);

INVx2_ASAP7_75t_SL g638 ( 
.A(n_474),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_481),
.B(n_378),
.Y(n_639)
);

INVx3_ASAP7_75t_L g640 ( 
.A(n_434),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_487),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_487),
.Y(n_642)
);

BUFx10_ASAP7_75t_L g643 ( 
.A(n_493),
.Y(n_643)
);

INVx2_ASAP7_75t_SL g644 ( 
.A(n_481),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_492),
.B(n_195),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_473),
.B(n_173),
.Y(n_646)
);

CKINVDCx20_ASAP7_75t_R g647 ( 
.A(n_460),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_476),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_476),
.Y(n_649)
);

INVx2_ASAP7_75t_SL g650 ( 
.A(n_473),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_487),
.Y(n_651)
);

INVx2_ASAP7_75t_SL g652 ( 
.A(n_473),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_504),
.B(n_386),
.Y(n_653)
);

INVx1_ASAP7_75t_SL g654 ( 
.A(n_460),
.Y(n_654)
);

CKINVDCx6p67_ASAP7_75t_R g655 ( 
.A(n_491),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_487),
.Y(n_656)
);

INVx3_ASAP7_75t_L g657 ( 
.A(n_461),
.Y(n_657)
);

AOI21xp5_ASAP7_75t_L g658 ( 
.A1(n_591),
.A2(n_470),
.B(n_439),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_579),
.B(n_449),
.Y(n_659)
);

AOI22xp33_ASAP7_75t_L g660 ( 
.A1(n_551),
.A2(n_480),
.B1(n_498),
.B2(n_507),
.Y(n_660)
);

OAI22xp5_ASAP7_75t_L g661 ( 
.A1(n_551),
.A2(n_283),
.B1(n_265),
.B2(n_198),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_509),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_532),
.Y(n_663)
);

AOI22xp33_ASAP7_75t_L g664 ( 
.A1(n_530),
.A2(n_498),
.B1(n_507),
.B2(n_501),
.Y(n_664)
);

BUFx5_ASAP7_75t_L g665 ( 
.A(n_643),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_545),
.B(n_449),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_509),
.B(n_227),
.Y(n_667)
);

OR2x2_ASAP7_75t_L g668 ( 
.A(n_512),
.B(n_462),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_644),
.B(n_449),
.Y(n_669)
);

OR2x6_ASAP7_75t_L g670 ( 
.A(n_529),
.B(n_600),
.Y(n_670)
);

NOR2x1p5_ASAP7_75t_L g671 ( 
.A(n_655),
.B(n_209),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_531),
.B(n_462),
.Y(n_672)
);

AOI22xp33_ASAP7_75t_L g673 ( 
.A1(n_530),
.A2(n_597),
.B1(n_622),
.B2(n_525),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_644),
.B(n_449),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_582),
.B(n_279),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_650),
.B(n_493),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_SL g677 ( 
.A(n_515),
.B(n_437),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_650),
.B(n_493),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_543),
.B(n_462),
.Y(n_679)
);

AOI22xp5_ASAP7_75t_L g680 ( 
.A1(n_525),
.A2(n_248),
.B1(n_493),
.B2(n_330),
.Y(n_680)
);

INVx2_ASAP7_75t_SL g681 ( 
.A(n_543),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_652),
.B(n_493),
.Y(n_682)
);

AND2x6_ASAP7_75t_SL g683 ( 
.A(n_633),
.B(n_403),
.Y(n_683)
);

INVx3_ASAP7_75t_L g684 ( 
.A(n_518),
.Y(n_684)
);

INVx8_ASAP7_75t_L g685 ( 
.A(n_630),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_652),
.B(n_493),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_522),
.B(n_493),
.Y(n_687)
);

BUFx6f_ASAP7_75t_L g688 ( 
.A(n_518),
.Y(n_688)
);

AOI22xp5_ASAP7_75t_L g689 ( 
.A1(n_559),
.A2(n_493),
.B1(n_302),
.B2(n_295),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_572),
.B(n_211),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_514),
.B(n_214),
.Y(n_691)
);

OAI22xp33_ASAP7_75t_L g692 ( 
.A1(n_622),
.A2(n_277),
.B1(n_333),
.B2(n_329),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_532),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_510),
.B(n_499),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_587),
.B(n_280),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_530),
.B(n_281),
.Y(n_696)
);

INVx8_ASAP7_75t_L g697 ( 
.A(n_630),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_511),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_511),
.B(n_499),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_593),
.B(n_571),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_523),
.B(n_246),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_537),
.Y(n_702)
);

OR2x2_ASAP7_75t_L g703 ( 
.A(n_512),
.B(n_492),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_517),
.B(n_524),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_524),
.B(n_499),
.Y(n_705)
);

INVxp67_ASAP7_75t_L g706 ( 
.A(n_639),
.Y(n_706)
);

OR2x6_ASAP7_75t_L g707 ( 
.A(n_529),
.B(n_218),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_570),
.Y(n_708)
);

INVx4_ASAP7_75t_L g709 ( 
.A(n_518),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_526),
.B(n_501),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_526),
.B(n_501),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_600),
.B(n_494),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_584),
.B(n_589),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_537),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_584),
.B(n_501),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_589),
.B(n_603),
.Y(n_716)
);

INVx2_ASAP7_75t_SL g717 ( 
.A(n_612),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_603),
.B(n_246),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_614),
.B(n_501),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_614),
.B(n_265),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_620),
.B(n_507),
.Y(n_721)
);

AOI22xp5_ASAP7_75t_L g722 ( 
.A1(n_620),
.A2(n_306),
.B1(n_291),
.B2(n_316),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_621),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_621),
.Y(n_724)
);

INVx3_ASAP7_75t_L g725 ( 
.A(n_567),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_627),
.B(n_507),
.Y(n_726)
);

AND2x2_ASAP7_75t_L g727 ( 
.A(n_608),
.B(n_495),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_558),
.B(n_289),
.Y(n_728)
);

AND2x2_ASAP7_75t_L g729 ( 
.A(n_608),
.B(n_495),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_597),
.B(n_292),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_541),
.Y(n_731)
);

INVxp67_ASAP7_75t_L g732 ( 
.A(n_645),
.Y(n_732)
);

INVx5_ASAP7_75t_L g733 ( 
.A(n_643),
.Y(n_733)
);

AOI22xp33_ASAP7_75t_L g734 ( 
.A1(n_653),
.A2(n_268),
.B1(n_205),
.B2(n_212),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_643),
.B(n_283),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_648),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_649),
.B(n_455),
.Y(n_737)
);

INVx2_ASAP7_75t_SL g738 ( 
.A(n_612),
.Y(n_738)
);

INVx2_ASAP7_75t_SL g739 ( 
.A(n_615),
.Y(n_739)
);

A2O1A1Ixp33_ASAP7_75t_L g740 ( 
.A1(n_635),
.A2(n_463),
.B(n_488),
.C(n_268),
.Y(n_740)
);

INVxp67_ASAP7_75t_L g741 ( 
.A(n_638),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_638),
.B(n_573),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_541),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_649),
.B(n_455),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_533),
.B(n_455),
.Y(n_745)
);

AOI22xp33_ASAP7_75t_L g746 ( 
.A1(n_653),
.A2(n_333),
.B1(n_212),
.B2(n_213),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_643),
.B(n_293),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_533),
.B(n_455),
.Y(n_748)
);

AND2x4_ASAP7_75t_L g749 ( 
.A(n_567),
.B(n_506),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_536),
.B(n_455),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_616),
.B(n_297),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_538),
.B(n_443),
.Y(n_752)
);

INVxp67_ASAP7_75t_L g753 ( 
.A(n_534),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_538),
.B(n_443),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_556),
.B(n_298),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_540),
.B(n_443),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_540),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_616),
.B(n_299),
.Y(n_758)
);

CKINVDCx16_ASAP7_75t_R g759 ( 
.A(n_566),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_542),
.B(n_443),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_542),
.B(n_196),
.Y(n_761)
);

INVxp67_ASAP7_75t_L g762 ( 
.A(n_534),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_548),
.B(n_213),
.Y(n_763)
);

AOI21xp5_ASAP7_75t_L g764 ( 
.A1(n_598),
.A2(n_439),
.B(n_435),
.Y(n_764)
);

CKINVDCx20_ASAP7_75t_R g765 ( 
.A(n_515),
.Y(n_765)
);

NOR2x1p5_ASAP7_75t_L g766 ( 
.A(n_655),
.B(n_220),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_548),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_550),
.Y(n_768)
);

A2O1A1Ixp33_ASAP7_75t_L g769 ( 
.A1(n_635),
.A2(n_463),
.B(n_488),
.C(n_217),
.Y(n_769)
);

INVxp33_ASAP7_75t_SL g770 ( 
.A(n_516),
.Y(n_770)
);

AND2x2_ASAP7_75t_L g771 ( 
.A(n_625),
.B(n_508),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_552),
.B(n_555),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_571),
.B(n_631),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_568),
.B(n_224),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_552),
.B(n_221),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_576),
.B(n_225),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_555),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_560),
.B(n_221),
.Y(n_778)
);

INVx3_ASAP7_75t_L g779 ( 
.A(n_567),
.Y(n_779)
);

HB1xp67_ASAP7_75t_L g780 ( 
.A(n_539),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_560),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_546),
.B(n_300),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_563),
.B(n_243),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_588),
.B(n_228),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_546),
.B(n_304),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_563),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_516),
.Y(n_787)
);

OAI22xp33_ASAP7_75t_L g788 ( 
.A1(n_610),
.A2(n_294),
.B1(n_321),
.B2(n_319),
.Y(n_788)
);

BUFx3_ASAP7_75t_L g789 ( 
.A(n_546),
.Y(n_789)
);

INVx2_ASAP7_75t_SL g790 ( 
.A(n_618),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_565),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_626),
.B(n_271),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_626),
.B(n_273),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_544),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_626),
.B(n_657),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_657),
.B(n_561),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_544),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_561),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_549),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_546),
.B(n_508),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_657),
.B(n_273),
.Y(n_801)
);

INVxp33_ASAP7_75t_SL g802 ( 
.A(n_547),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_562),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_646),
.B(n_229),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_619),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_619),
.Y(n_806)
);

BUFx3_ASAP7_75t_L g807 ( 
.A(n_647),
.Y(n_807)
);

AOI21xp5_ASAP7_75t_L g808 ( 
.A1(n_611),
.A2(n_451),
.B(n_448),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_623),
.Y(n_809)
);

NOR3xp33_ASAP7_75t_L g810 ( 
.A(n_610),
.B(n_277),
.C(n_284),
.Y(n_810)
);

INVxp67_ASAP7_75t_L g811 ( 
.A(n_577),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_617),
.B(n_632),
.Y(n_812)
);

BUFx5_ASAP7_75t_L g813 ( 
.A(n_513),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_623),
.B(n_307),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_L g815 ( 
.A(n_706),
.B(n_577),
.Y(n_815)
);

INVx2_ASAP7_75t_SL g816 ( 
.A(n_771),
.Y(n_816)
);

OR2x2_ASAP7_75t_L g817 ( 
.A(n_668),
.B(n_654),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_732),
.B(n_634),
.Y(n_818)
);

AOI22xp5_ASAP7_75t_L g819 ( 
.A1(n_700),
.A2(n_596),
.B1(n_527),
.B2(n_654),
.Y(n_819)
);

HB1xp67_ASAP7_75t_L g820 ( 
.A(n_670),
.Y(n_820)
);

INVxp67_ASAP7_75t_L g821 ( 
.A(n_780),
.Y(n_821)
);

INVx3_ASAP7_75t_L g822 ( 
.A(n_688),
.Y(n_822)
);

AOI22xp5_ASAP7_75t_L g823 ( 
.A1(n_700),
.A2(n_527),
.B1(n_651),
.B2(n_642),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_662),
.Y(n_824)
);

A2O1A1Ixp33_ASAP7_75t_L g825 ( 
.A1(n_784),
.A2(n_284),
.B(n_294),
.C(n_310),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_706),
.B(n_732),
.Y(n_826)
);

INVx3_ASAP7_75t_L g827 ( 
.A(n_688),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_813),
.B(n_624),
.Y(n_828)
);

OAI22xp5_ASAP7_75t_L g829 ( 
.A1(n_673),
.A2(n_656),
.B1(n_651),
.B2(n_642),
.Y(n_829)
);

BUFx6f_ASAP7_75t_L g830 ( 
.A(n_688),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_698),
.Y(n_831)
);

BUFx6f_ASAP7_75t_L g832 ( 
.A(n_688),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_663),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_693),
.Y(n_834)
);

INVx2_ASAP7_75t_SL g835 ( 
.A(n_670),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_753),
.B(n_618),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_708),
.Y(n_837)
);

INVx2_ASAP7_75t_SL g838 ( 
.A(n_670),
.Y(n_838)
);

AOI22xp33_ASAP7_75t_L g839 ( 
.A1(n_673),
.A2(n_746),
.B1(n_734),
.B2(n_692),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_659),
.B(n_519),
.Y(n_840)
);

OAI22xp5_ASAP7_75t_SL g841 ( 
.A1(n_802),
.A2(n_547),
.B1(n_328),
.B2(n_327),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_666),
.B(n_519),
.Y(n_842)
);

INVx2_ASAP7_75t_SL g843 ( 
.A(n_739),
.Y(n_843)
);

AOI22xp33_ASAP7_75t_L g844 ( 
.A1(n_734),
.A2(n_310),
.B1(n_319),
.B2(n_321),
.Y(n_844)
);

O2A1O1Ixp33_ASAP7_75t_L g845 ( 
.A1(n_692),
.A2(n_581),
.B(n_569),
.C(n_574),
.Y(n_845)
);

BUFx3_ASAP7_75t_L g846 ( 
.A(n_765),
.Y(n_846)
);

OAI21xp5_ASAP7_75t_L g847 ( 
.A1(n_658),
.A2(n_601),
.B(n_624),
.Y(n_847)
);

INVxp33_ASAP7_75t_L g848 ( 
.A(n_780),
.Y(n_848)
);

INVx3_ASAP7_75t_L g849 ( 
.A(n_709),
.Y(n_849)
);

OR2x6_ASAP7_75t_L g850 ( 
.A(n_685),
.B(n_592),
.Y(n_850)
);

INVx3_ASAP7_75t_L g851 ( 
.A(n_709),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_690),
.B(n_757),
.Y(n_852)
);

NOR2xp67_ASAP7_75t_L g853 ( 
.A(n_787),
.B(n_628),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_753),
.B(n_618),
.Y(n_854)
);

HB1xp67_ASAP7_75t_L g855 ( 
.A(n_741),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_690),
.B(n_520),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_741),
.B(n_618),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_723),
.Y(n_858)
);

OR2x6_ASAP7_75t_L g859 ( 
.A(n_685),
.B(n_592),
.Y(n_859)
);

AOI22xp5_ASAP7_75t_SL g860 ( 
.A1(n_784),
.A2(n_318),
.B1(n_230),
.B2(n_235),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_767),
.B(n_520),
.Y(n_861)
);

AOI22xp5_ASAP7_75t_L g862 ( 
.A1(n_773),
.A2(n_656),
.B1(n_641),
.B2(n_628),
.Y(n_862)
);

NOR2xp67_ASAP7_75t_L g863 ( 
.A(n_790),
.B(n_774),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_724),
.Y(n_864)
);

BUFx4f_ASAP7_75t_L g865 ( 
.A(n_685),
.Y(n_865)
);

INVx2_ASAP7_75t_SL g866 ( 
.A(n_703),
.Y(n_866)
);

INVx3_ASAP7_75t_L g867 ( 
.A(n_684),
.Y(n_867)
);

AOI22xp33_ASAP7_75t_SL g868 ( 
.A1(n_677),
.A2(n_259),
.B1(n_274),
.B2(n_332),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_SL g869 ( 
.A(n_813),
.B(n_637),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_736),
.Y(n_870)
);

AND2x4_ASAP7_75t_L g871 ( 
.A(n_717),
.B(n_404),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_749),
.Y(n_872)
);

NAND2x1_ASAP7_75t_L g873 ( 
.A(n_684),
.B(n_513),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_749),
.Y(n_874)
);

AOI22xp5_ASAP7_75t_L g875 ( 
.A1(n_812),
.A2(n_641),
.B1(n_637),
.B2(n_640),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_805),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_768),
.B(n_520),
.Y(n_877)
);

BUFx2_ASAP7_75t_L g878 ( 
.A(n_672),
.Y(n_878)
);

INVx3_ASAP7_75t_L g879 ( 
.A(n_725),
.Y(n_879)
);

CKINVDCx8_ASAP7_75t_R g880 ( 
.A(n_759),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_806),
.Y(n_881)
);

BUFx3_ASAP7_75t_L g882 ( 
.A(n_807),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_777),
.B(n_553),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_781),
.B(n_553),
.Y(n_884)
);

BUFx3_ASAP7_75t_L g885 ( 
.A(n_697),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_809),
.Y(n_886)
);

AOI22xp5_ASAP7_75t_L g887 ( 
.A1(n_691),
.A2(n_640),
.B1(n_557),
.B2(n_554),
.Y(n_887)
);

AOI22xp33_ASAP7_75t_L g888 ( 
.A1(n_746),
.A2(n_274),
.B1(n_259),
.B2(n_488),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_798),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_786),
.B(n_553),
.Y(n_890)
);

BUFx12f_ASAP7_75t_L g891 ( 
.A(n_683),
.Y(n_891)
);

BUFx3_ASAP7_75t_L g892 ( 
.A(n_697),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_SL g893 ( 
.A(n_800),
.B(n_308),
.Y(n_893)
);

INVx4_ASAP7_75t_L g894 ( 
.A(n_725),
.Y(n_894)
);

A2O1A1Ixp33_ASAP7_75t_L g895 ( 
.A1(n_691),
.A2(n_640),
.B(n_554),
.C(n_557),
.Y(n_895)
);

NAND3xp33_ASAP7_75t_SL g896 ( 
.A(n_774),
.B(n_315),
.C(n_311),
.Y(n_896)
);

NAND4xp25_ASAP7_75t_SL g897 ( 
.A(n_660),
.B(n_416),
.C(n_429),
.D(n_427),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_791),
.B(n_554),
.Y(n_898)
);

NOR2xp33_ASAP7_75t_SL g899 ( 
.A(n_770),
.B(n_197),
.Y(n_899)
);

NOR3xp33_ASAP7_75t_SL g900 ( 
.A(n_788),
.B(n_290),
.C(n_244),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_803),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_712),
.B(n_259),
.Y(n_902)
);

INVx3_ASAP7_75t_L g903 ( 
.A(n_779),
.Y(n_903)
);

AND2x4_ASAP7_75t_L g904 ( 
.A(n_738),
.B(n_404),
.Y(n_904)
);

AOI22xp33_ASAP7_75t_SL g905 ( 
.A1(n_776),
.A2(n_259),
.B1(n_274),
.B2(n_197),
.Y(n_905)
);

BUFx3_ASAP7_75t_L g906 ( 
.A(n_697),
.Y(n_906)
);

NOR2xp33_ASAP7_75t_L g907 ( 
.A(n_762),
.B(n_811),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_772),
.B(n_564),
.Y(n_908)
);

AND2x2_ASAP7_75t_L g909 ( 
.A(n_727),
.B(n_274),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_729),
.B(n_564),
.Y(n_910)
);

BUFx6f_ASAP7_75t_L g911 ( 
.A(n_779),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_L g912 ( 
.A(n_762),
.B(n_564),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_SL g913 ( 
.A(n_813),
.B(n_521),
.Y(n_913)
);

NOR2xp33_ASAP7_75t_L g914 ( 
.A(n_811),
.B(n_513),
.Y(n_914)
);

INVxp67_ASAP7_75t_SL g915 ( 
.A(n_713),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_716),
.Y(n_916)
);

AOI22xp5_ASAP7_75t_L g917 ( 
.A1(n_696),
.A2(n_758),
.B1(n_814),
.B2(n_751),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_679),
.B(n_406),
.Y(n_918)
);

AO22x1_ASAP7_75t_L g919 ( 
.A1(n_776),
.A2(n_287),
.B1(n_257),
.B2(n_261),
.Y(n_919)
);

AND2x4_ASAP7_75t_L g920 ( 
.A(n_789),
.B(n_406),
.Y(n_920)
);

INVx2_ASAP7_75t_SL g921 ( 
.A(n_681),
.Y(n_921)
);

NOR3xp33_ASAP7_75t_SL g922 ( 
.A(n_788),
.B(n_256),
.C(n_267),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_669),
.B(n_580),
.Y(n_923)
);

NOR2xp33_ASAP7_75t_L g924 ( 
.A(n_742),
.B(n_580),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_795),
.A2(n_580),
.B(n_629),
.Y(n_925)
);

AOI22xp33_ASAP7_75t_L g926 ( 
.A1(n_810),
.A2(n_578),
.B1(n_613),
.B2(n_609),
.Y(n_926)
);

AND2x4_ASAP7_75t_L g927 ( 
.A(n_707),
.B(n_412),
.Y(n_927)
);

AOI22xp33_ASAP7_75t_L g928 ( 
.A1(n_810),
.A2(n_578),
.B1(n_613),
.B2(n_609),
.Y(n_928)
);

NAND2x2_ASAP7_75t_L g929 ( 
.A(n_671),
.B(n_197),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_674),
.B(n_580),
.Y(n_930)
);

BUFx3_ASAP7_75t_L g931 ( 
.A(n_707),
.Y(n_931)
);

AND2x4_ASAP7_75t_L g932 ( 
.A(n_707),
.B(n_412),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_702),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_714),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_733),
.A2(n_711),
.B(n_710),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_728),
.B(n_629),
.Y(n_936)
);

OR2x6_ASAP7_75t_L g937 ( 
.A(n_766),
.B(n_782),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_664),
.B(n_629),
.Y(n_938)
);

HB1xp67_ASAP7_75t_L g939 ( 
.A(n_721),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_745),
.Y(n_940)
);

AND2x4_ASAP7_75t_L g941 ( 
.A(n_785),
.B(n_413),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_804),
.B(n_413),
.Y(n_942)
);

HB1xp67_ASAP7_75t_L g943 ( 
.A(n_726),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_748),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_SL g945 ( 
.A(n_813),
.B(n_521),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_750),
.Y(n_946)
);

INVxp67_ASAP7_75t_L g947 ( 
.A(n_804),
.Y(n_947)
);

NAND2x1_ASAP7_75t_L g948 ( 
.A(n_731),
.B(n_521),
.Y(n_948)
);

HB1xp67_ASAP7_75t_L g949 ( 
.A(n_715),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_660),
.B(n_416),
.Y(n_950)
);

INVx3_ASAP7_75t_L g951 ( 
.A(n_743),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_664),
.B(n_569),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_719),
.B(n_574),
.Y(n_953)
);

INVx2_ASAP7_75t_SL g954 ( 
.A(n_761),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_813),
.B(n_521),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_675),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_763),
.B(n_583),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_794),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_730),
.Y(n_959)
);

INVx1_ASAP7_75t_SL g960 ( 
.A(n_695),
.Y(n_960)
);

INVx4_ASAP7_75t_L g961 ( 
.A(n_733),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_752),
.Y(n_962)
);

BUFx2_ASAP7_75t_L g963 ( 
.A(n_792),
.Y(n_963)
);

OAI21xp33_ASAP7_75t_SL g964 ( 
.A1(n_718),
.A2(n_424),
.B(n_426),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_775),
.B(n_583),
.Y(n_965)
);

INVx1_ASAP7_75t_SL g966 ( 
.A(n_778),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_797),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_783),
.B(n_586),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_733),
.A2(n_699),
.B(n_694),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_754),
.Y(n_970)
);

BUFx2_ASAP7_75t_L g971 ( 
.A(n_793),
.Y(n_971)
);

AOI22xp33_ASAP7_75t_SL g972 ( 
.A1(n_661),
.A2(n_208),
.B1(n_276),
.B2(n_341),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_756),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_704),
.B(n_590),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_SL g975 ( 
.A(n_733),
.B(n_309),
.Y(n_975)
);

AND2x4_ASAP7_75t_L g976 ( 
.A(n_755),
.B(n_417),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_796),
.B(n_590),
.Y(n_977)
);

BUFx8_ASAP7_75t_L g978 ( 
.A(n_799),
.Y(n_978)
);

AND2x4_ASAP7_75t_L g979 ( 
.A(n_676),
.B(n_417),
.Y(n_979)
);

O2A1O1Ixp33_ASAP7_75t_L g980 ( 
.A1(n_740),
.A2(n_602),
.B(n_607),
.C(n_594),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_760),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_737),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_744),
.Y(n_983)
);

BUFx4f_ASAP7_75t_L g984 ( 
.A(n_680),
.Y(n_984)
);

BUFx6f_ASAP7_75t_L g985 ( 
.A(n_678),
.Y(n_985)
);

OR2x6_ASAP7_75t_L g986 ( 
.A(n_682),
.B(n_420),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_705),
.Y(n_987)
);

AND2x4_ASAP7_75t_L g988 ( 
.A(n_686),
.B(n_420),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_701),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_701),
.Y(n_990)
);

NOR2x2_ASAP7_75t_L g991 ( 
.A(n_722),
.B(n_208),
.Y(n_991)
);

CKINVDCx16_ASAP7_75t_R g992 ( 
.A(n_846),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_916),
.B(n_687),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_915),
.B(n_801),
.Y(n_994)
);

OAI22xp5_ASAP7_75t_L g995 ( 
.A1(n_839),
.A2(n_769),
.B1(n_720),
.B2(n_718),
.Y(n_995)
);

NOR3xp33_ASAP7_75t_L g996 ( 
.A(n_896),
.B(n_747),
.C(n_720),
.Y(n_996)
);

AND2x4_ASAP7_75t_L g997 ( 
.A(n_835),
.B(n_735),
.Y(n_997)
);

A2O1A1Ixp33_ASAP7_75t_L g998 ( 
.A1(n_984),
.A2(n_808),
.B(n_764),
.C(n_689),
.Y(n_998)
);

BUFx2_ASAP7_75t_R g999 ( 
.A(n_880),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_915),
.B(n_665),
.Y(n_1000)
);

BUFx6f_ASAP7_75t_L g1001 ( 
.A(n_830),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_833),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_834),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_L g1004 ( 
.A(n_826),
.B(n_735),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_923),
.A2(n_930),
.B(n_840),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_858),
.Y(n_1006)
);

OAI22xp5_ASAP7_75t_L g1007 ( 
.A1(n_839),
.A2(n_667),
.B1(n_270),
.B2(n_322),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_842),
.A2(n_665),
.B(n_585),
.Y(n_1008)
);

AND2x2_ASAP7_75t_L g1009 ( 
.A(n_878),
.B(n_422),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_913),
.A2(n_665),
.B(n_585),
.Y(n_1010)
);

A2O1A1Ixp33_ASAP7_75t_SL g1011 ( 
.A1(n_826),
.A2(n_595),
.B(n_599),
.C(n_594),
.Y(n_1011)
);

INVx3_ASAP7_75t_L g1012 ( 
.A(n_830),
.Y(n_1012)
);

AO32x2_ASAP7_75t_L g1013 ( 
.A1(n_829),
.A2(n_954),
.A3(n_894),
.B1(n_838),
.B2(n_866),
.Y(n_1013)
);

NAND2xp33_ASAP7_75t_SL g1014 ( 
.A(n_956),
.B(n_667),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_945),
.A2(n_665),
.B(n_636),
.Y(n_1015)
);

OAI21xp33_ASAP7_75t_L g1016 ( 
.A1(n_899),
.A2(n_334),
.B(n_338),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_945),
.A2(n_636),
.B(n_535),
.Y(n_1017)
);

OAI21x1_ASAP7_75t_L g1018 ( 
.A1(n_925),
.A2(n_602),
.B(n_606),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_864),
.Y(n_1019)
);

INVx2_ASAP7_75t_SL g1020 ( 
.A(n_843),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_942),
.B(n_599),
.Y(n_1021)
);

AOI21x1_ASAP7_75t_L g1022 ( 
.A1(n_935),
.A2(n_549),
.B(n_606),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_L g1023 ( 
.A(n_947),
.B(n_278),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_SL g1024 ( 
.A(n_947),
.B(n_312),
.Y(n_1024)
);

NAND2xp33_ASAP7_75t_L g1025 ( 
.A(n_852),
.B(n_342),
.Y(n_1025)
);

CKINVDCx11_ASAP7_75t_R g1026 ( 
.A(n_891),
.Y(n_1026)
);

HB1xp67_ASAP7_75t_L g1027 ( 
.A(n_821),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_966),
.B(n_604),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_955),
.A2(n_636),
.B(n_585),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_870),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_955),
.A2(n_636),
.B(n_585),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_939),
.B(n_604),
.Y(n_1032)
);

AND2x4_ASAP7_75t_L g1033 ( 
.A(n_853),
.B(n_872),
.Y(n_1033)
);

AND2x2_ASAP7_75t_L g1034 ( 
.A(n_918),
.B(n_424),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_856),
.A2(n_575),
.B(n_535),
.Y(n_1035)
);

A2O1A1Ixp33_ASAP7_75t_SL g1036 ( 
.A1(n_936),
.A2(n_605),
.B(n_431),
.C(n_426),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_935),
.A2(n_575),
.B(n_535),
.Y(n_1037)
);

AND2x2_ASAP7_75t_L g1038 ( 
.A(n_902),
.B(n_427),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_L g1039 ( 
.A(n_815),
.B(n_323),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_939),
.B(n_605),
.Y(n_1040)
);

NOR2xp33_ASAP7_75t_L g1041 ( 
.A(n_815),
.B(n_336),
.Y(n_1041)
);

NOR2xp33_ASAP7_75t_L g1042 ( 
.A(n_848),
.B(n_337),
.Y(n_1042)
);

INVx2_ASAP7_75t_SL g1043 ( 
.A(n_921),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_943),
.B(n_535),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_943),
.B(n_575),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_949),
.B(n_575),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_949),
.B(n_431),
.Y(n_1047)
);

NAND3xp33_ASAP7_75t_L g1048 ( 
.A(n_905),
.B(n_429),
.C(n_388),
.Y(n_1048)
);

NOR2xp33_ASAP7_75t_R g1049 ( 
.A(n_865),
.B(n_75),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_SL g1050 ( 
.A(n_819),
.B(n_208),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_837),
.Y(n_1051)
);

O2A1O1Ixp33_ASAP7_75t_L g1052 ( 
.A1(n_896),
.A2(n_388),
.B(n_393),
.C(n_394),
.Y(n_1052)
);

BUFx4f_ASAP7_75t_L g1053 ( 
.A(n_850),
.Y(n_1053)
);

AND2x2_ASAP7_75t_L g1054 ( 
.A(n_909),
.B(n_393),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_961),
.A2(n_528),
.B(n_451),
.Y(n_1055)
);

BUFx4f_ASAP7_75t_SL g1056 ( 
.A(n_885),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_824),
.Y(n_1057)
);

A2O1A1Ixp33_ASAP7_75t_L g1058 ( 
.A1(n_984),
.A2(n_394),
.B(n_451),
.C(n_448),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_SL g1059 ( 
.A(n_863),
.B(n_528),
.Y(n_1059)
);

AOI221x1_ASAP7_75t_L g1060 ( 
.A1(n_825),
.A2(n_454),
.B1(n_448),
.B2(n_439),
.C(n_435),
.Y(n_1060)
);

NOR2xp33_ASAP7_75t_L g1061 ( 
.A(n_817),
.B(n_1),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_982),
.B(n_528),
.Y(n_1062)
);

NOR2xp33_ASAP7_75t_L g1063 ( 
.A(n_821),
.B(n_818),
.Y(n_1063)
);

OAI22xp5_ASAP7_75t_L g1064 ( 
.A1(n_844),
.A2(n_454),
.B1(n_528),
.B2(n_448),
.Y(n_1064)
);

OAI22xp5_ASAP7_75t_SL g1065 ( 
.A1(n_905),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_983),
.B(n_987),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_979),
.B(n_454),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_963),
.B(n_971),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_SL g1069 ( 
.A(n_857),
.B(n_172),
.Y(n_1069)
);

INVx1_ASAP7_75t_SL g1070 ( 
.A(n_855),
.Y(n_1070)
);

INVx3_ASAP7_75t_L g1071 ( 
.A(n_830),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_950),
.B(n_5),
.Y(n_1072)
);

BUFx6f_ASAP7_75t_L g1073 ( 
.A(n_830),
.Y(n_1073)
);

BUFx2_ASAP7_75t_L g1074 ( 
.A(n_882),
.Y(n_1074)
);

OAI22xp5_ASAP7_75t_L g1075 ( 
.A1(n_844),
.A2(n_447),
.B1(n_9),
.B2(n_10),
.Y(n_1075)
);

AND2x2_ASAP7_75t_L g1076 ( 
.A(n_855),
.B(n_8),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_914),
.B(n_8),
.Y(n_1077)
);

AND3x2_ASAP7_75t_L g1078 ( 
.A(n_836),
.B(n_11),
.C(n_12),
.Y(n_1078)
);

BUFx3_ASAP7_75t_L g1079 ( 
.A(n_978),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_889),
.Y(n_1080)
);

CKINVDCx20_ASAP7_75t_R g1081 ( 
.A(n_892),
.Y(n_1081)
);

NOR3xp33_ASAP7_75t_SL g1082 ( 
.A(n_959),
.B(n_14),
.C(n_15),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_SL g1083 ( 
.A(n_874),
.B(n_71),
.Y(n_1083)
);

CKINVDCx11_ASAP7_75t_R g1084 ( 
.A(n_850),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_849),
.A2(n_447),
.B(n_67),
.Y(n_1085)
);

AO31x2_ASAP7_75t_L g1086 ( 
.A1(n_895),
.A2(n_15),
.A3(n_18),
.B(n_23),
.Y(n_1086)
);

AND2x2_ASAP7_75t_L g1087 ( 
.A(n_907),
.B(n_23),
.Y(n_1087)
);

A2O1A1Ixp33_ASAP7_75t_L g1088 ( 
.A1(n_917),
.A2(n_24),
.B(n_25),
.C(n_27),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_SL g1089 ( 
.A(n_941),
.B(n_96),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_901),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_849),
.A2(n_447),
.B(n_100),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_914),
.B(n_25),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_SL g1093 ( 
.A(n_941),
.B(n_102),
.Y(n_1093)
);

OR2x2_ASAP7_75t_SL g1094 ( 
.A(n_991),
.B(n_29),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_906),
.Y(n_1095)
);

AND2x2_ASAP7_75t_L g1096 ( 
.A(n_907),
.B(n_31),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_876),
.Y(n_1097)
);

AOI22xp33_ASAP7_75t_L g1098 ( 
.A1(n_976),
.A2(n_447),
.B1(n_35),
.B2(n_36),
.Y(n_1098)
);

NOR2xp33_ASAP7_75t_R g1099 ( 
.A(n_865),
.B(n_110),
.Y(n_1099)
);

BUFx3_ASAP7_75t_L g1100 ( 
.A(n_978),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_881),
.Y(n_1101)
);

O2A1O1Ixp5_ASAP7_75t_L g1102 ( 
.A1(n_936),
.A2(n_109),
.B(n_162),
.C(n_153),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_SL g1103 ( 
.A(n_960),
.B(n_92),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_851),
.A2(n_908),
.B(n_953),
.Y(n_1104)
);

CKINVDCx8_ASAP7_75t_R g1105 ( 
.A(n_850),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_851),
.A2(n_85),
.B(n_148),
.Y(n_1106)
);

INVxp33_ASAP7_75t_L g1107 ( 
.A(n_820),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_886),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_859),
.Y(n_1109)
);

BUFx2_ASAP7_75t_L g1110 ( 
.A(n_820),
.Y(n_1110)
);

BUFx6f_ASAP7_75t_L g1111 ( 
.A(n_832),
.Y(n_1111)
);

NAND3xp33_ASAP7_75t_SL g1112 ( 
.A(n_868),
.B(n_32),
.C(n_38),
.Y(n_1112)
);

NAND2x1p5_ASAP7_75t_L g1113 ( 
.A(n_832),
.B(n_111),
.Y(n_1113)
);

A2O1A1Ixp33_ASAP7_75t_L g1114 ( 
.A1(n_924),
.A2(n_32),
.B(n_42),
.C(n_48),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_979),
.B(n_116),
.Y(n_1115)
);

AOI22xp5_ASAP7_75t_L g1116 ( 
.A1(n_893),
.A2(n_163),
.B1(n_138),
.B2(n_128),
.Y(n_1116)
);

A2O1A1Ixp33_ASAP7_75t_L g1117 ( 
.A1(n_924),
.A2(n_42),
.B(n_48),
.C(n_50),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_988),
.B(n_126),
.Y(n_1118)
);

OAI22xp5_ASAP7_75t_SL g1119 ( 
.A1(n_841),
.A2(n_868),
.B1(n_937),
.B2(n_972),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_969),
.A2(n_50),
.B(n_55),
.Y(n_1120)
);

BUFx3_ASAP7_75t_L g1121 ( 
.A(n_931),
.Y(n_1121)
);

OR2x6_ASAP7_75t_L g1122 ( 
.A(n_859),
.B(n_55),
.Y(n_1122)
);

INVx4_ASAP7_75t_L g1123 ( 
.A(n_832),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_SL g1124 ( 
.A(n_836),
.B(n_57),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_969),
.A2(n_57),
.B(n_873),
.Y(n_1125)
);

NOR2xp33_ASAP7_75t_L g1126 ( 
.A(n_854),
.B(n_860),
.Y(n_1126)
);

NOR2xp33_ASAP7_75t_L g1127 ( 
.A(n_854),
.B(n_920),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_962),
.B(n_970),
.Y(n_1128)
);

NAND3xp33_ASAP7_75t_SL g1129 ( 
.A(n_972),
.B(n_900),
.C(n_922),
.Y(n_1129)
);

OR2x6_ASAP7_75t_L g1130 ( 
.A(n_859),
.B(n_937),
.Y(n_1130)
);

NAND2x1p5_ASAP7_75t_L g1131 ( 
.A(n_832),
.B(n_822),
.Y(n_1131)
);

OAI21x1_ASAP7_75t_L g1132 ( 
.A1(n_925),
.A2(n_980),
.B(n_847),
.Y(n_1132)
);

INVx1_ASAP7_75t_SL g1133 ( 
.A(n_920),
.Y(n_1133)
);

NOR3xp33_ASAP7_75t_L g1134 ( 
.A(n_919),
.B(n_897),
.C(n_927),
.Y(n_1134)
);

INVxp67_ASAP7_75t_L g1135 ( 
.A(n_927),
.Y(n_1135)
);

AO31x2_ASAP7_75t_L g1136 ( 
.A1(n_1060),
.A2(n_952),
.A3(n_938),
.B(n_912),
.Y(n_1136)
);

AOI221x1_ASAP7_75t_L g1137 ( 
.A1(n_1129),
.A2(n_946),
.B1(n_944),
.B2(n_940),
.C(n_973),
.Y(n_1137)
);

AOI21xp33_ASAP7_75t_L g1138 ( 
.A1(n_1039),
.A2(n_823),
.B(n_981),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_999),
.Y(n_1139)
);

INVx2_ASAP7_75t_SL g1140 ( 
.A(n_1074),
.Y(n_1140)
);

INVx2_ASAP7_75t_L g1141 ( 
.A(n_1003),
.Y(n_1141)
);

AO21x2_ASAP7_75t_L g1142 ( 
.A1(n_1132),
.A2(n_996),
.B(n_1036),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_1000),
.A2(n_957),
.B(n_968),
.Y(n_1143)
);

BUFx3_ASAP7_75t_L g1144 ( 
.A(n_1056),
.Y(n_1144)
);

AOI21x1_ASAP7_75t_L g1145 ( 
.A1(n_1005),
.A2(n_1104),
.B(n_1035),
.Y(n_1145)
);

CKINVDCx6p67_ASAP7_75t_R g1146 ( 
.A(n_1079),
.Y(n_1146)
);

OAI21x1_ASAP7_75t_L g1147 ( 
.A1(n_1010),
.A2(n_869),
.B(n_828),
.Y(n_1147)
);

OAI21x1_ASAP7_75t_L g1148 ( 
.A1(n_1015),
.A2(n_869),
.B(n_948),
.Y(n_1148)
);

AOI221xp5_ASAP7_75t_L g1149 ( 
.A1(n_1065),
.A2(n_1041),
.B1(n_1119),
.B2(n_1126),
.C(n_1112),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1006),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_994),
.A2(n_998),
.B(n_1008),
.Y(n_1151)
);

AO31x2_ASAP7_75t_L g1152 ( 
.A1(n_995),
.A2(n_965),
.A3(n_974),
.B(n_989),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_993),
.A2(n_977),
.B(n_910),
.Y(n_1153)
);

OAI21xp33_ASAP7_75t_SL g1154 ( 
.A1(n_1066),
.A2(n_990),
.B(n_888),
.Y(n_1154)
);

OAI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_995),
.A2(n_862),
.B(n_875),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1019),
.Y(n_1156)
);

AO31x2_ASAP7_75t_L g1157 ( 
.A1(n_1058),
.A2(n_898),
.A3(n_890),
.B(n_861),
.Y(n_1157)
);

INVx3_ASAP7_75t_L g1158 ( 
.A(n_1123),
.Y(n_1158)
);

OAI21x1_ASAP7_75t_L g1159 ( 
.A1(n_1017),
.A2(n_877),
.B(n_884),
.Y(n_1159)
);

OAI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_1004),
.A2(n_845),
.B(n_887),
.Y(n_1160)
);

OAI21x1_ASAP7_75t_L g1161 ( 
.A1(n_1029),
.A2(n_883),
.B(n_845),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_1030),
.Y(n_1162)
);

OAI21x1_ASAP7_75t_L g1163 ( 
.A1(n_1031),
.A2(n_879),
.B(n_903),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_1066),
.B(n_904),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_993),
.A2(n_1021),
.B(n_1128),
.Y(n_1165)
);

BUFx4_ASAP7_75t_SL g1166 ( 
.A(n_1081),
.Y(n_1166)
);

NOR2xp33_ASAP7_75t_SL g1167 ( 
.A(n_1105),
.B(n_937),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_1128),
.A2(n_975),
.B(n_867),
.Y(n_1168)
);

BUFx4f_ASAP7_75t_L g1169 ( 
.A(n_1130),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1063),
.B(n_1034),
.Y(n_1170)
);

BUFx6f_ASAP7_75t_L g1171 ( 
.A(n_1001),
.Y(n_1171)
);

O2A1O1Ixp33_ASAP7_75t_L g1172 ( 
.A1(n_1088),
.A2(n_900),
.B(n_922),
.C(n_964),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1032),
.B(n_871),
.Y(n_1173)
);

HB1xp67_ASAP7_75t_L g1174 ( 
.A(n_1070),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1032),
.B(n_871),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_SL g1176 ( 
.A(n_1068),
.B(n_932),
.Y(n_1176)
);

OAI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_1102),
.A2(n_928),
.B(n_926),
.Y(n_1177)
);

INVx2_ASAP7_75t_SL g1178 ( 
.A(n_1121),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_SL g1179 ( 
.A1(n_1115),
.A2(n_911),
.B(n_986),
.Y(n_1179)
);

AOI21x1_ASAP7_75t_L g1180 ( 
.A1(n_1125),
.A2(n_831),
.B(n_986),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1038),
.B(n_985),
.Y(n_1181)
);

AOI211x1_ASAP7_75t_L g1182 ( 
.A1(n_1072),
.A2(n_976),
.B(n_929),
.C(n_932),
.Y(n_1182)
);

OAI21xp33_ASAP7_75t_L g1183 ( 
.A1(n_1061),
.A2(n_888),
.B(n_933),
.Y(n_1183)
);

O2A1O1Ixp33_ASAP7_75t_SL g1184 ( 
.A1(n_1115),
.A2(n_934),
.B(n_967),
.C(n_958),
.Y(n_1184)
);

NAND3xp33_ASAP7_75t_L g1185 ( 
.A(n_1023),
.B(n_985),
.C(n_926),
.Y(n_1185)
);

BUFx3_ASAP7_75t_L g1186 ( 
.A(n_1110),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1080),
.Y(n_1187)
);

OAI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1077),
.A2(n_928),
.B(n_951),
.Y(n_1188)
);

AO31x2_ASAP7_75t_L g1189 ( 
.A1(n_1092),
.A2(n_985),
.A3(n_911),
.B(n_827),
.Y(n_1189)
);

OAI22xp5_ASAP7_75t_L g1190 ( 
.A1(n_1098),
.A2(n_1075),
.B1(n_1090),
.B2(n_1048),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_SL g1191 ( 
.A(n_1127),
.B(n_1133),
.Y(n_1191)
);

AO31x2_ASAP7_75t_L g1192 ( 
.A1(n_1114),
.A2(n_1117),
.A3(n_1120),
.B(n_1007),
.Y(n_1192)
);

A2O1A1Ixp33_ASAP7_75t_L g1193 ( 
.A1(n_1014),
.A2(n_1134),
.B(n_1118),
.C(n_1096),
.Y(n_1193)
);

OA21x2_ASAP7_75t_L g1194 ( 
.A1(n_1062),
.A2(n_1085),
.B(n_1091),
.Y(n_1194)
);

AO31x2_ASAP7_75t_L g1195 ( 
.A1(n_1007),
.A2(n_1118),
.A3(n_1064),
.B(n_1062),
.Y(n_1195)
);

INVx3_ASAP7_75t_L g1196 ( 
.A(n_1123),
.Y(n_1196)
);

O2A1O1Ixp5_ASAP7_75t_L g1197 ( 
.A1(n_1050),
.A2(n_1059),
.B(n_1124),
.C(n_1069),
.Y(n_1197)
);

INVx3_ASAP7_75t_L g1198 ( 
.A(n_1001),
.Y(n_1198)
);

OAI21x1_ASAP7_75t_L g1199 ( 
.A1(n_1055),
.A2(n_1067),
.B(n_1044),
.Y(n_1199)
);

AOI21x1_ASAP7_75t_L g1200 ( 
.A1(n_1040),
.A2(n_1044),
.B(n_1045),
.Y(n_1200)
);

INVx3_ASAP7_75t_L g1201 ( 
.A(n_1001),
.Y(n_1201)
);

AND2x4_ASAP7_75t_L g1202 ( 
.A(n_1033),
.B(n_1135),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_SL g1203 ( 
.A(n_1033),
.B(n_992),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_1095),
.Y(n_1204)
);

OAI21x1_ASAP7_75t_L g1205 ( 
.A1(n_1067),
.A2(n_1106),
.B(n_1046),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1051),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1047),
.B(n_1054),
.Y(n_1207)
);

BUFx6f_ASAP7_75t_L g1208 ( 
.A(n_1073),
.Y(n_1208)
);

AOI22xp5_ASAP7_75t_L g1209 ( 
.A1(n_1042),
.A2(n_1089),
.B1(n_1093),
.B2(n_1025),
.Y(n_1209)
);

AOI21x1_ASAP7_75t_L g1210 ( 
.A1(n_1024),
.A2(n_1083),
.B(n_1103),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1011),
.A2(n_1028),
.B(n_1108),
.Y(n_1211)
);

A2O1A1Ixp33_ASAP7_75t_L g1212 ( 
.A1(n_1087),
.A2(n_1016),
.B(n_1116),
.C(n_997),
.Y(n_1212)
);

AO31x2_ASAP7_75t_L g1213 ( 
.A1(n_1064),
.A2(n_1075),
.A3(n_1013),
.B(n_1101),
.Y(n_1213)
);

INVx2_ASAP7_75t_SL g1214 ( 
.A(n_1027),
.Y(n_1214)
);

AOI21xp5_ASAP7_75t_SL g1215 ( 
.A1(n_1113),
.A2(n_1111),
.B(n_1073),
.Y(n_1215)
);

BUFx2_ASAP7_75t_L g1216 ( 
.A(n_1009),
.Y(n_1216)
);

INVxp67_ASAP7_75t_SL g1217 ( 
.A(n_1073),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1097),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_997),
.A2(n_1131),
.B(n_1057),
.Y(n_1219)
);

AO21x2_ASAP7_75t_L g1220 ( 
.A1(n_1013),
.A2(n_1052),
.B(n_1099),
.Y(n_1220)
);

OAI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1113),
.A2(n_1076),
.B(n_1131),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1012),
.B(n_1071),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1012),
.B(n_1071),
.Y(n_1223)
);

BUFx2_ASAP7_75t_L g1224 ( 
.A(n_1020),
.Y(n_1224)
);

INVx4_ASAP7_75t_L g1225 ( 
.A(n_1111),
.Y(n_1225)
);

OAI21x1_ASAP7_75t_L g1226 ( 
.A1(n_1013),
.A2(n_1111),
.B(n_1086),
.Y(n_1226)
);

NOR2xp33_ASAP7_75t_L g1227 ( 
.A(n_1107),
.B(n_1043),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1086),
.B(n_1082),
.Y(n_1228)
);

OA21x2_ASAP7_75t_L g1229 ( 
.A1(n_1086),
.A2(n_1109),
.B(n_1078),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1053),
.A2(n_1130),
.B(n_1049),
.Y(n_1230)
);

OR2x2_ASAP7_75t_L g1231 ( 
.A(n_1130),
.B(n_1094),
.Y(n_1231)
);

OAI21x1_ASAP7_75t_L g1232 ( 
.A1(n_1053),
.A2(n_1084),
.B(n_1122),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_1026),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1122),
.B(n_1100),
.Y(n_1234)
);

AOI22xp33_ASAP7_75t_L g1235 ( 
.A1(n_1122),
.A2(n_1129),
.B1(n_984),
.B2(n_1119),
.Y(n_1235)
);

OAI22xp5_ASAP7_75t_L g1236 ( 
.A1(n_1066),
.A2(n_839),
.B1(n_844),
.B2(n_950),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_SL g1237 ( 
.A(n_1068),
.B(n_759),
.Y(n_1237)
);

A2O1A1Ixp33_ASAP7_75t_L g1238 ( 
.A1(n_1126),
.A2(n_947),
.B(n_984),
.C(n_691),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1066),
.B(n_916),
.Y(n_1239)
);

BUFx4_ASAP7_75t_SL g1240 ( 
.A(n_1081),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1066),
.B(n_916),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1002),
.Y(n_1242)
);

AO31x2_ASAP7_75t_L g1243 ( 
.A1(n_1060),
.A2(n_995),
.A3(n_998),
.B(n_895),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1066),
.B(n_916),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1000),
.A2(n_1005),
.B(n_733),
.Y(n_1245)
);

CKINVDCx5p33_ASAP7_75t_R g1246 ( 
.A(n_999),
.Y(n_1246)
);

NOR2xp33_ASAP7_75t_L g1247 ( 
.A(n_1063),
.B(n_706),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1002),
.Y(n_1248)
);

OAI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1005),
.A2(n_995),
.B(n_998),
.Y(n_1249)
);

AO31x2_ASAP7_75t_L g1250 ( 
.A1(n_1060),
.A2(n_995),
.A3(n_998),
.B(n_895),
.Y(n_1250)
);

INVx3_ASAP7_75t_L g1251 ( 
.A(n_1123),
.Y(n_1251)
);

BUFx6f_ASAP7_75t_L g1252 ( 
.A(n_1001),
.Y(n_1252)
);

AND2x4_ASAP7_75t_L g1253 ( 
.A(n_1033),
.B(n_1135),
.Y(n_1253)
);

INVx3_ASAP7_75t_L g1254 ( 
.A(n_1123),
.Y(n_1254)
);

INVx3_ASAP7_75t_L g1255 ( 
.A(n_1123),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1018),
.A2(n_1022),
.B(n_1037),
.Y(n_1256)
);

OAI22xp33_ASAP7_75t_L g1257 ( 
.A1(n_1126),
.A2(n_677),
.B1(n_438),
.B2(n_622),
.Y(n_1257)
);

OAI21x1_ASAP7_75t_L g1258 ( 
.A1(n_1018),
.A2(n_1022),
.B(n_1037),
.Y(n_1258)
);

OAI21x1_ASAP7_75t_L g1259 ( 
.A1(n_1018),
.A2(n_1022),
.B(n_1037),
.Y(n_1259)
);

BUFx6f_ASAP7_75t_L g1260 ( 
.A(n_1001),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1066),
.B(n_916),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1066),
.B(n_916),
.Y(n_1262)
);

AOI21xp33_ASAP7_75t_L g1263 ( 
.A1(n_1039),
.A2(n_1041),
.B(n_1126),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1066),
.B(n_916),
.Y(n_1264)
);

INVx5_ASAP7_75t_L g1265 ( 
.A(n_1001),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1066),
.B(n_916),
.Y(n_1266)
);

AND2x2_ASAP7_75t_L g1267 ( 
.A(n_1038),
.B(n_816),
.Y(n_1267)
);

BUFx2_ASAP7_75t_L g1268 ( 
.A(n_1074),
.Y(n_1268)
);

OAI21x1_ASAP7_75t_L g1269 ( 
.A1(n_1018),
.A2(n_1022),
.B(n_1037),
.Y(n_1269)
);

A2O1A1Ixp33_ASAP7_75t_L g1270 ( 
.A1(n_1126),
.A2(n_947),
.B(n_984),
.C(n_691),
.Y(n_1270)
);

INVx2_ASAP7_75t_L g1271 ( 
.A(n_1002),
.Y(n_1271)
);

NOR2xp33_ASAP7_75t_R g1272 ( 
.A(n_1081),
.B(n_787),
.Y(n_1272)
);

OR2x2_ASAP7_75t_L g1273 ( 
.A(n_1068),
.B(n_817),
.Y(n_1273)
);

AND2x2_ASAP7_75t_L g1274 ( 
.A(n_1038),
.B(n_816),
.Y(n_1274)
);

OAI22xp5_ASAP7_75t_L g1275 ( 
.A1(n_1066),
.A2(n_839),
.B1(n_844),
.B2(n_950),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1066),
.B(n_916),
.Y(n_1276)
);

AND2x4_ASAP7_75t_L g1277 ( 
.A(n_1033),
.B(n_1135),
.Y(n_1277)
);

AOI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1000),
.A2(n_1005),
.B(n_994),
.Y(n_1278)
);

OA21x2_ASAP7_75t_L g1279 ( 
.A1(n_1249),
.A2(n_1151),
.B(n_1256),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_1272),
.Y(n_1280)
);

NAND2x1p5_ASAP7_75t_L g1281 ( 
.A(n_1169),
.B(n_1265),
.Y(n_1281)
);

OAI21x1_ASAP7_75t_SL g1282 ( 
.A1(n_1210),
.A2(n_1221),
.B(n_1165),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1162),
.Y(n_1283)
);

OAI21x1_ASAP7_75t_L g1284 ( 
.A1(n_1258),
.A2(n_1269),
.B(n_1259),
.Y(n_1284)
);

BUFx6f_ASAP7_75t_L g1285 ( 
.A(n_1265),
.Y(n_1285)
);

AND2x4_ASAP7_75t_L g1286 ( 
.A(n_1230),
.B(n_1181),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1271),
.Y(n_1287)
);

OR2x2_ASAP7_75t_L g1288 ( 
.A(n_1170),
.B(n_1273),
.Y(n_1288)
);

INVx2_ASAP7_75t_SL g1289 ( 
.A(n_1166),
.Y(n_1289)
);

INVx4_ASAP7_75t_L g1290 ( 
.A(n_1265),
.Y(n_1290)
);

OAI21x1_ASAP7_75t_L g1291 ( 
.A1(n_1145),
.A2(n_1159),
.B(n_1148),
.Y(n_1291)
);

OAI21x1_ASAP7_75t_L g1292 ( 
.A1(n_1180),
.A2(n_1161),
.B(n_1199),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_1240),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_1139),
.Y(n_1294)
);

BUFx2_ASAP7_75t_L g1295 ( 
.A(n_1268),
.Y(n_1295)
);

OAI21x1_ASAP7_75t_L g1296 ( 
.A1(n_1205),
.A2(n_1147),
.B(n_1163),
.Y(n_1296)
);

BUFx3_ASAP7_75t_L g1297 ( 
.A(n_1144),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1150),
.Y(n_1298)
);

BUFx6f_ASAP7_75t_L g1299 ( 
.A(n_1265),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_1156),
.Y(n_1300)
);

NAND2x1p5_ASAP7_75t_L g1301 ( 
.A(n_1169),
.B(n_1203),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1247),
.B(n_1170),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1187),
.Y(n_1303)
);

OAI21x1_ASAP7_75t_L g1304 ( 
.A1(n_1143),
.A2(n_1153),
.B(n_1155),
.Y(n_1304)
);

OAI21x1_ASAP7_75t_L g1305 ( 
.A1(n_1226),
.A2(n_1155),
.B(n_1200),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_1246),
.Y(n_1306)
);

CKINVDCx5p33_ASAP7_75t_R g1307 ( 
.A(n_1204),
.Y(n_1307)
);

OAI22xp5_ASAP7_75t_SL g1308 ( 
.A1(n_1235),
.A2(n_1231),
.B1(n_1234),
.B2(n_1182),
.Y(n_1308)
);

AOI22xp33_ASAP7_75t_L g1309 ( 
.A1(n_1149),
.A2(n_1263),
.B1(n_1257),
.B2(n_1190),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_1233),
.Y(n_1310)
);

OAI21x1_ASAP7_75t_L g1311 ( 
.A1(n_1211),
.A2(n_1194),
.B(n_1177),
.Y(n_1311)
);

OA21x2_ASAP7_75t_L g1312 ( 
.A1(n_1137),
.A2(n_1177),
.B(n_1160),
.Y(n_1312)
);

INVx2_ASAP7_75t_L g1313 ( 
.A(n_1242),
.Y(n_1313)
);

AO31x2_ASAP7_75t_L g1314 ( 
.A1(n_1228),
.A2(n_1193),
.A3(n_1236),
.B(n_1275),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_1248),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1206),
.Y(n_1316)
);

AOI21x1_ASAP7_75t_L g1317 ( 
.A1(n_1228),
.A2(n_1160),
.B(n_1168),
.Y(n_1317)
);

OAI21x1_ASAP7_75t_L g1318 ( 
.A1(n_1194),
.A2(n_1221),
.B(n_1188),
.Y(n_1318)
);

OAI21x1_ASAP7_75t_L g1319 ( 
.A1(n_1188),
.A2(n_1219),
.B(n_1197),
.Y(n_1319)
);

INVxp67_ASAP7_75t_L g1320 ( 
.A(n_1174),
.Y(n_1320)
);

OR2x2_ASAP7_75t_L g1321 ( 
.A(n_1216),
.B(n_1207),
.Y(n_1321)
);

OR2x2_ASAP7_75t_L g1322 ( 
.A(n_1207),
.B(n_1164),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1218),
.Y(n_1323)
);

AO31x2_ASAP7_75t_L g1324 ( 
.A1(n_1236),
.A2(n_1275),
.A3(n_1190),
.B(n_1238),
.Y(n_1324)
);

BUFx4f_ASAP7_75t_L g1325 ( 
.A(n_1146),
.Y(n_1325)
);

BUFx2_ASAP7_75t_R g1326 ( 
.A(n_1234),
.Y(n_1326)
);

OAI21x1_ASAP7_75t_L g1327 ( 
.A1(n_1219),
.A2(n_1179),
.B(n_1172),
.Y(n_1327)
);

AO21x2_ASAP7_75t_L g1328 ( 
.A1(n_1142),
.A2(n_1220),
.B(n_1138),
.Y(n_1328)
);

OA21x2_ASAP7_75t_L g1329 ( 
.A1(n_1138),
.A2(n_1185),
.B(n_1183),
.Y(n_1329)
);

OAI21x1_ASAP7_75t_L g1330 ( 
.A1(n_1222),
.A2(n_1223),
.B(n_1215),
.Y(n_1330)
);

OR2x2_ASAP7_75t_L g1331 ( 
.A(n_1164),
.B(n_1237),
.Y(n_1331)
);

OAI21x1_ASAP7_75t_L g1332 ( 
.A1(n_1222),
.A2(n_1223),
.B(n_1181),
.Y(n_1332)
);

INVx2_ASAP7_75t_SL g1333 ( 
.A(n_1178),
.Y(n_1333)
);

AOI221x1_ASAP7_75t_L g1334 ( 
.A1(n_1263),
.A2(n_1270),
.B1(n_1212),
.B2(n_1264),
.C(n_1261),
.Y(n_1334)
);

OAI21x1_ASAP7_75t_L g1335 ( 
.A1(n_1173),
.A2(n_1175),
.B(n_1232),
.Y(n_1335)
);

OAI21x1_ASAP7_75t_L g1336 ( 
.A1(n_1173),
.A2(n_1175),
.B(n_1229),
.Y(n_1336)
);

OA21x2_ASAP7_75t_L g1337 ( 
.A1(n_1239),
.A2(n_1264),
.B(n_1276),
.Y(n_1337)
);

OAI21xp5_ASAP7_75t_L g1338 ( 
.A1(n_1149),
.A2(n_1154),
.B(n_1209),
.Y(n_1338)
);

AOI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1239),
.A2(n_1266),
.B(n_1276),
.Y(n_1339)
);

OAI21xp5_ASAP7_75t_L g1340 ( 
.A1(n_1241),
.A2(n_1244),
.B(n_1261),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_1241),
.Y(n_1341)
);

OAI21x1_ASAP7_75t_SL g1342 ( 
.A1(n_1244),
.A2(n_1262),
.B(n_1266),
.Y(n_1342)
);

AOI21xp5_ASAP7_75t_L g1343 ( 
.A1(n_1262),
.A2(n_1184),
.B(n_1142),
.Y(n_1343)
);

CKINVDCx16_ASAP7_75t_R g1344 ( 
.A(n_1186),
.Y(n_1344)
);

OAI21x1_ASAP7_75t_L g1345 ( 
.A1(n_1229),
.A2(n_1254),
.B(n_1251),
.Y(n_1345)
);

OAI21x1_ASAP7_75t_L g1346 ( 
.A1(n_1158),
.A2(n_1255),
.B(n_1254),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1189),
.Y(n_1347)
);

OAI21x1_ASAP7_75t_L g1348 ( 
.A1(n_1158),
.A2(n_1255),
.B(n_1251),
.Y(n_1348)
);

OAI22xp5_ASAP7_75t_L g1349 ( 
.A1(n_1191),
.A2(n_1214),
.B1(n_1176),
.B2(n_1253),
.Y(n_1349)
);

AOI22xp33_ASAP7_75t_L g1350 ( 
.A1(n_1167),
.A2(n_1267),
.B1(n_1274),
.B2(n_1202),
.Y(n_1350)
);

AO21x2_ASAP7_75t_L g1351 ( 
.A1(n_1152),
.A2(n_1250),
.B(n_1243),
.Y(n_1351)
);

INVx5_ASAP7_75t_L g1352 ( 
.A(n_1171),
.Y(n_1352)
);

INVx6_ASAP7_75t_L g1353 ( 
.A(n_1225),
.Y(n_1353)
);

OAI21x1_ASAP7_75t_L g1354 ( 
.A1(n_1196),
.A2(n_1198),
.B(n_1201),
.Y(n_1354)
);

BUFx2_ASAP7_75t_L g1355 ( 
.A(n_1224),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1202),
.B(n_1277),
.Y(n_1356)
);

OR2x2_ASAP7_75t_L g1357 ( 
.A(n_1253),
.B(n_1277),
.Y(n_1357)
);

AND2x4_ASAP7_75t_L g1358 ( 
.A(n_1198),
.B(n_1201),
.Y(n_1358)
);

NOR2xp33_ASAP7_75t_L g1359 ( 
.A(n_1167),
.B(n_1227),
.Y(n_1359)
);

OR2x6_ASAP7_75t_L g1360 ( 
.A(n_1140),
.B(n_1196),
.Y(n_1360)
);

CKINVDCx16_ASAP7_75t_R g1361 ( 
.A(n_1225),
.Y(n_1361)
);

OAI21x1_ASAP7_75t_L g1362 ( 
.A1(n_1243),
.A2(n_1250),
.B(n_1217),
.Y(n_1362)
);

BUFx10_ASAP7_75t_L g1363 ( 
.A(n_1171),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1189),
.Y(n_1364)
);

OA21x2_ASAP7_75t_L g1365 ( 
.A1(n_1243),
.A2(n_1250),
.B(n_1152),
.Y(n_1365)
);

OR2x2_ASAP7_75t_L g1366 ( 
.A(n_1171),
.B(n_1208),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1260),
.Y(n_1367)
);

BUFx8_ASAP7_75t_L g1368 ( 
.A(n_1208),
.Y(n_1368)
);

OAI21x1_ASAP7_75t_L g1369 ( 
.A1(n_1157),
.A2(n_1195),
.B(n_1192),
.Y(n_1369)
);

OAI21x1_ASAP7_75t_L g1370 ( 
.A1(n_1157),
.A2(n_1195),
.B(n_1136),
.Y(n_1370)
);

INVx8_ASAP7_75t_L g1371 ( 
.A(n_1252),
.Y(n_1371)
);

AOI22xp33_ASAP7_75t_L g1372 ( 
.A1(n_1192),
.A2(n_1213),
.B1(n_1136),
.B2(n_1157),
.Y(n_1372)
);

INVx3_ASAP7_75t_L g1373 ( 
.A(n_1213),
.Y(n_1373)
);

OR2x2_ASAP7_75t_L g1374 ( 
.A(n_1213),
.B(n_1136),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1247),
.B(n_1170),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1247),
.B(n_1170),
.Y(n_1376)
);

OAI21x1_ASAP7_75t_L g1377 ( 
.A1(n_1256),
.A2(n_1259),
.B(n_1258),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1141),
.Y(n_1378)
);

AOI22xp33_ASAP7_75t_SL g1379 ( 
.A1(n_1236),
.A2(n_438),
.B1(n_1065),
.B2(n_622),
.Y(n_1379)
);

A2O1A1Ixp33_ASAP7_75t_L g1380 ( 
.A1(n_1149),
.A2(n_839),
.B(n_1263),
.C(n_1249),
.Y(n_1380)
);

AOI22xp33_ASAP7_75t_L g1381 ( 
.A1(n_1149),
.A2(n_1263),
.B1(n_1065),
.B2(n_905),
.Y(n_1381)
);

AOI21xp5_ASAP7_75t_L g1382 ( 
.A1(n_1249),
.A2(n_1000),
.B(n_1278),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1141),
.Y(n_1383)
);

CKINVDCx5p33_ASAP7_75t_R g1384 ( 
.A(n_1272),
.Y(n_1384)
);

INVx3_ASAP7_75t_L g1385 ( 
.A(n_1158),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1247),
.B(n_1170),
.Y(n_1386)
);

OAI21xp5_ASAP7_75t_L g1387 ( 
.A1(n_1263),
.A2(n_947),
.B(n_706),
.Y(n_1387)
);

NOR2xp33_ASAP7_75t_SL g1388 ( 
.A(n_1139),
.B(n_770),
.Y(n_1388)
);

OAI21x1_ASAP7_75t_L g1389 ( 
.A1(n_1256),
.A2(n_1259),
.B(n_1258),
.Y(n_1389)
);

OR2x6_ASAP7_75t_L g1390 ( 
.A(n_1179),
.B(n_1230),
.Y(n_1390)
);

INVx3_ASAP7_75t_L g1391 ( 
.A(n_1158),
.Y(n_1391)
);

AOI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1180),
.A2(n_1022),
.B(n_1245),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1141),
.Y(n_1393)
);

AOI21xp5_ASAP7_75t_L g1394 ( 
.A1(n_1249),
.A2(n_1000),
.B(n_1278),
.Y(n_1394)
);

AO31x2_ASAP7_75t_L g1395 ( 
.A1(n_1137),
.A2(n_1151),
.A3(n_1060),
.B(n_1278),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1267),
.B(n_1274),
.Y(n_1396)
);

INVxp67_ASAP7_75t_SL g1397 ( 
.A(n_1278),
.Y(n_1397)
);

AOI22xp33_ASAP7_75t_SL g1398 ( 
.A1(n_1236),
.A2(n_438),
.B1(n_1065),
.B2(n_622),
.Y(n_1398)
);

AO21x1_ASAP7_75t_L g1399 ( 
.A1(n_1263),
.A2(n_1228),
.B(n_1092),
.Y(n_1399)
);

AO21x1_ASAP7_75t_L g1400 ( 
.A1(n_1263),
.A2(n_1228),
.B(n_1092),
.Y(n_1400)
);

AOI22xp33_ASAP7_75t_L g1401 ( 
.A1(n_1149),
.A2(n_1263),
.B1(n_1065),
.B2(n_905),
.Y(n_1401)
);

INVx2_ASAP7_75t_L g1402 ( 
.A(n_1141),
.Y(n_1402)
);

BUFx2_ASAP7_75t_L g1403 ( 
.A(n_1268),
.Y(n_1403)
);

INVx4_ASAP7_75t_SL g1404 ( 
.A(n_1192),
.Y(n_1404)
);

NAND3xp33_ASAP7_75t_L g1405 ( 
.A(n_1263),
.B(n_1149),
.C(n_1238),
.Y(n_1405)
);

AOI21xp33_ASAP7_75t_L g1406 ( 
.A1(n_1263),
.A2(n_691),
.B(n_1039),
.Y(n_1406)
);

NAND2x1p5_ASAP7_75t_L g1407 ( 
.A(n_1169),
.B(n_1265),
.Y(n_1407)
);

AOI22xp33_ASAP7_75t_L g1408 ( 
.A1(n_1149),
.A2(n_1263),
.B1(n_1065),
.B2(n_905),
.Y(n_1408)
);

AOI21xp5_ASAP7_75t_L g1409 ( 
.A1(n_1397),
.A2(n_1394),
.B(n_1382),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1396),
.B(n_1288),
.Y(n_1410)
);

OR2x6_ASAP7_75t_L g1411 ( 
.A(n_1390),
.B(n_1327),
.Y(n_1411)
);

OA21x2_ASAP7_75t_L g1412 ( 
.A1(n_1311),
.A2(n_1343),
.B(n_1305),
.Y(n_1412)
);

OR2x2_ASAP7_75t_L g1413 ( 
.A(n_1321),
.B(n_1331),
.Y(n_1413)
);

AOI21xp5_ASAP7_75t_SL g1414 ( 
.A1(n_1380),
.A2(n_1339),
.B(n_1337),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1341),
.B(n_1337),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1350),
.B(n_1387),
.Y(n_1416)
);

AOI21x1_ASAP7_75t_SL g1417 ( 
.A1(n_1302),
.A2(n_1376),
.B(n_1375),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1350),
.B(n_1357),
.Y(n_1418)
);

OR2x2_ASAP7_75t_L g1419 ( 
.A(n_1322),
.B(n_1300),
.Y(n_1419)
);

CKINVDCx12_ASAP7_75t_R g1420 ( 
.A(n_1366),
.Y(n_1420)
);

OR2x2_ASAP7_75t_L g1421 ( 
.A(n_1313),
.B(n_1315),
.Y(n_1421)
);

OA21x2_ASAP7_75t_L g1422 ( 
.A1(n_1292),
.A2(n_1369),
.B(n_1318),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1359),
.B(n_1356),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1359),
.B(n_1386),
.Y(n_1424)
);

NAND2x1p5_ASAP7_75t_L g1425 ( 
.A(n_1337),
.B(n_1345),
.Y(n_1425)
);

NAND2x1_ASAP7_75t_L g1426 ( 
.A(n_1390),
.B(n_1342),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1298),
.Y(n_1427)
);

BUFx3_ASAP7_75t_L g1428 ( 
.A(n_1297),
.Y(n_1428)
);

NOR2xp67_ASAP7_75t_L g1429 ( 
.A(n_1280),
.B(n_1384),
.Y(n_1429)
);

OA21x2_ASAP7_75t_L g1430 ( 
.A1(n_1370),
.A2(n_1319),
.B(n_1304),
.Y(n_1430)
);

OAI22xp5_ASAP7_75t_L g1431 ( 
.A1(n_1381),
.A2(n_1408),
.B1(n_1401),
.B2(n_1398),
.Y(n_1431)
);

A2O1A1Ixp33_ASAP7_75t_L g1432 ( 
.A1(n_1406),
.A2(n_1405),
.B(n_1380),
.C(n_1401),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1402),
.B(n_1309),
.Y(n_1433)
);

A2O1A1Ixp33_ASAP7_75t_L g1434 ( 
.A1(n_1381),
.A2(n_1408),
.B(n_1338),
.C(n_1309),
.Y(n_1434)
);

INVx1_ASAP7_75t_SL g1435 ( 
.A(n_1295),
.Y(n_1435)
);

CKINVDCx20_ASAP7_75t_R g1436 ( 
.A(n_1293),
.Y(n_1436)
);

INVxp33_ASAP7_75t_L g1437 ( 
.A(n_1388),
.Y(n_1437)
);

AND2x4_ASAP7_75t_L g1438 ( 
.A(n_1286),
.B(n_1358),
.Y(n_1438)
);

O2A1O1Ixp33_ASAP7_75t_L g1439 ( 
.A1(n_1349),
.A2(n_1320),
.B(n_1400),
.C(n_1399),
.Y(n_1439)
);

O2A1O1Ixp33_ASAP7_75t_L g1440 ( 
.A1(n_1320),
.A2(n_1340),
.B(n_1301),
.C(n_1282),
.Y(n_1440)
);

A2O1A1Ixp33_ASAP7_75t_L g1441 ( 
.A1(n_1379),
.A2(n_1398),
.B(n_1335),
.C(n_1336),
.Y(n_1441)
);

AOI221xp5_ASAP7_75t_L g1442 ( 
.A1(n_1379),
.A2(n_1308),
.B1(n_1341),
.B2(n_1372),
.C(n_1303),
.Y(n_1442)
);

O2A1O1Ixp33_ASAP7_75t_L g1443 ( 
.A1(n_1301),
.A2(n_1333),
.B(n_1316),
.C(n_1403),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1283),
.B(n_1287),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1323),
.Y(n_1445)
);

AOI21xp5_ASAP7_75t_SL g1446 ( 
.A1(n_1334),
.A2(n_1285),
.B(n_1299),
.Y(n_1446)
);

CKINVDCx5p33_ASAP7_75t_R g1447 ( 
.A(n_1307),
.Y(n_1447)
);

O2A1O1Ixp5_ASAP7_75t_L g1448 ( 
.A1(n_1317),
.A2(n_1364),
.B(n_1392),
.C(n_1347),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1314),
.B(n_1324),
.Y(n_1449)
);

AND2x2_ASAP7_75t_SL g1450 ( 
.A(n_1325),
.B(n_1312),
.Y(n_1450)
);

CKINVDCx5p33_ASAP7_75t_R g1451 ( 
.A(n_1307),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1314),
.B(n_1324),
.Y(n_1452)
);

O2A1O1Ixp33_ASAP7_75t_L g1453 ( 
.A1(n_1355),
.A2(n_1393),
.B(n_1383),
.C(n_1378),
.Y(n_1453)
);

OAI22xp5_ASAP7_75t_L g1454 ( 
.A1(n_1312),
.A2(n_1326),
.B1(n_1344),
.B2(n_1360),
.Y(n_1454)
);

O2A1O1Ixp33_ASAP7_75t_L g1455 ( 
.A1(n_1360),
.A2(n_1407),
.B(n_1281),
.C(n_1390),
.Y(n_1455)
);

AND2x4_ASAP7_75t_L g1456 ( 
.A(n_1360),
.B(n_1385),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1314),
.B(n_1324),
.Y(n_1457)
);

OR2x2_ASAP7_75t_L g1458 ( 
.A(n_1324),
.B(n_1314),
.Y(n_1458)
);

O2A1O1Ixp5_ASAP7_75t_L g1459 ( 
.A1(n_1347),
.A2(n_1373),
.B(n_1290),
.C(n_1374),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1312),
.B(n_1332),
.Y(n_1460)
);

AND2x4_ASAP7_75t_L g1461 ( 
.A(n_1385),
.B(n_1391),
.Y(n_1461)
);

OA21x2_ASAP7_75t_L g1462 ( 
.A1(n_1291),
.A2(n_1389),
.B(n_1296),
.Y(n_1462)
);

OAI22xp5_ASAP7_75t_SL g1463 ( 
.A1(n_1280),
.A2(n_1384),
.B1(n_1293),
.B2(n_1294),
.Y(n_1463)
);

INVxp67_ASAP7_75t_L g1464 ( 
.A(n_1367),
.Y(n_1464)
);

BUFx3_ASAP7_75t_L g1465 ( 
.A(n_1297),
.Y(n_1465)
);

OAI22xp5_ASAP7_75t_L g1466 ( 
.A1(n_1281),
.A2(n_1407),
.B1(n_1372),
.B2(n_1329),
.Y(n_1466)
);

INVx3_ASAP7_75t_L g1467 ( 
.A(n_1285),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1329),
.B(n_1351),
.Y(n_1468)
);

CKINVDCx20_ASAP7_75t_R g1469 ( 
.A(n_1310),
.Y(n_1469)
);

OR2x2_ASAP7_75t_L g1470 ( 
.A(n_1329),
.B(n_1289),
.Y(n_1470)
);

OR2x2_ASAP7_75t_L g1471 ( 
.A(n_1351),
.B(n_1361),
.Y(n_1471)
);

OAI22xp5_ASAP7_75t_L g1472 ( 
.A1(n_1352),
.A2(n_1299),
.B1(n_1285),
.B2(n_1353),
.Y(n_1472)
);

OAI22xp5_ASAP7_75t_L g1473 ( 
.A1(n_1352),
.A2(n_1299),
.B1(n_1353),
.B2(n_1365),
.Y(n_1473)
);

BUFx3_ASAP7_75t_L g1474 ( 
.A(n_1368),
.Y(n_1474)
);

OAI22xp5_ASAP7_75t_L g1475 ( 
.A1(n_1352),
.A2(n_1299),
.B1(n_1353),
.B2(n_1365),
.Y(n_1475)
);

NOR2xp67_ASAP7_75t_L g1476 ( 
.A(n_1310),
.B(n_1306),
.Y(n_1476)
);

BUFx3_ASAP7_75t_L g1477 ( 
.A(n_1368),
.Y(n_1477)
);

NOR2xp67_ASAP7_75t_L g1478 ( 
.A(n_1294),
.B(n_1306),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1404),
.B(n_1365),
.Y(n_1479)
);

O2A1O1Ixp33_ASAP7_75t_L g1480 ( 
.A1(n_1328),
.A2(n_1279),
.B(n_1404),
.C(n_1395),
.Y(n_1480)
);

OAI22xp5_ASAP7_75t_L g1481 ( 
.A1(n_1352),
.A2(n_1290),
.B1(n_1371),
.B2(n_1395),
.Y(n_1481)
);

A2O1A1Ixp33_ASAP7_75t_SL g1482 ( 
.A1(n_1404),
.A2(n_1330),
.B(n_1395),
.C(n_1362),
.Y(n_1482)
);

OAI22xp5_ASAP7_75t_L g1483 ( 
.A1(n_1371),
.A2(n_1395),
.B1(n_1368),
.B2(n_1363),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1354),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1346),
.Y(n_1485)
);

O2A1O1Ixp5_ASAP7_75t_L g1486 ( 
.A1(n_1348),
.A2(n_1263),
.B(n_1406),
.C(n_1338),
.Y(n_1486)
);

BUFx8_ASAP7_75t_L g1487 ( 
.A(n_1284),
.Y(n_1487)
);

NOR2xp67_ASAP7_75t_L g1488 ( 
.A(n_1377),
.B(n_1280),
.Y(n_1488)
);

OAI22xp5_ASAP7_75t_L g1489 ( 
.A1(n_1381),
.A2(n_839),
.B1(n_1408),
.B2(n_1401),
.Y(n_1489)
);

AOI21xp5_ASAP7_75t_L g1490 ( 
.A1(n_1397),
.A2(n_1249),
.B(n_1382),
.Y(n_1490)
);

O2A1O1Ixp5_ASAP7_75t_L g1491 ( 
.A1(n_1406),
.A2(n_1263),
.B(n_1338),
.C(n_1399),
.Y(n_1491)
);

OA21x2_ASAP7_75t_L g1492 ( 
.A1(n_1311),
.A2(n_1343),
.B(n_1305),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1396),
.B(n_1288),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1341),
.B(n_1337),
.Y(n_1494)
);

OAI211xp5_ASAP7_75t_L g1495 ( 
.A1(n_1408),
.A2(n_1263),
.B(n_905),
.C(n_1381),
.Y(n_1495)
);

BUFx6f_ASAP7_75t_L g1496 ( 
.A(n_1285),
.Y(n_1496)
);

AOI21xp5_ASAP7_75t_SL g1497 ( 
.A1(n_1380),
.A2(n_1275),
.B(n_1236),
.Y(n_1497)
);

NOR2xp67_ASAP7_75t_L g1498 ( 
.A(n_1280),
.B(n_1384),
.Y(n_1498)
);

OR2x2_ASAP7_75t_L g1499 ( 
.A(n_1288),
.B(n_1321),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1341),
.B(n_1337),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1396),
.B(n_1288),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1396),
.B(n_1288),
.Y(n_1502)
);

HB1xp67_ASAP7_75t_L g1503 ( 
.A(n_1321),
.Y(n_1503)
);

INVxp67_ASAP7_75t_L g1504 ( 
.A(n_1396),
.Y(n_1504)
);

INVx1_ASAP7_75t_SL g1505 ( 
.A(n_1321),
.Y(n_1505)
);

O2A1O1Ixp33_ASAP7_75t_L g1506 ( 
.A1(n_1406),
.A2(n_1263),
.B(n_1270),
.C(n_1238),
.Y(n_1506)
);

A2O1A1Ixp33_ASAP7_75t_L g1507 ( 
.A1(n_1406),
.A2(n_1263),
.B(n_1149),
.C(n_1126),
.Y(n_1507)
);

AOI21xp5_ASAP7_75t_SL g1508 ( 
.A1(n_1380),
.A2(n_1275),
.B(n_1236),
.Y(n_1508)
);

INVx3_ASAP7_75t_L g1509 ( 
.A(n_1358),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1415),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1438),
.B(n_1458),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1415),
.Y(n_1512)
);

INVx4_ASAP7_75t_SL g1513 ( 
.A(n_1411),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1438),
.B(n_1449),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1505),
.B(n_1503),
.Y(n_1515)
);

AOI221xp5_ASAP7_75t_L g1516 ( 
.A1(n_1431),
.A2(n_1507),
.B1(n_1489),
.B2(n_1495),
.C(n_1434),
.Y(n_1516)
);

OR2x2_ASAP7_75t_L g1517 ( 
.A(n_1494),
.B(n_1500),
.Y(n_1517)
);

INVx3_ASAP7_75t_L g1518 ( 
.A(n_1422),
.Y(n_1518)
);

OR2x2_ASAP7_75t_L g1519 ( 
.A(n_1494),
.B(n_1500),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1449),
.B(n_1452),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1452),
.B(n_1457),
.Y(n_1521)
);

BUFx2_ASAP7_75t_L g1522 ( 
.A(n_1487),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1484),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1457),
.B(n_1427),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1505),
.B(n_1499),
.Y(n_1525)
);

OR2x6_ASAP7_75t_L g1526 ( 
.A(n_1414),
.B(n_1411),
.Y(n_1526)
);

HB1xp67_ASAP7_75t_L g1527 ( 
.A(n_1419),
.Y(n_1527)
);

HB1xp67_ASAP7_75t_L g1528 ( 
.A(n_1470),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1445),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1424),
.B(n_1413),
.Y(n_1530)
);

INVx3_ASAP7_75t_L g1531 ( 
.A(n_1422),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1421),
.Y(n_1532)
);

BUFx3_ASAP7_75t_L g1533 ( 
.A(n_1487),
.Y(n_1533)
);

INVxp67_ASAP7_75t_SL g1534 ( 
.A(n_1453),
.Y(n_1534)
);

OR2x6_ASAP7_75t_L g1535 ( 
.A(n_1490),
.B(n_1409),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1423),
.B(n_1416),
.Y(n_1536)
);

OR2x6_ASAP7_75t_L g1537 ( 
.A(n_1455),
.B(n_1426),
.Y(n_1537)
);

OR2x2_ASAP7_75t_L g1538 ( 
.A(n_1460),
.B(n_1468),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1485),
.Y(n_1539)
);

OR2x2_ASAP7_75t_L g1540 ( 
.A(n_1460),
.B(n_1468),
.Y(n_1540)
);

AO21x2_ASAP7_75t_L g1541 ( 
.A1(n_1482),
.A2(n_1480),
.B(n_1441),
.Y(n_1541)
);

AND2x4_ASAP7_75t_L g1542 ( 
.A(n_1479),
.B(n_1509),
.Y(n_1542)
);

BUFx2_ASAP7_75t_L g1543 ( 
.A(n_1471),
.Y(n_1543)
);

INVx2_ASAP7_75t_SL g1544 ( 
.A(n_1456),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1418),
.B(n_1410),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1479),
.Y(n_1546)
);

AOI22xp33_ASAP7_75t_L g1547 ( 
.A1(n_1431),
.A2(n_1489),
.B1(n_1442),
.B2(n_1450),
.Y(n_1547)
);

OR2x2_ASAP7_75t_L g1548 ( 
.A(n_1425),
.B(n_1430),
.Y(n_1548)
);

AND2x4_ASAP7_75t_L g1549 ( 
.A(n_1509),
.B(n_1488),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_SL g1550 ( 
.A(n_1443),
.B(n_1432),
.Y(n_1550)
);

AOI21xp5_ASAP7_75t_L g1551 ( 
.A1(n_1497),
.A2(n_1508),
.B(n_1506),
.Y(n_1551)
);

HB1xp67_ASAP7_75t_L g1552 ( 
.A(n_1435),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1462),
.Y(n_1553)
);

HB1xp67_ASAP7_75t_L g1554 ( 
.A(n_1435),
.Y(n_1554)
);

BUFx6f_ASAP7_75t_SL g1555 ( 
.A(n_1474),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1493),
.B(n_1502),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1459),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1412),
.Y(n_1558)
);

OR2x6_ASAP7_75t_L g1559 ( 
.A(n_1466),
.B(n_1446),
.Y(n_1559)
);

OR2x2_ASAP7_75t_L g1560 ( 
.A(n_1466),
.B(n_1454),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1448),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1501),
.B(n_1433),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1444),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1492),
.Y(n_1564)
);

BUFx3_ASAP7_75t_L g1565 ( 
.A(n_1428),
.Y(n_1565)
);

OR2x2_ASAP7_75t_L g1566 ( 
.A(n_1454),
.B(n_1504),
.Y(n_1566)
);

HB1xp67_ASAP7_75t_L g1567 ( 
.A(n_1528),
.Y(n_1567)
);

NAND3xp33_ASAP7_75t_L g1568 ( 
.A(n_1516),
.B(n_1491),
.C(n_1442),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1535),
.B(n_1486),
.Y(n_1569)
);

OAI22xp5_ASAP7_75t_L g1570 ( 
.A1(n_1547),
.A2(n_1439),
.B1(n_1472),
.B2(n_1464),
.Y(n_1570)
);

NOR2x1_ASAP7_75t_L g1571 ( 
.A(n_1526),
.B(n_1473),
.Y(n_1571)
);

INVxp67_ASAP7_75t_SL g1572 ( 
.A(n_1523),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1535),
.B(n_1475),
.Y(n_1573)
);

HB1xp67_ASAP7_75t_L g1574 ( 
.A(n_1512),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1535),
.B(n_1481),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1535),
.B(n_1483),
.Y(n_1576)
);

NOR2x1_ASAP7_75t_L g1577 ( 
.A(n_1526),
.B(n_1440),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1512),
.B(n_1461),
.Y(n_1578)
);

AND2x4_ASAP7_75t_L g1579 ( 
.A(n_1513),
.B(n_1461),
.Y(n_1579)
);

OAI211xp5_ASAP7_75t_SL g1580 ( 
.A1(n_1551),
.A2(n_1417),
.B(n_1472),
.C(n_1467),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1553),
.B(n_1465),
.Y(n_1581)
);

BUFx2_ASAP7_75t_L g1582 ( 
.A(n_1548),
.Y(n_1582)
);

BUFx3_ASAP7_75t_L g1583 ( 
.A(n_1533),
.Y(n_1583)
);

HB1xp67_ASAP7_75t_L g1584 ( 
.A(n_1510),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_1518),
.Y(n_1585)
);

OR2x2_ASAP7_75t_L g1586 ( 
.A(n_1538),
.B(n_1496),
.Y(n_1586)
);

OAI22xp5_ASAP7_75t_L g1587 ( 
.A1(n_1550),
.A2(n_1534),
.B1(n_1559),
.B2(n_1560),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1531),
.B(n_1496),
.Y(n_1588)
);

NOR2x1p5_ASAP7_75t_L g1589 ( 
.A(n_1533),
.B(n_1477),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1539),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1531),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1539),
.Y(n_1592)
);

INVx1_ASAP7_75t_SL g1593 ( 
.A(n_1517),
.Y(n_1593)
);

BUFx2_ASAP7_75t_L g1594 ( 
.A(n_1583),
.Y(n_1594)
);

OAI221xp5_ASAP7_75t_L g1595 ( 
.A1(n_1568),
.A2(n_1559),
.B1(n_1522),
.B2(n_1526),
.C(n_1560),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1590),
.Y(n_1596)
);

NAND4xp25_ASAP7_75t_L g1597 ( 
.A(n_1568),
.B(n_1515),
.C(n_1557),
.D(n_1566),
.Y(n_1597)
);

OAI211xp5_ASAP7_75t_L g1598 ( 
.A1(n_1568),
.A2(n_1566),
.B(n_1557),
.C(n_1552),
.Y(n_1598)
);

OAI22xp5_ASAP7_75t_L g1599 ( 
.A1(n_1587),
.A2(n_1559),
.B1(n_1522),
.B2(n_1533),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1590),
.Y(n_1600)
);

A2O1A1Ixp33_ASAP7_75t_L g1601 ( 
.A1(n_1587),
.A2(n_1437),
.B(n_1554),
.C(n_1536),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1593),
.B(n_1543),
.Y(n_1602)
);

AOI22xp33_ASAP7_75t_L g1603 ( 
.A1(n_1570),
.A2(n_1559),
.B1(n_1525),
.B2(n_1526),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1593),
.B(n_1543),
.Y(n_1604)
);

AOI21xp5_ASAP7_75t_L g1605 ( 
.A1(n_1587),
.A2(n_1537),
.B(n_1541),
.Y(n_1605)
);

NAND2x1_ASAP7_75t_L g1606 ( 
.A(n_1577),
.B(n_1537),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1582),
.B(n_1514),
.Y(n_1607)
);

CKINVDCx16_ASAP7_75t_R g1608 ( 
.A(n_1583),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_SL g1609 ( 
.A(n_1577),
.B(n_1549),
.Y(n_1609)
);

AOI222xp33_ASAP7_75t_L g1610 ( 
.A1(n_1570),
.A2(n_1530),
.B1(n_1545),
.B2(n_1556),
.C1(n_1521),
.C2(n_1520),
.Y(n_1610)
);

AOI33xp33_ASAP7_75t_L g1611 ( 
.A1(n_1569),
.A2(n_1561),
.A3(n_1546),
.B1(n_1510),
.B2(n_1529),
.B3(n_1563),
.Y(n_1611)
);

OAI221xp5_ASAP7_75t_SL g1612 ( 
.A1(n_1569),
.A2(n_1537),
.B1(n_1561),
.B2(n_1545),
.C(n_1517),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1590),
.Y(n_1613)
);

BUFx6f_ASAP7_75t_L g1614 ( 
.A(n_1583),
.Y(n_1614)
);

HB1xp67_ASAP7_75t_L g1615 ( 
.A(n_1567),
.Y(n_1615)
);

OR2x2_ASAP7_75t_L g1616 ( 
.A(n_1567),
.B(n_1519),
.Y(n_1616)
);

OAI221xp5_ASAP7_75t_L g1617 ( 
.A1(n_1577),
.A2(n_1537),
.B1(n_1544),
.B2(n_1565),
.C(n_1546),
.Y(n_1617)
);

OAI211xp5_ASAP7_75t_L g1618 ( 
.A1(n_1570),
.A2(n_1540),
.B(n_1538),
.C(n_1529),
.Y(n_1618)
);

AOI221xp5_ASAP7_75t_L g1619 ( 
.A1(n_1569),
.A2(n_1556),
.B1(n_1562),
.B2(n_1532),
.C(n_1524),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1592),
.Y(n_1620)
);

OAI22xp5_ASAP7_75t_L g1621 ( 
.A1(n_1583),
.A2(n_1537),
.B1(n_1565),
.B2(n_1544),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1592),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1592),
.Y(n_1623)
);

OR2x2_ASAP7_75t_L g1624 ( 
.A(n_1582),
.B(n_1540),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1584),
.Y(n_1625)
);

OR2x2_ASAP7_75t_L g1626 ( 
.A(n_1582),
.B(n_1527),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1584),
.Y(n_1627)
);

BUFx2_ASAP7_75t_L g1628 ( 
.A(n_1583),
.Y(n_1628)
);

AND2x4_ASAP7_75t_L g1629 ( 
.A(n_1579),
.B(n_1513),
.Y(n_1629)
);

AOI22xp5_ASAP7_75t_L g1630 ( 
.A1(n_1580),
.A2(n_1555),
.B1(n_1511),
.B2(n_1514),
.Y(n_1630)
);

OA21x2_ASAP7_75t_L g1631 ( 
.A1(n_1585),
.A2(n_1558),
.B(n_1564),
.Y(n_1631)
);

INVxp67_ASAP7_75t_SL g1632 ( 
.A(n_1574),
.Y(n_1632)
);

AOI22xp5_ASAP7_75t_L g1633 ( 
.A1(n_1580),
.A2(n_1555),
.B1(n_1511),
.B2(n_1420),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1578),
.B(n_1542),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1596),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1631),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1610),
.B(n_1578),
.Y(n_1637)
);

INVx1_ASAP7_75t_SL g1638 ( 
.A(n_1626),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1600),
.Y(n_1639)
);

INVx2_ASAP7_75t_L g1640 ( 
.A(n_1631),
.Y(n_1640)
);

HB1xp67_ASAP7_75t_L g1641 ( 
.A(n_1615),
.Y(n_1641)
);

INVx1_ASAP7_75t_SL g1642 ( 
.A(n_1626),
.Y(n_1642)
);

INVx4_ASAP7_75t_SL g1643 ( 
.A(n_1614),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1613),
.Y(n_1644)
);

NOR2xp33_ASAP7_75t_L g1645 ( 
.A(n_1597),
.B(n_1555),
.Y(n_1645)
);

HB1xp67_ASAP7_75t_L g1646 ( 
.A(n_1602),
.Y(n_1646)
);

BUFx2_ASAP7_75t_L g1647 ( 
.A(n_1629),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1619),
.B(n_1578),
.Y(n_1648)
);

INVx2_ASAP7_75t_SL g1649 ( 
.A(n_1614),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1620),
.Y(n_1650)
);

INVx4_ASAP7_75t_L g1651 ( 
.A(n_1614),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1622),
.Y(n_1652)
);

INVxp67_ASAP7_75t_SL g1653 ( 
.A(n_1609),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1623),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1625),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1607),
.B(n_1634),
.Y(n_1656)
);

AO21x1_ASAP7_75t_L g1657 ( 
.A1(n_1605),
.A2(n_1569),
.B(n_1572),
.Y(n_1657)
);

INVx4_ASAP7_75t_SL g1658 ( 
.A(n_1614),
.Y(n_1658)
);

BUFx8_ASAP7_75t_L g1659 ( 
.A(n_1598),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1627),
.Y(n_1660)
);

NAND3xp33_ASAP7_75t_SL g1661 ( 
.A(n_1618),
.B(n_1575),
.C(n_1573),
.Y(n_1661)
);

INVx4_ASAP7_75t_SL g1662 ( 
.A(n_1629),
.Y(n_1662)
);

HB1xp67_ASAP7_75t_L g1663 ( 
.A(n_1602),
.Y(n_1663)
);

OA21x2_ASAP7_75t_L g1664 ( 
.A1(n_1609),
.A2(n_1591),
.B(n_1585),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_SL g1665 ( 
.A(n_1630),
.B(n_1579),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1632),
.Y(n_1666)
);

NOR2xp33_ASAP7_75t_L g1667 ( 
.A(n_1633),
.B(n_1555),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1624),
.Y(n_1668)
);

BUFx6f_ASAP7_75t_L g1669 ( 
.A(n_1606),
.Y(n_1669)
);

BUFx3_ASAP7_75t_L g1670 ( 
.A(n_1594),
.Y(n_1670)
);

HB1xp67_ASAP7_75t_L g1671 ( 
.A(n_1604),
.Y(n_1671)
);

INVxp67_ASAP7_75t_SL g1672 ( 
.A(n_1624),
.Y(n_1672)
);

INVx2_ASAP7_75t_SL g1673 ( 
.A(n_1662),
.Y(n_1673)
);

BUFx3_ASAP7_75t_L g1674 ( 
.A(n_1670),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1662),
.B(n_1629),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1639),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1662),
.B(n_1607),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1662),
.B(n_1634),
.Y(n_1678)
);

OR2x2_ASAP7_75t_L g1679 ( 
.A(n_1668),
.B(n_1616),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1647),
.B(n_1628),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1645),
.B(n_1611),
.Y(n_1681)
);

HB1xp67_ASAP7_75t_L g1682 ( 
.A(n_1641),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1639),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1644),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1647),
.B(n_1604),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1644),
.Y(n_1686)
);

OR2x2_ASAP7_75t_L g1687 ( 
.A(n_1672),
.B(n_1586),
.Y(n_1687)
);

AOI22xp33_ASAP7_75t_L g1688 ( 
.A1(n_1659),
.A2(n_1603),
.B1(n_1595),
.B2(n_1599),
.Y(n_1688)
);

NAND3xp33_ASAP7_75t_L g1689 ( 
.A(n_1659),
.B(n_1601),
.C(n_1603),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1652),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1652),
.Y(n_1691)
);

AND2x4_ASAP7_75t_L g1692 ( 
.A(n_1643),
.B(n_1589),
.Y(n_1692)
);

OR2x6_ASAP7_75t_L g1693 ( 
.A(n_1669),
.B(n_1589),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1654),
.Y(n_1694)
);

HB1xp67_ASAP7_75t_L g1695 ( 
.A(n_1646),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1653),
.B(n_1608),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1643),
.B(n_1575),
.Y(n_1697)
);

AOI322xp5_ASAP7_75t_L g1698 ( 
.A1(n_1661),
.A2(n_1601),
.A3(n_1571),
.B1(n_1575),
.B2(n_1573),
.C1(n_1576),
.C2(n_1562),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1654),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1643),
.B(n_1575),
.Y(n_1700)
);

OR2x2_ASAP7_75t_L g1701 ( 
.A(n_1638),
.B(n_1642),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1635),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1650),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1655),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1655),
.Y(n_1705)
);

OR2x2_ASAP7_75t_L g1706 ( 
.A(n_1666),
.B(n_1663),
.Y(n_1706)
);

CKINVDCx20_ASAP7_75t_R g1707 ( 
.A(n_1659),
.Y(n_1707)
);

OR2x2_ASAP7_75t_L g1708 ( 
.A(n_1666),
.B(n_1586),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1660),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1664),
.Y(n_1710)
);

NAND3xp33_ASAP7_75t_L g1711 ( 
.A(n_1669),
.B(n_1612),
.C(n_1611),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1660),
.Y(n_1712)
);

HB1xp67_ASAP7_75t_L g1713 ( 
.A(n_1671),
.Y(n_1713)
);

OR2x2_ASAP7_75t_L g1714 ( 
.A(n_1637),
.B(n_1586),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1690),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1675),
.B(n_1643),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1690),
.Y(n_1717)
);

INVx2_ASAP7_75t_SL g1718 ( 
.A(n_1692),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1680),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1691),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1675),
.B(n_1658),
.Y(n_1721)
);

INVxp67_ASAP7_75t_L g1722 ( 
.A(n_1674),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1693),
.B(n_1658),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1691),
.Y(n_1724)
);

NAND2x1_ASAP7_75t_SL g1725 ( 
.A(n_1692),
.B(n_1651),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1676),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1683),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1693),
.B(n_1658),
.Y(n_1728)
);

INVx2_ASAP7_75t_SL g1729 ( 
.A(n_1692),
.Y(n_1729)
);

NOR2xp33_ASAP7_75t_L g1730 ( 
.A(n_1707),
.B(n_1436),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1682),
.B(n_1656),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1684),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1686),
.Y(n_1733)
);

OR2x2_ASAP7_75t_L g1734 ( 
.A(n_1706),
.B(n_1648),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1681),
.B(n_1656),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1674),
.B(n_1649),
.Y(n_1736)
);

INVx1_ASAP7_75t_SL g1737 ( 
.A(n_1707),
.Y(n_1737)
);

AND2x2_ASAP7_75t_SL g1738 ( 
.A(n_1688),
.B(n_1669),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1698),
.B(n_1649),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1680),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1714),
.B(n_1670),
.Y(n_1741)
);

INVx2_ASAP7_75t_SL g1742 ( 
.A(n_1673),
.Y(n_1742)
);

AOI22xp5_ASAP7_75t_L g1743 ( 
.A1(n_1689),
.A2(n_1665),
.B1(n_1657),
.B2(n_1667),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1693),
.B(n_1658),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1694),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1714),
.B(n_1651),
.Y(n_1746)
);

INVx2_ASAP7_75t_SL g1747 ( 
.A(n_1673),
.Y(n_1747)
);

INVx1_ASAP7_75t_SL g1748 ( 
.A(n_1701),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1696),
.B(n_1651),
.Y(n_1749)
);

AND2x4_ASAP7_75t_L g1750 ( 
.A(n_1693),
.B(n_1669),
.Y(n_1750)
);

AOI22xp33_ASAP7_75t_L g1751 ( 
.A1(n_1738),
.A2(n_1711),
.B1(n_1657),
.B2(n_1696),
.Y(n_1751)
);

OR2x2_ASAP7_75t_L g1752 ( 
.A(n_1748),
.B(n_1701),
.Y(n_1752)
);

INVx1_ASAP7_75t_SL g1753 ( 
.A(n_1737),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1717),
.Y(n_1754)
);

INVxp67_ASAP7_75t_L g1755 ( 
.A(n_1749),
.Y(n_1755)
);

NOR2x1_ASAP7_75t_L g1756 ( 
.A(n_1723),
.B(n_1697),
.Y(n_1756)
);

AND2x4_ASAP7_75t_L g1757 ( 
.A(n_1716),
.B(n_1677),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1717),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1716),
.B(n_1677),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1722),
.B(n_1695),
.Y(n_1760)
);

INVx1_ASAP7_75t_SL g1761 ( 
.A(n_1721),
.Y(n_1761)
);

INVx5_ASAP7_75t_L g1762 ( 
.A(n_1723),
.Y(n_1762)
);

INVx1_ASAP7_75t_SL g1763 ( 
.A(n_1721),
.Y(n_1763)
);

INVx1_ASAP7_75t_SL g1764 ( 
.A(n_1725),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1728),
.B(n_1744),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1724),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1724),
.Y(n_1767)
);

NOR2xp33_ASAP7_75t_L g1768 ( 
.A(n_1730),
.B(n_1669),
.Y(n_1768)
);

INVx1_ASAP7_75t_SL g1769 ( 
.A(n_1725),
.Y(n_1769)
);

AND2x2_ASAP7_75t_L g1770 ( 
.A(n_1728),
.B(n_1697),
.Y(n_1770)
);

AND2x4_ASAP7_75t_L g1771 ( 
.A(n_1718),
.B(n_1678),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1715),
.Y(n_1772)
);

INVx1_ASAP7_75t_SL g1773 ( 
.A(n_1744),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1720),
.Y(n_1774)
);

OR2x2_ASAP7_75t_L g1775 ( 
.A(n_1731),
.B(n_1706),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1726),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1753),
.B(n_1719),
.Y(n_1777)
);

OAI221xp5_ASAP7_75t_L g1778 ( 
.A1(n_1751),
.A2(n_1743),
.B1(n_1739),
.B2(n_1729),
.C(n_1718),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1754),
.Y(n_1779)
);

NOR3xp33_ASAP7_75t_L g1780 ( 
.A(n_1773),
.B(n_1747),
.C(n_1742),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1758),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1761),
.B(n_1719),
.Y(n_1782)
);

NOR2xp33_ASAP7_75t_L g1783 ( 
.A(n_1768),
.B(n_1738),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1766),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1763),
.B(n_1740),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1767),
.Y(n_1786)
);

INVx1_ASAP7_75t_SL g1787 ( 
.A(n_1759),
.Y(n_1787)
);

NAND2xp33_ASAP7_75t_SL g1788 ( 
.A(n_1751),
.B(n_1729),
.Y(n_1788)
);

INVx2_ASAP7_75t_SL g1789 ( 
.A(n_1762),
.Y(n_1789)
);

OAI221xp5_ASAP7_75t_SL g1790 ( 
.A1(n_1752),
.A2(n_1734),
.B1(n_1735),
.B2(n_1746),
.C(n_1741),
.Y(n_1790)
);

AOI21xp33_ASAP7_75t_L g1791 ( 
.A1(n_1768),
.A2(n_1750),
.B(n_1747),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_1757),
.Y(n_1792)
);

AOI22xp5_ASAP7_75t_L g1793 ( 
.A1(n_1757),
.A2(n_1750),
.B1(n_1740),
.B2(n_1736),
.Y(n_1793)
);

OR2x2_ASAP7_75t_L g1794 ( 
.A(n_1760),
.B(n_1734),
.Y(n_1794)
);

AOI22xp5_ASAP7_75t_L g1795 ( 
.A1(n_1757),
.A2(n_1750),
.B1(n_1700),
.B2(n_1742),
.Y(n_1795)
);

INVx2_ASAP7_75t_L g1796 ( 
.A(n_1759),
.Y(n_1796)
);

AND2x4_ASAP7_75t_SL g1797 ( 
.A(n_1792),
.B(n_1765),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1787),
.B(n_1755),
.Y(n_1798)
);

INVxp67_ASAP7_75t_L g1799 ( 
.A(n_1783),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1796),
.Y(n_1800)
);

NOR3xp33_ASAP7_75t_L g1801 ( 
.A(n_1788),
.B(n_1765),
.C(n_1764),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1780),
.B(n_1762),
.Y(n_1802)
);

INVx2_ASAP7_75t_L g1803 ( 
.A(n_1789),
.Y(n_1803)
);

INVx2_ASAP7_75t_L g1804 ( 
.A(n_1777),
.Y(n_1804)
);

NAND3xp33_ASAP7_75t_L g1805 ( 
.A(n_1778),
.B(n_1762),
.C(n_1776),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1795),
.B(n_1770),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1782),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_SL g1808 ( 
.A(n_1783),
.B(n_1762),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_L g1809 ( 
.A(n_1780),
.B(n_1770),
.Y(n_1809)
);

OAI211xp5_ASAP7_75t_SL g1810 ( 
.A1(n_1805),
.A2(n_1791),
.B(n_1793),
.C(n_1794),
.Y(n_1810)
);

AOI211xp5_ASAP7_75t_SL g1811 ( 
.A1(n_1801),
.A2(n_1802),
.B(n_1799),
.C(n_1809),
.Y(n_1811)
);

NOR4xp25_ASAP7_75t_L g1812 ( 
.A(n_1805),
.B(n_1790),
.C(n_1786),
.D(n_1779),
.Y(n_1812)
);

AOI221xp5_ASAP7_75t_L g1813 ( 
.A1(n_1808),
.A2(n_1790),
.B1(n_1785),
.B2(n_1784),
.C(n_1781),
.Y(n_1813)
);

NAND5xp2_ASAP7_75t_SL g1814 ( 
.A(n_1806),
.B(n_1769),
.C(n_1756),
.D(n_1700),
.E(n_1447),
.Y(n_1814)
);

NAND3xp33_ASAP7_75t_L g1815 ( 
.A(n_1803),
.B(n_1771),
.C(n_1772),
.Y(n_1815)
);

A2O1A1Ixp33_ASAP7_75t_L g1816 ( 
.A1(n_1797),
.A2(n_1771),
.B(n_1775),
.C(n_1774),
.Y(n_1816)
);

NOR2xp33_ASAP7_75t_R g1817 ( 
.A(n_1807),
.B(n_1469),
.Y(n_1817)
);

OAI322xp33_ASAP7_75t_L g1818 ( 
.A1(n_1798),
.A2(n_1726),
.A3(n_1727),
.B1(n_1733),
.B2(n_1732),
.C1(n_1745),
.C2(n_1710),
.Y(n_1818)
);

O2A1O1Ixp5_ASAP7_75t_L g1819 ( 
.A1(n_1798),
.A2(n_1771),
.B(n_1727),
.C(n_1710),
.Y(n_1819)
);

OA21x2_ASAP7_75t_L g1820 ( 
.A1(n_1819),
.A2(n_1800),
.B(n_1804),
.Y(n_1820)
);

AND2x2_ASAP7_75t_SL g1821 ( 
.A(n_1812),
.B(n_1713),
.Y(n_1821)
);

INVx1_ASAP7_75t_SL g1822 ( 
.A(n_1817),
.Y(n_1822)
);

OAI22xp33_ASAP7_75t_L g1823 ( 
.A1(n_1811),
.A2(n_1617),
.B1(n_1687),
.B2(n_1709),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1815),
.Y(n_1824)
);

INVxp33_ASAP7_75t_SL g1825 ( 
.A(n_1822),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1820),
.Y(n_1826)
);

OR2x2_ASAP7_75t_L g1827 ( 
.A(n_1824),
.B(n_1816),
.Y(n_1827)
);

NAND3xp33_ASAP7_75t_L g1828 ( 
.A(n_1821),
.B(n_1813),
.C(n_1810),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1820),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1822),
.Y(n_1830)
);

OAI22xp5_ASAP7_75t_L g1831 ( 
.A1(n_1828),
.A2(n_1823),
.B1(n_1705),
.B2(n_1712),
.Y(n_1831)
);

AOI222xp33_ASAP7_75t_L g1832 ( 
.A1(n_1826),
.A2(n_1814),
.B1(n_1818),
.B2(n_1704),
.C1(n_1685),
.C2(n_1703),
.Y(n_1832)
);

AOI21xp33_ASAP7_75t_SL g1833 ( 
.A1(n_1825),
.A2(n_1451),
.B(n_1463),
.Y(n_1833)
);

NOR3xp33_ASAP7_75t_L g1834 ( 
.A(n_1830),
.B(n_1476),
.C(n_1478),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1829),
.Y(n_1835)
);

AND3x4_ASAP7_75t_L g1836 ( 
.A(n_1834),
.B(n_1429),
.C(n_1498),
.Y(n_1836)
);

NOR2x1_ASAP7_75t_L g1837 ( 
.A(n_1835),
.B(n_1827),
.Y(n_1837)
);

INVx2_ASAP7_75t_L g1838 ( 
.A(n_1831),
.Y(n_1838)
);

AND2x4_ASAP7_75t_L g1839 ( 
.A(n_1837),
.B(n_1685),
.Y(n_1839)
);

AOI31xp33_ASAP7_75t_L g1840 ( 
.A1(n_1839),
.A2(n_1838),
.A3(n_1833),
.B(n_1832),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1840),
.Y(n_1841)
);

BUFx6f_ASAP7_75t_L g1842 ( 
.A(n_1840),
.Y(n_1842)
);

NAND2x1p5_ASAP7_75t_L g1843 ( 
.A(n_1842),
.B(n_1836),
.Y(n_1843)
);

NAND2x1p5_ASAP7_75t_L g1844 ( 
.A(n_1842),
.B(n_1589),
.Y(n_1844)
);

AOI21xp5_ASAP7_75t_L g1845 ( 
.A1(n_1844),
.A2(n_1841),
.B(n_1702),
.Y(n_1845)
);

CKINVDCx20_ASAP7_75t_R g1846 ( 
.A(n_1845),
.Y(n_1846)
);

AOI22xp33_ASAP7_75t_SL g1847 ( 
.A1(n_1846),
.A2(n_1843),
.B1(n_1699),
.B2(n_1678),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1847),
.B(n_1708),
.Y(n_1848)
);

AOI322xp5_ASAP7_75t_L g1849 ( 
.A1(n_1848),
.A2(n_1636),
.A3(n_1640),
.B1(n_1571),
.B2(n_1565),
.C1(n_1581),
.C2(n_1588),
.Y(n_1849)
);

AOI22xp5_ASAP7_75t_L g1850 ( 
.A1(n_1849),
.A2(n_1708),
.B1(n_1687),
.B2(n_1679),
.Y(n_1850)
);

AOI211xp5_ASAP7_75t_L g1851 ( 
.A1(n_1850),
.A2(n_1580),
.B(n_1496),
.C(n_1621),
.Y(n_1851)
);


endmodule