module fake_jpeg_18516_n_164 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_164);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_164;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_122;
wire n_75;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_30),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_46),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_7),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_12),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_7),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_14),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_23),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_13),
.Y(n_68)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_2),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_31),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_0),
.Y(n_72)
);

INVx6_ASAP7_75t_SL g73 ( 
.A(n_40),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_24),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_17),
.Y(n_76)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_79),
.Y(n_87)
);

BUFx16f_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_81),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_54),
.B(n_1),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_51),
.B(n_1),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_72),
.Y(n_93)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_83),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_78),
.A2(n_70),
.B1(n_76),
.B2(n_69),
.Y(n_84)
);

AO22x1_ASAP7_75t_SL g100 ( 
.A1(n_84),
.A2(n_64),
.B1(n_71),
.B2(n_68),
.Y(n_100)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_80),
.Y(n_85)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_83),
.A2(n_76),
.B1(n_62),
.B2(n_73),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_89),
.B(n_67),
.Y(n_99)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_77),
.Y(n_92)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_92),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_93),
.B(n_94),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_79),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_84),
.A2(n_49),
.B1(n_56),
.B2(n_64),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_96),
.A2(n_99),
.B1(n_71),
.B2(n_49),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_91),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_97),
.B(n_102),
.Y(n_114)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_86),
.Y(n_98)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_98),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_100),
.A2(n_88),
.B1(n_87),
.B2(n_68),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_86),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_85),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_103),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_90),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_SL g111 ( 
.A(n_104),
.B(n_101),
.C(n_53),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_93),
.B(n_80),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_106),
.A2(n_60),
.B(n_52),
.Y(n_117)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_107),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_107),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_108),
.B(n_115),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_111),
.A2(n_116),
.B(n_117),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_112),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_105),
.Y(n_115)
);

NAND3xp33_ASAP7_75t_L g116 ( 
.A(n_106),
.B(n_50),
.C(n_74),
.Y(n_116)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_100),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_118),
.Y(n_132)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_95),
.Y(n_119)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_119),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_120),
.A2(n_55),
.B1(n_5),
.B2(n_6),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_95),
.A2(n_66),
.B(n_65),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_121),
.B(n_122),
.Y(n_134)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_107),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_101),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_123),
.A2(n_124),
.B1(n_59),
.B2(n_58),
.Y(n_129)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_107),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_116),
.B(n_48),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_125),
.B(n_127),
.Y(n_147)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_114),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_113),
.B(n_63),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_128),
.B(n_133),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_129),
.Y(n_143)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_109),
.Y(n_130)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_130),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_110),
.B(n_75),
.C(n_61),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_135),
.A2(n_138),
.B1(n_4),
.B2(n_5),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_123),
.B(n_3),
.Y(n_137)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_137),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_134),
.B(n_124),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_139),
.B(n_126),
.C(n_132),
.Y(n_148)
);

OR2x2_ASAP7_75t_L g141 ( 
.A(n_136),
.B(n_122),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_141),
.A2(n_145),
.B1(n_146),
.B2(n_6),
.Y(n_151)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_136),
.Y(n_146)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_148),
.Y(n_152)
);

OAI21xp33_ASAP7_75t_SL g149 ( 
.A1(n_141),
.A2(n_132),
.B(n_131),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_144),
.B(n_27),
.C(n_45),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_150),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_143),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_151),
.C(n_149),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_155),
.A2(n_140),
.B1(n_147),
.B2(n_142),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_156),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_32),
.C(n_11),
.Y(n_158)
);

NOR2xp67_ASAP7_75t_SL g159 ( 
.A(n_158),
.B(n_33),
.Y(n_159)
);

NOR2x1_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_29),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_160),
.B(n_37),
.C(n_16),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_161),
.A2(n_41),
.B(n_18),
.Y(n_162)
);

FAx1_ASAP7_75t_SL g163 ( 
.A(n_162),
.B(n_20),
.CI(n_26),
.CON(n_163),
.SN(n_163)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_42),
.Y(n_164)
);


endmodule