module fake_jpeg_15130_n_212 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_212);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_212;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_0),
.Y(n_13)
);

INVx5_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx2_ASAP7_75t_SL g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx8_ASAP7_75t_SL g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_10),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_27),
.B(n_12),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_28),
.B(n_32),
.Y(n_50)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

CKINVDCx6p67_ASAP7_75t_R g41 ( 
.A(n_30),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_6),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_35),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_37),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_37),
.B(n_25),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_38),
.B(n_16),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_34),
.A2(n_15),
.B1(n_23),
.B2(n_14),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_45),
.A2(n_27),
.B1(n_20),
.B2(n_35),
.Y(n_72)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_29),
.A2(n_22),
.B1(n_14),
.B2(n_24),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_47),
.A2(n_15),
.B1(n_34),
.B2(n_20),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_28),
.B(n_23),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_49),
.B(n_50),
.Y(n_59)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_51),
.B(n_62),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_46),
.B(n_28),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_52),
.B(n_53),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_50),
.B(n_37),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_47),
.A2(n_14),
.B1(n_34),
.B2(n_24),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_54),
.A2(n_57),
.B1(n_70),
.B2(n_75),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_37),
.Y(n_55)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_32),
.Y(n_56)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_42),
.A2(n_34),
.B1(n_15),
.B2(n_29),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_29),
.C(n_33),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_58),
.B(n_67),
.C(n_31),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_45),
.A2(n_15),
.B1(n_27),
.B2(n_20),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_60),
.A2(n_30),
.B(n_31),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_49),
.B(n_26),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_16),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_65),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_16),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_69),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_36),
.C(n_33),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_47),
.B(n_21),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_41),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_71),
.B(n_77),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_72),
.A2(n_73),
.B1(n_40),
.B2(n_71),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_40),
.A2(n_35),
.B1(n_13),
.B2(n_26),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_48),
.B(n_21),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_74),
.B(n_13),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_48),
.A2(n_35),
.B1(n_36),
.B2(n_33),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_39),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_41),
.Y(n_77)
);

AO21x1_ASAP7_75t_L g113 ( 
.A1(n_78),
.A2(n_97),
.B(n_41),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_83),
.B(n_88),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_74),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_85),
.B(n_94),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_87),
.B(n_69),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_64),
.B(n_36),
.Y(n_88)
);

MAJx2_ASAP7_75t_L g91 ( 
.A(n_55),
.B(n_31),
.C(n_30),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_91),
.B(n_60),
.C(n_70),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_66),
.B(n_36),
.Y(n_94)
);

OAI21xp33_ASAP7_75t_L g95 ( 
.A1(n_56),
.A2(n_53),
.B(n_52),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_95),
.A2(n_98),
.B(n_101),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_65),
.B(n_33),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_30),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_58),
.B(n_31),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_61),
.B(n_59),
.Y(n_100)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_100),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_67),
.B(n_31),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_104),
.A2(n_110),
.B1(n_113),
.B2(n_101),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_84),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_105),
.B(n_108),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_106),
.B(n_80),
.C(n_81),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_98),
.A2(n_65),
.B1(n_61),
.B2(n_51),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_107),
.A2(n_112),
.B1(n_120),
.B2(n_97),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_82),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_82),
.B(n_62),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g125 ( 
.A(n_109),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_79),
.A2(n_75),
.B1(n_59),
.B2(n_76),
.Y(n_110)
);

NOR2xp67_ASAP7_75t_R g111 ( 
.A(n_99),
.B(n_30),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_111),
.A2(n_94),
.B(n_96),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_79),
.A2(n_77),
.B1(n_68),
.B2(n_63),
.Y(n_112)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_86),
.Y(n_114)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_114),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_92),
.B(n_17),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_116),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_117),
.B(n_89),
.Y(n_135)
);

AO22x1_ASAP7_75t_SL g118 ( 
.A1(n_91),
.A2(n_41),
.B1(n_35),
.B2(n_17),
.Y(n_118)
);

AO22x1_ASAP7_75t_SL g145 ( 
.A1(n_118),
.A2(n_41),
.B1(n_86),
.B2(n_4),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_84),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_119),
.B(n_121),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_87),
.A2(n_41),
.B1(n_17),
.B2(n_18),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_92),
.B(n_18),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_1),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_122),
.B(n_124),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_88),
.B(n_1),
.Y(n_124)
);

NAND3xp33_ASAP7_75t_L g127 ( 
.A(n_108),
.B(n_80),
.C(n_85),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_127),
.B(n_142),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_128),
.A2(n_142),
.B1(n_132),
.B2(n_140),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_129),
.A2(n_104),
.B1(n_113),
.B2(n_118),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_130),
.A2(n_111),
.B(n_117),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_110),
.A2(n_101),
.B1(n_98),
.B2(n_89),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_132),
.A2(n_105),
.B1(n_118),
.B2(n_103),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_135),
.B(n_145),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_136),
.B(n_140),
.C(n_141),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_123),
.B(n_81),
.Y(n_137)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_137),
.Y(n_147)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_114),
.Y(n_139)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_139),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_115),
.B(n_91),
.C(n_99),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_115),
.B(n_83),
.C(n_90),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_120),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_102),
.Y(n_143)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_143),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_103),
.B(n_93),
.Y(n_144)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_144),
.Y(n_160)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_112),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_146),
.B(n_2),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_148),
.A2(n_131),
.B(n_5),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_146),
.A2(n_106),
.B1(n_113),
.B2(n_119),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_150),
.A2(n_156),
.B1(n_141),
.B2(n_130),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_136),
.B(n_104),
.C(n_107),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_153),
.B(n_162),
.C(n_139),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_155),
.A2(n_157),
.B1(n_2),
.B2(n_5),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_126),
.B(n_102),
.Y(n_159)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_159),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_133),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_161),
.B(n_125),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_128),
.B(n_1),
.C(n_2),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_163),
.A2(n_144),
.B(n_135),
.Y(n_165)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_152),
.Y(n_164)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_164),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_165),
.Y(n_177)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_152),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_166),
.B(n_172),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_167),
.B(n_171),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_158),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_168),
.B(n_174),
.Y(n_185)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_169),
.Y(n_180)
);

OAI322xp33_ASAP7_75t_L g170 ( 
.A1(n_147),
.A2(n_137),
.A3(n_143),
.B1(n_134),
.B2(n_129),
.C1(n_145),
.C2(n_138),
.Y(n_170)
);

NOR4xp25_ASAP7_75t_L g179 ( 
.A(n_170),
.B(n_157),
.C(n_154),
.D(n_151),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_149),
.B(n_131),
.C(n_145),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_173),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_165),
.A2(n_154),
.B(n_156),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_178),
.A2(n_148),
.B(n_153),
.Y(n_190)
);

OAI31xp33_ASAP7_75t_L g193 ( 
.A1(n_179),
.A2(n_6),
.A3(n_7),
.B(n_8),
.Y(n_193)
);

NOR3xp33_ASAP7_75t_SL g181 ( 
.A(n_175),
.B(n_159),
.C(n_162),
.Y(n_181)
);

AOI31xp67_ASAP7_75t_L g187 ( 
.A1(n_181),
.A2(n_173),
.A3(n_163),
.B(n_160),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_164),
.B(n_160),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g195 ( 
.A(n_183),
.Y(n_195)
);

NAND3xp33_ASAP7_75t_SL g196 ( 
.A(n_187),
.B(n_188),
.C(n_184),
.Y(n_196)
);

NAND4xp25_ASAP7_75t_L g188 ( 
.A(n_181),
.B(n_172),
.C(n_171),
.D(n_174),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_177),
.A2(n_147),
.B1(n_158),
.B2(n_150),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_189),
.A2(n_191),
.B1(n_192),
.B2(n_183),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_190),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_186),
.B(n_182),
.C(n_149),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_186),
.B(n_5),
.C(n_6),
.Y(n_192)
);

NAND3xp33_ASAP7_75t_L g201 ( 
.A(n_193),
.B(n_194),
.C(n_7),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_178),
.B(n_7),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_196),
.B(n_197),
.Y(n_202)
);

INVxp33_ASAP7_75t_L g197 ( 
.A(n_195),
.Y(n_197)
);

AOI31xp33_ASAP7_75t_L g198 ( 
.A1(n_194),
.A2(n_180),
.A3(n_185),
.B(n_176),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_198),
.B(n_9),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_200),
.B(n_192),
.C(n_191),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_201),
.B(n_9),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_203),
.B(n_204),
.C(n_197),
.Y(n_207)
);

AND2x4_ASAP7_75t_L g205 ( 
.A(n_199),
.B(n_9),
.Y(n_205)
);

NAND3xp33_ASAP7_75t_L g209 ( 
.A(n_205),
.B(n_206),
.C(n_11),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_207),
.B(n_208),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_202),
.B(n_11),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_209),
.A2(n_205),
.B(n_11),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_211),
.B(n_210),
.Y(n_212)
);


endmodule