module fake_netlist_5_1675_n_1774 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1774);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1774;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_156;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_157;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_1723;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1097;
wire n_1036;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_290;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_433;
wire n_368;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_1757;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1363;
wire n_1301;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_1722;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_172;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_1771;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_159;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_1747;
wire n_714;
wire n_1683;
wire n_909;
wire n_1530;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_158;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_41),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_44),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g158 ( 
.A(n_5),
.Y(n_158)
);

BUFx10_ASAP7_75t_L g159 ( 
.A(n_3),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_13),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_63),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_67),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_20),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_153),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_105),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_19),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_9),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_98),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_66),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_104),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_34),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_116),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_44),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_70),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_136),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_130),
.Y(n_176)
);

INVx2_ASAP7_75t_SL g177 ( 
.A(n_76),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_23),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_73),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_55),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_74),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_75),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_7),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_61),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_93),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_145),
.Y(n_186)
);

BUFx2_ASAP7_75t_L g187 ( 
.A(n_154),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_26),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_135),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_31),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_29),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_131),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_59),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_83),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_77),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_82),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_134),
.Y(n_197)
);

BUFx5_ASAP7_75t_L g198 ( 
.A(n_117),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_60),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_39),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_5),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_123),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_121),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_109),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_65),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_18),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_3),
.Y(n_207)
);

INVx2_ASAP7_75t_SL g208 ( 
.A(n_155),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_11),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_133),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_81),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_84),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_1),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_49),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_21),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_112),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_48),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_10),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_13),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_32),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_89),
.Y(n_221)
);

BUFx10_ASAP7_75t_L g222 ( 
.A(n_107),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_8),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_54),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_38),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_96),
.Y(n_226)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_62),
.Y(n_227)
);

BUFx10_ASAP7_75t_L g228 ( 
.A(n_33),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_78),
.Y(n_229)
);

BUFx2_ASAP7_75t_L g230 ( 
.A(n_97),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_80),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_106),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_122),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_102),
.Y(n_234)
);

BUFx8_ASAP7_75t_SL g235 ( 
.A(n_24),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_147),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_57),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_12),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_144),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_1),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_15),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_113),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_15),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_0),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_100),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_69),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_36),
.Y(n_247)
);

INVx2_ASAP7_75t_SL g248 ( 
.A(n_53),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_141),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_17),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_88),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_132),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_17),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_32),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_26),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_150),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_125),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_0),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_25),
.Y(n_259)
);

INVx2_ASAP7_75t_SL g260 ( 
.A(n_101),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_8),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_4),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_91),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_40),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_94),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_124),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_86),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_33),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_71),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_146),
.Y(n_270)
);

BUFx10_ASAP7_75t_L g271 ( 
.A(n_108),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_46),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_21),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_128),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g275 ( 
.A(n_9),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_85),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_4),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_79),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_35),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_126),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_111),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_10),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_50),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_139),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_2),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_56),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_14),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_152),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_36),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_149),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_34),
.Y(n_291)
);

BUFx10_ASAP7_75t_L g292 ( 
.A(n_22),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_45),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_35),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_6),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_99),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_64),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_90),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_27),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_72),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_2),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_40),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_29),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_6),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_52),
.Y(n_305)
);

BUFx10_ASAP7_75t_L g306 ( 
.A(n_7),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_148),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_18),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_183),
.Y(n_309)
);

CKINVDCx14_ASAP7_75t_R g310 ( 
.A(n_227),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_235),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_183),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_183),
.Y(n_313)
);

HB1xp67_ASAP7_75t_L g314 ( 
.A(n_295),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_168),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_159),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_183),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_219),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_219),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_219),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_159),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_219),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_166),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_168),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_166),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_159),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_244),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_198),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_244),
.Y(n_329)
);

INVxp33_ASAP7_75t_SL g330 ( 
.A(n_171),
.Y(n_330)
);

CKINVDCx16_ASAP7_75t_R g331 ( 
.A(n_256),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_161),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_193),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_162),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_193),
.Y(n_335)
);

HB1xp67_ASAP7_75t_L g336 ( 
.A(n_171),
.Y(n_336)
);

INVx1_ASAP7_75t_SL g337 ( 
.A(n_228),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_188),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_164),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_169),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_201),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_195),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_206),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_215),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_308),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_198),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_238),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_243),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_181),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_250),
.Y(n_350)
);

BUFx3_ASAP7_75t_L g351 ( 
.A(n_170),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_182),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_253),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_255),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_189),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_195),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_259),
.Y(n_357)
);

INVxp67_ASAP7_75t_SL g358 ( 
.A(n_187),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_268),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_279),
.Y(n_360)
);

INVx3_ASAP7_75t_L g361 ( 
.A(n_170),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_216),
.Y(n_362)
);

CKINVDCx14_ASAP7_75t_R g363 ( 
.A(n_230),
.Y(n_363)
);

INVxp67_ASAP7_75t_SL g364 ( 
.A(n_179),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_216),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_287),
.Y(n_366)
);

INVxp33_ASAP7_75t_SL g367 ( 
.A(n_178),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_293),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_194),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_304),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_199),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_242),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_186),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_204),
.Y(n_374)
);

INVxp33_ASAP7_75t_SL g375 ( 
.A(n_178),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_186),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_205),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_203),
.Y(n_378)
);

INVxp33_ASAP7_75t_SL g379 ( 
.A(n_299),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_332),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_328),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_309),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_328),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_346),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_346),
.Y(n_385)
);

INVx3_ASAP7_75t_L g386 ( 
.A(n_309),
.Y(n_386)
);

INVx3_ASAP7_75t_L g387 ( 
.A(n_312),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_361),
.B(n_364),
.Y(n_388)
);

INVx4_ASAP7_75t_L g389 ( 
.A(n_361),
.Y(n_389)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_312),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_313),
.Y(n_391)
);

BUFx12f_ASAP7_75t_L g392 ( 
.A(n_311),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_313),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_361),
.B(n_177),
.Y(n_394)
);

AND2x4_ASAP7_75t_L g395 ( 
.A(n_373),
.B(n_179),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_317),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_373),
.Y(n_397)
);

NAND2xp33_ASAP7_75t_R g398 ( 
.A(n_330),
.B(n_299),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_317),
.Y(n_399)
);

INVxp33_ASAP7_75t_SL g400 ( 
.A(n_314),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_376),
.Y(n_401)
);

BUFx3_ASAP7_75t_L g402 ( 
.A(n_318),
.Y(n_402)
);

BUFx8_ASAP7_75t_L g403 ( 
.A(n_351),
.Y(n_403)
);

OA21x2_ASAP7_75t_L g404 ( 
.A1(n_376),
.A2(n_203),
.B(n_174),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_334),
.Y(n_405)
);

INVx2_ASAP7_75t_SL g406 ( 
.A(n_351),
.Y(n_406)
);

AND2x4_ASAP7_75t_L g407 ( 
.A(n_378),
.B(n_232),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_318),
.Y(n_408)
);

BUFx3_ASAP7_75t_L g409 ( 
.A(n_319),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_319),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_320),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_339),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_320),
.B(n_177),
.Y(n_413)
);

CKINVDCx16_ASAP7_75t_R g414 ( 
.A(n_331),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_322),
.Y(n_415)
);

HB1xp67_ASAP7_75t_L g416 ( 
.A(n_336),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_337),
.A2(n_303),
.B1(n_200),
.B2(n_254),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_322),
.Y(n_418)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_378),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_344),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_344),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_323),
.B(n_232),
.Y(n_422)
);

BUFx3_ASAP7_75t_L g423 ( 
.A(n_338),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_341),
.B(n_208),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_345),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_340),
.Y(n_426)
);

HB1xp67_ASAP7_75t_L g427 ( 
.A(n_316),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_323),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_325),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_315),
.Y(n_430)
);

INVx1_ASAP7_75t_SL g431 ( 
.A(n_324),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_358),
.B(n_208),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_367),
.B(n_248),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_345),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_325),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_349),
.Y(n_436)
);

AND2x4_ASAP7_75t_L g437 ( 
.A(n_327),
.B(n_274),
.Y(n_437)
);

INVx3_ASAP7_75t_L g438 ( 
.A(n_327),
.Y(n_438)
);

BUFx2_ASAP7_75t_L g439 ( 
.A(n_310),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_347),
.Y(n_440)
);

OR2x2_ASAP7_75t_L g441 ( 
.A(n_321),
.B(n_326),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_343),
.B(n_248),
.Y(n_442)
);

OA21x2_ASAP7_75t_L g443 ( 
.A1(n_329),
.A2(n_175),
.B(n_165),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_347),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_433),
.B(n_352),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_381),
.Y(n_446)
);

NOR3xp33_ASAP7_75t_L g447 ( 
.A(n_417),
.B(n_433),
.C(n_414),
.Y(n_447)
);

HB1xp67_ASAP7_75t_L g448 ( 
.A(n_406),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g449 ( 
.A(n_422),
.B(n_329),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_381),
.Y(n_450)
);

BUFx3_ASAP7_75t_L g451 ( 
.A(n_406),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_381),
.Y(n_452)
);

AO21x2_ASAP7_75t_L g453 ( 
.A1(n_388),
.A2(n_192),
.B(n_184),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_383),
.Y(n_454)
);

CKINVDCx11_ASAP7_75t_R g455 ( 
.A(n_392),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_389),
.B(n_355),
.Y(n_456)
);

OAI21xp33_ASAP7_75t_SL g457 ( 
.A1(n_432),
.A2(n_260),
.B(n_348),
.Y(n_457)
);

INVx6_ASAP7_75t_L g458 ( 
.A(n_389),
.Y(n_458)
);

AND2x6_ASAP7_75t_L g459 ( 
.A(n_432),
.B(n_269),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_383),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_383),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_380),
.B(n_369),
.Y(n_462)
);

NAND2xp33_ASAP7_75t_L g463 ( 
.A(n_406),
.B(n_371),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_384),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_389),
.B(n_374),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_398),
.A2(n_249),
.B1(n_242),
.B2(n_303),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_384),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_384),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_408),
.Y(n_469)
);

INVx2_ASAP7_75t_SL g470 ( 
.A(n_388),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_408),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_405),
.B(n_377),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_408),
.Y(n_473)
);

INVx3_ASAP7_75t_L g474 ( 
.A(n_385),
.Y(n_474)
);

BUFx2_ASAP7_75t_L g475 ( 
.A(n_427),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_422),
.B(n_348),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_402),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_412),
.B(n_375),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_408),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_426),
.B(n_379),
.Y(n_480)
);

BUFx10_ASAP7_75t_L g481 ( 
.A(n_436),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_402),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_402),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_410),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_403),
.B(n_249),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_410),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_402),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_400),
.B(n_363),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_409),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_410),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_389),
.B(n_260),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_403),
.B(n_222),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_410),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_389),
.B(n_274),
.Y(n_494)
);

INVxp67_ASAP7_75t_SL g495 ( 
.A(n_385),
.Y(n_495)
);

OR2x2_ASAP7_75t_L g496 ( 
.A(n_441),
.B(n_158),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_411),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_411),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_400),
.B(n_333),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_395),
.B(n_185),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_392),
.Y(n_501)
);

HB1xp67_ASAP7_75t_L g502 ( 
.A(n_416),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_403),
.B(n_441),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_392),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_403),
.B(n_222),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_411),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_411),
.Y(n_507)
);

INVx2_ASAP7_75t_SL g508 ( 
.A(n_441),
.Y(n_508)
);

BUFx2_ASAP7_75t_L g509 ( 
.A(n_427),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_385),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_422),
.B(n_350),
.Y(n_511)
);

INVxp67_ASAP7_75t_SL g512 ( 
.A(n_385),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_430),
.Y(n_513)
);

INVxp67_ASAP7_75t_SL g514 ( 
.A(n_385),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_409),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_428),
.Y(n_516)
);

INVx3_ASAP7_75t_L g517 ( 
.A(n_385),
.Y(n_517)
);

AOI21x1_ASAP7_75t_L g518 ( 
.A1(n_394),
.A2(n_197),
.B(n_196),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_395),
.B(n_211),
.Y(n_519)
);

AOI22xp33_ASAP7_75t_L g520 ( 
.A1(n_395),
.A2(n_269),
.B1(n_370),
.B2(n_368),
.Y(n_520)
);

AND2x2_ASAP7_75t_SL g521 ( 
.A(n_404),
.B(n_269),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_428),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_403),
.B(n_222),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_428),
.Y(n_524)
);

NOR2x1p5_ASAP7_75t_L g525 ( 
.A(n_424),
.B(n_156),
.Y(n_525)
);

INVx2_ASAP7_75t_SL g526 ( 
.A(n_416),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_395),
.B(n_229),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_428),
.Y(n_528)
);

OR2x2_ASAP7_75t_SL g529 ( 
.A(n_414),
.B(n_398),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_439),
.B(n_271),
.Y(n_530)
);

INVx2_ASAP7_75t_SL g531 ( 
.A(n_395),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_437),
.B(n_350),
.Y(n_532)
);

OR2x2_ASAP7_75t_L g533 ( 
.A(n_417),
.B(n_275),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_385),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_437),
.B(n_353),
.Y(n_535)
);

INVx2_ASAP7_75t_SL g536 ( 
.A(n_407),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_407),
.B(n_212),
.Y(n_537)
);

INVx2_ASAP7_75t_SL g538 ( 
.A(n_407),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_385),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_409),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_409),
.Y(n_541)
);

AO22x2_ASAP7_75t_L g542 ( 
.A1(n_394),
.A2(n_245),
.B1(n_239),
.B2(n_233),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_439),
.B(n_271),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_386),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_386),
.Y(n_545)
);

OAI21xp5_ASAP7_75t_L g546 ( 
.A1(n_404),
.A2(n_297),
.B(n_210),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_386),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_386),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_386),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_382),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_387),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_423),
.B(n_335),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_435),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_382),
.Y(n_554)
);

AOI22xp33_ASAP7_75t_L g555 ( 
.A1(n_407),
.A2(n_269),
.B1(n_370),
.B2(n_368),
.Y(n_555)
);

INVx2_ASAP7_75t_SL g556 ( 
.A(n_407),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_391),
.Y(n_557)
);

INVx2_ASAP7_75t_SL g558 ( 
.A(n_437),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_437),
.B(n_214),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_435),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_437),
.B(n_221),
.Y(n_561)
);

AND3x2_ASAP7_75t_L g562 ( 
.A(n_439),
.B(n_173),
.C(n_224),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_423),
.B(n_226),
.Y(n_563)
);

NOR2x1p5_ASAP7_75t_L g564 ( 
.A(n_424),
.B(n_157),
.Y(n_564)
);

BUFx3_ASAP7_75t_L g565 ( 
.A(n_423),
.Y(n_565)
);

INVx3_ASAP7_75t_L g566 ( 
.A(n_397),
.Y(n_566)
);

INVxp67_ASAP7_75t_L g567 ( 
.A(n_442),
.Y(n_567)
);

INVx3_ASAP7_75t_L g568 ( 
.A(n_397),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_391),
.Y(n_569)
);

INVx3_ASAP7_75t_L g570 ( 
.A(n_397),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_423),
.B(n_393),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_393),
.B(n_231),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_387),
.Y(n_573)
);

BUFx6f_ASAP7_75t_L g574 ( 
.A(n_397),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_387),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_387),
.Y(n_576)
);

OR2x2_ASAP7_75t_L g577 ( 
.A(n_442),
.B(n_431),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_387),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_420),
.B(n_271),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_420),
.B(n_342),
.Y(n_580)
);

AND2x2_ASAP7_75t_SL g581 ( 
.A(n_404),
.B(n_202),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_396),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_396),
.B(n_234),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_399),
.B(n_236),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_390),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_399),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_397),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_421),
.B(n_172),
.Y(n_588)
);

OAI22xp5_ASAP7_75t_L g589 ( 
.A1(n_421),
.A2(n_218),
.B1(n_223),
.B2(n_213),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_415),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_390),
.Y(n_591)
);

HB1xp67_ASAP7_75t_L g592 ( 
.A(n_431),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_470),
.B(n_443),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_470),
.B(n_443),
.Y(n_594)
);

AOI22xp33_ASAP7_75t_L g595 ( 
.A1(n_581),
.A2(n_443),
.B1(n_404),
.B2(n_247),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_567),
.B(n_443),
.Y(n_596)
);

O2A1O1Ixp33_ASAP7_75t_L g597 ( 
.A1(n_457),
.A2(n_413),
.B(n_444),
.C(n_440),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_477),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_481),
.Y(n_599)
);

HB1xp67_ASAP7_75t_L g600 ( 
.A(n_526),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_477),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_577),
.B(n_172),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_446),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_482),
.Y(n_604)
);

OR2x2_ASAP7_75t_L g605 ( 
.A(n_577),
.B(n_425),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_451),
.B(n_448),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_482),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_508),
.B(n_176),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_483),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_451),
.B(n_443),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_508),
.B(n_176),
.Y(n_611)
);

OAI22xp33_ASAP7_75t_L g612 ( 
.A1(n_466),
.A2(n_240),
.B1(n_247),
.B2(n_200),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_483),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_446),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_487),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_451),
.B(n_443),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_532),
.B(n_535),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_445),
.B(n_496),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_476),
.B(n_180),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_487),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_532),
.B(n_419),
.Y(n_621)
);

OAI22xp5_ASAP7_75t_L g622 ( 
.A1(n_531),
.A2(n_283),
.B1(n_286),
.B2(n_276),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_535),
.B(n_419),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_531),
.B(n_419),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_476),
.B(n_180),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_489),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_511),
.B(n_296),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_536),
.B(n_419),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_489),
.Y(n_629)
);

INVx2_ASAP7_75t_SL g630 ( 
.A(n_511),
.Y(n_630)
);

INVx1_ASAP7_75t_SL g631 ( 
.A(n_592),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_526),
.B(n_296),
.Y(n_632)
);

AOI22xp33_ASAP7_75t_L g633 ( 
.A1(n_581),
.A2(n_404),
.B1(n_282),
.B2(n_254),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_515),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_515),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_536),
.B(n_419),
.Y(n_636)
);

NOR2xp67_ASAP7_75t_SL g637 ( 
.A(n_458),
.B(n_492),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_446),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_500),
.B(n_298),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_540),
.Y(n_640)
);

NOR2x1p5_ASAP7_75t_L g641 ( 
.A(n_501),
.B(n_160),
.Y(n_641)
);

BUFx5_ASAP7_75t_L g642 ( 
.A(n_521),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_SL g643 ( 
.A(n_481),
.B(n_240),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_538),
.B(n_438),
.Y(n_644)
);

NOR2x1p5_ASAP7_75t_L g645 ( 
.A(n_504),
.B(n_163),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_540),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_538),
.B(n_438),
.Y(n_647)
);

AOI22xp33_ASAP7_75t_L g648 ( 
.A1(n_581),
.A2(n_404),
.B1(n_282),
.B2(n_267),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_541),
.Y(n_649)
);

AOI22xp33_ASAP7_75t_L g650 ( 
.A1(n_546),
.A2(n_217),
.B1(n_265),
.B2(n_444),
.Y(n_650)
);

INVx8_ASAP7_75t_L g651 ( 
.A(n_459),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_496),
.B(n_298),
.Y(n_652)
);

AOI22xp33_ASAP7_75t_L g653 ( 
.A1(n_453),
.A2(n_440),
.B1(n_425),
.B2(n_434),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_468),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_519),
.B(n_300),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_556),
.B(n_438),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_541),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_556),
.B(n_438),
.Y(n_658)
);

AOI22xp33_ASAP7_75t_L g659 ( 
.A1(n_453),
.A2(n_434),
.B1(n_198),
.B2(n_438),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_558),
.B(n_390),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_550),
.Y(n_661)
);

AOI22xp5_ASAP7_75t_L g662 ( 
.A1(n_558),
.A2(n_356),
.B1(n_362),
.B2(n_365),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_527),
.B(n_300),
.Y(n_663)
);

NAND3xp33_ASAP7_75t_SL g664 ( 
.A(n_466),
.B(n_372),
.C(n_430),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_462),
.B(n_167),
.Y(n_665)
);

INVx3_ASAP7_75t_L g666 ( 
.A(n_565),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_480),
.B(n_237),
.Y(n_667)
);

INVxp67_ASAP7_75t_SL g668 ( 
.A(n_449),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_468),
.Y(n_669)
);

AOI22xp5_ASAP7_75t_L g670 ( 
.A1(n_447),
.A2(n_305),
.B1(n_246),
.B2(n_251),
.Y(n_670)
);

BUFx3_ASAP7_75t_L g671 ( 
.A(n_513),
.Y(n_671)
);

INVx2_ASAP7_75t_SL g672 ( 
.A(n_525),
.Y(n_672)
);

NAND2xp33_ASAP7_75t_L g673 ( 
.A(n_459),
.B(n_198),
.Y(n_673)
);

BUFx3_ASAP7_75t_L g674 ( 
.A(n_481),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_468),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_472),
.B(n_190),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_550),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_521),
.B(n_390),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_521),
.B(n_390),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_452),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_572),
.B(n_191),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_571),
.B(n_415),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_583),
.B(n_207),
.Y(n_683)
);

AOI21xp5_ASAP7_75t_L g684 ( 
.A1(n_495),
.A2(n_413),
.B(n_435),
.Y(n_684)
);

OR2x2_ASAP7_75t_L g685 ( 
.A(n_475),
.B(n_353),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_452),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_475),
.B(n_228),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_580),
.B(n_252),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_456),
.B(n_418),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_554),
.Y(n_690)
);

INVx2_ASAP7_75t_SL g691 ( 
.A(n_525),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_465),
.B(n_418),
.Y(n_692)
);

NOR2xp67_ASAP7_75t_SL g693 ( 
.A(n_458),
.B(n_257),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_488),
.B(n_263),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_460),
.Y(n_695)
);

BUFx3_ASAP7_75t_L g696 ( 
.A(n_481),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_460),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_565),
.B(n_397),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_554),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_552),
.B(n_266),
.Y(n_700)
);

BUFx6f_ASAP7_75t_L g701 ( 
.A(n_565),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_557),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_557),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_458),
.B(n_397),
.Y(n_704)
);

AOI22xp5_ASAP7_75t_L g705 ( 
.A1(n_564),
.A2(n_281),
.B1(n_290),
.B2(n_270),
.Y(n_705)
);

OR2x6_ASAP7_75t_L g706 ( 
.A(n_485),
.B(n_354),
.Y(n_706)
);

BUFx5_ASAP7_75t_L g707 ( 
.A(n_450),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_458),
.B(n_397),
.Y(n_708)
);

OR2x2_ASAP7_75t_L g709 ( 
.A(n_509),
.B(n_354),
.Y(n_709)
);

OAI21xp5_ASAP7_75t_L g710 ( 
.A1(n_512),
.A2(n_435),
.B(n_429),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_584),
.B(n_209),
.Y(n_711)
);

INVx8_ASAP7_75t_L g712 ( 
.A(n_459),
.Y(n_712)
);

BUFx3_ASAP7_75t_L g713 ( 
.A(n_529),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_569),
.B(n_401),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_569),
.B(n_582),
.Y(n_715)
);

OR2x2_ASAP7_75t_L g716 ( 
.A(n_509),
.B(n_357),
.Y(n_716)
);

BUFx6f_ASAP7_75t_L g717 ( 
.A(n_574),
.Y(n_717)
);

INVx2_ASAP7_75t_SL g718 ( 
.A(n_564),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_582),
.Y(n_719)
);

NOR3xp33_ASAP7_75t_L g720 ( 
.A(n_457),
.B(n_357),
.C(n_366),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_R g721 ( 
.A(n_455),
.B(n_278),
.Y(n_721)
);

BUFx3_ASAP7_75t_L g722 ( 
.A(n_529),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_563),
.B(n_280),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_586),
.B(n_401),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_537),
.B(n_284),
.Y(n_725)
);

OR2x6_ASAP7_75t_L g726 ( 
.A(n_503),
.B(n_359),
.Y(n_726)
);

A2O1A1Ixp33_ASAP7_75t_L g727 ( 
.A1(n_586),
.A2(n_429),
.B(n_359),
.C(n_366),
.Y(n_727)
);

NAND2xp33_ASAP7_75t_L g728 ( 
.A(n_459),
.B(n_198),
.Y(n_728)
);

INVx3_ASAP7_75t_L g729 ( 
.A(n_544),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_590),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_530),
.B(n_220),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_590),
.B(n_514),
.Y(n_732)
);

OAI221xp5_ASAP7_75t_L g733 ( 
.A1(n_533),
.A2(n_360),
.B1(n_241),
.B2(n_225),
.C(n_258),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_543),
.B(n_261),
.Y(n_734)
);

AOI22xp33_ASAP7_75t_L g735 ( 
.A1(n_453),
.A2(n_198),
.B1(n_228),
.B2(n_292),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_544),
.Y(n_736)
);

BUFx4f_ASAP7_75t_L g737 ( 
.A(n_459),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_559),
.B(n_288),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_561),
.B(n_307),
.Y(n_739)
);

NAND2xp33_ASAP7_75t_L g740 ( 
.A(n_459),
.B(n_198),
.Y(n_740)
);

BUFx3_ASAP7_75t_L g741 ( 
.A(n_502),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_478),
.B(n_292),
.Y(n_742)
);

O2A1O1Ixp33_ASAP7_75t_L g743 ( 
.A1(n_588),
.A2(n_360),
.B(n_429),
.C(n_306),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_544),
.Y(n_744)
);

AOI22xp33_ASAP7_75t_L g745 ( 
.A1(n_542),
.A2(n_292),
.B1(n_306),
.B2(n_302),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_505),
.B(n_285),
.Y(n_746)
);

NAND2x1p5_ASAP7_75t_L g747 ( 
.A(n_523),
.B(n_401),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_545),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_545),
.Y(n_749)
);

NAND3xp33_ASAP7_75t_L g750 ( 
.A(n_463),
.B(n_589),
.C(n_579),
.Y(n_750)
);

AND2x2_ASAP7_75t_L g751 ( 
.A(n_499),
.B(n_306),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_510),
.B(n_401),
.Y(n_752)
);

AOI22xp33_ASAP7_75t_L g753 ( 
.A1(n_542),
.A2(n_277),
.B1(n_301),
.B2(n_294),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_461),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_510),
.B(n_401),
.Y(n_755)
);

BUFx3_ASAP7_75t_L g756 ( 
.A(n_545),
.Y(n_756)
);

BUFx3_ASAP7_75t_L g757 ( 
.A(n_547),
.Y(n_757)
);

AOI22xp33_ASAP7_75t_L g758 ( 
.A1(n_542),
.A2(n_291),
.B1(n_289),
.B2(n_273),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_547),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_494),
.B(n_262),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_491),
.B(n_264),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_510),
.B(n_401),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_534),
.B(n_401),
.Y(n_763)
);

AO22x1_ASAP7_75t_L g764 ( 
.A1(n_731),
.A2(n_459),
.B1(n_272),
.B2(n_533),
.Y(n_764)
);

BUFx6f_ASAP7_75t_L g765 ( 
.A(n_701),
.Y(n_765)
);

AND2x2_ASAP7_75t_L g766 ( 
.A(n_600),
.B(n_562),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_598),
.Y(n_767)
);

OAI21xp33_ASAP7_75t_L g768 ( 
.A1(n_652),
.A2(n_542),
.B(n_520),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_599),
.Y(n_769)
);

BUFx3_ASAP7_75t_L g770 ( 
.A(n_671),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_601),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_604),
.Y(n_772)
);

INVx4_ASAP7_75t_L g773 ( 
.A(n_701),
.Y(n_773)
);

AOI22xp33_ASAP7_75t_L g774 ( 
.A1(n_648),
.A2(n_555),
.B1(n_454),
.B2(n_464),
.Y(n_774)
);

NOR2x1p5_ASAP7_75t_L g775 ( 
.A(n_674),
.B(n_518),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_756),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_607),
.Y(n_777)
);

BUFx8_ASAP7_75t_L g778 ( 
.A(n_741),
.Y(n_778)
);

AND2x6_ASAP7_75t_L g779 ( 
.A(n_610),
.B(n_534),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_668),
.B(n_474),
.Y(n_780)
);

AOI22xp5_ASAP7_75t_L g781 ( 
.A1(n_618),
.A2(n_517),
.B1(n_474),
.B2(n_539),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_642),
.B(n_534),
.Y(n_782)
);

OAI22xp5_ASAP7_75t_SL g783 ( 
.A1(n_662),
.A2(n_618),
.B1(n_631),
.B2(n_633),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_696),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_L g785 ( 
.A(n_600),
.B(n_474),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_668),
.B(n_474),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_609),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_757),
.Y(n_788)
);

NOR3xp33_ASAP7_75t_SL g789 ( 
.A(n_612),
.B(n_450),
.C(n_454),
.Y(n_789)
);

AND2x4_ASAP7_75t_L g790 ( 
.A(n_630),
.B(n_539),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_613),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_602),
.B(n_461),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_729),
.Y(n_793)
);

NAND2x2_ASAP7_75t_L g794 ( 
.A(n_641),
.B(n_645),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_642),
.B(n_539),
.Y(n_795)
);

AOI22xp5_ASAP7_75t_L g796 ( 
.A1(n_642),
.A2(n_517),
.B1(n_547),
.B2(n_585),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_721),
.Y(n_797)
);

INVxp67_ASAP7_75t_L g798 ( 
.A(n_605),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_595),
.B(n_517),
.Y(n_799)
);

INVx1_ASAP7_75t_SL g800 ( 
.A(n_685),
.Y(n_800)
);

INVx2_ASAP7_75t_SL g801 ( 
.A(n_709),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_602),
.B(n_517),
.Y(n_802)
);

INVx2_ASAP7_75t_SL g803 ( 
.A(n_716),
.Y(n_803)
);

AOI22xp33_ASAP7_75t_SL g804 ( 
.A1(n_643),
.A2(n_11),
.B1(n_12),
.B2(n_14),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_595),
.B(n_464),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_729),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_648),
.B(n_467),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_652),
.B(n_548),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_615),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_687),
.B(n_518),
.Y(n_810)
);

INVx2_ASAP7_75t_SL g811 ( 
.A(n_713),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_736),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_642),
.B(n_633),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_642),
.B(n_548),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_744),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_620),
.Y(n_816)
);

AND2x6_ASAP7_75t_L g817 ( 
.A(n_616),
.B(n_548),
.Y(n_817)
);

NOR2xp33_ASAP7_75t_R g818 ( 
.A(n_664),
.B(n_47),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_606),
.B(n_467),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_642),
.B(n_549),
.Y(n_820)
);

BUFx6f_ASAP7_75t_L g821 ( 
.A(n_701),
.Y(n_821)
);

OAI22xp5_ASAP7_75t_L g822 ( 
.A1(n_650),
.A2(n_591),
.B1(n_551),
.B2(n_585),
.Y(n_822)
);

INVx4_ASAP7_75t_L g823 ( 
.A(n_701),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_626),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_629),
.Y(n_825)
);

AOI22xp5_ASAP7_75t_L g826 ( 
.A1(n_681),
.A2(n_591),
.B1(n_551),
.B2(n_585),
.Y(n_826)
);

INVx1_ASAP7_75t_SL g827 ( 
.A(n_722),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_650),
.B(n_591),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_760),
.B(n_549),
.Y(n_829)
);

INVxp67_ASAP7_75t_L g830 ( 
.A(n_611),
.Y(n_830)
);

INVx3_ASAP7_75t_L g831 ( 
.A(n_666),
.Y(n_831)
);

BUFx3_ASAP7_75t_L g832 ( 
.A(n_672),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_634),
.Y(n_833)
);

BUFx3_ASAP7_75t_L g834 ( 
.A(n_691),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_617),
.B(n_549),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_621),
.B(n_551),
.Y(n_836)
);

INVx5_ASAP7_75t_L g837 ( 
.A(n_651),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_760),
.B(n_573),
.Y(n_838)
);

NAND2xp33_ASAP7_75t_L g839 ( 
.A(n_651),
.B(n_573),
.Y(n_839)
);

AOI22xp33_ASAP7_75t_L g840 ( 
.A1(n_753),
.A2(n_758),
.B1(n_735),
.B2(n_594),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_681),
.B(n_573),
.Y(n_841)
);

AOI22xp33_ASAP7_75t_L g842 ( 
.A1(n_753),
.A2(n_516),
.B1(n_522),
.B2(n_524),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_683),
.B(n_575),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_748),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_683),
.B(n_575),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_635),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_SL g847 ( 
.A(n_623),
.B(n_575),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_711),
.B(n_576),
.Y(n_848)
);

AOI22xp33_ASAP7_75t_L g849 ( 
.A1(n_758),
.A2(n_524),
.B1(n_560),
.B2(n_553),
.Y(n_849)
);

BUFx6f_ASAP7_75t_L g850 ( 
.A(n_717),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_721),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_711),
.B(n_576),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_655),
.B(n_576),
.Y(n_853)
);

OAI22xp33_ASAP7_75t_L g854 ( 
.A1(n_726),
.A2(n_578),
.B1(n_522),
.B2(n_516),
.Y(n_854)
);

BUFx2_ASAP7_75t_L g855 ( 
.A(n_706),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_751),
.B(n_578),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_749),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_640),
.Y(n_858)
);

AOI22xp33_ASAP7_75t_L g859 ( 
.A1(n_735),
.A2(n_528),
.B1(n_553),
.B2(n_560),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_646),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_649),
.Y(n_861)
);

HB1xp67_ASAP7_75t_L g862 ( 
.A(n_706),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_SL g863 ( 
.A(n_612),
.B(n_578),
.Y(n_863)
);

AND2x4_ASAP7_75t_L g864 ( 
.A(n_718),
.B(n_587),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_657),
.Y(n_865)
);

AOI21x1_ASAP7_75t_L g866 ( 
.A1(n_593),
.A2(n_528),
.B(n_469),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_655),
.B(n_587),
.Y(n_867)
);

INVx3_ASAP7_75t_L g868 ( 
.A(n_666),
.Y(n_868)
);

AND2x6_ASAP7_75t_L g869 ( 
.A(n_678),
.B(n_587),
.Y(n_869)
);

HB1xp67_ASAP7_75t_L g870 ( 
.A(n_661),
.Y(n_870)
);

INVx5_ASAP7_75t_L g871 ( 
.A(n_651),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_759),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_677),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_690),
.B(n_587),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_680),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_699),
.B(n_566),
.Y(n_876)
);

INVx5_ASAP7_75t_L g877 ( 
.A(n_712),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_702),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_703),
.B(n_566),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_719),
.Y(n_880)
);

AOI22xp33_ASAP7_75t_L g881 ( 
.A1(n_596),
.A2(n_493),
.B1(n_471),
.B2(n_473),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_730),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_761),
.B(n_715),
.Y(n_883)
);

HB1xp67_ASAP7_75t_L g884 ( 
.A(n_726),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_761),
.B(n_566),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_686),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_750),
.B(n_574),
.Y(n_887)
);

INVx3_ASAP7_75t_L g888 ( 
.A(n_717),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_689),
.B(n_566),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_695),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_697),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_754),
.Y(n_892)
);

AOI22xp33_ASAP7_75t_L g893 ( 
.A1(n_659),
.A2(n_490),
.B1(n_471),
.B2(n_473),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_714),
.Y(n_894)
);

AOI22xp5_ASAP7_75t_L g895 ( 
.A1(n_665),
.A2(n_676),
.B1(n_726),
.B2(n_637),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_SL g896 ( 
.A(n_665),
.B(n_574),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_724),
.Y(n_897)
);

OAI22xp5_ASAP7_75t_SL g898 ( 
.A1(n_733),
.A2(n_16),
.B1(n_19),
.B2(n_20),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_SL g899 ( 
.A(n_707),
.B(n_570),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_676),
.B(n_574),
.Y(n_900)
);

AND2x6_ASAP7_75t_SL g901 ( 
.A(n_731),
.B(n_734),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_603),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_L g903 ( 
.A(n_611),
.B(n_568),
.Y(n_903)
);

NOR2xp33_ASAP7_75t_L g904 ( 
.A(n_608),
.B(n_568),
.Y(n_904)
);

NAND2x1p5_ASAP7_75t_L g905 ( 
.A(n_717),
.B(n_570),
.Y(n_905)
);

OAI22xp5_ASAP7_75t_L g906 ( 
.A1(n_679),
.A2(n_692),
.B1(n_732),
.B2(n_659),
.Y(n_906)
);

BUFx8_ASAP7_75t_L g907 ( 
.A(n_742),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_653),
.B(n_568),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_614),
.Y(n_909)
);

NOR2xp33_ASAP7_75t_L g910 ( 
.A(n_734),
.B(n_568),
.Y(n_910)
);

INVx5_ASAP7_75t_L g911 ( 
.A(n_712),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_632),
.B(n_619),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_653),
.B(n_570),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_638),
.Y(n_914)
);

NOR2xp33_ASAP7_75t_R g915 ( 
.A(n_712),
.B(n_115),
.Y(n_915)
);

AOI22xp33_ASAP7_75t_L g916 ( 
.A1(n_745),
.A2(n_490),
.B1(n_471),
.B2(n_507),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_682),
.B(n_570),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_654),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_L g919 ( 
.A(n_625),
.B(n_16),
.Y(n_919)
);

INVx3_ASAP7_75t_L g920 ( 
.A(n_717),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_597),
.B(n_490),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_707),
.B(n_486),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_669),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_707),
.B(n_486),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_707),
.B(n_486),
.Y(n_925)
);

BUFx2_ASAP7_75t_L g926 ( 
.A(n_670),
.Y(n_926)
);

AND2x6_ASAP7_75t_L g927 ( 
.A(n_704),
.B(n_574),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_708),
.A2(n_710),
.B(n_737),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_675),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_707),
.B(n_493),
.Y(n_930)
);

BUFx3_ASAP7_75t_L g931 ( 
.A(n_705),
.Y(n_931)
);

BUFx12f_ASAP7_75t_L g932 ( 
.A(n_747),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_707),
.B(n_493),
.Y(n_933)
);

CKINVDCx11_ASAP7_75t_R g934 ( 
.A(n_622),
.Y(n_934)
);

AOI22xp33_ASAP7_75t_L g935 ( 
.A1(n_745),
.A2(n_484),
.B1(n_507),
.B2(n_506),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_624),
.Y(n_936)
);

OAI21xp5_ASAP7_75t_L g937 ( 
.A1(n_628),
.A2(n_484),
.B(n_507),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_667),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_684),
.B(n_484),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_752),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_694),
.Y(n_941)
);

NAND3xp33_ASAP7_75t_SL g942 ( 
.A(n_743),
.B(n_469),
.C(n_473),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_639),
.B(n_663),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_752),
.Y(n_944)
);

BUFx3_ASAP7_75t_L g945 ( 
.A(n_747),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_636),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_627),
.B(n_469),
.Y(n_947)
);

A2O1A1Ixp33_ASAP7_75t_L g948 ( 
.A1(n_644),
.A2(n_506),
.B(n_498),
.C(n_497),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_SL g949 ( 
.A(n_737),
.B(n_574),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_647),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_812),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_928),
.A2(n_658),
.B(n_656),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_883),
.B(n_688),
.Y(n_953)
);

OAI22xp5_ASAP7_75t_L g954 ( 
.A1(n_840),
.A2(n_746),
.B1(n_720),
.B2(n_700),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_830),
.B(n_739),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_815),
.Y(n_956)
);

BUFx4f_ASAP7_75t_L g957 ( 
.A(n_811),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_808),
.B(n_720),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_L g959 ( 
.A(n_830),
.B(n_725),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_808),
.B(n_660),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_L g961 ( 
.A(n_800),
.B(n_738),
.Y(n_961)
);

A2O1A1Ixp33_ASAP7_75t_L g962 ( 
.A1(n_895),
.A2(n_698),
.B(n_723),
.C(n_740),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_SL g963 ( 
.A(n_938),
.B(n_763),
.Y(n_963)
);

INVxp67_ASAP7_75t_L g964 ( 
.A(n_801),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_870),
.Y(n_965)
);

NAND2x1_ASAP7_75t_L g966 ( 
.A(n_773),
.B(n_693),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_SL g967 ( 
.A(n_941),
.B(n_763),
.Y(n_967)
);

OR2x2_ASAP7_75t_L g968 ( 
.A(n_803),
.B(n_727),
.Y(n_968)
);

NOR3xp33_ASAP7_75t_SL g969 ( 
.A(n_898),
.B(n_762),
.C(n_755),
.Y(n_969)
);

AO22x1_ASAP7_75t_L g970 ( 
.A1(n_919),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_970)
);

A2O1A1Ixp33_ASAP7_75t_L g971 ( 
.A1(n_919),
.A2(n_728),
.B(n_673),
.C(n_762),
.Y(n_971)
);

O2A1O1Ixp33_ASAP7_75t_L g972 ( 
.A1(n_798),
.A2(n_755),
.B(n_506),
.C(n_498),
.Y(n_972)
);

O2A1O1Ixp33_ASAP7_75t_SL g973 ( 
.A1(n_949),
.A2(n_498),
.B(n_497),
.C(n_479),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_870),
.Y(n_974)
);

O2A1O1Ixp33_ASAP7_75t_L g975 ( 
.A1(n_798),
.A2(n_497),
.B(n_479),
.C(n_28),
.Y(n_975)
);

A2O1A1Ixp33_ASAP7_75t_L g976 ( 
.A1(n_768),
.A2(n_479),
.B(n_401),
.C(n_28),
.Y(n_976)
);

NAND3xp33_ASAP7_75t_SL g977 ( 
.A(n_818),
.B(n_25),
.C(n_27),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_873),
.Y(n_978)
);

NOR3xp33_ASAP7_75t_L g979 ( 
.A(n_783),
.B(n_30),
.C(n_31),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_926),
.B(n_95),
.Y(n_980)
);

BUFx12f_ASAP7_75t_L g981 ( 
.A(n_778),
.Y(n_981)
);

O2A1O1Ixp33_ASAP7_75t_L g982 ( 
.A1(n_943),
.A2(n_30),
.B(n_37),
.C(n_38),
.Y(n_982)
);

BUFx6f_ASAP7_75t_L g983 ( 
.A(n_850),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_792),
.B(n_37),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_912),
.B(n_39),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_931),
.B(n_114),
.Y(n_986)
);

AND2x4_ASAP7_75t_L g987 ( 
.A(n_832),
.B(n_834),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_844),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_878),
.Y(n_989)
);

NAND2x1p5_ASAP7_75t_L g990 ( 
.A(n_837),
.B(n_110),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_880),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_856),
.B(n_41),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_839),
.A2(n_118),
.B(n_143),
.Y(n_993)
);

AOI22xp33_ASAP7_75t_L g994 ( 
.A1(n_813),
.A2(n_42),
.B1(n_43),
.B2(n_45),
.Y(n_994)
);

BUFx8_ASAP7_75t_L g995 ( 
.A(n_766),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_882),
.Y(n_996)
);

AOI22xp5_ASAP7_75t_L g997 ( 
.A1(n_813),
.A2(n_863),
.B1(n_810),
.B2(n_884),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_857),
.Y(n_998)
);

NOR2x1_ASAP7_75t_R g999 ( 
.A(n_797),
.B(n_851),
.Y(n_999)
);

NOR2xp67_ASAP7_75t_L g1000 ( 
.A(n_769),
.B(n_119),
.Y(n_1000)
);

BUFx12f_ASAP7_75t_L g1001 ( 
.A(n_778),
.Y(n_1001)
);

OAI22x1_ASAP7_75t_L g1002 ( 
.A1(n_855),
.A2(n_42),
.B1(n_43),
.B2(n_46),
.Y(n_1002)
);

BUFx4f_ASAP7_75t_L g1003 ( 
.A(n_932),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_L g1004 ( 
.A(n_901),
.B(n_51),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_L g1005 ( 
.A(n_827),
.B(n_58),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_841),
.A2(n_68),
.B(n_87),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_784),
.Y(n_1007)
);

INVx6_ASAP7_75t_L g1008 ( 
.A(n_907),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_843),
.A2(n_92),
.B(n_103),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_936),
.B(n_120),
.Y(n_1010)
);

INVx4_ASAP7_75t_L g1011 ( 
.A(n_765),
.Y(n_1011)
);

BUFx6f_ASAP7_75t_SL g1012 ( 
.A(n_770),
.Y(n_1012)
);

O2A1O1Ixp33_ASAP7_75t_L g1013 ( 
.A1(n_789),
.A2(n_127),
.B(n_129),
.C(n_137),
.Y(n_1013)
);

INVxp67_ASAP7_75t_SL g1014 ( 
.A(n_765),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_946),
.B(n_138),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_950),
.B(n_140),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_767),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_845),
.A2(n_142),
.B(n_151),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_848),
.A2(n_900),
.B(n_896),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_835),
.B(n_894),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_835),
.B(n_897),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_829),
.A2(n_838),
.B(n_885),
.Y(n_1022)
);

O2A1O1Ixp33_ASAP7_75t_L g1023 ( 
.A1(n_789),
.A2(n_862),
.B(n_906),
.C(n_887),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_922),
.A2(n_930),
.B(n_933),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_771),
.Y(n_1025)
);

O2A1O1Ixp33_ASAP7_75t_L g1026 ( 
.A1(n_862),
.A2(n_884),
.B(n_861),
.C(n_772),
.Y(n_1026)
);

A2O1A1Ixp33_ASAP7_75t_SL g1027 ( 
.A1(n_802),
.A2(n_910),
.B(n_903),
.C(n_904),
.Y(n_1027)
);

NAND2xp33_ASAP7_75t_SL g1028 ( 
.A(n_915),
.B(n_818),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_777),
.Y(n_1029)
);

AOI21x1_ASAP7_75t_L g1030 ( 
.A1(n_866),
.A2(n_921),
.B(n_852),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_787),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_924),
.A2(n_925),
.B(n_889),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_872),
.Y(n_1033)
);

OAI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_840),
.A2(n_828),
.B(n_847),
.Y(n_1034)
);

AO21x1_ASAP7_75t_L g1035 ( 
.A1(n_910),
.A2(n_802),
.B(n_903),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_SL g1036 ( 
.A(n_776),
.B(n_788),
.Y(n_1036)
);

O2A1O1Ixp33_ASAP7_75t_SL g1037 ( 
.A1(n_949),
.A2(n_814),
.B(n_795),
.C(n_820),
.Y(n_1037)
);

NOR2xp33_ASAP7_75t_L g1038 ( 
.A(n_791),
.B(n_809),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_816),
.B(n_824),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_917),
.A2(n_786),
.B(n_780),
.Y(n_1040)
);

BUFx2_ASAP7_75t_L g1041 ( 
.A(n_907),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_785),
.B(n_853),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_785),
.B(n_819),
.Y(n_1043)
);

NOR3xp33_ASAP7_75t_SL g1044 ( 
.A(n_825),
.B(n_860),
.C(n_865),
.Y(n_1044)
);

NOR2xp33_ASAP7_75t_L g1045 ( 
.A(n_833),
.B(n_846),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_858),
.Y(n_1046)
);

AOI22x1_ASAP7_75t_L g1047 ( 
.A1(n_775),
.A2(n_940),
.B1(n_944),
.B2(n_947),
.Y(n_1047)
);

O2A1O1Ixp33_ASAP7_75t_L g1048 ( 
.A1(n_854),
.A2(n_867),
.B(n_904),
.C(n_892),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_793),
.Y(n_1049)
);

BUFx12f_ASAP7_75t_L g1050 ( 
.A(n_934),
.Y(n_1050)
);

AND2x2_ASAP7_75t_L g1051 ( 
.A(n_790),
.B(n_764),
.Y(n_1051)
);

BUFx6f_ASAP7_75t_L g1052 ( 
.A(n_850),
.Y(n_1052)
);

INVx2_ASAP7_75t_SL g1053 ( 
.A(n_864),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_806),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_899),
.A2(n_908),
.B(n_913),
.Y(n_1055)
);

A2O1A1Ixp33_ASAP7_75t_L g1056 ( 
.A1(n_807),
.A2(n_805),
.B(n_799),
.C(n_826),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_914),
.Y(n_1057)
);

NAND2xp33_ASAP7_75t_SL g1058 ( 
.A(n_915),
.B(n_850),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_790),
.B(n_774),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_L g1060 ( 
.A(n_864),
.B(n_795),
.Y(n_1060)
);

A2O1A1Ixp33_ASAP7_75t_SL g1061 ( 
.A1(n_937),
.A2(n_888),
.B(n_920),
.C(n_868),
.Y(n_1061)
);

INVx6_ASAP7_75t_L g1062 ( 
.A(n_794),
.Y(n_1062)
);

OAI22xp5_ASAP7_75t_L g1063 ( 
.A1(n_774),
.A2(n_804),
.B1(n_893),
.B2(n_859),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_SL g1064 ( 
.A(n_765),
.B(n_821),
.Y(n_1064)
);

INVx1_ASAP7_75t_SL g1065 ( 
.A(n_765),
.Y(n_1065)
);

HB1xp67_ASAP7_75t_L g1066 ( 
.A(n_821),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_831),
.B(n_868),
.Y(n_1067)
);

NOR2xp33_ASAP7_75t_L g1068 ( 
.A(n_831),
.B(n_814),
.Y(n_1068)
);

INVxp67_ASAP7_75t_SL g1069 ( 
.A(n_821),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_899),
.A2(n_939),
.B(n_837),
.Y(n_1070)
);

O2A1O1Ixp33_ASAP7_75t_L g1071 ( 
.A1(n_854),
.A2(n_876),
.B(n_879),
.C(n_874),
.Y(n_1071)
);

OAI21xp33_ASAP7_75t_L g1072 ( 
.A1(n_804),
.A2(n_842),
.B(n_849),
.Y(n_1072)
);

A2O1A1Ixp33_ASAP7_75t_L g1073 ( 
.A1(n_781),
.A2(n_796),
.B(n_945),
.C(n_886),
.Y(n_1073)
);

O2A1O1Ixp33_ASAP7_75t_SL g1074 ( 
.A1(n_782),
.A2(n_847),
.B(n_836),
.C(n_948),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_837),
.A2(n_871),
.B(n_911),
.Y(n_1075)
);

AOI21x1_ASAP7_75t_L g1076 ( 
.A1(n_836),
.A2(n_822),
.B(n_929),
.Y(n_1076)
);

AOI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_794),
.A2(n_869),
.B1(n_817),
.B2(n_779),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_902),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_817),
.B(n_891),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_SL g1080 ( 
.A(n_821),
.B(n_871),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_817),
.B(n_890),
.Y(n_1081)
);

BUFx2_ASAP7_75t_L g1082 ( 
.A(n_875),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_817),
.B(n_773),
.Y(n_1083)
);

NOR2x1_ASAP7_75t_L g1084 ( 
.A(n_823),
.B(n_888),
.Y(n_1084)
);

AOI22xp5_ASAP7_75t_L g1085 ( 
.A1(n_869),
.A2(n_817),
.B1(n_779),
.B2(n_918),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_SL g1086 ( 
.A(n_837),
.B(n_877),
.Y(n_1086)
);

AOI22xp5_ASAP7_75t_L g1087 ( 
.A1(n_869),
.A2(n_779),
.B1(n_823),
.B2(n_923),
.Y(n_1087)
);

AO21x1_ASAP7_75t_L g1088 ( 
.A1(n_905),
.A2(n_909),
.B(n_869),
.Y(n_1088)
);

NAND2xp33_ASAP7_75t_SL g1089 ( 
.A(n_850),
.B(n_920),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_905),
.Y(n_1090)
);

INVx2_ASAP7_75t_SL g1091 ( 
.A(n_869),
.Y(n_1091)
);

INVx3_ASAP7_75t_L g1092 ( 
.A(n_871),
.Y(n_1092)
);

OAI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_881),
.A2(n_779),
.B(n_893),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_779),
.B(n_881),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_871),
.A2(n_911),
.B(n_877),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_916),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_L g1097 ( 
.A(n_942),
.B(n_842),
.Y(n_1097)
);

NOR2xp33_ASAP7_75t_SL g1098 ( 
.A(n_1007),
.B(n_877),
.Y(n_1098)
);

OAI21x1_ASAP7_75t_L g1099 ( 
.A1(n_1070),
.A2(n_942),
.B(n_916),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_1022),
.A2(n_877),
.B(n_911),
.Y(n_1100)
);

INVx4_ASAP7_75t_SL g1101 ( 
.A(n_983),
.Y(n_1101)
);

INVxp67_ASAP7_75t_SL g1102 ( 
.A(n_964),
.Y(n_1102)
);

OAI22x1_ASAP7_75t_L g1103 ( 
.A1(n_959),
.A2(n_911),
.B1(n_935),
.B2(n_849),
.Y(n_1103)
);

INVx3_ASAP7_75t_L g1104 ( 
.A(n_1092),
.Y(n_1104)
);

OAI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_1097),
.A2(n_859),
.B(n_935),
.Y(n_1105)
);

OA21x2_ASAP7_75t_L g1106 ( 
.A1(n_1034),
.A2(n_927),
.B(n_1019),
.Y(n_1106)
);

OAI21x1_ASAP7_75t_L g1107 ( 
.A1(n_952),
.A2(n_927),
.B(n_1076),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_1020),
.B(n_927),
.Y(n_1108)
);

NAND2xp33_ASAP7_75t_L g1109 ( 
.A(n_969),
.B(n_953),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_978),
.Y(n_1110)
);

AND2x4_ASAP7_75t_L g1111 ( 
.A(n_987),
.B(n_927),
.Y(n_1111)
);

INVxp67_ASAP7_75t_SL g1112 ( 
.A(n_965),
.Y(n_1112)
);

OAI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_1034),
.A2(n_927),
.B(n_1056),
.Y(n_1113)
);

AND2x2_ASAP7_75t_L g1114 ( 
.A(n_985),
.B(n_1082),
.Y(n_1114)
);

AND2x2_ASAP7_75t_L g1115 ( 
.A(n_961),
.B(n_974),
.Y(n_1115)
);

AO31x2_ASAP7_75t_L g1116 ( 
.A1(n_1035),
.A2(n_1088),
.A3(n_954),
.B(n_1063),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_989),
.Y(n_1117)
);

OAI21x1_ASAP7_75t_L g1118 ( 
.A1(n_1024),
.A2(n_1030),
.B(n_1032),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_1093),
.A2(n_1040),
.B(n_1027),
.Y(n_1119)
);

BUFx2_ASAP7_75t_L g1120 ( 
.A(n_987),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_1020),
.B(n_1021),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_1093),
.A2(n_960),
.B(n_1021),
.Y(n_1122)
);

OR2x2_ASAP7_75t_L g1123 ( 
.A(n_984),
.B(n_1039),
.Y(n_1123)
);

AOI22xp33_ASAP7_75t_L g1124 ( 
.A1(n_979),
.A2(n_954),
.B1(n_1072),
.B2(n_977),
.Y(n_1124)
);

OAI21x1_ASAP7_75t_L g1125 ( 
.A1(n_1055),
.A2(n_1047),
.B(n_1079),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_960),
.A2(n_962),
.B(n_1063),
.Y(n_1126)
);

OAI21x1_ASAP7_75t_L g1127 ( 
.A1(n_1081),
.A2(n_1095),
.B(n_1075),
.Y(n_1127)
);

OAI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_958),
.A2(n_1023),
.B(n_1094),
.Y(n_1128)
);

AOI21x1_ASAP7_75t_L g1129 ( 
.A1(n_1083),
.A2(n_1042),
.B(n_966),
.Y(n_1129)
);

AOI22xp5_ASAP7_75t_L g1130 ( 
.A1(n_1028),
.A2(n_980),
.B1(n_955),
.B2(n_1051),
.Y(n_1130)
);

NOR2xp33_ASAP7_75t_L g1131 ( 
.A(n_963),
.B(n_967),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_958),
.B(n_1043),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_SL g1133 ( 
.A(n_957),
.B(n_1038),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_1042),
.A2(n_1048),
.B(n_1043),
.Y(n_1134)
);

OAI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_1094),
.A2(n_997),
.B(n_971),
.Y(n_1135)
);

BUFx12f_ASAP7_75t_L g1136 ( 
.A(n_981),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_1071),
.A2(n_1037),
.B(n_1074),
.Y(n_1137)
);

OA21x2_ASAP7_75t_L g1138 ( 
.A1(n_1085),
.A2(n_1073),
.B(n_976),
.Y(n_1138)
);

AO31x2_ASAP7_75t_L g1139 ( 
.A1(n_1096),
.A2(n_1068),
.A3(n_1060),
.B(n_1059),
.Y(n_1139)
);

OAI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_1013),
.A2(n_972),
.B(n_1087),
.Y(n_1140)
);

INVx3_ASAP7_75t_L g1141 ( 
.A(n_1092),
.Y(n_1141)
);

HB1xp67_ASAP7_75t_L g1142 ( 
.A(n_1066),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_991),
.Y(n_1143)
);

AO31x2_ASAP7_75t_L g1144 ( 
.A1(n_1010),
.A2(n_1016),
.A3(n_1015),
.B(n_1006),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_1045),
.B(n_996),
.Y(n_1145)
);

AOI21x1_ASAP7_75t_L g1146 ( 
.A1(n_992),
.A2(n_1064),
.B(n_1091),
.Y(n_1146)
);

OAI21x1_ASAP7_75t_L g1147 ( 
.A1(n_1086),
.A2(n_1077),
.B(n_993),
.Y(n_1147)
);

AO31x2_ASAP7_75t_L g1148 ( 
.A1(n_1009),
.A2(n_1018),
.A3(n_1067),
.B(n_1002),
.Y(n_1148)
);

OAI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_1061),
.A2(n_975),
.B(n_973),
.Y(n_1149)
);

BUFx2_ASAP7_75t_L g1150 ( 
.A(n_995),
.Y(n_1150)
);

OAI21x1_ASAP7_75t_L g1151 ( 
.A1(n_1080),
.A2(n_990),
.B(n_1084),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1017),
.B(n_1025),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1029),
.Y(n_1153)
);

INVxp67_ASAP7_75t_SL g1154 ( 
.A(n_983),
.Y(n_1154)
);

AND2x4_ASAP7_75t_L g1155 ( 
.A(n_1053),
.B(n_1044),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_1058),
.A2(n_1089),
.B(n_1069),
.Y(n_1156)
);

BUFx3_ASAP7_75t_L g1157 ( 
.A(n_1062),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_SL g1158 ( 
.A1(n_990),
.A2(n_986),
.B(n_1014),
.Y(n_1158)
);

OR2x2_ASAP7_75t_L g1159 ( 
.A(n_1031),
.B(n_1046),
.Y(n_1159)
);

INVx2_ASAP7_75t_SL g1160 ( 
.A(n_957),
.Y(n_1160)
);

OAI21xp5_ASAP7_75t_SL g1161 ( 
.A1(n_1004),
.A2(n_994),
.B(n_982),
.Y(n_1161)
);

OAI22xp5_ASAP7_75t_L g1162 ( 
.A1(n_968),
.A2(n_1057),
.B1(n_956),
.B2(n_1033),
.Y(n_1162)
);

NAND3x1_ASAP7_75t_L g1163 ( 
.A(n_1005),
.B(n_1001),
.C(n_970),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1065),
.A2(n_951),
.B(n_988),
.Y(n_1164)
);

OAI21x1_ASAP7_75t_L g1165 ( 
.A1(n_1026),
.A2(n_1090),
.B(n_998),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_SL g1166 ( 
.A1(n_983),
.A2(n_1052),
.B(n_1011),
.Y(n_1166)
);

OAI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_1078),
.A2(n_1003),
.B1(n_1065),
.B2(n_1000),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_1036),
.A2(n_1011),
.B(n_1052),
.Y(n_1168)
);

BUFx2_ASAP7_75t_L g1169 ( 
.A(n_995),
.Y(n_1169)
);

NAND2x1p5_ASAP7_75t_L g1170 ( 
.A(n_1052),
.B(n_1003),
.Y(n_1170)
);

AO21x2_ASAP7_75t_L g1171 ( 
.A1(n_1049),
.A2(n_1054),
.B(n_999),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_SL g1172 ( 
.A(n_1050),
.B(n_1041),
.Y(n_1172)
);

OAI21x1_ASAP7_75t_SL g1173 ( 
.A1(n_1062),
.A2(n_1012),
.B(n_1008),
.Y(n_1173)
);

NAND3xp33_ASAP7_75t_SL g1174 ( 
.A(n_1012),
.B(n_643),
.C(n_895),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1008),
.Y(n_1175)
);

OAI21x1_ASAP7_75t_L g1176 ( 
.A1(n_1070),
.A2(n_866),
.B(n_952),
.Y(n_1176)
);

NAND2xp33_ASAP7_75t_L g1177 ( 
.A(n_969),
.B(n_642),
.Y(n_1177)
);

O2A1O1Ixp5_ASAP7_75t_SL g1178 ( 
.A1(n_954),
.A2(n_887),
.B(n_505),
.C(n_523),
.Y(n_1178)
);

OA22x2_ASAP7_75t_L g1179 ( 
.A1(n_1002),
.A2(n_466),
.B1(n_898),
.B2(n_417),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1020),
.B(n_1021),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1020),
.B(n_1021),
.Y(n_1181)
);

OAI21x1_ASAP7_75t_L g1182 ( 
.A1(n_1070),
.A2(n_866),
.B(n_952),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_978),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_978),
.Y(n_1184)
);

OAI21xp5_ASAP7_75t_SL g1185 ( 
.A1(n_979),
.A2(n_466),
.B(n_612),
.Y(n_1185)
);

HB1xp67_ASAP7_75t_L g1186 ( 
.A(n_964),
.Y(n_1186)
);

BUFx4f_ASAP7_75t_SL g1187 ( 
.A(n_981),
.Y(n_1187)
);

BUFx2_ASAP7_75t_L g1188 ( 
.A(n_964),
.Y(n_1188)
);

NAND2x1p5_ASAP7_75t_L g1189 ( 
.A(n_1011),
.B(n_773),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_978),
.Y(n_1190)
);

OAI21x1_ASAP7_75t_L g1191 ( 
.A1(n_1070),
.A2(n_866),
.B(n_952),
.Y(n_1191)
);

OR2x2_ASAP7_75t_L g1192 ( 
.A(n_965),
.B(n_800),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_SL g1193 ( 
.A(n_961),
.B(n_643),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1020),
.B(n_1021),
.Y(n_1194)
);

AOI21x1_ASAP7_75t_L g1195 ( 
.A1(n_1030),
.A2(n_1076),
.B(n_1070),
.Y(n_1195)
);

O2A1O1Ixp5_ASAP7_75t_L g1196 ( 
.A1(n_1035),
.A2(n_954),
.B(n_637),
.C(n_1097),
.Y(n_1196)
);

AOI21x1_ASAP7_75t_SL g1197 ( 
.A1(n_958),
.A2(n_953),
.B(n_984),
.Y(n_1197)
);

OAI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1097),
.A2(n_1034),
.B(n_1056),
.Y(n_1198)
);

BUFx2_ASAP7_75t_L g1199 ( 
.A(n_964),
.Y(n_1199)
);

OA21x2_ASAP7_75t_L g1200 ( 
.A1(n_1034),
.A2(n_1019),
.B(n_1093),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1020),
.B(n_1021),
.Y(n_1201)
);

AOI21x1_ASAP7_75t_SL g1202 ( 
.A1(n_958),
.A2(n_953),
.B(n_984),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_978),
.Y(n_1203)
);

OR2x2_ASAP7_75t_L g1204 ( 
.A(n_965),
.B(n_800),
.Y(n_1204)
);

OAI21x1_ASAP7_75t_L g1205 ( 
.A1(n_1070),
.A2(n_866),
.B(n_952),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_978),
.Y(n_1206)
);

OR2x2_ASAP7_75t_L g1207 ( 
.A(n_965),
.B(n_800),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1020),
.B(n_1021),
.Y(n_1208)
);

AND2x4_ASAP7_75t_L g1209 ( 
.A(n_987),
.B(n_811),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_978),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1022),
.A2(n_883),
.B(n_1019),
.Y(n_1211)
);

NAND3xp33_ASAP7_75t_L g1212 ( 
.A(n_979),
.B(n_895),
.C(n_499),
.Y(n_1212)
);

AO31x2_ASAP7_75t_L g1213 ( 
.A1(n_1035),
.A2(n_1088),
.A3(n_1097),
.B(n_954),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1020),
.B(n_1021),
.Y(n_1214)
);

HB1xp67_ASAP7_75t_L g1215 ( 
.A(n_964),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_L g1216 ( 
.A1(n_1070),
.A2(n_866),
.B(n_952),
.Y(n_1216)
);

NAND3x1_ASAP7_75t_L g1217 ( 
.A(n_979),
.B(n_466),
.C(n_1004),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1022),
.A2(n_1040),
.B(n_737),
.Y(n_1218)
);

NOR2xp33_ASAP7_75t_L g1219 ( 
.A(n_959),
.B(n_315),
.Y(n_1219)
);

INVx3_ASAP7_75t_L g1220 ( 
.A(n_1092),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1020),
.B(n_1021),
.Y(n_1221)
);

OAI21x1_ASAP7_75t_L g1222 ( 
.A1(n_1070),
.A2(n_866),
.B(n_952),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_SL g1223 ( 
.A(n_961),
.B(n_643),
.Y(n_1223)
);

OAI21x1_ASAP7_75t_L g1224 ( 
.A1(n_1070),
.A2(n_866),
.B(n_952),
.Y(n_1224)
);

OAI21x1_ASAP7_75t_L g1225 ( 
.A1(n_1070),
.A2(n_866),
.B(n_952),
.Y(n_1225)
);

NAND2x1p5_ASAP7_75t_L g1226 ( 
.A(n_1011),
.B(n_773),
.Y(n_1226)
);

OAI22xp5_ASAP7_75t_L g1227 ( 
.A1(n_1063),
.A2(n_633),
.B1(n_648),
.B2(n_840),
.Y(n_1227)
);

INVxp67_ASAP7_75t_SL g1228 ( 
.A(n_964),
.Y(n_1228)
);

XOR2xp5_ASAP7_75t_L g1229 ( 
.A(n_1007),
.B(n_513),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1020),
.B(n_1021),
.Y(n_1230)
);

A2O1A1Ixp33_ASAP7_75t_L g1231 ( 
.A1(n_1072),
.A2(n_895),
.B(n_618),
.C(n_954),
.Y(n_1231)
);

AOI211x1_ASAP7_75t_L g1232 ( 
.A1(n_970),
.A2(n_612),
.B(n_1072),
.C(n_733),
.Y(n_1232)
);

NOR2xp67_ASAP7_75t_L g1233 ( 
.A(n_1007),
.B(n_769),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_978),
.Y(n_1234)
);

A2O1A1Ixp33_ASAP7_75t_L g1235 ( 
.A1(n_1072),
.A2(n_895),
.B(n_618),
.C(n_954),
.Y(n_1235)
);

AOI21xp5_ASAP7_75t_SL g1236 ( 
.A1(n_1063),
.A2(n_813),
.B(n_1093),
.Y(n_1236)
);

HB1xp67_ASAP7_75t_L g1237 ( 
.A(n_964),
.Y(n_1237)
);

NOR4xp25_ASAP7_75t_L g1238 ( 
.A(n_977),
.B(n_982),
.C(n_612),
.D(n_1072),
.Y(n_1238)
);

OAI21x1_ASAP7_75t_L g1239 ( 
.A1(n_1107),
.A2(n_1182),
.B(n_1176),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1159),
.Y(n_1240)
);

OAI22xp33_ASAP7_75t_L g1241 ( 
.A1(n_1227),
.A2(n_1185),
.B1(n_1179),
.B2(n_1212),
.Y(n_1241)
);

O2A1O1Ixp33_ASAP7_75t_L g1242 ( 
.A1(n_1231),
.A2(n_1235),
.B(n_1161),
.C(n_1193),
.Y(n_1242)
);

BUFx2_ASAP7_75t_L g1243 ( 
.A(n_1188),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1152),
.Y(n_1244)
);

OR2x6_ASAP7_75t_L g1245 ( 
.A(n_1158),
.B(n_1236),
.Y(n_1245)
);

INVx2_ASAP7_75t_L g1246 ( 
.A(n_1110),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1152),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1132),
.B(n_1121),
.Y(n_1248)
);

O2A1O1Ixp33_ASAP7_75t_SL g1249 ( 
.A1(n_1227),
.A2(n_1105),
.B(n_1132),
.C(n_1108),
.Y(n_1249)
);

INVx3_ASAP7_75t_L g1250 ( 
.A(n_1111),
.Y(n_1250)
);

OA21x2_ASAP7_75t_L g1251 ( 
.A1(n_1196),
.A2(n_1119),
.B(n_1137),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1143),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_1190),
.Y(n_1253)
);

AND2x4_ASAP7_75t_L g1254 ( 
.A(n_1111),
.B(n_1155),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1206),
.Y(n_1255)
);

O2A1O1Ixp33_ASAP7_75t_SL g1256 ( 
.A1(n_1105),
.A2(n_1108),
.B(n_1181),
.C(n_1194),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_1117),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_1153),
.Y(n_1258)
);

OAI21x1_ASAP7_75t_L g1259 ( 
.A1(n_1191),
.A2(n_1222),
.B(n_1216),
.Y(n_1259)
);

AND2x2_ASAP7_75t_L g1260 ( 
.A(n_1114),
.B(n_1115),
.Y(n_1260)
);

AOI22xp33_ASAP7_75t_L g1261 ( 
.A1(n_1124),
.A2(n_1179),
.B1(n_1198),
.B2(n_1109),
.Y(n_1261)
);

AND2x4_ASAP7_75t_L g1262 ( 
.A(n_1155),
.B(n_1104),
.Y(n_1262)
);

BUFx12f_ASAP7_75t_L g1263 ( 
.A(n_1136),
.Y(n_1263)
);

OA21x2_ASAP7_75t_L g1264 ( 
.A1(n_1119),
.A2(n_1137),
.B(n_1140),
.Y(n_1264)
);

AOI22xp5_ASAP7_75t_L g1265 ( 
.A1(n_1219),
.A2(n_1217),
.B1(n_1174),
.B2(n_1223),
.Y(n_1265)
);

NAND2x1p5_ASAP7_75t_L g1266 ( 
.A(n_1104),
.B(n_1141),
.Y(n_1266)
);

INVx2_ASAP7_75t_SL g1267 ( 
.A(n_1157),
.Y(n_1267)
);

OAI21x1_ASAP7_75t_L g1268 ( 
.A1(n_1205),
.A2(n_1225),
.B(n_1224),
.Y(n_1268)
);

NOR2xp33_ASAP7_75t_L g1269 ( 
.A(n_1131),
.B(n_1123),
.Y(n_1269)
);

AOI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1211),
.A2(n_1218),
.B(n_1100),
.Y(n_1270)
);

AND2x4_ASAP7_75t_L g1271 ( 
.A(n_1141),
.B(n_1220),
.Y(n_1271)
);

NOR2xp67_ASAP7_75t_L g1272 ( 
.A(n_1186),
.B(n_1215),
.Y(n_1272)
);

HB1xp67_ASAP7_75t_L g1273 ( 
.A(n_1237),
.Y(n_1273)
);

OAI21x1_ASAP7_75t_SL g1274 ( 
.A1(n_1130),
.A2(n_1128),
.B(n_1167),
.Y(n_1274)
);

INVx5_ASAP7_75t_L g1275 ( 
.A(n_1220),
.Y(n_1275)
);

BUFx8_ASAP7_75t_SL g1276 ( 
.A(n_1150),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_1187),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_1183),
.Y(n_1278)
);

OA21x2_ASAP7_75t_L g1279 ( 
.A1(n_1140),
.A2(n_1118),
.B(n_1211),
.Y(n_1279)
);

OAI21x1_ASAP7_75t_L g1280 ( 
.A1(n_1195),
.A2(n_1125),
.B(n_1100),
.Y(n_1280)
);

AND2x4_ASAP7_75t_L g1281 ( 
.A(n_1171),
.B(n_1184),
.Y(n_1281)
);

OAI21x1_ASAP7_75t_L g1282 ( 
.A1(n_1127),
.A2(n_1099),
.B(n_1147),
.Y(n_1282)
);

OAI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1134),
.A2(n_1178),
.B(n_1122),
.Y(n_1283)
);

AOI221xp5_ASAP7_75t_L g1284 ( 
.A1(n_1238),
.A2(n_1232),
.B1(n_1198),
.B2(n_1126),
.C(n_1128),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1203),
.Y(n_1285)
);

OAI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1134),
.A2(n_1122),
.B(n_1126),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1210),
.Y(n_1287)
);

NOR2x1_ASAP7_75t_R g1288 ( 
.A(n_1169),
.B(n_1120),
.Y(n_1288)
);

CKINVDCx20_ASAP7_75t_R g1289 ( 
.A(n_1229),
.Y(n_1289)
);

OAI21x1_ASAP7_75t_L g1290 ( 
.A1(n_1129),
.A2(n_1113),
.B(n_1146),
.Y(n_1290)
);

INVx2_ASAP7_75t_L g1291 ( 
.A(n_1234),
.Y(n_1291)
);

BUFx3_ASAP7_75t_L g1292 ( 
.A(n_1199),
.Y(n_1292)
);

AO21x2_ASAP7_75t_L g1293 ( 
.A1(n_1113),
.A2(n_1149),
.B(n_1135),
.Y(n_1293)
);

HB1xp67_ASAP7_75t_L g1294 ( 
.A(n_1192),
.Y(n_1294)
);

INVxp67_ASAP7_75t_L g1295 ( 
.A(n_1204),
.Y(n_1295)
);

AO22x2_ASAP7_75t_L g1296 ( 
.A1(n_1162),
.A2(n_1230),
.B1(n_1208),
.B2(n_1201),
.Y(n_1296)
);

OAI21x1_ASAP7_75t_L g1297 ( 
.A1(n_1197),
.A2(n_1202),
.B(n_1164),
.Y(n_1297)
);

NOR2xp33_ASAP7_75t_L g1298 ( 
.A(n_1180),
.B(n_1208),
.Y(n_1298)
);

BUFx3_ASAP7_75t_L g1299 ( 
.A(n_1209),
.Y(n_1299)
);

AO31x2_ASAP7_75t_L g1300 ( 
.A1(n_1103),
.A2(n_1164),
.A3(n_1181),
.B(n_1230),
.Y(n_1300)
);

INVx1_ASAP7_75t_SL g1301 ( 
.A(n_1207),
.Y(n_1301)
);

OAI21x1_ASAP7_75t_L g1302 ( 
.A1(n_1151),
.A2(n_1165),
.B(n_1106),
.Y(n_1302)
);

BUFx2_ASAP7_75t_L g1303 ( 
.A(n_1102),
.Y(n_1303)
);

AND2x2_ASAP7_75t_L g1304 ( 
.A(n_1142),
.B(n_1209),
.Y(n_1304)
);

AND2x4_ASAP7_75t_L g1305 ( 
.A(n_1171),
.B(n_1101),
.Y(n_1305)
);

BUFx6f_ASAP7_75t_L g1306 ( 
.A(n_1170),
.Y(n_1306)
);

AOI22xp33_ASAP7_75t_L g1307 ( 
.A1(n_1138),
.A2(n_1221),
.B1(n_1201),
.B2(n_1194),
.Y(n_1307)
);

OR2x6_ASAP7_75t_L g1308 ( 
.A(n_1156),
.B(n_1173),
.Y(n_1308)
);

CKINVDCx11_ASAP7_75t_R g1309 ( 
.A(n_1175),
.Y(n_1309)
);

AO22x1_ASAP7_75t_L g1310 ( 
.A1(n_1228),
.A2(n_1145),
.B1(n_1112),
.B2(n_1160),
.Y(n_1310)
);

OAI21x1_ASAP7_75t_L g1311 ( 
.A1(n_1106),
.A2(n_1200),
.B(n_1138),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1133),
.B(n_1233),
.Y(n_1312)
);

BUFx4f_ASAP7_75t_SL g1313 ( 
.A(n_1172),
.Y(n_1313)
);

INVx3_ASAP7_75t_L g1314 ( 
.A(n_1189),
.Y(n_1314)
);

INVx4_ASAP7_75t_L g1315 ( 
.A(n_1101),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1214),
.A2(n_1221),
.B1(n_1200),
.B2(n_1177),
.Y(n_1316)
);

OAI21x1_ASAP7_75t_L g1317 ( 
.A1(n_1168),
.A2(n_1189),
.B(n_1226),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1214),
.Y(n_1318)
);

INVx1_ASAP7_75t_SL g1319 ( 
.A(n_1101),
.Y(n_1319)
);

NOR2xp33_ASAP7_75t_L g1320 ( 
.A(n_1098),
.B(n_1154),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1139),
.Y(n_1321)
);

OR2x2_ASAP7_75t_L g1322 ( 
.A(n_1213),
.B(n_1116),
.Y(n_1322)
);

NOR2xp33_ASAP7_75t_L g1323 ( 
.A(n_1226),
.B(n_1166),
.Y(n_1323)
);

OAI21x1_ASAP7_75t_L g1324 ( 
.A1(n_1163),
.A2(n_1144),
.B(n_1116),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1148),
.Y(n_1325)
);

O2A1O1Ixp33_ASAP7_75t_L g1326 ( 
.A1(n_1144),
.A2(n_1235),
.B(n_1231),
.C(n_1161),
.Y(n_1326)
);

HB1xp67_ASAP7_75t_L g1327 ( 
.A(n_1186),
.Y(n_1327)
);

BUFx3_ASAP7_75t_L g1328 ( 
.A(n_1120),
.Y(n_1328)
);

AND2x2_ASAP7_75t_L g1329 ( 
.A(n_1114),
.B(n_713),
.Y(n_1329)
);

OAI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1231),
.A2(n_1235),
.B(n_895),
.Y(n_1330)
);

BUFx2_ASAP7_75t_SL g1331 ( 
.A(n_1233),
.Y(n_1331)
);

OAI21x1_ASAP7_75t_L g1332 ( 
.A1(n_1107),
.A2(n_1182),
.B(n_1176),
.Y(n_1332)
);

NOR2xp33_ASAP7_75t_L g1333 ( 
.A(n_1219),
.B(n_315),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1159),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_1110),
.Y(n_1335)
);

OAI21x1_ASAP7_75t_SL g1336 ( 
.A1(n_1130),
.A2(n_1023),
.B(n_1124),
.Y(n_1336)
);

AO31x2_ASAP7_75t_L g1337 ( 
.A1(n_1119),
.A2(n_1035),
.A3(n_1227),
.B(n_1231),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1159),
.Y(n_1338)
);

HB1xp67_ASAP7_75t_L g1339 ( 
.A(n_1186),
.Y(n_1339)
);

AOI22xp33_ASAP7_75t_L g1340 ( 
.A1(n_1227),
.A2(n_979),
.B1(n_1124),
.B2(n_1179),
.Y(n_1340)
);

AND2x4_ASAP7_75t_L g1341 ( 
.A(n_1111),
.B(n_1155),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1114),
.B(n_713),
.Y(n_1342)
);

INVx2_ASAP7_75t_SL g1343 ( 
.A(n_1157),
.Y(n_1343)
);

OAI21x1_ASAP7_75t_L g1344 ( 
.A1(n_1107),
.A2(n_1182),
.B(n_1176),
.Y(n_1344)
);

CKINVDCx11_ASAP7_75t_R g1345 ( 
.A(n_1136),
.Y(n_1345)
);

BUFx3_ASAP7_75t_L g1346 ( 
.A(n_1120),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1110),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1159),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1114),
.B(n_713),
.Y(n_1349)
);

AO21x2_ASAP7_75t_L g1350 ( 
.A1(n_1119),
.A2(n_1140),
.B(n_1137),
.Y(n_1350)
);

OR2x6_ASAP7_75t_L g1351 ( 
.A(n_1158),
.B(n_1236),
.Y(n_1351)
);

BUFx3_ASAP7_75t_L g1352 ( 
.A(n_1120),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1110),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1114),
.B(n_713),
.Y(n_1354)
);

OA21x2_ASAP7_75t_L g1355 ( 
.A1(n_1196),
.A2(n_1119),
.B(n_1137),
.Y(n_1355)
);

AOI22xp33_ASAP7_75t_L g1356 ( 
.A1(n_1227),
.A2(n_979),
.B1(n_1124),
.B2(n_1179),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1132),
.B(n_1121),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_SL g1358 ( 
.A(n_1227),
.B(n_895),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_1114),
.B(n_713),
.Y(n_1359)
);

INVx3_ASAP7_75t_L g1360 ( 
.A(n_1111),
.Y(n_1360)
);

OAI21x1_ASAP7_75t_L g1361 ( 
.A1(n_1107),
.A2(n_1182),
.B(n_1176),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_1110),
.Y(n_1362)
);

OAI21xp5_ASAP7_75t_L g1363 ( 
.A1(n_1231),
.A2(n_1235),
.B(n_895),
.Y(n_1363)
);

OAI21xp5_ASAP7_75t_L g1364 ( 
.A1(n_1231),
.A2(n_1235),
.B(n_895),
.Y(n_1364)
);

AND2x4_ASAP7_75t_L g1365 ( 
.A(n_1111),
.B(n_1155),
.Y(n_1365)
);

OAI21x1_ASAP7_75t_L g1366 ( 
.A1(n_1107),
.A2(n_1182),
.B(n_1176),
.Y(n_1366)
);

OAI22xp33_ASAP7_75t_L g1367 ( 
.A1(n_1227),
.A2(n_643),
.B1(n_1185),
.B2(n_1179),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1269),
.B(n_1298),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1260),
.B(n_1269),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1298),
.B(n_1248),
.Y(n_1370)
);

AOI21x1_ASAP7_75t_SL g1371 ( 
.A1(n_1305),
.A2(n_1312),
.B(n_1281),
.Y(n_1371)
);

OA21x2_ASAP7_75t_L g1372 ( 
.A1(n_1283),
.A2(n_1270),
.B(n_1286),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1254),
.B(n_1341),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1357),
.B(n_1318),
.Y(n_1374)
);

CKINVDCx20_ASAP7_75t_R g1375 ( 
.A(n_1345),
.Y(n_1375)
);

NOR2xp33_ASAP7_75t_L g1376 ( 
.A(n_1241),
.B(n_1367),
.Y(n_1376)
);

AOI211xp5_ASAP7_75t_L g1377 ( 
.A1(n_1367),
.A2(n_1241),
.B(n_1242),
.C(n_1265),
.Y(n_1377)
);

BUFx8_ASAP7_75t_SL g1378 ( 
.A(n_1263),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1258),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1278),
.Y(n_1380)
);

AOI21xp5_ASAP7_75t_SL g1381 ( 
.A1(n_1245),
.A2(n_1351),
.B(n_1363),
.Y(n_1381)
);

AND2x4_ASAP7_75t_L g1382 ( 
.A(n_1281),
.B(n_1305),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1365),
.B(n_1329),
.Y(n_1383)
);

AOI21xp5_ASAP7_75t_L g1384 ( 
.A1(n_1245),
.A2(n_1351),
.B(n_1330),
.Y(n_1384)
);

O2A1O1Ixp33_ASAP7_75t_L g1385 ( 
.A1(n_1336),
.A2(n_1358),
.B(n_1364),
.C(n_1326),
.Y(n_1385)
);

AOI221x1_ASAP7_75t_SL g1386 ( 
.A1(n_1272),
.A2(n_1333),
.B1(n_1240),
.B2(n_1338),
.C(n_1334),
.Y(n_1386)
);

AOI21xp5_ASAP7_75t_SL g1387 ( 
.A1(n_1245),
.A2(n_1351),
.B(n_1323),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1301),
.B(n_1244),
.Y(n_1388)
);

A2O1A1Ixp33_ASAP7_75t_L g1389 ( 
.A1(n_1261),
.A2(n_1356),
.B(n_1340),
.C(n_1284),
.Y(n_1389)
);

AOI221x1_ASAP7_75t_SL g1390 ( 
.A1(n_1333),
.A2(n_1348),
.B1(n_1247),
.B2(n_1285),
.C(n_1287),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1295),
.B(n_1261),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1293),
.B(n_1296),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1340),
.B(n_1356),
.Y(n_1393)
);

OR2x2_ASAP7_75t_L g1394 ( 
.A(n_1358),
.B(n_1303),
.Y(n_1394)
);

OR2x2_ASAP7_75t_L g1395 ( 
.A(n_1273),
.B(n_1327),
.Y(n_1395)
);

AND2x4_ASAP7_75t_L g1396 ( 
.A(n_1291),
.B(n_1262),
.Y(n_1396)
);

OAI22xp5_ASAP7_75t_L g1397 ( 
.A1(n_1313),
.A2(n_1292),
.B1(n_1307),
.B2(n_1243),
.Y(n_1397)
);

OA21x2_ASAP7_75t_L g1398 ( 
.A1(n_1290),
.A2(n_1280),
.B(n_1297),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1339),
.B(n_1246),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1365),
.B(n_1342),
.Y(n_1400)
);

AOI21xp5_ASAP7_75t_L g1401 ( 
.A1(n_1350),
.A2(n_1264),
.B(n_1293),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1349),
.B(n_1354),
.Y(n_1402)
);

A2O1A1Ixp33_ASAP7_75t_L g1403 ( 
.A1(n_1307),
.A2(n_1324),
.B(n_1316),
.C(n_1323),
.Y(n_1403)
);

O2A1O1Ixp5_ASAP7_75t_L g1404 ( 
.A1(n_1310),
.A2(n_1325),
.B(n_1321),
.C(n_1320),
.Y(n_1404)
);

OR2x2_ASAP7_75t_L g1405 ( 
.A(n_1253),
.B(n_1335),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1359),
.B(n_1304),
.Y(n_1406)
);

A2O1A1Ixp33_ASAP7_75t_L g1407 ( 
.A1(n_1324),
.A2(n_1316),
.B(n_1290),
.C(n_1297),
.Y(n_1407)
);

AOI21xp5_ASAP7_75t_L g1408 ( 
.A1(n_1350),
.A2(n_1264),
.B(n_1279),
.Y(n_1408)
);

AOI21xp5_ASAP7_75t_SL g1409 ( 
.A1(n_1315),
.A2(n_1264),
.B(n_1308),
.Y(n_1409)
);

NOR2xp67_ASAP7_75t_L g1410 ( 
.A(n_1252),
.B(n_1255),
.Y(n_1410)
);

OAI22xp5_ASAP7_75t_L g1411 ( 
.A1(n_1313),
.A2(n_1299),
.B1(n_1352),
.B2(n_1346),
.Y(n_1411)
);

OR2x2_ASAP7_75t_L g1412 ( 
.A(n_1347),
.B(n_1353),
.Y(n_1412)
);

O2A1O1Ixp5_ASAP7_75t_L g1413 ( 
.A1(n_1320),
.A2(n_1322),
.B(n_1314),
.C(n_1271),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1347),
.B(n_1362),
.Y(n_1414)
);

AOI21xp5_ASAP7_75t_SL g1415 ( 
.A1(n_1315),
.A2(n_1308),
.B(n_1279),
.Y(n_1415)
);

AND2x4_ASAP7_75t_L g1416 ( 
.A(n_1308),
.B(n_1271),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1328),
.B(n_1352),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1296),
.Y(n_1418)
);

AOI21xp5_ASAP7_75t_SL g1419 ( 
.A1(n_1315),
.A2(n_1279),
.B(n_1355),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1300),
.Y(n_1420)
);

OAI22xp5_ASAP7_75t_L g1421 ( 
.A1(n_1289),
.A2(n_1331),
.B1(n_1360),
.B2(n_1250),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1271),
.B(n_1306),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1249),
.B(n_1256),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1306),
.B(n_1266),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1249),
.B(n_1256),
.Y(n_1425)
);

AOI21xp5_ASAP7_75t_L g1426 ( 
.A1(n_1251),
.A2(n_1355),
.B(n_1259),
.Y(n_1426)
);

AOI21x1_ASAP7_75t_SL g1427 ( 
.A1(n_1309),
.A2(n_1288),
.B(n_1276),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1274),
.B(n_1337),
.Y(n_1428)
);

OAI211xp5_ASAP7_75t_L g1429 ( 
.A1(n_1251),
.A2(n_1355),
.B(n_1345),
.C(n_1267),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1314),
.B(n_1337),
.Y(n_1430)
);

HB1xp67_ASAP7_75t_L g1431 ( 
.A(n_1251),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1337),
.B(n_1289),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1275),
.B(n_1319),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1275),
.B(n_1343),
.Y(n_1434)
);

BUFx12f_ASAP7_75t_L g1435 ( 
.A(n_1277),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1275),
.B(n_1311),
.Y(n_1436)
);

O2A1O1Ixp5_ASAP7_75t_L g1437 ( 
.A1(n_1302),
.A2(n_1282),
.B(n_1317),
.C(n_1280),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_1239),
.Y(n_1438)
);

AND2x4_ASAP7_75t_L g1439 ( 
.A(n_1239),
.B(n_1366),
.Y(n_1439)
);

HB1xp67_ASAP7_75t_L g1440 ( 
.A(n_1332),
.Y(n_1440)
);

OR2x2_ASAP7_75t_L g1441 ( 
.A(n_1332),
.B(n_1366),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1344),
.B(n_1361),
.Y(n_1442)
);

O2A1O1Ixp5_ASAP7_75t_L g1443 ( 
.A1(n_1344),
.A2(n_1361),
.B(n_1268),
.C(n_1263),
.Y(n_1443)
);

AOI21xp5_ASAP7_75t_SL g1444 ( 
.A1(n_1277),
.A2(n_1227),
.B(n_1231),
.Y(n_1444)
);

OR2x2_ASAP7_75t_L g1445 ( 
.A(n_1301),
.B(n_1294),
.Y(n_1445)
);

OR2x2_ASAP7_75t_L g1446 ( 
.A(n_1301),
.B(n_1294),
.Y(n_1446)
);

AOI21x1_ASAP7_75t_SL g1447 ( 
.A1(n_1305),
.A2(n_1312),
.B(n_1281),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1257),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1260),
.B(n_1269),
.Y(n_1449)
);

OAI22xp5_ASAP7_75t_L g1450 ( 
.A1(n_1340),
.A2(n_1356),
.B1(n_1124),
.B2(n_1261),
.Y(n_1450)
);

NAND2xp33_ASAP7_75t_SL g1451 ( 
.A(n_1315),
.B(n_1227),
.Y(n_1451)
);

BUFx6f_ASAP7_75t_L g1452 ( 
.A(n_1315),
.Y(n_1452)
);

O2A1O1Ixp5_ASAP7_75t_L g1453 ( 
.A1(n_1358),
.A2(n_1227),
.B(n_1363),
.C(n_1330),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1368),
.B(n_1370),
.Y(n_1454)
);

AO21x2_ASAP7_75t_L g1455 ( 
.A1(n_1426),
.A2(n_1408),
.B(n_1401),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_1438),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1392),
.B(n_1418),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1420),
.Y(n_1458)
);

AO21x2_ASAP7_75t_L g1459 ( 
.A1(n_1407),
.A2(n_1419),
.B(n_1429),
.Y(n_1459)
);

OR2x2_ASAP7_75t_L g1460 ( 
.A(n_1392),
.B(n_1428),
.Y(n_1460)
);

INVx3_ASAP7_75t_L g1461 ( 
.A(n_1439),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1430),
.B(n_1372),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1374),
.B(n_1376),
.Y(n_1463)
);

OA21x2_ASAP7_75t_L g1464 ( 
.A1(n_1437),
.A2(n_1431),
.B(n_1403),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1372),
.B(n_1431),
.Y(n_1465)
);

HB1xp67_ASAP7_75t_L g1466 ( 
.A(n_1436),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1376),
.B(n_1432),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_SL g1468 ( 
.A(n_1385),
.B(n_1377),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1372),
.B(n_1382),
.Y(n_1469)
);

INVx2_ASAP7_75t_SL g1470 ( 
.A(n_1439),
.Y(n_1470)
);

BUFx2_ASAP7_75t_L g1471 ( 
.A(n_1440),
.Y(n_1471)
);

AO21x2_ASAP7_75t_L g1472 ( 
.A1(n_1403),
.A2(n_1423),
.B(n_1425),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1379),
.Y(n_1473)
);

AO21x2_ASAP7_75t_L g1474 ( 
.A1(n_1384),
.A2(n_1415),
.B(n_1409),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1441),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1442),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1380),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1394),
.B(n_1448),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1442),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1398),
.Y(n_1480)
);

AO21x2_ASAP7_75t_L g1481 ( 
.A1(n_1389),
.A2(n_1381),
.B(n_1450),
.Y(n_1481)
);

AO21x2_ASAP7_75t_L g1482 ( 
.A1(n_1389),
.A2(n_1381),
.B(n_1410),
.Y(n_1482)
);

NOR3xp33_ASAP7_75t_L g1483 ( 
.A(n_1453),
.B(n_1393),
.C(n_1397),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1398),
.Y(n_1484)
);

OAI21xp5_ASAP7_75t_L g1485 ( 
.A1(n_1444),
.A2(n_1404),
.B(n_1413),
.Y(n_1485)
);

INVx2_ASAP7_75t_SL g1486 ( 
.A(n_1416),
.Y(n_1486)
);

AOI22xp33_ASAP7_75t_L g1487 ( 
.A1(n_1451),
.A2(n_1391),
.B1(n_1449),
.B2(n_1369),
.Y(n_1487)
);

NAND2x1p5_ASAP7_75t_L g1488 ( 
.A(n_1416),
.B(n_1396),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1443),
.Y(n_1489)
);

AOI21x1_ASAP7_75t_L g1490 ( 
.A1(n_1421),
.A2(n_1414),
.B(n_1416),
.Y(n_1490)
);

AO21x2_ASAP7_75t_L g1491 ( 
.A1(n_1387),
.A2(n_1444),
.B(n_1399),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1405),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1422),
.B(n_1412),
.Y(n_1493)
);

OR2x2_ASAP7_75t_L g1494 ( 
.A(n_1395),
.B(n_1445),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1424),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1451),
.Y(n_1496)
);

INVx3_ASAP7_75t_L g1497 ( 
.A(n_1452),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1390),
.Y(n_1498)
);

OAI21xp5_ASAP7_75t_L g1499 ( 
.A1(n_1485),
.A2(n_1388),
.B(n_1411),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1476),
.B(n_1406),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1458),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1456),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1458),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1462),
.B(n_1465),
.Y(n_1504)
);

INVx1_ASAP7_75t_SL g1505 ( 
.A(n_1471),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1458),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1479),
.B(n_1373),
.Y(n_1507)
);

NOR2x1p5_ASAP7_75t_L g1508 ( 
.A(n_1498),
.B(n_1452),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1462),
.B(n_1465),
.Y(n_1509)
);

INVx3_ASAP7_75t_L g1510 ( 
.A(n_1461),
.Y(n_1510)
);

AO21x2_ASAP7_75t_L g1511 ( 
.A1(n_1455),
.A2(n_1434),
.B(n_1417),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1492),
.B(n_1386),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1462),
.B(n_1402),
.Y(n_1513)
);

AOI22xp33_ASAP7_75t_SL g1514 ( 
.A1(n_1481),
.A2(n_1375),
.B1(n_1383),
.B2(n_1400),
.Y(n_1514)
);

BUFx2_ASAP7_75t_L g1515 ( 
.A(n_1461),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1469),
.B(n_1446),
.Y(n_1516)
);

AOI22xp33_ASAP7_75t_L g1517 ( 
.A1(n_1468),
.A2(n_1375),
.B1(n_1378),
.B2(n_1435),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1469),
.B(n_1433),
.Y(n_1518)
);

AND2x4_ASAP7_75t_L g1519 ( 
.A(n_1461),
.B(n_1452),
.Y(n_1519)
);

OA21x2_ASAP7_75t_L g1520 ( 
.A1(n_1489),
.A2(n_1371),
.B(n_1447),
.Y(n_1520)
);

OR2x2_ASAP7_75t_L g1521 ( 
.A(n_1460),
.B(n_1452),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1469),
.B(n_1461),
.Y(n_1522)
);

AOI22xp33_ASAP7_75t_L g1523 ( 
.A1(n_1514),
.A2(n_1481),
.B1(n_1468),
.B2(n_1483),
.Y(n_1523)
);

AOI22xp33_ASAP7_75t_L g1524 ( 
.A1(n_1514),
.A2(n_1481),
.B1(n_1483),
.B2(n_1482),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1502),
.Y(n_1525)
);

AOI221xp5_ASAP7_75t_L g1526 ( 
.A1(n_1512),
.A2(n_1498),
.B1(n_1467),
.B2(n_1485),
.C(n_1463),
.Y(n_1526)
);

AND2x4_ASAP7_75t_L g1527 ( 
.A(n_1519),
.B(n_1470),
.Y(n_1527)
);

AOI22xp33_ASAP7_75t_L g1528 ( 
.A1(n_1499),
.A2(n_1481),
.B1(n_1482),
.B2(n_1498),
.Y(n_1528)
);

OAI211xp5_ASAP7_75t_SL g1529 ( 
.A1(n_1512),
.A2(n_1463),
.B(n_1454),
.C(n_1467),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1501),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1501),
.Y(n_1531)
);

AOI22xp5_ASAP7_75t_L g1532 ( 
.A1(n_1499),
.A2(n_1481),
.B1(n_1482),
.B2(n_1491),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1502),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1516),
.B(n_1494),
.Y(n_1534)
);

BUFx3_ASAP7_75t_L g1535 ( 
.A(n_1521),
.Y(n_1535)
);

OAI221xp5_ASAP7_75t_L g1536 ( 
.A1(n_1499),
.A2(n_1487),
.B1(n_1454),
.B2(n_1494),
.C(n_1478),
.Y(n_1536)
);

AOI22xp33_ASAP7_75t_L g1537 ( 
.A1(n_1508),
.A2(n_1482),
.B1(n_1491),
.B2(n_1487),
.Y(n_1537)
);

AOI221xp5_ASAP7_75t_L g1538 ( 
.A1(n_1516),
.A2(n_1457),
.B1(n_1478),
.B2(n_1492),
.C(n_1472),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1501),
.Y(n_1539)
);

AND2x4_ASAP7_75t_L g1540 ( 
.A(n_1519),
.B(n_1470),
.Y(n_1540)
);

OAI221xp5_ASAP7_75t_L g1541 ( 
.A1(n_1517),
.A2(n_1494),
.B1(n_1486),
.B2(n_1460),
.C(n_1488),
.Y(n_1541)
);

INVx3_ASAP7_75t_L g1542 ( 
.A(n_1510),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1513),
.B(n_1466),
.Y(n_1543)
);

BUFx3_ASAP7_75t_L g1544 ( 
.A(n_1521),
.Y(n_1544)
);

AOI221xp5_ASAP7_75t_L g1545 ( 
.A1(n_1516),
.A2(n_1457),
.B1(n_1492),
.B2(n_1472),
.C(n_1496),
.Y(n_1545)
);

NAND2xp33_ASAP7_75t_SL g1546 ( 
.A(n_1508),
.B(n_1482),
.Y(n_1546)
);

AND2x4_ASAP7_75t_L g1547 ( 
.A(n_1519),
.B(n_1470),
.Y(n_1547)
);

OAI22xp5_ASAP7_75t_L g1548 ( 
.A1(n_1517),
.A2(n_1496),
.B1(n_1486),
.B2(n_1488),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1503),
.Y(n_1549)
);

NOR2xp33_ASAP7_75t_L g1550 ( 
.A(n_1516),
.B(n_1495),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1513),
.B(n_1466),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1513),
.B(n_1457),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1503),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1513),
.B(n_1500),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1503),
.Y(n_1555)
);

AOI22xp5_ASAP7_75t_L g1556 ( 
.A1(n_1519),
.A2(n_1491),
.B1(n_1474),
.B2(n_1486),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1506),
.Y(n_1557)
);

NAND3xp33_ASAP7_75t_L g1558 ( 
.A(n_1520),
.B(n_1489),
.C(n_1496),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1500),
.B(n_1493),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1522),
.B(n_1470),
.Y(n_1560)
);

NAND2xp33_ASAP7_75t_R g1561 ( 
.A(n_1520),
.B(n_1464),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1506),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1500),
.B(n_1493),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1500),
.B(n_1493),
.Y(n_1564)
);

NOR2x1_ASAP7_75t_SL g1565 ( 
.A(n_1511),
.B(n_1474),
.Y(n_1565)
);

AOI33xp33_ASAP7_75t_L g1566 ( 
.A1(n_1505),
.A2(n_1465),
.A3(n_1489),
.B1(n_1475),
.B2(n_1477),
.B3(n_1473),
.Y(n_1566)
);

OR2x2_ASAP7_75t_L g1567 ( 
.A(n_1554),
.B(n_1504),
.Y(n_1567)
);

INVx3_ASAP7_75t_L g1568 ( 
.A(n_1542),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1525),
.Y(n_1569)
);

AOI21xp5_ASAP7_75t_L g1570 ( 
.A1(n_1532),
.A2(n_1474),
.B(n_1524),
.Y(n_1570)
);

INVx2_ASAP7_75t_SL g1571 ( 
.A(n_1542),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1530),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1531),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1560),
.B(n_1522),
.Y(n_1574)
);

INVxp67_ASAP7_75t_SL g1575 ( 
.A(n_1558),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1539),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1552),
.B(n_1522),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1552),
.B(n_1504),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1538),
.B(n_1504),
.Y(n_1579)
);

NAND3xp33_ASAP7_75t_SL g1580 ( 
.A(n_1526),
.B(n_1505),
.C(n_1521),
.Y(n_1580)
);

OA21x2_ASAP7_75t_L g1581 ( 
.A1(n_1556),
.A2(n_1484),
.B(n_1480),
.Y(n_1581)
);

HB1xp67_ASAP7_75t_L g1582 ( 
.A(n_1549),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_SL g1583 ( 
.A(n_1523),
.B(n_1486),
.Y(n_1583)
);

INVx2_ASAP7_75t_L g1584 ( 
.A(n_1525),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_1533),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1533),
.Y(n_1586)
);

INVxp67_ASAP7_75t_L g1587 ( 
.A(n_1536),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1553),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1543),
.B(n_1509),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1566),
.B(n_1509),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1555),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1557),
.Y(n_1592)
);

OR2x2_ASAP7_75t_L g1593 ( 
.A(n_1534),
.B(n_1509),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1562),
.Y(n_1594)
);

BUFx2_ASAP7_75t_L g1595 ( 
.A(n_1546),
.Y(n_1595)
);

AND2x4_ASAP7_75t_L g1596 ( 
.A(n_1527),
.B(n_1515),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1543),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1535),
.Y(n_1598)
);

AOI21xp33_ASAP7_75t_L g1599 ( 
.A1(n_1529),
.A2(n_1528),
.B(n_1561),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1551),
.Y(n_1600)
);

INVx4_ASAP7_75t_L g1601 ( 
.A(n_1598),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1578),
.B(n_1551),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1587),
.B(n_1545),
.Y(n_1603)
);

OR2x2_ASAP7_75t_L g1604 ( 
.A(n_1590),
.B(n_1559),
.Y(n_1604)
);

NAND3xp33_ASAP7_75t_L g1605 ( 
.A(n_1570),
.B(n_1561),
.C(n_1537),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1578),
.B(n_1535),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1587),
.B(n_1544),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1590),
.B(n_1544),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1578),
.B(n_1527),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1577),
.B(n_1527),
.Y(n_1610)
);

NOR2x1_ASAP7_75t_L g1611 ( 
.A(n_1580),
.B(n_1541),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1582),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1582),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1577),
.B(n_1540),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1579),
.B(n_1566),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1572),
.Y(n_1616)
);

OR2x2_ASAP7_75t_L g1617 ( 
.A(n_1593),
.B(n_1563),
.Y(n_1617)
);

OR2x2_ASAP7_75t_L g1618 ( 
.A(n_1593),
.B(n_1564),
.Y(n_1618)
);

AND2x4_ASAP7_75t_L g1619 ( 
.A(n_1598),
.B(n_1540),
.Y(n_1619)
);

NAND2x1_ASAP7_75t_L g1620 ( 
.A(n_1595),
.B(n_1540),
.Y(n_1620)
);

AND2x4_ASAP7_75t_L g1621 ( 
.A(n_1598),
.B(n_1547),
.Y(n_1621)
);

INVxp67_ASAP7_75t_L g1622 ( 
.A(n_1583),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1577),
.B(n_1547),
.Y(n_1623)
);

NAND3xp33_ASAP7_75t_L g1624 ( 
.A(n_1570),
.B(n_1548),
.C(n_1546),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1572),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1569),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1569),
.Y(n_1627)
);

OR2x2_ASAP7_75t_L g1628 ( 
.A(n_1593),
.B(n_1460),
.Y(n_1628)
);

INVx1_ASAP7_75t_SL g1629 ( 
.A(n_1595),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1589),
.B(n_1547),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1573),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1589),
.B(n_1518),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1589),
.B(n_1574),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1569),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1574),
.B(n_1518),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1579),
.B(n_1550),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1574),
.B(n_1518),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1573),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1576),
.Y(n_1639)
);

NOR3xp33_ASAP7_75t_L g1640 ( 
.A(n_1580),
.B(n_1490),
.C(n_1497),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1576),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1599),
.B(n_1507),
.Y(n_1642)
);

OR2x2_ASAP7_75t_L g1643 ( 
.A(n_1607),
.B(n_1583),
.Y(n_1643)
);

AND2x4_ASAP7_75t_L g1644 ( 
.A(n_1601),
.B(n_1575),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1603),
.B(n_1622),
.Y(n_1645)
);

NAND4xp25_ASAP7_75t_L g1646 ( 
.A(n_1611),
.B(n_1599),
.C(n_1595),
.D(n_1521),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1601),
.Y(n_1647)
);

OR2x2_ASAP7_75t_L g1648 ( 
.A(n_1608),
.B(n_1567),
.Y(n_1648)
);

OR2x2_ASAP7_75t_L g1649 ( 
.A(n_1604),
.B(n_1567),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1616),
.Y(n_1650)
);

INVx2_ASAP7_75t_SL g1651 ( 
.A(n_1620),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1619),
.B(n_1596),
.Y(n_1652)
);

OR2x2_ASAP7_75t_L g1653 ( 
.A(n_1604),
.B(n_1575),
.Y(n_1653)
);

NOR2xp33_ASAP7_75t_L g1654 ( 
.A(n_1636),
.B(n_1378),
.Y(n_1654)
);

AOI22xp33_ASAP7_75t_L g1655 ( 
.A1(n_1605),
.A2(n_1491),
.B1(n_1474),
.B2(n_1459),
.Y(n_1655)
);

NOR2xp33_ASAP7_75t_L g1656 ( 
.A(n_1615),
.B(n_1435),
.Y(n_1656)
);

INVxp67_ASAP7_75t_L g1657 ( 
.A(n_1642),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1619),
.B(n_1596),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1619),
.B(n_1596),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1616),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1625),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1640),
.B(n_1606),
.Y(n_1662)
);

HB1xp67_ASAP7_75t_L g1663 ( 
.A(n_1612),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1625),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1631),
.Y(n_1665)
);

AND2x4_ASAP7_75t_L g1666 ( 
.A(n_1601),
.B(n_1596),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1621),
.B(n_1596),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1633),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1631),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1638),
.Y(n_1670)
);

NAND2xp67_ASAP7_75t_L g1671 ( 
.A(n_1606),
.B(n_1584),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1602),
.B(n_1597),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1638),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_1633),
.Y(n_1674)
);

AOI22xp33_ASAP7_75t_SL g1675 ( 
.A1(n_1624),
.A2(n_1565),
.B1(n_1459),
.B2(n_1581),
.Y(n_1675)
);

NOR2xp67_ASAP7_75t_L g1676 ( 
.A(n_1612),
.B(n_1597),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1602),
.B(n_1600),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1663),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_1651),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1645),
.B(n_1629),
.Y(n_1680)
);

INVx1_ASAP7_75t_SL g1681 ( 
.A(n_1643),
.Y(n_1681)
);

CKINVDCx16_ASAP7_75t_R g1682 ( 
.A(n_1654),
.Y(n_1682)
);

HB1xp67_ASAP7_75t_L g1683 ( 
.A(n_1644),
.Y(n_1683)
);

OR2x6_ASAP7_75t_L g1684 ( 
.A(n_1647),
.B(n_1620),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1650),
.Y(n_1685)
);

OR2x2_ASAP7_75t_L g1686 ( 
.A(n_1648),
.B(n_1617),
.Y(n_1686)
);

OAI22xp5_ASAP7_75t_L g1687 ( 
.A1(n_1655),
.A2(n_1628),
.B1(n_1618),
.B2(n_1617),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1654),
.B(n_1632),
.Y(n_1688)
);

OR2x2_ASAP7_75t_L g1689 ( 
.A(n_1657),
.B(n_1618),
.Y(n_1689)
);

INVx1_ASAP7_75t_SL g1690 ( 
.A(n_1653),
.Y(n_1690)
);

OR2x2_ASAP7_75t_L g1691 ( 
.A(n_1653),
.B(n_1628),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1652),
.B(n_1621),
.Y(n_1692)
);

HB1xp67_ASAP7_75t_L g1693 ( 
.A(n_1644),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1652),
.B(n_1658),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1660),
.Y(n_1695)
);

INVxp67_ASAP7_75t_SL g1696 ( 
.A(n_1651),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1661),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1664),
.Y(n_1698)
);

NOR2xp33_ASAP7_75t_L g1699 ( 
.A(n_1656),
.B(n_1621),
.Y(n_1699)
);

OR2x2_ASAP7_75t_L g1700 ( 
.A(n_1646),
.B(n_1662),
.Y(n_1700)
);

OAI22xp5_ASAP7_75t_L g1701 ( 
.A1(n_1655),
.A2(n_1567),
.B1(n_1600),
.B2(n_1632),
.Y(n_1701)
);

INVx1_ASAP7_75t_SL g1702 ( 
.A(n_1666),
.Y(n_1702)
);

OAI22xp5_ASAP7_75t_L g1703 ( 
.A1(n_1700),
.A2(n_1675),
.B1(n_1656),
.B2(n_1674),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1690),
.B(n_1644),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1694),
.B(n_1658),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1683),
.Y(n_1706)
);

OAI21xp33_ASAP7_75t_L g1707 ( 
.A1(n_1688),
.A2(n_1671),
.B(n_1674),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1683),
.B(n_1647),
.Y(n_1708)
);

NOR2xp33_ASAP7_75t_L g1709 ( 
.A(n_1682),
.B(n_1649),
.Y(n_1709)
);

OAI21xp5_ASAP7_75t_L g1710 ( 
.A1(n_1681),
.A2(n_1676),
.B(n_1665),
.Y(n_1710)
);

NAND3xp33_ASAP7_75t_SL g1711 ( 
.A(n_1702),
.B(n_1668),
.C(n_1673),
.Y(n_1711)
);

OAI21xp5_ASAP7_75t_SL g1712 ( 
.A1(n_1699),
.A2(n_1668),
.B(n_1666),
.Y(n_1712)
);

AOI21xp5_ASAP7_75t_L g1713 ( 
.A1(n_1680),
.A2(n_1666),
.B(n_1670),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1693),
.B(n_1669),
.Y(n_1714)
);

NAND3xp33_ASAP7_75t_L g1715 ( 
.A(n_1693),
.B(n_1613),
.C(n_1672),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1678),
.B(n_1659),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1696),
.B(n_1694),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1692),
.B(n_1699),
.Y(n_1718)
);

NAND2x1_ASAP7_75t_L g1719 ( 
.A(n_1684),
.B(n_1659),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1679),
.B(n_1667),
.Y(n_1720)
);

AOI21xp33_ASAP7_75t_SL g1721 ( 
.A1(n_1687),
.A2(n_1613),
.B(n_1667),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1685),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1709),
.B(n_1679),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1706),
.Y(n_1724)
);

INVx1_ASAP7_75t_SL g1725 ( 
.A(n_1717),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1718),
.B(n_1692),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1704),
.B(n_1695),
.Y(n_1727)
);

NOR2xp33_ASAP7_75t_L g1728 ( 
.A(n_1716),
.B(n_1689),
.Y(n_1728)
);

AOI22xp33_ASAP7_75t_SL g1729 ( 
.A1(n_1703),
.A2(n_1701),
.B1(n_1565),
.B2(n_1686),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1714),
.Y(n_1730)
);

AOI22xp33_ASAP7_75t_L g1731 ( 
.A1(n_1705),
.A2(n_1691),
.B1(n_1684),
.B2(n_1697),
.Y(n_1731)
);

NAND2x1_ASAP7_75t_L g1732 ( 
.A(n_1710),
.B(n_1684),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1713),
.B(n_1698),
.Y(n_1733)
);

AOI221xp5_ASAP7_75t_L g1734 ( 
.A1(n_1733),
.A2(n_1721),
.B1(n_1711),
.B2(n_1715),
.C(n_1710),
.Y(n_1734)
);

OAI211xp5_ASAP7_75t_L g1735 ( 
.A1(n_1732),
.A2(n_1719),
.B(n_1712),
.C(n_1708),
.Y(n_1735)
);

NAND3xp33_ASAP7_75t_L g1736 ( 
.A(n_1729),
.B(n_1722),
.C(n_1720),
.Y(n_1736)
);

NOR2xp33_ASAP7_75t_L g1737 ( 
.A(n_1723),
.B(n_1707),
.Y(n_1737)
);

AOI22xp33_ASAP7_75t_SL g1738 ( 
.A1(n_1725),
.A2(n_1728),
.B1(n_1726),
.B2(n_1730),
.Y(n_1738)
);

NOR3xp33_ASAP7_75t_L g1739 ( 
.A(n_1727),
.B(n_1677),
.C(n_1634),
.Y(n_1739)
);

O2A1O1Ixp5_ASAP7_75t_L g1740 ( 
.A1(n_1724),
.A2(n_1626),
.B(n_1627),
.C(n_1634),
.Y(n_1740)
);

AOI221xp5_ASAP7_75t_L g1741 ( 
.A1(n_1731),
.A2(n_1641),
.B1(n_1639),
.B2(n_1626),
.C(n_1627),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1724),
.Y(n_1742)
);

OAI21xp33_ASAP7_75t_SL g1743 ( 
.A1(n_1734),
.A2(n_1684),
.B(n_1610),
.Y(n_1743)
);

INVxp67_ASAP7_75t_L g1744 ( 
.A(n_1737),
.Y(n_1744)
);

O2A1O1Ixp33_ASAP7_75t_L g1745 ( 
.A1(n_1735),
.A2(n_1641),
.B(n_1639),
.C(n_1571),
.Y(n_1745)
);

AOI22xp5_ASAP7_75t_L g1746 ( 
.A1(n_1736),
.A2(n_1614),
.B1(n_1623),
.B2(n_1610),
.Y(n_1746)
);

O2A1O1Ixp5_ASAP7_75t_L g1747 ( 
.A1(n_1742),
.A2(n_1568),
.B(n_1569),
.C(n_1584),
.Y(n_1747)
);

OAI21xp5_ASAP7_75t_L g1748 ( 
.A1(n_1743),
.A2(n_1738),
.B(n_1741),
.Y(n_1748)
);

INVx1_ASAP7_75t_SL g1749 ( 
.A(n_1746),
.Y(n_1749)
);

CKINVDCx5p33_ASAP7_75t_R g1750 ( 
.A(n_1744),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1745),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1747),
.B(n_1739),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1744),
.Y(n_1753)
);

NOR2x1_ASAP7_75t_L g1754 ( 
.A(n_1753),
.B(n_1751),
.Y(n_1754)
);

CKINVDCx5p33_ASAP7_75t_R g1755 ( 
.A(n_1750),
.Y(n_1755)
);

INVx3_ASAP7_75t_SL g1756 ( 
.A(n_1750),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1752),
.Y(n_1757)
);

AOI21xp5_ASAP7_75t_L g1758 ( 
.A1(n_1748),
.A2(n_1740),
.B(n_1571),
.Y(n_1758)
);

NOR3xp33_ASAP7_75t_L g1759 ( 
.A(n_1755),
.B(n_1749),
.C(n_1752),
.Y(n_1759)
);

NOR2x1_ASAP7_75t_L g1760 ( 
.A(n_1757),
.B(n_1568),
.Y(n_1760)
);

OAI211xp5_ASAP7_75t_SL g1761 ( 
.A1(n_1754),
.A2(n_1427),
.B(n_1568),
.C(n_1594),
.Y(n_1761)
);

NOR3xp33_ASAP7_75t_SL g1762 ( 
.A(n_1761),
.B(n_1758),
.C(n_1756),
.Y(n_1762)
);

INVx2_ASAP7_75t_L g1763 ( 
.A(n_1762),
.Y(n_1763)
);

XOR2xp5_ASAP7_75t_L g1764 ( 
.A(n_1763),
.B(n_1760),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1764),
.B(n_1759),
.Y(n_1765)
);

AO22x1_ASAP7_75t_L g1766 ( 
.A1(n_1765),
.A2(n_1568),
.B1(n_1571),
.B2(n_1614),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1766),
.Y(n_1767)
);

AOI21xp5_ASAP7_75t_L g1768 ( 
.A1(n_1767),
.A2(n_1609),
.B(n_1630),
.Y(n_1768)
);

OAI21x1_ASAP7_75t_L g1769 ( 
.A1(n_1768),
.A2(n_1623),
.B(n_1609),
.Y(n_1769)
);

AND3x1_ASAP7_75t_L g1770 ( 
.A(n_1768),
.B(n_1568),
.C(n_1630),
.Y(n_1770)
);

AOI22xp33_ASAP7_75t_L g1771 ( 
.A1(n_1769),
.A2(n_1585),
.B1(n_1586),
.B2(n_1584),
.Y(n_1771)
);

AOI22xp33_ASAP7_75t_SL g1772 ( 
.A1(n_1770),
.A2(n_1637),
.B1(n_1635),
.B2(n_1594),
.Y(n_1772)
);

OAI22xp5_ASAP7_75t_L g1773 ( 
.A1(n_1772),
.A2(n_1771),
.B1(n_1637),
.B2(n_1635),
.Y(n_1773)
);

AOI211xp5_ASAP7_75t_L g1774 ( 
.A1(n_1773),
.A2(n_1592),
.B(n_1591),
.C(n_1588),
.Y(n_1774)
);


endmodule