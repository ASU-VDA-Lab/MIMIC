module fake_jpeg_16072_n_177 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_177);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_177;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g50 ( 
.A(n_10),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

BUFx16f_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

BUFx4f_ASAP7_75t_L g54 ( 
.A(n_13),
.Y(n_54)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_42),
.Y(n_57)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_22),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_11),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_17),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_49),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_12),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_32),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_77),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_79),
.Y(n_86)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_82),
.Y(n_87)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_78),
.Y(n_84)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_84),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_77),
.A2(n_58),
.B1(n_55),
.B2(n_53),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_88),
.A2(n_50),
.B1(n_73),
.B2(n_66),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_63),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_89),
.B(n_99),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_76),
.A2(n_54),
.B1(n_55),
.B2(n_70),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_90),
.A2(n_97),
.B1(n_74),
.B2(n_67),
.Y(n_121)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_75),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_93),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_82),
.B(n_56),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_94),
.B(n_95),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_56),
.C(n_70),
.Y(n_95)
);

OA22x2_ASAP7_75t_L g97 ( 
.A1(n_79),
.A2(n_54),
.B1(n_69),
.B2(n_73),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_96),
.Y(n_100)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_100),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_103),
.B(n_106),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_88),
.B(n_51),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_104),
.B(n_0),
.Y(n_127)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_98),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_98),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_107),
.A2(n_110),
.B1(n_118),
.B2(n_119),
.Y(n_128)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_85),
.Y(n_108)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_108),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_83),
.A2(n_57),
.B1(n_61),
.B2(n_68),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_97),
.A2(n_92),
.B1(n_90),
.B2(n_87),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_111),
.A2(n_121),
.B1(n_0),
.B2(n_1),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_97),
.B(n_59),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_112),
.B(n_104),
.Y(n_130)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_91),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_114),
.Y(n_125)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_92),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_115),
.A2(n_117),
.B1(n_120),
.B2(n_101),
.Y(n_131)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_91),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_116),
.Y(n_132)
);

HB1xp67_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_84),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_84),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_124),
.A2(n_133),
.B1(n_134),
.B2(n_62),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_127),
.B(n_130),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_131),
.Y(n_137)
);

OAI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_111),
.A2(n_102),
.B1(n_117),
.B2(n_109),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_102),
.A2(n_23),
.B1(n_48),
.B2(n_47),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_125),
.Y(n_135)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_135),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_129),
.B(n_113),
.Y(n_138)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_138),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_129),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_139),
.B(n_140),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_134),
.B(n_64),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_127),
.A2(n_72),
.B(n_71),
.Y(n_141)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_141),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_142),
.A2(n_128),
.B1(n_124),
.B2(n_126),
.Y(n_145)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_122),
.Y(n_143)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_143),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_145),
.A2(n_150),
.B1(n_123),
.B2(n_60),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_137),
.A2(n_123),
.B1(n_132),
.B2(n_126),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_148),
.B(n_140),
.C(n_145),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_151),
.B(n_36),
.C(n_35),
.Y(n_160)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_144),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_152),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_150),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_153),
.A2(n_154),
.B1(n_155),
.B2(n_156),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_146),
.B(n_135),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_147),
.A2(n_142),
.B1(n_149),
.B2(n_136),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_153),
.A2(n_39),
.B1(n_38),
.B2(n_37),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_158),
.A2(n_160),
.B(n_151),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_159),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_161),
.B(n_162),
.C(n_157),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_160),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_163),
.A2(n_164),
.B1(n_30),
.B2(n_28),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_27),
.C(n_26),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_166),
.A2(n_24),
.B1(n_16),
.B2(n_15),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_167),
.A2(n_14),
.B1(n_2),
.B2(n_3),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_1),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_169),
.B(n_3),
.Y(n_170)
);

OAI321xp33_ASAP7_75t_L g171 ( 
.A1(n_170),
.A2(n_4),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C(n_8),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_171),
.A2(n_4),
.B(n_5),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_172),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_173),
.B(n_6),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_7),
.C(n_8),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_175),
.B(n_9),
.C(n_10),
.Y(n_176)
);

FAx1_ASAP7_75t_SL g177 ( 
.A(n_176),
.B(n_9),
.CI(n_11),
.CON(n_177),
.SN(n_177)
);


endmodule