module fake_netlist_1_9459_n_43 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_14, n_7, n_15, n_10, n_8, n_0, n_43);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_14;
input n_7;
input n_15;
input n_10;
input n_8;
input n_0;
output n_43;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_17;
wire n_42;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_40;
wire n_27;
wire n_39;
INVx1_ASAP7_75t_L g16 ( .A(n_0), .Y(n_16) );
CKINVDCx20_ASAP7_75t_R g17 ( .A(n_9), .Y(n_17) );
OAI21x1_ASAP7_75t_L g18 ( .A1(n_7), .A2(n_14), .B(n_13), .Y(n_18) );
OA21x2_ASAP7_75t_L g19 ( .A1(n_4), .A2(n_1), .B(n_6), .Y(n_19) );
CKINVDCx5p33_ASAP7_75t_R g20 ( .A(n_10), .Y(n_20) );
CKINVDCx5p33_ASAP7_75t_R g21 ( .A(n_5), .Y(n_21) );
CKINVDCx5p33_ASAP7_75t_R g22 ( .A(n_12), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_0), .Y(n_23) );
NOR2xp33_ASAP7_75t_R g24 ( .A(n_21), .B(n_8), .Y(n_24) );
NOR3xp33_ASAP7_75t_SL g25 ( .A(n_16), .B(n_1), .C(n_2), .Y(n_25) );
INVx1_ASAP7_75t_L g26 ( .A(n_23), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_26), .Y(n_27) );
O2A1O1Ixp5_ASAP7_75t_L g28 ( .A1(n_26), .A2(n_24), .B(n_25), .C(n_18), .Y(n_28) );
OAI31xp33_ASAP7_75t_L g29 ( .A1(n_27), .A2(n_17), .A3(n_3), .B(n_4), .Y(n_29) );
OAI22xp33_ASAP7_75t_L g30 ( .A1(n_27), .A2(n_22), .B1(n_20), .B2(n_19), .Y(n_30) );
AND2x2_ASAP7_75t_L g31 ( .A(n_29), .B(n_28), .Y(n_31) );
NOR2xp33_ASAP7_75t_L g32 ( .A(n_30), .B(n_22), .Y(n_32) );
NOR3xp33_ASAP7_75t_SL g33 ( .A(n_32), .B(n_29), .C(n_20), .Y(n_33) );
INVx1_ASAP7_75t_L g34 ( .A(n_31), .Y(n_34) );
AOI22xp5_ASAP7_75t_L g35 ( .A1(n_33), .A2(n_19), .B1(n_18), .B2(n_3), .Y(n_35) );
NAND2xp5_ASAP7_75t_L g36 ( .A(n_34), .B(n_2), .Y(n_36) );
AND2x2_ASAP7_75t_L g37 ( .A(n_33), .B(n_19), .Y(n_37) );
AOI221xp5_ASAP7_75t_SL g38 ( .A1(n_37), .A2(n_11), .B1(n_15), .B2(n_36), .C(n_35), .Y(n_38) );
INVxp67_ASAP7_75t_SL g39 ( .A(n_36), .Y(n_39) );
INVx1_ASAP7_75t_L g40 ( .A(n_36), .Y(n_40) );
HB1xp67_ASAP7_75t_L g41 ( .A(n_39), .Y(n_41) );
INVx1_ASAP7_75t_L g42 ( .A(n_40), .Y(n_42) );
NAND3xp33_ASAP7_75t_L g43 ( .A(n_41), .B(n_38), .C(n_42), .Y(n_43) );
endmodule