module fake_jpeg_24813_n_306 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_306);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_306;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_181;
wire n_38;
wire n_26;
wire n_28;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_288;
wire n_272;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_303;
wire n_90;
wire n_304;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_300;
wire n_211;
wire n_299;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_93;
wire n_91;
wire n_54;
wire n_227;
wire n_305;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_282;
wire n_96;

INVx6_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_13),
.B(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_16),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_14),
.B(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx24_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_25),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_37),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_22),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

BUFx10_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_42),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_46),
.Y(n_58)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g50 ( 
.A(n_44),
.Y(n_50)
);

BUFx16f_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_22),
.Y(n_46)
);

AOI21xp33_ASAP7_75t_L g47 ( 
.A1(n_36),
.A2(n_33),
.B(n_25),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_47),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_44),
.A2(n_17),
.B1(n_23),
.B2(n_20),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_48),
.A2(n_52),
.B1(n_62),
.B2(n_63),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_44),
.A2(n_17),
.B1(n_23),
.B2(n_20),
.Y(n_52)
);

AO22x1_ASAP7_75t_SL g53 ( 
.A1(n_39),
.A2(n_18),
.B1(n_19),
.B2(n_17),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_53),
.A2(n_60),
.B1(n_64),
.B2(n_67),
.Y(n_71)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_56),
.B(n_57),
.Y(n_78)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_59),
.B(n_61),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_40),
.A2(n_17),
.B1(n_20),
.B2(n_23),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_44),
.A2(n_26),
.B1(n_18),
.B2(n_27),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_44),
.A2(n_26),
.B1(n_18),
.B2(n_27),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_40),
.A2(n_26),
.B1(n_18),
.B2(n_30),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_36),
.B(n_29),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_66),
.B(n_37),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_40),
.A2(n_29),
.B1(n_34),
.B2(n_27),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_39),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_49),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_70),
.B(n_81),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_64),
.A2(n_19),
.B1(n_43),
.B2(n_42),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_72),
.A2(n_74),
.B1(n_80),
.B2(n_59),
.Y(n_120)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_73),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_L g74 ( 
.A1(n_53),
.A2(n_19),
.B1(n_35),
.B2(n_39),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_58),
.B(n_46),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_75),
.B(n_83),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_77),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_48),
.A2(n_43),
.B1(n_42),
.B2(n_34),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_82),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_58),
.B(n_49),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_84),
.B(n_90),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_47),
.B(n_46),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_85),
.B(n_87),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_53),
.A2(n_60),
.B1(n_43),
.B2(n_42),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_86),
.A2(n_93),
.B1(n_94),
.B2(n_97),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_55),
.B(n_46),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_53),
.B(n_39),
.C(n_45),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_89),
.B(n_41),
.Y(n_108)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_67),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_91),
.B(n_92),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_65),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_53),
.A2(n_39),
.B1(n_29),
.B2(n_30),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_62),
.A2(n_39),
.B1(n_30),
.B2(n_32),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_51),
.B(n_37),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_95),
.B(n_96),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_52),
.A2(n_35),
.B1(n_32),
.B2(n_34),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_65),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_98),
.B(n_99),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_65),
.Y(n_99)
);

BUFx24_ASAP7_75t_SL g103 ( 
.A(n_70),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_103),
.B(n_123),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_83),
.B(n_63),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_105),
.B(n_118),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_108),
.B(n_111),
.C(n_127),
.Y(n_137)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_95),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_110),
.B(n_128),
.Y(n_146)
);

AND2x6_ASAP7_75t_L g111 ( 
.A(n_76),
.B(n_11),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_89),
.B(n_50),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_112),
.A2(n_121),
.B(n_124),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_76),
.A2(n_50),
.B1(n_69),
.B2(n_61),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_113),
.A2(n_117),
.B1(n_125),
.B2(n_73),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_90),
.A2(n_61),
.B1(n_59),
.B2(n_57),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_114),
.A2(n_99),
.B1(n_98),
.B2(n_91),
.Y(n_157)
);

AO22x2_ASAP7_75t_L g117 ( 
.A1(n_71),
.A2(n_41),
.B1(n_56),
.B2(n_45),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_75),
.B(n_45),
.Y(n_118)
);

A2O1A1Ixp33_ASAP7_75t_SL g156 ( 
.A1(n_120),
.A2(n_97),
.B(n_35),
.C(n_73),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_89),
.B(n_0),
.Y(n_121)
);

INVx13_ASAP7_75t_L g123 ( 
.A(n_77),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_96),
.B(n_0),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_88),
.A2(n_69),
.B1(n_68),
.B2(n_56),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_88),
.A2(n_68),
.B1(n_69),
.B2(n_32),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_126),
.A2(n_94),
.B1(n_93),
.B2(n_84),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_85),
.A2(n_54),
.B(n_41),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_78),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_102),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_129),
.B(n_136),
.Y(n_176)
);

AOI22x1_ASAP7_75t_SL g131 ( 
.A1(n_117),
.A2(n_71),
.B1(n_72),
.B2(n_94),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_131),
.A2(n_125),
.B1(n_106),
.B2(n_121),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_102),
.B(n_81),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_132),
.B(n_143),
.Y(n_183)
);

BUFx4f_ASAP7_75t_L g134 ( 
.A(n_107),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_134),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_115),
.B(n_87),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_135),
.B(n_150),
.Y(n_172)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_122),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_138),
.A2(n_139),
.B1(n_147),
.B2(n_148),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_117),
.A2(n_105),
.B1(n_127),
.B2(n_116),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_122),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_140),
.B(n_141),
.Y(n_179)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_119),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_113),
.B(n_86),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_142),
.A2(n_121),
.B(n_100),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_115),
.B(n_93),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_119),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_144),
.B(n_145),
.Y(n_184)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_104),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_117),
.A2(n_116),
.B1(n_120),
.B2(n_106),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_101),
.B(n_78),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_104),
.B(n_79),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_151),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_108),
.B(n_82),
.C(n_92),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_152),
.B(n_159),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_110),
.B(n_79),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_153),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_101),
.B(n_80),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_154),
.B(n_124),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_123),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_155),
.B(n_158),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_156),
.A2(n_123),
.B1(n_109),
.B2(n_100),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_157),
.A2(n_117),
.B1(n_109),
.B2(n_126),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_128),
.B(n_22),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g159 ( 
.A(n_112),
.B(n_21),
.Y(n_159)
);

NOR4xp25_ASAP7_75t_L g160 ( 
.A(n_149),
.B(n_118),
.C(n_112),
.D(n_111),
.Y(n_160)
);

A2O1A1O1Ixp25_ASAP7_75t_L g202 ( 
.A1(n_160),
.A2(n_156),
.B(n_142),
.C(n_136),
.D(n_144),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_161),
.A2(n_147),
.B1(n_156),
.B2(n_145),
.Y(n_203)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_146),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_162),
.B(n_166),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_165),
.A2(n_168),
.B1(n_192),
.B2(n_41),
.Y(n_216)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_146),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_134),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_167),
.B(n_170),
.Y(n_214)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_134),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_134),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_171),
.B(n_175),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_150),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_177),
.A2(n_178),
.B(n_181),
.Y(n_219)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_132),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_180),
.B(n_185),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_143),
.A2(n_124),
.B(n_33),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_139),
.B(n_21),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_182),
.B(n_28),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_135),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_154),
.B(n_77),
.Y(n_186)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_186),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_149),
.B(n_77),
.Y(n_188)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_188),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_130),
.B(n_54),
.Y(n_189)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_189),
.Y(n_217)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_157),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_190),
.B(n_191),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_141),
.B(n_37),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_148),
.A2(n_24),
.B1(n_33),
.B2(n_25),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_164),
.A2(n_137),
.B1(n_131),
.B2(n_156),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_194),
.A2(n_216),
.B1(n_54),
.B2(n_24),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_189),
.B(n_152),
.C(n_137),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_195),
.B(n_196),
.C(n_220),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_175),
.B(n_159),
.C(n_130),
.Y(n_196)
);

AND2x2_ASAP7_75t_SL g198 ( 
.A(n_185),
.B(n_140),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_198),
.A2(n_179),
.B(n_184),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_180),
.B(n_133),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_199),
.B(n_205),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_202),
.B(n_179),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_172),
.B(n_45),
.Y(n_204)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_204),
.Y(n_224)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_184),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_161),
.A2(n_164),
.B1(n_186),
.B2(n_165),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_207),
.A2(n_211),
.B1(n_188),
.B2(n_177),
.Y(n_221)
);

NAND3xp33_ASAP7_75t_L g208 ( 
.A(n_162),
.B(n_12),
.C(n_16),
.Y(n_208)
);

OA21x2_ASAP7_75t_SL g225 ( 
.A1(n_208),
.A2(n_215),
.B(n_15),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_163),
.Y(n_210)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_210),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_160),
.A2(n_24),
.B1(n_54),
.B2(n_35),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_172),
.B(n_45),
.Y(n_212)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_212),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_213),
.B(n_28),
.Y(n_235)
);

NAND3xp33_ASAP7_75t_L g215 ( 
.A(n_166),
.B(n_11),
.C(n_16),
.Y(n_215)
);

OAI22x1_ASAP7_75t_SL g218 ( 
.A1(n_168),
.A2(n_192),
.B1(n_178),
.B2(n_182),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_174),
.B(n_54),
.C(n_155),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_221),
.B(n_225),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_214),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_226),
.B(n_234),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_227),
.A2(n_236),
.B(n_217),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_195),
.B(n_174),
.C(n_183),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_228),
.B(n_243),
.C(n_196),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_200),
.B(n_176),
.Y(n_229)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_229),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_218),
.A2(n_169),
.B1(n_176),
.B2(n_173),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_230),
.A2(n_231),
.B1(n_238),
.B2(n_201),
.Y(n_253)
);

OAI22x1_ASAP7_75t_SL g231 ( 
.A1(n_203),
.A2(n_169),
.B1(n_181),
.B2(n_187),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_207),
.A2(n_191),
.B1(n_171),
.B2(n_170),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_233),
.B(n_241),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_198),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_235),
.B(n_213),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_217),
.A2(n_167),
.B(n_54),
.Y(n_236)
);

AOI322xp5_ASAP7_75t_L g240 ( 
.A1(n_219),
.A2(n_155),
.A3(n_15),
.B1(n_14),
.B2(n_13),
.C1(n_12),
.C2(n_11),
.Y(n_240)
);

BUFx24_ASAP7_75t_SL g259 ( 
.A(n_240),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_197),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_197),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_242),
.B(n_209),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_220),
.B(n_0),
.C(n_1),
.Y(n_243)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_245),
.Y(n_263)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_229),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_246),
.B(n_251),
.Y(n_264)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_248),
.Y(n_266)
);

AOI21x1_ASAP7_75t_L g249 ( 
.A1(n_234),
.A2(n_198),
.B(n_201),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g273 ( 
.A(n_249),
.B(n_194),
.Y(n_273)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_227),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_236),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_252),
.B(n_206),
.Y(n_268)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_253),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_254),
.B(n_255),
.C(n_222),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_241),
.A2(n_200),
.B(n_206),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_256),
.A2(n_239),
.B1(n_224),
.B2(n_204),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_230),
.B(n_193),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_257),
.B(n_221),
.Y(n_262)
);

BUFx12_ASAP7_75t_L g260 ( 
.A(n_231),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_260),
.B(n_238),
.Y(n_272)
);

FAx1_ASAP7_75t_L g261 ( 
.A(n_223),
.B(n_242),
.CI(n_212),
.CON(n_261),
.SN(n_261)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_261),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_262),
.B(n_270),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_267),
.A2(n_269),
.B(n_271),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_268),
.A2(n_272),
.B(n_274),
.Y(n_278)
);

OAI321xp33_ASAP7_75t_L g269 ( 
.A1(n_256),
.A2(n_248),
.A3(n_247),
.B1(n_246),
.B2(n_202),
.C(n_258),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_255),
.B(n_222),
.C(n_228),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_251),
.B(n_224),
.C(n_239),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_273),
.B(n_276),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_244),
.B(n_209),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_266),
.A2(n_275),
.B1(n_265),
.B2(n_252),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_281),
.A2(n_280),
.B1(n_235),
.B2(n_259),
.Y(n_291)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_263),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_282),
.B(n_253),
.Y(n_288)
);

OAI21xp33_ASAP7_75t_L g283 ( 
.A1(n_264),
.A2(n_274),
.B(n_268),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_266),
.A2(n_249),
.B(n_250),
.Y(n_284)
);

OR2x2_ASAP7_75t_L g285 ( 
.A(n_283),
.B(n_264),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_285),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_279),
.B(n_270),
.C(n_267),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_286),
.B(n_287),
.C(n_12),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_277),
.B(n_245),
.C(n_232),
.Y(n_287)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_288),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_278),
.B(n_237),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_289),
.B(n_290),
.Y(n_293)
);

OR2x2_ASAP7_75t_L g290 ( 
.A(n_278),
.B(n_284),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_291),
.B(n_292),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_281),
.B(n_13),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_SL g298 ( 
.A(n_294),
.B(n_286),
.C(n_6),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_298),
.A2(n_300),
.B(n_297),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_293),
.Y(n_299)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_299),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_296),
.A2(n_5),
.B(n_6),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_298),
.B(n_295),
.C(n_293),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_301),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_304),
.B(n_302),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_305),
.B(n_303),
.Y(n_306)
);


endmodule