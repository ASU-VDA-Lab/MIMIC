module fake_jpeg_30492_n_228 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_228);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_228;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx11_ASAP7_75t_SL g26 ( 
.A(n_4),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_13),
.B(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_29),
.B(n_0),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_34),
.B(n_36),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_35),
.B(n_39),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_2),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_21),
.B(n_2),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

CKINVDCx5p33_ASAP7_75t_R g42 ( 
.A(n_26),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_44),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_26),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_43),
.Y(n_45)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_40),
.A2(n_27),
.B1(n_32),
.B2(n_24),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_47),
.A2(n_48),
.B1(n_69),
.B2(n_44),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_40),
.A2(n_27),
.B1(n_32),
.B2(n_24),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_25),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_49),
.B(n_65),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_38),
.A2(n_32),
.B1(n_24),
.B2(n_20),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_50),
.Y(n_103)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_38),
.A2(n_32),
.B1(n_24),
.B2(n_20),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_53),
.Y(n_81)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_56),
.Y(n_93)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_58),
.B(n_71),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_34),
.B(n_23),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_60),
.B(n_61),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_34),
.B(n_35),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

CKINVDCx14_ASAP7_75t_R g86 ( 
.A(n_62),
.Y(n_86)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_36),
.B(n_16),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_66),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_37),
.A2(n_17),
.B1(n_25),
.B2(n_19),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_67),
.A2(n_73),
.B1(n_44),
.B2(n_33),
.Y(n_91)
);

BUFx10_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_68),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_41),
.A2(n_16),
.B1(n_25),
.B2(n_19),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_39),
.B(n_18),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_37),
.A2(n_16),
.B1(n_19),
.B2(n_23),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_74),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_71),
.B(n_31),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_75),
.B(n_85),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_49),
.A2(n_18),
.B(n_23),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_76),
.A2(n_46),
.B(n_62),
.Y(n_122)
);

OAI22x1_ASAP7_75t_SL g78 ( 
.A1(n_64),
.A2(n_65),
.B1(n_42),
.B2(n_68),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_78),
.A2(n_70),
.B1(n_62),
.B2(n_8),
.Y(n_125)
);

A2O1A1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_64),
.A2(n_18),
.B(n_31),
.C(n_30),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_80),
.B(n_87),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_54),
.B(n_30),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_68),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_88),
.B(n_72),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_68),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_89),
.B(n_96),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_91),
.A2(n_45),
.B1(n_63),
.B2(n_59),
.Y(n_119)
);

OAI32xp33_ASAP7_75t_L g92 ( 
.A1(n_64),
.A2(n_28),
.A3(n_22),
.B1(n_21),
.B2(n_7),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_98),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_57),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_57),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_70),
.Y(n_99)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_99),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_54),
.B(n_28),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_100),
.B(n_102),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_61),
.A2(n_22),
.B1(n_5),
.B2(n_6),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_101),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_60),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_95),
.B(n_52),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_104),
.B(n_80),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_95),
.B(n_66),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_107),
.B(n_114),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_77),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_111),
.B(n_112),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_77),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_81),
.A2(n_58),
.B1(n_55),
.B2(n_51),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_113),
.A2(n_83),
.B(n_74),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_56),
.Y(n_114)
);

NOR3xp33_ASAP7_75t_SL g115 ( 
.A(n_78),
.B(n_45),
.C(n_46),
.Y(n_115)
);

NOR3xp33_ASAP7_75t_L g148 ( 
.A(n_115),
.B(n_86),
.C(n_83),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_90),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_116),
.B(n_120),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_117),
.A2(n_88),
.B1(n_111),
.B2(n_119),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_118),
.A2(n_76),
.B1(n_103),
.B2(n_101),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_119),
.A2(n_89),
.B1(n_87),
.B2(n_82),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_90),
.B(n_72),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_94),
.B(n_59),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_121),
.B(n_130),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_122),
.B(n_125),
.Y(n_139)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_97),
.Y(n_124)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_124),
.Y(n_140)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_97),
.Y(n_126)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_126),
.Y(n_147)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_93),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_128),
.Y(n_155)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_93),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_129),
.B(n_3),
.Y(n_152)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_79),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_90),
.B(n_62),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_131),
.B(n_9),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_123),
.B(n_94),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_134),
.B(n_142),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_135),
.B(n_141),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_136),
.B(n_131),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_105),
.A2(n_92),
.B(n_91),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_137),
.A2(n_149),
.B(n_120),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_127),
.B(n_82),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_144),
.A2(n_145),
.B1(n_153),
.B2(n_122),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_117),
.A2(n_115),
.B1(n_104),
.B2(n_107),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_109),
.B(n_79),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_146),
.B(n_118),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_148),
.B(n_150),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_117),
.A2(n_99),
.B1(n_84),
.B2(n_8),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_116),
.A2(n_84),
.B1(n_6),
.B2(n_8),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_151),
.B(n_154),
.Y(n_166)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_152),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_114),
.A2(n_3),
.B1(n_9),
.B2(n_11),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_156),
.B(n_171),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_133),
.B(n_108),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_157),
.B(n_161),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_160),
.A2(n_139),
.B(n_144),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_163),
.A2(n_139),
.B1(n_135),
.B2(n_141),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_143),
.B(n_129),
.C(n_106),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_165),
.B(n_167),
.C(n_147),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_143),
.B(n_106),
.C(n_124),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_132),
.Y(n_168)
);

INVx3_ASAP7_75t_SL g187 ( 
.A(n_168),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_138),
.B(n_126),
.Y(n_169)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_169),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_151),
.B(n_110),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_170),
.Y(n_185)
);

MAJx2_ASAP7_75t_L g171 ( 
.A(n_138),
.B(n_14),
.C(n_15),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_136),
.B(n_110),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_172),
.A2(n_158),
.B1(n_166),
.B2(n_168),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_140),
.Y(n_173)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_173),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_175),
.B(n_186),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_156),
.B(n_145),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_176),
.B(n_180),
.C(n_163),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_177),
.Y(n_191)
);

NOR2xp67_ASAP7_75t_SL g178 ( 
.A(n_160),
.B(n_149),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_178),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_158),
.B(n_154),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_181),
.B(n_188),
.Y(n_189)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_169),
.Y(n_184)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_184),
.Y(n_200)
);

OA21x2_ASAP7_75t_SL g186 ( 
.A1(n_159),
.A2(n_137),
.B(n_139),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_181),
.B(n_167),
.C(n_165),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_190),
.B(n_194),
.Y(n_202)
);

AOI21xp33_ASAP7_75t_L g192 ( 
.A1(n_183),
.A2(n_162),
.B(n_164),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_192),
.A2(n_187),
.B(n_179),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_174),
.B(n_164),
.C(n_171),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_195),
.B(n_180),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_174),
.B(n_173),
.C(n_162),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_196),
.B(n_198),
.C(n_182),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_176),
.B(n_166),
.C(n_155),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_185),
.A2(n_150),
.B1(n_155),
.B2(n_153),
.Y(n_199)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_199),
.Y(n_205)
);

OAI21x1_ASAP7_75t_L g201 ( 
.A1(n_197),
.A2(n_187),
.B(n_178),
.Y(n_201)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_201),
.Y(n_214)
);

AOI31xp67_ASAP7_75t_L g203 ( 
.A1(n_191),
.A2(n_187),
.A3(n_175),
.B(n_177),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_203),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_204),
.A2(n_206),
.B(n_207),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_189),
.B(n_184),
.C(n_179),
.Y(n_207)
);

AOI21x1_ASAP7_75t_L g216 ( 
.A1(n_208),
.A2(n_193),
.B(n_189),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_191),
.A2(n_182),
.B1(n_140),
.B2(n_147),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_209),
.A2(n_210),
.B1(n_193),
.B2(n_195),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_200),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_211),
.B(n_213),
.Y(n_219)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_205),
.Y(n_213)
);

NAND2xp33_ASAP7_75t_SL g220 ( 
.A(n_216),
.B(n_209),
.Y(n_220)
);

MAJx2_ASAP7_75t_L g217 ( 
.A(n_214),
.B(n_202),
.C(n_206),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_217),
.A2(n_218),
.B(n_220),
.Y(n_223)
);

OAI21xp33_ASAP7_75t_L g218 ( 
.A1(n_212),
.A2(n_207),
.B(n_204),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_219),
.B(n_211),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_221),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_219),
.B(n_213),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_222),
.A2(n_210),
.B(n_215),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_225),
.B(n_12),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_224),
.A2(n_223),
.B(n_12),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_226),
.B(n_227),
.Y(n_228)
);


endmodule