module fake_jpeg_27860_n_255 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_255);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_255;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_15),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_21),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_34),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g34 ( 
.A(n_17),
.Y(n_34)
);

INVx6_ASAP7_75t_SL g35 ( 
.A(n_24),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_16),
.B(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_43),
.Y(n_56)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_21),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_39),
.A2(n_22),
.B1(n_20),
.B2(n_19),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_44),
.A2(n_50),
.B1(n_53),
.B2(n_34),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_25),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_45),
.B(n_47),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_40),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_39),
.A2(n_22),
.B1(n_32),
.B2(n_27),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_34),
.A2(n_22),
.B1(n_20),
.B2(n_19),
.Y(n_53)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_55),
.B(n_63),
.Y(n_67)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_17),
.C(n_18),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_58),
.B(n_37),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_33),
.B(n_25),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_16),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_43),
.B(n_23),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_61),
.B(n_64),
.Y(n_88)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_23),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_38),
.A2(n_32),
.B1(n_27),
.B2(n_30),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_65),
.A2(n_34),
.B1(n_32),
.B2(n_27),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_64),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_69),
.B(n_71),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_48),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_61),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_72),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_73),
.B(n_75),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_48),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_74),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_26),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_56),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_46),
.Y(n_93)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_54),
.B(n_26),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_78),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_55),
.A2(n_30),
.B1(n_29),
.B2(n_28),
.Y(n_79)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_79),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_80),
.A2(n_85),
.B1(n_35),
.B2(n_38),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_59),
.Y(n_100)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_83),
.Y(n_112)
);

CKINVDCx12_ASAP7_75t_R g84 ( 
.A(n_46),
.Y(n_84)
);

NAND3xp33_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_41),
.C(n_57),
.Y(n_102)
);

OA22x2_ASAP7_75t_L g85 ( 
.A1(n_58),
.A2(n_38),
.B1(n_41),
.B2(n_37),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_86),
.A2(n_63),
.B(n_52),
.Y(n_95)
);

AND2x6_ASAP7_75t_L g89 ( 
.A(n_86),
.B(n_15),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_89),
.B(n_102),
.Y(n_128)
);

OR2x4_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_71),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_92),
.A2(n_108),
.B(n_54),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_93),
.B(n_104),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_85),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_74),
.B(n_59),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_103),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_98),
.A2(n_105),
.B1(n_82),
.B2(n_84),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_100),
.A2(n_81),
.B1(n_69),
.B2(n_85),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_67),
.B(n_59),
.Y(n_103)
);

OAI211xp5_ASAP7_75t_L g104 ( 
.A1(n_70),
.A2(n_16),
.B(n_26),
.C(n_31),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_77),
.A2(n_49),
.B1(n_62),
.B2(n_35),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_87),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_106),
.B(n_110),
.Y(n_114)
);

AOI32xp33_ASAP7_75t_L g108 ( 
.A1(n_86),
.A2(n_52),
.A3(n_42),
.B1(n_36),
.B2(n_37),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_67),
.B(n_49),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_109),
.B(n_79),
.Y(n_118)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_68),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_113),
.A2(n_133),
.B1(n_112),
.B2(n_110),
.Y(n_145)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_97),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_118),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_116),
.B(n_129),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_119),
.A2(n_107),
.B1(n_96),
.B2(n_99),
.Y(n_138)
);

CKINVDCx14_ASAP7_75t_R g120 ( 
.A(n_93),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_120),
.B(n_121),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_94),
.B(n_72),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_94),
.B(n_88),
.Y(n_123)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_123),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_88),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_124),
.B(n_126),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_103),
.B(n_109),
.Y(n_125)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_125),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_91),
.B(n_88),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_91),
.B(n_85),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_131),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_129),
.A2(n_29),
.B(n_28),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_92),
.B(n_87),
.Y(n_130)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_130),
.Y(n_147)
);

INVx1_ASAP7_75t_SL g131 ( 
.A(n_100),
.Y(n_131)
);

O2A1O1Ixp33_ASAP7_75t_L g132 ( 
.A1(n_90),
.A2(n_51),
.B(n_68),
.C(n_37),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_132),
.A2(n_68),
.B(n_83),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_98),
.A2(n_51),
.B1(n_83),
.B2(n_37),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_105),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_134),
.B(n_68),
.Y(n_153)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_106),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_135),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_138),
.A2(n_142),
.B(n_145),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_119),
.A2(n_107),
.B1(n_96),
.B2(n_99),
.Y(n_140)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_140),
.Y(n_161)
);

OAI22x1_ASAP7_75t_L g142 ( 
.A1(n_131),
.A2(n_108),
.B1(n_89),
.B2(n_95),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_143),
.B(n_154),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_127),
.A2(n_112),
.B(n_111),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_146),
.B(n_149),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_114),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_150),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_123),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_151),
.Y(n_180)
);

INVx11_ASAP7_75t_L g152 ( 
.A(n_132),
.Y(n_152)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_152),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_153),
.B(n_155),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_116),
.B(n_24),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_130),
.B(n_66),
.C(n_42),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_115),
.B(n_66),
.C(n_42),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_157),
.B(n_158),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_117),
.B(n_24),
.C(n_31),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_159),
.B(n_133),
.Y(n_175)
);

NOR3xp33_ASAP7_75t_L g160 ( 
.A(n_142),
.B(n_126),
.C(n_128),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_160),
.B(n_165),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_139),
.B(n_118),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_164),
.B(n_168),
.Y(n_189)
);

NAND3xp33_ASAP7_75t_L g165 ( 
.A(n_137),
.B(n_122),
.C(n_128),
.Y(n_165)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_137),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_167),
.B(n_176),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_150),
.B(n_122),
.Y(n_168)
);

BUFx12_ASAP7_75t_L g170 ( 
.A(n_156),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_170),
.B(n_175),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_136),
.B(n_117),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_172),
.B(n_173),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_138),
.B(n_113),
.Y(n_173)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_157),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_141),
.B(n_125),
.Y(n_177)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_177),
.Y(n_181)
);

INVx2_ASAP7_75t_SL g178 ( 
.A(n_149),
.Y(n_178)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_178),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_174),
.B(n_143),
.C(n_154),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_182),
.B(n_183),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_174),
.B(n_144),
.C(n_141),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_178),
.A2(n_147),
.B1(n_146),
.B2(n_134),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_184),
.A2(n_166),
.B(n_163),
.Y(n_213)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_179),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_186),
.B(n_187),
.Y(n_209)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_179),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_161),
.A2(n_147),
.B1(n_140),
.B2(n_144),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_188),
.A2(n_161),
.B1(n_169),
.B2(n_178),
.Y(n_199)
);

BUFx12f_ASAP7_75t_L g190 ( 
.A(n_170),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_190),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_162),
.B(n_159),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_191),
.B(n_195),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_176),
.B(n_155),
.C(n_148),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_171),
.Y(n_197)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_197),
.Y(n_200)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_171),
.Y(n_198)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_198),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_199),
.A2(n_208),
.B1(n_209),
.B2(n_213),
.Y(n_225)
);

NOR2xp67_ASAP7_75t_R g201 ( 
.A(n_184),
.B(n_166),
.Y(n_201)
);

OR2x2_ASAP7_75t_L g217 ( 
.A(n_201),
.B(n_191),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_194),
.A2(n_180),
.B1(n_169),
.B2(n_167),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_204),
.A2(n_181),
.B1(n_188),
.B2(n_152),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_189),
.B(n_180),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_205),
.B(n_207),
.Y(n_215)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_192),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_185),
.A2(n_166),
.B(n_162),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_208),
.B(n_210),
.Y(n_219)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_192),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_196),
.Y(n_211)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_211),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_213),
.B(n_190),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_216),
.B(n_218),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_217),
.B(n_220),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_201),
.A2(n_207),
.B1(n_202),
.B2(n_200),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_206),
.B(n_195),
.C(n_183),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_212),
.A2(n_193),
.B1(n_158),
.B2(n_182),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_221),
.B(n_222),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_206),
.B(n_190),
.C(n_170),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_223),
.B(n_31),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_203),
.B(n_24),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_224),
.B(n_24),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_225),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_215),
.A2(n_209),
.B(n_199),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_226),
.B(n_230),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_228),
.B(n_223),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_229),
.B(n_231),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_219),
.B(n_14),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_224),
.B(n_13),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_234),
.B(n_12),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_236),
.B(n_237),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_227),
.B(n_220),
.C(n_222),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_233),
.A2(n_214),
.B(n_217),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_238),
.A2(n_1),
.B(n_2),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_232),
.Y(n_240)
);

OR2x2_ASAP7_75t_L g246 ( 
.A(n_240),
.B(n_241),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_240),
.A2(n_231),
.B1(n_229),
.B2(n_3),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_242),
.B(n_243),
.C(n_235),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_239),
.B(n_1),
.Y(n_243)
);

AOI322xp5_ASAP7_75t_L g248 ( 
.A1(n_244),
.A2(n_2),
.A3(n_3),
.B1(n_4),
.B2(n_6),
.C1(n_7),
.C2(n_8),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_247),
.B(n_248),
.C(n_249),
.Y(n_251)
);

AOI322xp5_ASAP7_75t_L g249 ( 
.A1(n_245),
.A2(n_4),
.A3(n_6),
.B1(n_9),
.B2(n_10),
.C1(n_11),
.C2(n_246),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_246),
.B(n_243),
.C(n_10),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_250),
.B(n_9),
.C(n_11),
.Y(n_252)
);

BUFx24_ASAP7_75t_SL g253 ( 
.A(n_252),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_253),
.B(n_251),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_254),
.B(n_11),
.Y(n_255)
);


endmodule