module real_jpeg_2813_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_202;
wire n_128;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_215;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_1),
.A2(n_62),
.B1(n_63),
.B2(n_75),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_1),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_1),
.A2(n_69),
.B1(n_71),
.B2(n_75),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_1),
.A2(n_46),
.B1(n_48),
.B2(n_75),
.Y(n_157)
);

OAI22xp33_ASAP7_75t_L g202 ( 
.A1(n_1),
.A2(n_34),
.B1(n_41),
.B2(n_75),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_2),
.A2(n_62),
.B1(n_63),
.B2(n_185),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_2),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_2),
.A2(n_69),
.B1(n_71),
.B2(n_185),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_2),
.A2(n_46),
.B1(n_48),
.B2(n_185),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_2),
.A2(n_34),
.B1(n_41),
.B2(n_185),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_3),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_4),
.A2(n_46),
.B1(n_48),
.B2(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_4),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_4),
.A2(n_55),
.B1(n_69),
.B2(n_71),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_4),
.A2(n_34),
.B1(n_41),
.B2(n_55),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_4),
.A2(n_55),
.B1(n_62),
.B2(n_63),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_6),
.B(n_62),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_6),
.B(n_166),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_6),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_6),
.A2(n_62),
.B(n_175),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_6),
.B(n_84),
.Y(n_237)
);

AOI21xp33_ASAP7_75t_L g244 ( 
.A1(n_6),
.A2(n_71),
.B(n_245),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_6),
.B(n_34),
.C(n_51),
.Y(n_253)
);

OAI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_6),
.A2(n_46),
.B1(n_48),
.B2(n_211),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_6),
.B(n_37),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_6),
.B(n_56),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_7),
.A2(n_62),
.B1(n_63),
.B2(n_131),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_7),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_7),
.A2(n_69),
.B1(n_71),
.B2(n_131),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_7),
.A2(n_46),
.B1(n_48),
.B2(n_131),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_7),
.A2(n_34),
.B1(n_41),
.B2(n_131),
.Y(n_239)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_8),
.Y(n_333)
);

BUFx8_ASAP7_75t_L g64 ( 
.A(n_9),
.Y(n_64)
);

BUFx16f_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_11),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_12),
.A2(n_21),
.B(n_332),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_12),
.B(n_333),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_13),
.A2(n_62),
.B1(n_63),
.B2(n_165),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_13),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_13),
.A2(n_69),
.B1(n_71),
.B2(n_165),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_13),
.A2(n_46),
.B1(n_48),
.B2(n_165),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_13),
.A2(n_34),
.B1(n_41),
.B2(n_165),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_14),
.A2(n_45),
.B1(n_46),
.B2(n_48),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_14),
.A2(n_45),
.B1(n_69),
.B2(n_71),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_14),
.A2(n_45),
.B1(n_62),
.B2(n_63),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_14),
.A2(n_34),
.B1(n_41),
.B2(n_45),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_15),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_16),
.A2(n_62),
.B1(n_63),
.B2(n_73),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_16),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_16),
.A2(n_69),
.B1(n_71),
.B2(n_73),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_16),
.A2(n_46),
.B1(n_48),
.B2(n_73),
.Y(n_207)
);

OAI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_16),
.A2(n_34),
.B1(n_41),
.B2(n_73),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_17),
.A2(n_69),
.B1(n_71),
.B2(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_17),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_17),
.A2(n_62),
.B1(n_63),
.B2(n_81),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_17),
.A2(n_46),
.B1(n_48),
.B2(n_81),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_17),
.A2(n_34),
.B1(n_41),
.B2(n_81),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_18),
.A2(n_34),
.B1(n_40),
.B2(n_41),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_18),
.A2(n_40),
.B1(n_46),
.B2(n_48),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_18),
.A2(n_40),
.B1(n_69),
.B2(n_71),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_18),
.A2(n_40),
.B1(n_62),
.B2(n_63),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

AOI21xp33_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_327),
.B(n_330),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_319),
.B(n_323),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_306),
.B(n_318),
.Y(n_23)
);

AO21x1_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_145),
.B(n_303),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_132),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_105),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_27),
.B(n_105),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_76),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_28),
.B(n_91),
.C(n_103),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_57),
.B(n_58),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_29),
.A2(n_30),
.B1(n_108),
.B2(n_109),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_42),
.Y(n_30)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_31),
.A2(n_57),
.B1(n_58),
.B2(n_110),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_31),
.A2(n_42),
.B1(n_43),
.B2(n_57),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_36),
.B(n_38),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_32),
.A2(n_36),
.B1(n_119),
.B2(n_160),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_32),
.A2(n_36),
.B1(n_214),
.B2(n_216),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_32),
.A2(n_36),
.B1(n_273),
.B2(n_274),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_33),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_33),
.A2(n_37),
.B1(n_39),
.B2(n_118),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_33),
.A2(n_37),
.B1(n_178),
.B2(n_179),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_33),
.A2(n_37),
.B1(n_178),
.B2(n_202),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_33),
.A2(n_37),
.B1(n_215),
.B2(n_239),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_33),
.A2(n_37),
.B1(n_211),
.B2(n_265),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_33),
.A2(n_37),
.B1(n_265),
.B2(n_269),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_36),
.Y(n_33)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

OA22x2_ASAP7_75t_L g53 ( 
.A1(n_34),
.A2(n_41),
.B1(n_51),
.B2(n_52),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_34),
.B(n_263),
.Y(n_262)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_49),
.B1(n_54),
.B2(n_56),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_44),
.A2(n_49),
.B1(n_56),
.B2(n_122),
.Y(n_121)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_46),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_L g50 ( 
.A1(n_46),
.A2(n_48),
.B1(n_51),
.B2(n_52),
.Y(n_50)
);

AO22x2_ASAP7_75t_SL g84 ( 
.A1(n_46),
.A2(n_48),
.B1(n_85),
.B2(n_86),
.Y(n_84)
);

OAI32xp33_ASAP7_75t_L g209 ( 
.A1(n_46),
.A2(n_71),
.A3(n_85),
.B1(n_210),
.B2(n_212),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_46),
.B(n_253),
.Y(n_252)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_48),
.B(n_86),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_49),
.A2(n_54),
.B1(n_56),
.B2(n_90),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_49),
.A2(n_56),
.B(n_90),
.Y(n_97)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_49),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_49),
.A2(n_56),
.B1(n_205),
.B2(n_207),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_49),
.A2(n_56),
.B1(n_207),
.B2(n_227),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_49),
.A2(n_56),
.B1(n_235),
.B2(n_236),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_49),
.A2(n_56),
.B1(n_235),
.B2(n_256),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_53),
.Y(n_49)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_51),
.Y(n_52)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_53),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_53),
.A2(n_123),
.B1(n_157),
.B2(n_158),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_53),
.A2(n_158),
.B1(n_206),
.B2(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_58),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_68),
.B1(n_72),
.B2(n_74),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_59),
.A2(n_68),
.B1(n_74),
.B2(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_59),
.A2(n_68),
.B1(n_72),
.B2(n_129),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_59),
.A2(n_68),
.B1(n_94),
.B2(n_142),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_59),
.A2(n_68),
.B1(n_184),
.B2(n_186),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_59),
.A2(n_68),
.B1(n_184),
.B2(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_60),
.A2(n_130),
.B1(n_164),
.B2(n_166),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_60),
.A2(n_166),
.B1(n_313),
.B2(n_314),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_60),
.A2(n_166),
.B1(n_314),
.B2(n_321),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_60),
.A2(n_166),
.B(n_321),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_68),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_63),
.B1(n_65),
.B2(n_67),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AOI32xp33_ASAP7_75t_L g174 ( 
.A1(n_63),
.A2(n_67),
.A3(n_71),
.B1(n_175),
.B2(n_176),
.Y(n_174)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx6_ASAP7_75t_SL g67 ( 
.A(n_65),
.Y(n_67)
);

OA22x2_ASAP7_75t_L g68 ( 
.A1(n_65),
.A2(n_67),
.B1(n_69),
.B2(n_71),
.Y(n_68)
);

NAND2xp33_ASAP7_75t_SL g176 ( 
.A(n_65),
.B(n_69),
.Y(n_176)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_68),
.Y(n_166)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_69),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_69),
.A2(n_71),
.B1(n_85),
.B2(n_86),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_69),
.B(n_211),
.Y(n_210)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_91),
.B1(n_103),
.B2(n_104),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_77),
.Y(n_103)
);

OAI21xp33_ASAP7_75t_L g112 ( 
.A1(n_77),
.A2(n_78),
.B(n_89),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_89),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_82),
.B1(n_84),
.B2(n_88),
.Y(n_78)
);

INVxp33_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_80),
.A2(n_83),
.B1(n_125),
.B2(n_127),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_82),
.A2(n_84),
.B1(n_88),
.B2(n_100),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_82),
.A2(n_84),
.B1(n_126),
.B2(n_162),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_82),
.A2(n_84),
.B(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_83),
.A2(n_101),
.B1(n_127),
.B2(n_140),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_83),
.A2(n_127),
.B1(n_181),
.B2(n_182),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_83),
.A2(n_127),
.B1(n_196),
.B2(n_197),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_83),
.A2(n_127),
.B1(n_181),
.B2(n_197),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_83),
.A2(n_127),
.B1(n_196),
.B2(n_244),
.Y(n_243)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_87),
.Y(n_83)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_84),
.Y(n_127)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_85),
.Y(n_86)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_91),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_93),
.B1(n_95),
.B2(n_96),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_92),
.A2(n_93),
.B1(n_135),
.B2(n_136),
.Y(n_134)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_93),
.B(n_97),
.C(n_99),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_93),
.B(n_136),
.C(n_143),
.Y(n_307)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_98),
.B1(n_99),
.B2(n_102),
.Y(n_96)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_97),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_97),
.A2(n_102),
.B1(n_138),
.B2(n_139),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_97),
.B(n_139),
.C(n_141),
.Y(n_317)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_111),
.C(n_113),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_106),
.A2(n_107),
.B1(n_111),
.B2(n_112),
.Y(n_148)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_113),
.B(n_148),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_124),
.C(n_128),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_114),
.A2(n_115),
.B1(n_151),
.B2(n_152),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_120),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_116),
.A2(n_117),
.B1(n_120),
.B2(n_121),
.Y(n_187)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_124),
.B(n_128),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_132),
.A2(n_304),
.B(n_305),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_133),
.B(n_144),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_133),
.B(n_144),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_143),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_141),
.Y(n_136)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g311 ( 
.A(n_140),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_142),
.Y(n_313)
);

AO21x1_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_167),
.B(n_302),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_147),
.B(n_149),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_147),
.B(n_149),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_153),
.C(n_154),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_150),
.B(n_153),
.Y(n_189)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_151),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_154),
.B(n_189),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_161),
.C(n_163),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_155),
.B(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_156),
.B(n_159),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_156),
.B(n_159),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_157),
.Y(n_227)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_160),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_161),
.B(n_163),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_162),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_164),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_190),
.B(n_301),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_188),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_169),
.B(n_188),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_172),
.C(n_187),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_170),
.B(n_187),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_172),
.B(n_288),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_180),
.C(n_183),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_SL g290 ( 
.A(n_173),
.B(n_291),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_177),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_174),
.B(n_177),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_180),
.B(n_183),
.Y(n_291)
);

AOI31xp33_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_285),
.A3(n_294),
.B(n_298),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_230),
.B(n_284),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_217),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_193),
.B(n_217),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_204),
.C(n_208),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_194),
.B(n_281),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_198),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_195),
.B(n_199),
.C(n_203),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_200),
.B1(n_201),
.B2(n_203),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_201),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_202),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_204),
.B(n_208),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_213),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_209),
.B(n_213),
.Y(n_241)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_210),
.Y(n_245)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_221),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_219),
.B(n_220),
.C(n_221),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_224),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_222),
.B(n_225),
.C(n_229),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_226),
.B1(n_228),
.B2(n_229),
.Y(n_224)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_225),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_226),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_231),
.A2(n_279),
.B(n_283),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_248),
.B(n_278),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_240),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_233),
.B(n_240),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_237),
.C(n_238),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_234),
.B(n_237),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_236),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_238),
.B(n_258),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_239),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_241),
.B(n_243),
.C(n_246),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_246),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_259),
.B(n_277),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_257),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_250),
.B(n_257),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_254),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_251),
.A2(n_252),
.B1(n_254),
.B2(n_255),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_260),
.A2(n_271),
.B(n_276),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_261),
.A2(n_266),
.B(n_270),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_264),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_267),
.B(n_268),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_269),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_275),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_272),
.B(n_275),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_280),
.B(n_282),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_280),
.B(n_282),
.Y(n_283)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_286),
.A2(n_299),
.B(n_300),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_287),
.B(n_289),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_287),
.B(n_289),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_292),
.C(n_293),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_290),
.B(n_297),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_292),
.B(n_293),
.Y(n_297)
);

OR2x2_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_295),
.B(n_296),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_307),
.B(n_308),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_307),
.B(n_308),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_317),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_310),
.A2(n_312),
.B1(n_315),
.B2(n_316),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_310),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_312),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_312),
.B(n_315),
.C(n_317),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_322),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_320),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_320),
.B(n_328),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g326 ( 
.A(n_322),
.Y(n_326)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_326),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_325),
.B(n_329),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_329),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_331),
.Y(n_330)
);


endmodule