module fake_jpeg_23334_n_267 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_267);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_267;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_96;

INVx2_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_19),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_37),
.A2(n_19),
.B1(n_31),
.B2(n_30),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_0),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_47),
.Y(n_55)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_39),
.Y(n_85)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_31),
.B(n_1),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_36),
.Y(n_54)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g44 ( 
.A(n_24),
.Y(n_44)
);

INVx3_ASAP7_75t_SL g82 ( 
.A(n_44),
.Y(n_82)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_30),
.B(n_36),
.Y(n_47)
);

INVx4_ASAP7_75t_SL g48 ( 
.A(n_35),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_48),
.B(n_49),
.Y(n_50)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_52),
.A2(n_57),
.B1(n_73),
.B2(n_83),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_23),
.Y(n_53)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_53),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_54),
.B(n_69),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_43),
.A2(n_17),
.B1(n_27),
.B2(n_35),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

CKINVDCx14_ASAP7_75t_R g114 ( 
.A(n_58),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_47),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_59),
.B(n_63),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_38),
.B(n_23),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_60),
.B(n_66),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_62),
.Y(n_98)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_28),
.Y(n_64)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_64),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_38),
.B(n_25),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_41),
.B(n_26),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_67),
.B(n_88),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_45),
.A2(n_26),
.B1(n_33),
.B2(n_29),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_68),
.A2(n_71),
.B1(n_89),
.B2(n_39),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_41),
.B(n_25),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_70),
.B(n_72),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_45),
.A2(n_20),
.B1(n_33),
.B2(n_29),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_74),
.Y(n_104)
);

CKINVDCx12_ASAP7_75t_R g75 ( 
.A(n_46),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_75),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_40),
.B(n_28),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_76),
.B(n_77),
.Y(n_108)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

CKINVDCx12_ASAP7_75t_R g78 ( 
.A(n_48),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_78),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_37),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_79),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_49),
.B(n_34),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_87),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_48),
.A2(n_17),
.B1(n_27),
.B2(n_35),
.Y(n_83)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_84),
.B(n_86),
.Y(n_109)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_49),
.B(n_34),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_39),
.A2(n_21),
.B1(n_22),
.B2(n_20),
.Y(n_89)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_91),
.B(n_94),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_54),
.B(n_22),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_93),
.B(n_106),
.Y(n_121)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_61),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_55),
.B(n_49),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_99),
.B(n_106),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_55),
.A2(n_39),
.B1(n_21),
.B2(n_34),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_100),
.A2(n_56),
.B1(n_84),
.B2(n_65),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_55),
.B(n_2),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_81),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_107),
.B(n_110),
.Y(n_137)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_58),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_111),
.B(n_118),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_89),
.B(n_2),
.Y(n_115)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_115),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_87),
.A2(n_3),
.B(n_4),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_116),
.B(n_7),
.C(n_8),
.Y(n_132)
);

A2O1A1Ixp33_ASAP7_75t_L g117 ( 
.A1(n_50),
.A2(n_4),
.B(n_7),
.C(n_8),
.Y(n_117)
);

OAI21xp33_ASAP7_75t_L g125 ( 
.A1(n_117),
.A2(n_7),
.B(n_8),
.Y(n_125)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_61),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_102),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_120),
.B(n_124),
.Y(n_152)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_101),
.B(n_82),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_122),
.B(n_134),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_123),
.B(n_125),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_109),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_99),
.B(n_82),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_126),
.B(n_132),
.C(n_114),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_90),
.B(n_80),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_130),
.A2(n_105),
.B(n_111),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_90),
.B(n_77),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_131),
.B(n_133),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_107),
.B(n_72),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_108),
.B(n_85),
.Y(n_134)
);

AOI32xp33_ASAP7_75t_L g135 ( 
.A1(n_97),
.A2(n_85),
.A3(n_70),
.B1(n_63),
.B2(n_80),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_135),
.B(n_138),
.Y(n_154)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_96),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_136),
.B(n_141),
.Y(n_157)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_98),
.Y(n_138)
);

INVx3_ASAP7_75t_SL g139 ( 
.A(n_102),
.Y(n_139)
);

HB1xp67_ASAP7_75t_L g164 ( 
.A(n_139),
.Y(n_164)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_94),
.Y(n_140)
);

INVx13_ASAP7_75t_L g156 ( 
.A(n_140),
.Y(n_156)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_96),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_108),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_142),
.Y(n_160)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_109),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_143),
.B(n_149),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_103),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_144),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_97),
.A2(n_73),
.B1(n_65),
.B2(n_51),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_145),
.A2(n_148),
.B1(n_98),
.B2(n_104),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_146),
.A2(n_115),
.B1(n_144),
.B2(n_149),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_117),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_147),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_110),
.A2(n_51),
.B1(n_56),
.B2(n_62),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_112),
.B(n_74),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_93),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_150),
.B(n_92),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_155),
.A2(n_161),
.B1(n_165),
.B2(n_169),
.Y(n_198)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_131),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_158),
.B(n_166),
.Y(n_187)
);

AO22x1_ASAP7_75t_L g163 ( 
.A1(n_146),
.A2(n_100),
.B1(n_116),
.B2(n_118),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_163),
.A2(n_172),
.B(n_113),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_137),
.A2(n_104),
.B1(n_98),
.B2(n_112),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_133),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_128),
.Y(n_167)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_167),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_127),
.A2(n_104),
.B1(n_112),
.B2(n_105),
.Y(n_169)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_140),
.Y(n_171)
);

INVx2_ASAP7_75t_SL g185 ( 
.A(n_171),
.Y(n_185)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_129),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_173),
.B(n_177),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_174),
.B(n_176),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_175),
.B(n_122),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_130),
.A2(n_92),
.B1(n_95),
.B2(n_119),
.Y(n_176)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_176),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_130),
.B(n_119),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_126),
.B(n_95),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_178),
.B(n_150),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_172),
.A2(n_123),
.B(n_136),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_179),
.B(n_189),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_178),
.B(n_143),
.C(n_148),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_183),
.B(n_186),
.C(n_190),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_157),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_184),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_175),
.B(n_132),
.C(n_145),
.Y(n_186)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_162),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_188),
.B(n_192),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_162),
.B(n_121),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_191),
.B(n_194),
.Y(n_202)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_168),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_158),
.B(n_120),
.Y(n_193)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_193),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_166),
.B(n_91),
.C(n_138),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_195),
.A2(n_167),
.B1(n_152),
.B2(n_160),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_174),
.B(n_13),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_196),
.B(n_199),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_168),
.B(n_9),
.Y(n_197)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_197),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_197),
.B(n_159),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_203),
.B(n_211),
.Y(n_217)
);

AOI322xp5_ASAP7_75t_L g204 ( 
.A1(n_179),
.A2(n_154),
.A3(n_177),
.B1(n_163),
.B2(n_153),
.C1(n_170),
.C2(n_155),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_204),
.B(n_212),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_198),
.A2(n_163),
.B1(n_165),
.B2(n_151),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_206),
.A2(n_208),
.B1(n_210),
.B2(n_180),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_181),
.A2(n_161),
.B1(n_151),
.B2(n_159),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_181),
.A2(n_192),
.B1(n_188),
.B2(n_198),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_193),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_189),
.B(n_169),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_214),
.A2(n_206),
.B1(n_205),
.B2(n_200),
.Y(n_223)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_187),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_216),
.B(n_173),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_218),
.A2(n_222),
.B1(n_223),
.B2(n_211),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_209),
.B(n_186),
.C(n_183),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_219),
.B(n_221),
.C(n_224),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g220 ( 
.A(n_216),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_220),
.B(n_228),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_209),
.B(n_195),
.C(n_180),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_200),
.A2(n_185),
.B1(n_171),
.B2(n_156),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_212),
.B(n_194),
.C(n_191),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_225),
.B(n_226),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_208),
.Y(n_226)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_202),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_201),
.B(n_182),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_229),
.B(n_230),
.Y(n_240)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_210),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_224),
.B(n_213),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_232),
.B(n_236),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_233),
.B(n_234),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_217),
.B(n_215),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_218),
.A2(n_202),
.B1(n_207),
.B2(n_213),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_226),
.A2(n_207),
.B(n_164),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_237),
.A2(n_238),
.B(n_11),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_221),
.A2(n_185),
.B1(n_156),
.B2(n_139),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_219),
.B(n_190),
.C(n_185),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_241),
.B(n_227),
.C(n_220),
.Y(n_245)
);

OA21x2_ASAP7_75t_SL g242 ( 
.A1(n_227),
.A2(n_13),
.B(n_14),
.Y(n_242)
);

FAx1_ASAP7_75t_SL g243 ( 
.A(n_242),
.B(n_14),
.CI(n_15),
.CON(n_243),
.SN(n_243)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_243),
.B(n_12),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_245),
.B(n_246),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_239),
.B(n_9),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_239),
.B(n_9),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_247),
.B(n_248),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_232),
.B(n_10),
.Y(n_248)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_249),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_250),
.A2(n_235),
.B(n_238),
.Y(n_253)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_253),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_244),
.A2(n_237),
.B(n_231),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_254),
.B(n_255),
.Y(n_258)
);

AOI21x1_ASAP7_75t_L g257 ( 
.A1(n_252),
.A2(n_240),
.B(n_244),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_257),
.A2(n_236),
.B1(n_255),
.B2(n_241),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_251),
.B(n_246),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_259),
.B(n_248),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_258),
.B(n_245),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_261),
.B(n_262),
.C(n_263),
.Y(n_265)
);

A2O1A1O1Ixp25_ASAP7_75t_L g264 ( 
.A1(n_262),
.A2(n_260),
.B(n_247),
.C(n_256),
.D(n_243),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_264),
.B(n_261),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_266),
.B(n_265),
.Y(n_267)
);


endmodule