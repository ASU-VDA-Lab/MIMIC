module real_jpeg_33073_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_216;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_470;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_17;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_487;
wire n_93;
wire n_493;
wire n_242;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_508;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_537;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_534;
wire n_358;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_519;
wire n_205;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_0),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_1),
.B(n_526),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_2),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_L g540 ( 
.A1(n_2),
.A2(n_528),
.B1(n_537),
.B2(n_541),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_3),
.A2(n_49),
.B1(n_53),
.B2(n_54),
.Y(n_48)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_3),
.A2(n_53),
.B1(n_126),
.B2(n_128),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g246 ( 
.A1(n_3),
.A2(n_53),
.B1(n_247),
.B2(n_248),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_3),
.A2(n_53),
.B1(n_340),
.B2(n_341),
.Y(n_339)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_4),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_4),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_4),
.Y(n_119)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_5),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_5),
.Y(n_164)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_6),
.Y(n_379)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_6),
.Y(n_388)
);

AO22x1_ASAP7_75t_SL g36 ( 
.A1(n_7),
.A2(n_37),
.B1(n_41),
.B2(n_43),
.Y(n_36)
);

INVx2_ASAP7_75t_SL g43 ( 
.A(n_7),
.Y(n_43)
);

OAI22x1_ASAP7_75t_SL g172 ( 
.A1(n_7),
.A2(n_43),
.B1(n_173),
.B2(n_175),
.Y(n_172)
);

AOI22x1_ASAP7_75t_SL g215 ( 
.A1(n_7),
.A2(n_43),
.B1(n_216),
.B2(n_218),
.Y(n_215)
);

NAND2xp33_ASAP7_75t_SL g299 ( 
.A(n_7),
.B(n_300),
.Y(n_299)
);

OAI32xp33_ASAP7_75t_L g372 ( 
.A1(n_7),
.A2(n_373),
.A3(n_380),
.B1(n_383),
.B2(n_389),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_7),
.B(n_132),
.Y(n_408)
);

OAI22x1_ASAP7_75t_R g84 ( 
.A1(n_8),
.A2(n_50),
.B1(n_85),
.B2(n_88),
.Y(n_84)
);

INVx2_ASAP7_75t_SL g88 ( 
.A(n_8),
.Y(n_88)
);

AO22x2_ASAP7_75t_SL g148 ( 
.A1(n_8),
.A2(n_88),
.B1(n_149),
.B2(n_152),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_8),
.A2(n_88),
.B1(n_185),
.B2(n_187),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_8),
.A2(n_88),
.B1(n_209),
.B2(n_210),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_9),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_9),
.Y(n_87)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_9),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_10),
.Y(n_97)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_10),
.Y(n_111)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_11),
.Y(n_67)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_11),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_12),
.Y(n_105)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_12),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_12),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_12),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_13),
.A2(n_225),
.B1(n_228),
.B2(n_229),
.Y(n_224)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_13),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_13),
.A2(n_152),
.B1(n_228),
.B2(n_284),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_13),
.A2(n_228),
.B1(n_305),
.B2(n_307),
.Y(n_304)
);

OAI22xp33_ASAP7_75t_SL g400 ( 
.A1(n_13),
.A2(n_228),
.B1(n_401),
.B2(n_404),
.Y(n_400)
);

OAI21xp33_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_511),
.B(n_535),
.Y(n_14)
);

AOI211xp5_ASAP7_75t_L g535 ( 
.A1(n_15),
.A2(n_536),
.B(n_539),
.C(n_540),
.Y(n_535)
);

AOI21xp5_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_263),
.B(n_508),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_239),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_197),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_18),
.B(n_197),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_120),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_19),
.B(n_121),
.C(n_180),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_44),
.B(n_89),
.Y(n_19)
);

INVx1_ASAP7_75t_SL g45 ( 
.A(n_20),
.Y(n_45)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_20),
.B(n_90),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_20),
.B(n_290),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_20),
.A2(n_45),
.B1(n_290),
.B2(n_364),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_20),
.A2(n_45),
.B1(n_486),
.B2(n_487),
.Y(n_485)
);

AO21x2_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_25),
.B(n_35),
.Y(n_20)
);

CKINVDCx5p33_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g458 ( 
.A1(n_25),
.A2(n_273),
.B(n_339),
.Y(n_458)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_26),
.B(n_208),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_26),
.B(n_36),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_26),
.B(n_400),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_31),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_30),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_30),
.Y(n_338)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_31),
.Y(n_340)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g422 ( 
.A(n_32),
.Y(n_422)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_34),
.Y(n_79)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_36),
.B(n_203),
.Y(n_202)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_40),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_40),
.Y(n_403)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_42),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_43),
.A2(n_114),
.B(n_115),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_43),
.B(n_116),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_43),
.B(n_190),
.Y(n_277)
);

AOI32xp33_ASAP7_75t_L g290 ( 
.A1(n_43),
.A2(n_291),
.A3(n_294),
.B1(n_298),
.B2(n_299),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_43),
.B(n_384),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_R g413 ( 
.A(n_43),
.B(n_73),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_43),
.B(n_275),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_44),
.B(n_238),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_46),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g487 ( 
.A(n_46),
.Y(n_487)
);

OAI21xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_57),
.B(n_82),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_48),
.B(n_83),
.Y(n_200)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_52),
.Y(n_56)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_52),
.Y(n_306)
);

INVx4_ASAP7_75t_SL g54 ( 
.A(n_55),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_58),
.B(n_84),
.Y(n_178)
);

OA21x2_ASAP7_75t_L g196 ( 
.A1(n_58),
.A2(n_83),
.B(n_172),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_58),
.B(n_304),
.Y(n_303)
);

NAND2x1_ASAP7_75t_L g396 ( 
.A(n_58),
.B(n_172),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_73),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_63),
.B1(n_68),
.B2(n_70),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_61),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_62),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_62),
.Y(n_293)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_67),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_69),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g393 ( 
.A(n_70),
.Y(n_393)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

OA22x2_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_76),
.B1(n_78),
.B2(n_80),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_75),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_79),
.Y(n_211)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_82),
.B(n_303),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_82),
.B(n_396),
.Y(n_459)
);

NAND2x1p5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_84),
.Y(n_82)
);

NAND2xp33_ASAP7_75t_SL g171 ( 
.A(n_83),
.B(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_83),
.B(n_304),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_87),
.Y(n_391)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_91),
.A2(n_112),
.B(n_113),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_91),
.B(n_113),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_91),
.B(n_224),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_91),
.B(n_184),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g521 ( 
.A(n_91),
.Y(n_521)
);

NOR2x1p5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_102),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_95),
.B1(n_98),
.B2(n_101),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_97),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_97),
.Y(n_329)
);

INVx3_ASAP7_75t_SL g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g250 ( 
.A(n_99),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_100),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_100),
.Y(n_227)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_100),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_100),
.Y(n_324)
);

AO22x2_ASAP7_75t_L g102 ( 
.A1(n_101),
.A2(n_103),
.B1(n_106),
.B2(n_109),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g320 ( 
.A(n_101),
.Y(n_320)
);

HB1xp67_ASAP7_75t_L g112 ( 
.A(n_102),
.Y(n_112)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_102),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_102),
.B(n_224),
.Y(n_347)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g220 ( 
.A(n_105),
.Y(n_220)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_107),
.Y(n_127)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_107),
.Y(n_160)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_107),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g131 ( 
.A(n_108),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_108),
.Y(n_155)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_112),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_113),
.B(n_189),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_115),
.Y(n_334)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_117),
.Y(n_186)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_117),
.Y(n_188)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_122),
.B1(n_179),
.B2(n_180),
.Y(n_120)
);

INVxp67_ASAP7_75t_SL g121 ( 
.A(n_122),
.Y(n_121)
);

OAI21x1_ASAP7_75t_SL g234 ( 
.A1(n_122),
.A2(n_123),
.B(n_170),
.Y(n_234)
);

NAND2x1p5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_170),
.Y(n_122)
);

AOI21x1_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_132),
.B(n_146),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_125),
.A2(n_157),
.B(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_132),
.B(n_259),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_132),
.B(n_283),
.Y(n_350)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_133),
.Y(n_195)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

AO21x2_ASAP7_75t_L g157 ( 
.A1(n_134),
.A2(n_158),
.B(n_165),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_138),
.B1(n_142),
.B2(n_145),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_137),
.Y(n_144)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_140),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_141),
.Y(n_169)
);

INVx2_ASAP7_75t_SL g142 ( 
.A(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

NOR2x1_ASAP7_75t_L g256 ( 
.A(n_146),
.B(n_257),
.Y(n_256)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_147),
.B(n_350),
.Y(n_349)
);

NAND2x1_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_156),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_148),
.B(n_195),
.Y(n_194)
);

BUFx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_150),
.Y(n_166)
);

INVx5_ASAP7_75t_L g317 ( 
.A(n_150),
.Y(n_317)
);

INVx8_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_151),
.Y(n_217)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_155),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_156),
.B(n_283),
.Y(n_282)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

NOR2x1_ASAP7_75t_L g214 ( 
.A(n_157),
.B(n_215),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g454 ( 
.A1(n_157),
.A2(n_215),
.B(n_455),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_159),
.B(n_161),
.Y(n_158)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVxp33_ASAP7_75t_L g298 ( 
.A(n_165),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_167),
.Y(n_165)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_178),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_171),
.B(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_SL g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_178),
.A2(n_200),
.B(n_201),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_178),
.B(n_357),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_178),
.B(n_200),
.Y(n_451)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

XNOR2x1_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_191),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_181),
.B(n_192),
.C(n_196),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_181),
.A2(n_244),
.B1(n_261),
.B2(n_262),
.Y(n_243)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_181),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_182),
.B(n_347),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_183),
.B(n_223),
.Y(n_447)
);

OAI21xp5_ASAP7_75t_L g520 ( 
.A1(n_183),
.A2(n_246),
.B(n_521),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_189),
.Y(n_183)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_185),
.Y(n_247)
);

INVx3_ASAP7_75t_SL g185 ( 
.A(n_186),
.Y(n_185)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_196),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_193),
.B(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

NOR2x1p5_ASAP7_75t_SL g213 ( 
.A(n_194),
.B(n_214),
.Y(n_213)
);

INVxp67_ASAP7_75t_SL g455 ( 
.A(n_195),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_196),
.A2(n_255),
.B1(n_256),
.B2(n_260),
.Y(n_254)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_196),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_196),
.A2(n_260),
.B1(n_349),
.B2(n_351),
.Y(n_348)
);

MAJx2_ASAP7_75t_L g465 ( 
.A(n_196),
.B(n_346),
.C(n_349),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_196),
.B(n_256),
.C(n_519),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_233),
.C(n_235),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_198),
.B(n_493),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_212),
.C(n_221),
.Y(n_198)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_199),
.Y(n_489)
);

XOR2x2_ASAP7_75t_SL g450 ( 
.A(n_201),
.B(n_451),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_207),
.Y(n_201)
);

AND2x4_ASAP7_75t_SL g398 ( 
.A(n_202),
.B(n_399),
.Y(n_398)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx2_ASAP7_75t_SL g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_206),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_L g335 ( 
.A1(n_207),
.A2(n_336),
.B(n_339),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_207),
.B(n_417),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_208),
.B(n_274),
.Y(n_273)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVxp33_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_213),
.B(n_222),
.Y(n_490)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_214),
.Y(n_361)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_215),
.Y(n_259)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_232),
.Y(n_222)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_232),
.B(n_252),
.Y(n_516)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_234),
.B(n_237),
.Y(n_493)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g508 ( 
.A1(n_239),
.A2(n_509),
.B(n_510),
.Y(n_508)
);

NOR2xp67_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_240),
.B(n_241),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

INVxp67_ASAP7_75t_SL g534 ( 
.A(n_242),
.Y(n_534)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_244),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g533 ( 
.A(n_244),
.Y(n_533)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_254),
.Y(n_244)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_245),
.Y(n_519)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_246),
.A2(n_251),
.B(n_252),
.Y(n_245)
);

INVx4_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx11_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_253),
.B(n_347),
.Y(n_456)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_258),
.B(n_282),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_261),
.B(n_533),
.C(n_534),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_499),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_265),
.A2(n_439),
.B(n_498),
.Y(n_264)
);

AO21x1_ASAP7_75t_L g265 ( 
.A1(n_266),
.A2(n_352),
.B(n_438),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_309),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_267),
.B(n_309),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_288),
.C(n_302),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_268),
.B(n_366),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_280),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_277),
.B1(n_278),
.B2(n_279),
.Y(n_269)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_270),
.Y(n_279)
);

NOR2xp67_ASAP7_75t_SL g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g420 ( 
.A(n_271),
.Y(n_420)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_273),
.B(n_399),
.Y(n_414)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_277),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_277),
.B(n_279),
.C(n_281),
.Y(n_311)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx8_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_289),
.B(n_302),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_290),
.Y(n_364)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_293),
.Y(n_301)
);

INVx5_ASAP7_75t_L g308 ( 
.A(n_293),
.Y(n_308)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVxp67_ASAP7_75t_SL g305 ( 
.A(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_306),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_345),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_311),
.A2(n_312),
.B1(n_313),
.B2(n_344),
.Y(n_310)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_311),
.Y(n_344)
);

HB1xp67_ASAP7_75t_L g471 ( 
.A(n_311),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_312),
.B(n_469),
.C(n_470),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_312),
.B(n_469),
.C(n_470),
.Y(n_503)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_335),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_314),
.B(n_335),
.Y(n_448)
);

OAI31xp33_ASAP7_75t_L g314 ( 
.A1(n_315),
.A2(n_318),
.A3(n_321),
.B(n_325),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_326),
.A2(n_330),
.B(n_334),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_SL g336 ( 
.A(n_337),
.Y(n_336)
);

BUFx2_ASAP7_75t_R g337 ( 
.A(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_345),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_348),
.Y(n_345)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_349),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_350),
.B(n_361),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_L g352 ( 
.A1(n_353),
.A2(n_367),
.B(n_437),
.Y(n_352)
);

NOR2x1_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_365),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_354),
.B(n_365),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_358),
.C(n_362),
.Y(n_354)
);

OAI22xp33_ASAP7_75t_L g435 ( 
.A1(n_355),
.A2(n_356),
.B1(n_359),
.B2(n_360),
.Y(n_435)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_357),
.B(n_396),
.Y(n_395)
);

HB1xp67_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVxp67_ASAP7_75t_SL g362 ( 
.A(n_363),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_363),
.B(n_435),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_L g367 ( 
.A1(n_368),
.A2(n_430),
.B(n_436),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_L g368 ( 
.A1(n_369),
.A2(n_410),
.B(n_429),
.Y(n_368)
);

NOR2x1_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_397),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_370),
.B(n_397),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_394),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_371),
.A2(n_372),
.B1(n_394),
.B2(n_395),
.Y(n_427)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

BUFx4f_ASAP7_75t_SL g381 ( 
.A(n_382),
.Y(n_381)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_392),
.Y(n_389)
);

BUFx2_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_407),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_398),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_400),
.B(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx4_ASAP7_75t_L g406 ( 
.A(n_403),
.Y(n_406)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_409),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_408),
.B(n_432),
.C(n_433),
.Y(n_431)
);

HB1xp67_ASAP7_75t_L g433 ( 
.A(n_409),
.Y(n_433)
);

AOI21x1_ASAP7_75t_L g410 ( 
.A1(n_411),
.A2(n_425),
.B(n_428),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_SL g411 ( 
.A1(n_412),
.A2(n_415),
.B(n_424),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_413),
.B(n_414),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_413),
.B(n_414),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_416),
.B(n_421),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_420),
.Y(n_416)
);

BUFx2_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_422),
.B(n_423),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_427),
.Y(n_425)
);

NOR2x1_ASAP7_75t_L g428 ( 
.A(n_426),
.B(n_427),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_431),
.B(n_434),
.Y(n_430)
);

NOR2xp67_ASAP7_75t_L g436 ( 
.A(n_431),
.B(n_434),
.Y(n_436)
);

NOR3xp33_ASAP7_75t_L g439 ( 
.A(n_440),
.B(n_474),
.C(n_491),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_441),
.B(n_467),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_441),
.B(n_502),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_460),
.Y(n_441)
);

OR2x2_ASAP7_75t_L g505 ( 
.A(n_442),
.B(n_460),
.Y(n_505)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_443),
.B(n_449),
.Y(n_442)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_443),
.Y(n_476)
);

MAJx2_ASAP7_75t_L g443 ( 
.A(n_444),
.B(n_446),
.C(n_448),
.Y(n_443)
);

INVxp67_ASAP7_75t_SL g444 ( 
.A(n_445),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_L g462 ( 
.A1(n_445),
.A2(n_446),
.B(n_463),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_445),
.B(n_464),
.Y(n_463)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_447),
.Y(n_464)
);

XNOR2x1_ASAP7_75t_L g461 ( 
.A(n_448),
.B(n_462),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_452),
.Y(n_449)
);

INVxp33_ASAP7_75t_SL g477 ( 
.A(n_450),
.Y(n_477)
);

HB1xp67_ASAP7_75t_L g478 ( 
.A(n_452),
.Y(n_478)
);

XNOR2x1_ASAP7_75t_L g452 ( 
.A(n_453),
.B(n_457),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_454),
.B(n_456),
.Y(n_453)
);

HB1xp67_ASAP7_75t_L g483 ( 
.A(n_454),
.Y(n_483)
);

HB1xp67_ASAP7_75t_L g482 ( 
.A(n_456),
.Y(n_482)
);

HB1xp67_ASAP7_75t_L g481 ( 
.A(n_457),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_458),
.B(n_459),
.Y(n_457)
);

XOR2x2_ASAP7_75t_L g466 ( 
.A(n_458),
.B(n_459),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_465),
.C(n_466),
.Y(n_460)
);

XNOR2x1_ASAP7_75t_L g472 ( 
.A(n_461),
.B(n_473),
.Y(n_472)
);

XOR2x1_ASAP7_75t_SL g473 ( 
.A(n_465),
.B(n_466),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_468),
.B(n_472),
.Y(n_467)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_472),
.B(n_503),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_474),
.B(n_504),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_475),
.B(n_479),
.Y(n_474)
);

OR2x2_ASAP7_75t_L g504 ( 
.A(n_475),
.B(n_479),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_476),
.B(n_477),
.C(n_478),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_480),
.B(n_484),
.Y(n_479)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_480),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_481),
.B(n_482),
.C(n_483),
.Y(n_480)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_483),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_L g530 ( 
.A1(n_483),
.A2(n_520),
.B1(n_522),
.B2(n_531),
.Y(n_530)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_485),
.B(n_488),
.Y(n_484)
);

INVxp67_ASAP7_75t_SL g496 ( 
.A(n_485),
.Y(n_496)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

INVxp33_ASAP7_75t_L g495 ( 
.A(n_488),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_489),
.B(n_490),
.Y(n_488)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_491),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_492),
.B(n_494),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_492),
.B(n_494),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_495),
.B(n_496),
.C(n_497),
.Y(n_494)
);

NAND3xp33_ASAP7_75t_L g499 ( 
.A(n_500),
.B(n_506),
.C(n_507),
.Y(n_499)
);

NAND3xp33_ASAP7_75t_L g500 ( 
.A(n_501),
.B(n_504),
.C(n_505),
.Y(n_500)
);

OR2x2_ASAP7_75t_L g511 ( 
.A(n_512),
.B(n_527),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_SL g539 ( 
.A(n_512),
.B(n_538),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_513),
.B(n_525),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

NAND3xp33_ASAP7_75t_L g537 ( 
.A(n_514),
.B(n_525),
.C(n_538),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_515),
.B(n_523),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_516),
.B(n_517),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_516),
.B(n_517),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_518),
.B(n_520),
.C(n_522),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_L g529 ( 
.A(n_518),
.B(n_530),
.Y(n_529)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_520),
.Y(n_531)
);

INVxp67_ASAP7_75t_L g523 ( 
.A(n_524),
.Y(n_523)
);

INVxp67_ASAP7_75t_L g541 ( 
.A(n_525),
.Y(n_541)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_528),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_529),
.B(n_532),
.Y(n_528)
);

OR2x2_ASAP7_75t_L g538 ( 
.A(n_529),
.B(n_532),
.Y(n_538)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_537),
.Y(n_536)
);


endmodule