module fake_jpeg_15003_n_44 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_44);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_44;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_25;
wire n_17;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_32;
wire n_15;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_12),
.B(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx4f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_15),
.B(n_0),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_22),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_15),
.B(n_0),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_19),
.B(n_1),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_23),
.B(n_4),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g24 ( 
.A1(n_20),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g29 ( 
.A1(n_24),
.A2(n_25),
.B(n_20),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_SL g25 ( 
.A1(n_19),
.A2(n_4),
.B(n_5),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_24),
.B(n_17),
.C(n_20),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_27),
.C(n_31),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_29),
.A2(n_16),
.B1(n_7),
.B2(n_8),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_18),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_30),
.Y(n_33)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

HB1xp67_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_17),
.C(n_16),
.Y(n_35)
);

XOR2xp5_ASAP7_75t_L g39 ( 
.A(n_35),
.B(n_17),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g37 ( 
.A1(n_36),
.A2(n_6),
.B(n_7),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_SL g41 ( 
.A1(n_37),
.A2(n_33),
.B(n_8),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_39),
.B(n_34),
.Y(n_40)
);

AO21x1_ASAP7_75t_L g42 ( 
.A1(n_40),
.A2(n_41),
.B(n_32),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_42),
.B(n_38),
.Y(n_43)
);

AOI31xp67_ASAP7_75t_SL g44 ( 
.A1(n_43),
.A2(n_6),
.A3(n_11),
.B(n_10),
.Y(n_44)
);


endmodule