module real_jpeg_4813_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_216;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_215;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx5_ASAP7_75t_L g173 ( 
.A(n_0),
.Y(n_173)
);

INVx8_ASAP7_75t_L g179 ( 
.A(n_0),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_0),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_0),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_0),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_1),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_1),
.Y(n_59)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_1),
.Y(n_148)
);

BUFx5_ASAP7_75t_L g237 ( 
.A(n_1),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_1),
.Y(n_239)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_1),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_2),
.A2(n_236),
.B1(n_238),
.B2(n_239),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_2),
.Y(n_238)
);

OAI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_2),
.A2(n_238),
.B1(n_270),
.B2(n_273),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g337 ( 
.A1(n_2),
.A2(n_238),
.B1(n_338),
.B2(n_340),
.Y(n_337)
);

AOI22xp33_ASAP7_75t_L g424 ( 
.A1(n_2),
.A2(n_139),
.B1(n_238),
.B2(n_425),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_3),
.Y(n_504)
);

AOI22xp33_ASAP7_75t_L g290 ( 
.A1(n_4),
.A2(n_291),
.B1(n_293),
.B2(n_294),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_4),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_4),
.A2(n_293),
.B1(n_312),
.B2(n_313),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g372 ( 
.A1(n_4),
.A2(n_122),
.B1(n_293),
.B2(n_373),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_4),
.A2(n_51),
.B1(n_293),
.B2(n_451),
.Y(n_450)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g400 ( 
.A(n_5),
.Y(n_400)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_6),
.Y(n_500)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_7),
.A2(n_122),
.B1(n_126),
.B2(n_128),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_7),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_7),
.A2(n_128),
.B1(n_157),
.B2(n_158),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_7),
.A2(n_128),
.B1(n_216),
.B2(n_220),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_8),
.A2(n_194),
.B1(n_195),
.B2(n_196),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_8),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_8),
.A2(n_88),
.B1(n_194),
.B2(n_258),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_L g278 ( 
.A1(n_8),
.A2(n_194),
.B1(n_279),
.B2(n_283),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_8),
.A2(n_126),
.B1(n_194),
.B2(n_348),
.Y(n_347)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_9),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_9),
.Y(n_75)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_9),
.Y(n_80)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_10),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_11),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_11),
.Y(n_85)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_11),
.Y(n_177)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_12),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_13),
.A2(n_252),
.B1(n_253),
.B2(n_255),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_13),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_13),
.B(n_75),
.C(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_13),
.B(n_107),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_13),
.B(n_173),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_13),
.B(n_160),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_13),
.B(n_127),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_14),
.A2(n_56),
.B1(n_59),
.B2(n_60),
.Y(n_55)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_14),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_14),
.A2(n_60),
.B1(n_166),
.B2(n_167),
.Y(n_165)
);

OAI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_14),
.A2(n_60),
.B1(n_227),
.B2(n_228),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g381 ( 
.A1(n_14),
.A2(n_60),
.B1(n_304),
.B2(n_382),
.Y(n_381)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_15),
.A2(n_87),
.B1(n_89),
.B2(n_91),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_15),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_15),
.A2(n_91),
.B1(n_137),
.B2(n_139),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_15),
.A2(n_91),
.B1(n_181),
.B2(n_182),
.Y(n_180)
);

OAI22xp33_ASAP7_75t_L g49 ( 
.A1(n_16),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_16),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_16),
.A2(n_50),
.B1(n_231),
.B2(n_233),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_L g352 ( 
.A1(n_16),
.A2(n_50),
.B1(n_271),
.B2(n_312),
.Y(n_352)
);

AOI22xp33_ASAP7_75t_SL g429 ( 
.A1(n_16),
.A2(n_50),
.B1(n_188),
.B2(n_430),
.Y(n_429)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_18),
.A2(n_115),
.B1(n_119),
.B2(n_120),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_18),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_18),
.A2(n_51),
.B1(n_119),
.B2(n_144),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_18),
.A2(n_119),
.B1(n_186),
.B2(n_188),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g411 ( 
.A1(n_18),
.A2(n_81),
.B1(n_119),
.B2(n_183),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_499),
.B(n_501),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_200),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_199),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_150),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_24),
.B(n_150),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_129),
.B2(n_130),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_61),
.C(n_92),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_27),
.A2(n_131),
.B1(n_132),
.B2(n_149),
.Y(n_130)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_27),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_27),
.A2(n_149),
.B1(n_152),
.B2(n_153),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_28),
.A2(n_48),
.B1(n_53),
.B2(n_55),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_28),
.A2(n_53),
.B1(n_55),
.B2(n_143),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_28),
.A2(n_235),
.B(n_240),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_28),
.A2(n_53),
.B1(n_235),
.B2(n_450),
.Y(n_449)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_29),
.B(n_193),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g417 ( 
.A1(n_29),
.A2(n_418),
.B(n_421),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_39),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_33),
.B1(n_35),
.B2(n_36),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_32),
.Y(n_397)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_35),
.Y(n_195)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_41),
.B1(n_45),
.B2(n_47),
.Y(n_39)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g396 ( 
.A(n_42),
.Y(n_396)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g166 ( 
.A(n_43),
.Y(n_166)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_43),
.Y(n_375)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_44),
.Y(n_118)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_44),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_44),
.Y(n_127)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_44),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_46),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_46),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_46),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_49),
.B(n_54),
.Y(n_191)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_51),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_51),
.B(n_255),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_53),
.B(n_255),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_L g468 ( 
.A1(n_53),
.A2(n_192),
.B(n_450),
.Y(n_468)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_54),
.B(n_193),
.Y(n_240)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_61),
.A2(n_62),
.B1(n_134),
.B2(n_135),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_61),
.A2(n_62),
.B1(n_92),
.B2(n_93),
.Y(n_152)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_SL g62 ( 
.A1(n_63),
.A2(n_77),
.B(n_86),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_63),
.A2(n_251),
.B(n_256),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_63),
.A2(n_77),
.B1(n_290),
.B2(n_337),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g368 ( 
.A1(n_63),
.A2(n_256),
.B(n_337),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_63),
.A2(n_77),
.B1(n_429),
.B2(n_444),
.Y(n_443)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_64),
.A2(n_156),
.B1(n_160),
.B2(n_161),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_64),
.A2(n_156),
.B1(n_160),
.B2(n_185),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_64),
.A2(n_160),
.B1(n_185),
.B2(n_226),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_64),
.B(n_257),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_77),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_71),
.B1(n_74),
.B2(n_76),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

INVx5_ASAP7_75t_L g340 ( 
.A(n_68),
.Y(n_340)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_69),
.Y(n_157)
);

INVx5_ASAP7_75t_L g187 ( 
.A(n_69),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_69),
.Y(n_296)
);

INVx6_ASAP7_75t_L g431 ( 
.A(n_69),
.Y(n_431)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_70),
.Y(n_110)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_70),
.Y(n_159)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_70),
.Y(n_254)
);

BUFx3_ASAP7_75t_L g260 ( 
.A(n_70),
.Y(n_260)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

AOI22x1_ASAP7_75t_L g77 ( 
.A1(n_74),
.A2(n_78),
.B1(n_81),
.B2(n_84),
.Y(n_77)
);

INVx4_ASAP7_75t_SL g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_77),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_77),
.A2(n_290),
.B(n_297),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g428 ( 
.A1(n_77),
.A2(n_297),
.B(n_429),
.Y(n_428)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_83),
.Y(n_219)
);

BUFx5_ASAP7_75t_L g272 ( 
.A(n_83),
.Y(n_272)
);

BUFx8_ASAP7_75t_L g306 ( 
.A(n_83),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_85),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_85),
.Y(n_183)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_85),
.Y(n_266)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_85),
.Y(n_286)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_86),
.Y(n_161)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

AO22x2_ASAP7_75t_L g107 ( 
.A1(n_88),
.A2(n_108),
.B1(n_109),
.B2(n_111),
.Y(n_107)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_90),
.Y(n_227)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_94),
.A2(n_113),
.B1(n_124),
.B2(n_125),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_94),
.A2(n_124),
.B1(n_125),
.B2(n_136),
.Y(n_135)
);

INVx2_ASAP7_75t_SL g163 ( 
.A(n_94),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_94),
.A2(n_124),
.B1(n_165),
.B2(n_230),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_94),
.A2(n_124),
.B1(n_372),
.B2(n_424),
.Y(n_423)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_107),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_100),
.B1(n_102),
.B2(n_105),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_98),
.Y(n_356)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_99),
.Y(n_104)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_99),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx5_ASAP7_75t_L g427 ( 
.A(n_101),
.Y(n_427)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_104),
.Y(n_112)
);

INVx4_ASAP7_75t_L g361 ( 
.A(n_104),
.Y(n_361)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_SL g124 ( 
.A(n_107),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_107),
.A2(n_114),
.B1(n_163),
.B2(n_164),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_107),
.A2(n_163),
.B1(n_377),
.B2(n_455),
.Y(n_454)
);

INVx4_ASAP7_75t_L g263 ( 
.A(n_109),
.Y(n_263)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_109),
.Y(n_292)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g339 ( 
.A(n_110),
.Y(n_339)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

OAI21xp33_ASAP7_75t_SL g343 ( 
.A1(n_115),
.A2(n_255),
.B(n_344),
.Y(n_343)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_118),
.Y(n_141)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_118),
.Y(n_167)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_118),
.Y(n_232)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_124),
.B(n_347),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_124),
.A2(n_372),
.B(n_376),
.Y(n_371)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_SL g132 ( 
.A(n_133),
.B(n_142),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_137),
.Y(n_233)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_139),
.Y(n_348)
);

AOI32xp33_ASAP7_75t_L g353 ( 
.A1(n_139),
.A2(n_338),
.A3(n_345),
.B1(n_354),
.B2(n_357),
.Y(n_353)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_148),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_154),
.C(n_168),
.Y(n_150)
);

FAx1_ASAP7_75t_SL g202 ( 
.A(n_151),
.B(n_154),
.CI(n_168),
.CON(n_202),
.SN(n_202)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_152),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_154),
.A2(n_210),
.B(n_211),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_162),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_155),
.Y(n_211)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_160),
.B(n_257),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_162),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_163),
.A2(n_343),
.B(n_346),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_163),
.B(n_377),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_163),
.A2(n_346),
.B(n_471),
.Y(n_470)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_170),
.B(n_190),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_169),
.B(n_206),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_184),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_170),
.A2(n_190),
.B1(n_207),
.B2(n_208),
.Y(n_206)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_170),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_170),
.A2(n_184),
.B1(n_208),
.B2(n_440),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_171),
.A2(n_178),
.B(n_180),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_171),
.A2(n_180),
.B1(n_215),
.B2(n_223),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_171),
.A2(n_269),
.B(n_276),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_171),
.A2(n_255),
.B(n_276),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_171),
.A2(n_407),
.B1(n_408),
.B2(n_410),
.Y(n_406)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_172),
.B(n_278),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_172),
.A2(n_323),
.B1(n_324),
.B2(n_325),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_172),
.A2(n_352),
.B1(n_381),
.B2(n_383),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_172),
.A2(n_411),
.B1(n_446),
.B2(n_447),
.Y(n_445)
);

OR2x2_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_174),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_175),
.Y(n_174)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_177),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_177),
.Y(n_282)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_178),
.Y(n_277)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g440 ( 
.A(n_184),
.Y(n_440)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_186),
.Y(n_252)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx5_ASAP7_75t_L g189 ( 
.A(n_187),
.Y(n_189)
);

BUFx2_ASAP7_75t_L g228 ( 
.A(n_187),
.Y(n_228)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_190),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_192),
.Y(n_190)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_241),
.B(n_498),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_202),
.B(n_203),
.Y(n_498)
);

BUFx24_ASAP7_75t_SL g505 ( 
.A(n_202),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_209),
.C(n_212),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_204),
.A2(n_205),
.B1(n_209),
.B2(n_458),
.Y(n_457)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_209),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_212),
.B(n_457),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_229),
.C(n_234),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_213),
.B(n_438),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_225),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_214),
.B(n_225),
.Y(n_465)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_215),
.Y(n_446)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_219),
.Y(n_275)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_220),
.Y(n_312)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx8_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g326 ( 
.A(n_223),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g350 ( 
.A1(n_223),
.A2(n_318),
.B(n_351),
.Y(n_350)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_223),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_224),
.Y(n_409)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_226),
.Y(n_444)
);

NAND2xp33_ASAP7_75t_SL g357 ( 
.A(n_227),
.B(n_358),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_229),
.B(n_234),
.Y(n_438)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_230),
.Y(n_455)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

OAI32xp33_ASAP7_75t_L g393 ( 
.A1(n_236),
.A2(n_394),
.A3(n_397),
.B1(n_398),
.B2(n_404),
.Y(n_393)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx8_ASAP7_75t_L g453 ( 
.A(n_239),
.Y(n_453)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_240),
.Y(n_421)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

OAI311xp33_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_434),
.A3(n_474),
.B1(n_492),
.C1(n_497),
.Y(n_243)
);

AOI21x1_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_387),
.B(n_433),
.Y(n_244)
);

AO21x1_ASAP7_75t_SL g245 ( 
.A1(n_246),
.A2(n_363),
.B(n_386),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_247),
.A2(n_331),
.B(n_362),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_300),
.B(n_330),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_267),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_249),
.B(n_267),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_250),
.B(n_261),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_250),
.A2(n_261),
.B1(n_262),
.B2(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_250),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

OAI21xp33_ASAP7_75t_SL g418 ( 
.A1(n_255),
.A2(n_404),
.B(n_419),
.Y(n_418)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_259),
.Y(n_258)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_262),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_287),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_268),
.B(n_288),
.C(n_299),
.Y(n_332)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_269),
.Y(n_324)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_271),
.Y(n_270)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_280),
.Y(n_382)
);

INVx6_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_282),
.Y(n_314)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx6_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_288),
.A2(n_289),
.B1(n_298),
.B2(n_299),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx4_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_301),
.A2(n_321),
.B(n_329),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_302),
.A2(n_309),
.B(n_320),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_308),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_307),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx8_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_310),
.B(n_319),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_310),
.B(n_319),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_311),
.A2(n_315),
.B(n_318),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_311),
.Y(n_323)
);

INVx4_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx4_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx4_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_327),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_322),
.B(n_327),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_326),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_333),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_332),
.B(n_333),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_349),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_335),
.A2(n_336),
.B1(n_341),
.B2(n_342),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_336),
.B(n_341),
.C(n_349),
.Y(n_364)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVxp33_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_347),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_353),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_350),
.B(n_353),
.Y(n_369)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

CKINVDCx14_ASAP7_75t_R g354 ( 
.A(n_355),
.Y(n_354)
);

BUFx3_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx4_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx8_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_365),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_SL g386 ( 
.A(n_364),
.B(n_365),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_366),
.A2(n_367),
.B1(n_370),
.B2(n_385),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_SL g367 ( 
.A(n_368),
.B(n_369),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_368),
.B(n_369),
.C(n_385),
.Y(n_388)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_370),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_SL g370 ( 
.A(n_371),
.B(n_378),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_371),
.B(n_379),
.C(n_380),
.Y(n_412)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_380),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_381),
.Y(n_407)
);

INVx3_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_389),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_SL g433 ( 
.A(n_388),
.B(n_389),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_415),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_391),
.A2(n_412),
.B1(n_413),
.B2(n_414),
.Y(n_390)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_391),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_392),
.A2(n_393),
.B1(n_405),
.B2(n_406),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_393),
.B(n_405),
.Y(n_469)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx3_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_401),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx3_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

BUFx12f_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_412),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_412),
.B(n_413),
.C(n_415),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_416),
.A2(n_417),
.B1(n_422),
.B2(n_432),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_416),
.B(n_423),
.C(n_428),
.Y(n_483)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_422),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_SL g422 ( 
.A(n_423),
.B(n_428),
.Y(n_422)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_424),
.Y(n_471)
);

INVx3_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

INVx6_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

INVx8_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

NAND2xp33_ASAP7_75t_SL g434 ( 
.A(n_435),
.B(n_459),
.Y(n_434)
);

A2O1A1Ixp33_ASAP7_75t_SL g492 ( 
.A1(n_435),
.A2(n_459),
.B(n_493),
.C(n_496),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_436),
.B(n_456),
.Y(n_435)
);

OR2x2_ASAP7_75t_L g497 ( 
.A(n_436),
.B(n_456),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_437),
.B(n_439),
.C(n_441),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_437),
.B(n_439),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_441),
.B(n_473),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_448),
.C(n_454),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_442),
.B(n_463),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_443),
.B(n_445),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_443),
.B(n_445),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_448),
.A2(n_449),
.B1(n_454),
.B2(n_464),
.Y(n_463)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

INVx3_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_454),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_460),
.B(n_472),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_460),
.B(n_472),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_465),
.C(n_466),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_461),
.A2(n_462),
.B1(n_465),
.B2(n_486),
.Y(n_485)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_465),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_466),
.B(n_485),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_467),
.B(n_469),
.C(n_470),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_467),
.A2(n_468),
.B1(n_470),
.B2(n_480),
.Y(n_479)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_469),
.B(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_470),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_475),
.B(n_487),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

OAI21xp5_ASAP7_75t_L g493 ( 
.A1(n_476),
.A2(n_494),
.B(n_495),
.Y(n_493)
);

NOR2x1_ASAP7_75t_L g476 ( 
.A(n_477),
.B(n_484),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_477),
.B(n_484),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_478),
.B(n_481),
.C(n_483),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_478),
.B(n_490),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_481),
.A2(n_482),
.B1(n_483),
.B2(n_491),
.Y(n_490)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_483),
.Y(n_491)
);

OR2x2_ASAP7_75t_L g487 ( 
.A(n_488),
.B(n_489),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_488),
.B(n_489),
.Y(n_494)
);

INVx6_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

INVx13_ASAP7_75t_L g503 ( 
.A(n_500),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_502),
.B(n_504),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);


endmodule