module fake_jpeg_17497_n_191 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_191);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_191;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

CKINVDCx16_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_35),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_19),
.Y(n_61)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_24),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_39),
.A2(n_21),
.B1(n_1),
.B2(n_4),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_38),
.A2(n_31),
.B1(n_24),
.B2(n_20),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_43),
.A2(n_54),
.B1(n_59),
.B2(n_18),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_38),
.A2(n_20),
.B1(n_21),
.B2(n_23),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_44),
.A2(n_22),
.B1(n_21),
.B2(n_17),
.Y(n_77)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_22),
.Y(n_48)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_48),
.B(n_17),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_28),
.Y(n_52)
);

OAI21xp33_ASAP7_75t_L g72 ( 
.A1(n_52),
.A2(n_53),
.B(n_18),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_28),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_33),
.A2(n_20),
.B1(n_36),
.B2(n_41),
.Y(n_54)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_34),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_58),
.B(n_30),
.Y(n_79)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_59),
.A2(n_41),
.B1(n_36),
.B2(n_33),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_62),
.A2(n_68),
.B1(n_77),
.B2(n_27),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_52),
.B(n_40),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_63),
.B(n_73),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_53),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_65),
.B(n_66),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_53),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_50),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_67),
.B(n_76),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_69),
.B(n_27),
.Y(n_95)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_72),
.B(n_74),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_52),
.B(n_40),
.Y(n_73)
);

OA22x2_ASAP7_75t_L g74 ( 
.A1(n_49),
.A2(n_47),
.B1(n_56),
.B2(n_57),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_78),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_79),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_44),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_47),
.Y(n_94)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_60),
.C(n_37),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_83),
.B(n_88),
.Y(n_109)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_90),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_71),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_97),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_93),
.A2(n_94),
.B1(n_102),
.B2(n_29),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_95),
.B(n_29),
.Y(n_106)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_69),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_73),
.B(n_55),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_99),
.B(n_100),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_80),
.B(n_45),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_101),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_75),
.A2(n_77),
.B1(n_25),
.B2(n_56),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_98),
.A2(n_75),
.B(n_64),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_104),
.A2(n_98),
.B(n_87),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_106),
.B(n_116),
.Y(n_127)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_96),
.Y(n_107)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_107),
.Y(n_123)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_96),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_108),
.B(n_111),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_97),
.B(n_64),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_101),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_112),
.B(n_117),
.Y(n_136)
);

CKINVDCx14_ASAP7_75t_R g114 ( 
.A(n_89),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_114),
.B(n_119),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_82),
.B(n_78),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_84),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_100),
.A2(n_74),
.B(n_23),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_118),
.A2(n_16),
.B(n_74),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_90),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_120),
.A2(n_25),
.B1(n_98),
.B2(n_16),
.Y(n_124)
);

XNOR2x2_ASAP7_75t_SL g139 ( 
.A(n_121),
.B(n_133),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_103),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_122),
.B(n_124),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_109),
.B(n_83),
.C(n_86),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_125),
.B(n_126),
.C(n_128),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_104),
.B(n_86),
.C(n_99),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_91),
.C(n_85),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_118),
.A2(n_51),
.B1(n_85),
.B2(n_91),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_130),
.A2(n_134),
.B1(n_119),
.B2(n_113),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_115),
.B(n_74),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_SL g145 ( 
.A(n_131),
.B(n_137),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_105),
.A2(n_112),
.B1(n_108),
.B2(n_107),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_132),
.A2(n_129),
.B1(n_134),
.B2(n_128),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_105),
.A2(n_51),
.B1(n_88),
.B2(n_58),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_103),
.B(n_60),
.C(n_35),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_136),
.Y(n_138)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_138),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_140),
.A2(n_141),
.B1(n_143),
.B2(n_34),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_135),
.A2(n_113),
.B1(n_117),
.B2(n_40),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_123),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_142),
.B(n_144),
.Y(n_158)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_130),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_127),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_146),
.A2(n_147),
.B1(n_10),
.B2(n_12),
.Y(n_157)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_131),
.Y(n_147)
);

NAND3xp33_ASAP7_75t_L g150 ( 
.A(n_124),
.B(n_11),
.C(n_14),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_150),
.B(n_151),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_126),
.B(n_19),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_149),
.B(n_125),
.C(n_137),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_152),
.B(n_149),
.C(n_140),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_139),
.A2(n_15),
.B1(n_30),
.B2(n_4),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_154),
.B(n_159),
.Y(n_164)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_155),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_157),
.B(n_148),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_SL g159 ( 
.A(n_145),
.B(n_30),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_143),
.A2(n_7),
.B1(n_9),
.B2(n_6),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_160),
.B(n_162),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_145),
.B(n_35),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_161),
.B(n_139),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g162 ( 
.A(n_141),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_163),
.B(n_167),
.C(n_153),
.Y(n_174)
);

INVxp33_ASAP7_75t_L g165 ( 
.A(n_158),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_165),
.B(n_154),
.Y(n_171)
);

BUFx24_ASAP7_75t_SL g166 ( 
.A(n_156),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_166),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_169),
.B(n_161),
.Y(n_176)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_171),
.Y(n_181)
);

INVxp67_ASAP7_75t_SL g172 ( 
.A(n_165),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_172),
.B(n_173),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_168),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_174),
.B(n_177),
.C(n_170),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_176),
.B(n_15),
.C(n_6),
.Y(n_180)
);

MAJx2_ASAP7_75t_L g177 ( 
.A(n_164),
.B(n_159),
.C(n_152),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_178),
.B(n_179),
.C(n_180),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_171),
.B(n_162),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_182),
.B(n_175),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_183),
.B(n_185),
.Y(n_187)
);

MAJx2_ASAP7_75t_L g185 ( 
.A(n_181),
.B(n_7),
.C(n_1),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_184),
.B(n_182),
.Y(n_186)
);

OR2x2_ASAP7_75t_L g188 ( 
.A(n_186),
.B(n_19),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_188),
.B(n_187),
.Y(n_189)
);

AO21x2_ASAP7_75t_L g190 ( 
.A1(n_189),
.A2(n_0),
.B(n_5),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_190),
.B(n_5),
.Y(n_191)
);


endmodule