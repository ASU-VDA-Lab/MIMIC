module real_jpeg_4403_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_455;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_438;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g61 ( 
.A(n_0),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_1),
.A2(n_141),
.B1(n_143),
.B2(n_144),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_1),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_1),
.A2(n_143),
.B1(n_248),
.B2(n_249),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g324 ( 
.A1(n_1),
.A2(n_143),
.B1(n_325),
.B2(n_327),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_1),
.A2(n_143),
.B1(n_391),
.B2(n_396),
.Y(n_390)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_2),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_3),
.A2(n_45),
.B1(n_47),
.B2(n_50),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_3),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_3),
.A2(n_50),
.B1(n_127),
.B2(n_149),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_3),
.A2(n_50),
.B1(n_196),
.B2(n_197),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_3),
.A2(n_50),
.B1(n_88),
.B2(n_219),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_4),
.A2(n_185),
.B1(n_189),
.B2(n_190),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_4),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_4),
.A2(n_189),
.B1(n_320),
.B2(n_321),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_L g335 ( 
.A1(n_4),
.A2(n_33),
.B1(n_189),
.B2(n_336),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_4),
.A2(n_189),
.B1(n_375),
.B2(n_407),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_5),
.B(n_270),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_5),
.B(n_47),
.C(n_298),
.Y(n_297)
);

OAI22xp33_ASAP7_75t_L g301 ( 
.A1(n_5),
.A2(n_302),
.B1(n_303),
.B2(n_305),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_5),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_5),
.B(n_203),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_5),
.A2(n_26),
.B1(n_346),
.B2(n_349),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_5),
.B(n_150),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g437 ( 
.A1(n_5),
.A2(n_269),
.B(n_438),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_6),
.A2(n_258),
.B1(n_282),
.B2(n_285),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_6),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_6),
.A2(n_285),
.B1(n_309),
.B2(n_312),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_6),
.A2(n_285),
.B1(n_330),
.B2(n_347),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_6),
.A2(n_285),
.B1(n_386),
.B2(n_387),
.Y(n_385)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_7),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g157 ( 
.A(n_8),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_8),
.Y(n_178)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_8),
.Y(n_351)
);

INVx8_ASAP7_75t_L g359 ( 
.A(n_8),
.Y(n_359)
);

AOI22xp33_ASAP7_75t_L g32 ( 
.A1(n_9),
.A2(n_33),
.B1(n_38),
.B2(n_39),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_9),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_9),
.A2(n_38),
.B1(n_107),
.B2(n_122),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_9),
.A2(n_38),
.B1(n_163),
.B2(n_166),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g229 ( 
.A1(n_9),
.A2(n_38),
.B1(n_192),
.B2(n_230),
.Y(n_229)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_10),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g129 ( 
.A(n_11),
.Y(n_129)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_11),
.Y(n_134)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_11),
.Y(n_137)
);

BUFx5_ASAP7_75t_L g139 ( 
.A(n_11),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_11),
.Y(n_264)
);

BUFx5_ASAP7_75t_L g127 ( 
.A(n_12),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_12),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_12),
.Y(n_142)
);

BUFx5_ASAP7_75t_L g146 ( 
.A(n_12),
.Y(n_146)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_12),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_12),
.Y(n_192)
);

INVx6_ASAP7_75t_L g260 ( 
.A(n_12),
.Y(n_260)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_12),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_13),
.A2(n_86),
.B1(n_87),
.B2(n_90),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_13),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_13),
.A2(n_86),
.B1(n_173),
.B2(n_176),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_13),
.A2(n_86),
.B1(n_210),
.B2(n_214),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_14),
.Y(n_70)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_14),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_14),
.Y(n_78)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_14),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_15),
.A2(n_58),
.B1(n_62),
.B2(n_63),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_15),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_15),
.A2(n_62),
.B1(n_104),
.B2(n_107),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_15),
.A2(n_34),
.B1(n_62),
.B2(n_276),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_234),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_232),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_204),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_19),
.B(n_204),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_153),
.C(n_168),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_20),
.A2(n_21),
.B1(n_153),
.B2(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_93),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_22),
.B(n_123),
.C(n_152),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_54),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_23),
.A2(n_54),
.B1(n_55),
.B2(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_23),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_42),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g413 ( 
.A1(n_25),
.A2(n_275),
.B(n_414),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_32),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_26),
.A2(n_44),
.B(n_156),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_26),
.A2(n_172),
.B(n_177),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_26),
.A2(n_172),
.B1(n_274),
.B2(n_279),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_26),
.A2(n_42),
.B(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_26),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_26),
.A2(n_335),
.B1(n_346),
.B2(n_349),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_L g381 ( 
.A1(n_26),
.A2(n_44),
.B(n_177),
.Y(n_381)
);

OR2x2_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_30),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx8_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_31),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_32),
.Y(n_179)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx4_ASAP7_75t_L g348 ( 
.A(n_35),
.Y(n_348)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_36),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_37),
.Y(n_175)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g354 ( 
.A(n_40),
.B(n_355),
.Y(n_354)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_43),
.B(n_51),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_48),
.A2(n_78),
.B1(n_79),
.B2(n_81),
.Y(n_77)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_53),
.Y(n_279)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_66),
.B1(n_83),
.B2(n_85),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_57),
.A2(n_84),
.B1(n_160),
.B2(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_60),
.Y(n_166)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g304 ( 
.A(n_61),
.Y(n_304)
);

INVx3_ASAP7_75t_L g307 ( 
.A(n_61),
.Y(n_307)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_66),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_66),
.A2(n_83),
.B1(n_301),
.B2(n_308),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_66),
.A2(n_83),
.B1(n_308),
.B2(n_319),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_66),
.A2(n_83),
.B1(n_319),
.B2(n_390),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_77),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_69),
.B1(n_71),
.B2(n_74),
.Y(n_67)
);

INVx5_ASAP7_75t_L g296 ( 
.A(n_68),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_74),
.Y(n_313)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_75),
.Y(n_311)
);

INVx6_ASAP7_75t_L g372 ( 
.A(n_75),
.Y(n_372)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_76),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_76),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_76),
.Y(n_395)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_77),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx5_ASAP7_75t_L g176 ( 
.A(n_80),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_80),
.Y(n_326)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_80),
.Y(n_330)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_82),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_83),
.B(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_84),
.B(n_218),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_84),
.B(n_302),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_85),
.Y(n_159)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

OA22x2_ASAP7_75t_L g95 ( 
.A1(n_92),
.A2(n_96),
.B1(n_98),
.B2(n_101),
.Y(n_95)
);

INVx5_ASAP7_75t_L g220 ( 
.A(n_92),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_94),
.A2(n_123),
.B1(n_124),
.B2(n_152),
.Y(n_93)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_94),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_103),
.B(n_108),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_95),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_95),
.B(n_195),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_95),
.A2(n_201),
.B1(n_405),
.B2(n_406),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_95),
.A2(n_201),
.B1(n_406),
.B2(n_434),
.Y(n_433)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx6_ASAP7_75t_L g373 ( 
.A(n_98),
.Y(n_373)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_99),
.Y(n_120)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_100),
.Y(n_102)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_100),
.Y(n_116)
);

INVx3_ASAP7_75t_L g380 ( 
.A(n_100),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_103),
.Y(n_208)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_104),
.Y(n_107)
);

INVx5_ASAP7_75t_L g248 ( 
.A(n_104),
.Y(n_248)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_106),
.Y(n_113)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_106),
.Y(n_119)
);

BUFx5_ASAP7_75t_L g200 ( 
.A(n_106),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_106),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_106),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_109),
.B(n_121),
.Y(n_108)
);

INVx2_ASAP7_75t_SL g201 ( 
.A(n_109),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_109),
.A2(n_203),
.B1(n_208),
.B2(n_209),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_109),
.A2(n_247),
.B(n_252),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_109),
.A2(n_203),
.B1(n_384),
.B2(n_385),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_111),
.A2(n_114),
.B1(n_117),
.B2(n_120),
.Y(n_110)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_112),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_113),
.Y(n_136)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_113),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_113),
.Y(n_257)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_119),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_121),
.B(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_140),
.B(n_147),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_125),
.A2(n_140),
.B1(n_151),
.B2(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_125),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g436 ( 
.A1(n_125),
.A2(n_151),
.B1(n_437),
.B2(n_440),
.Y(n_436)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_135),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_128),
.B1(n_130),
.B2(n_132),
.Y(n_126)
);

INVx8_ASAP7_75t_L g149 ( 
.A(n_127),
.Y(n_149)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_134),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g151 ( 
.A(n_135),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_137),
.B1(n_138),
.B2(n_139),
.Y(n_135)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_150),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_148),
.A2(n_227),
.B(n_228),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_150),
.A2(n_227),
.B1(n_281),
.B2(n_286),
.Y(n_280)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_151),
.B(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_153),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_155),
.B1(n_158),
.B2(n_167),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_154),
.A2(n_155),
.B1(n_226),
.B2(n_231),
.Y(n_225)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_155),
.B(n_158),
.Y(n_224)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_158),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_160),
.B(n_161),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_160),
.B(n_181),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g420 ( 
.A1(n_160),
.A2(n_421),
.B(n_422),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_L g435 ( 
.A1(n_160),
.A2(n_161),
.B(n_218),
.Y(n_435)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_162),
.Y(n_181)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g320 ( 
.A(n_165),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_168),
.B(n_238),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_182),
.C(n_193),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_170),
.B(n_242),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_180),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_171),
.B(n_180),
.Y(n_450)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx8_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_182),
.A2(n_183),
.B1(n_193),
.B2(n_194),
.Y(n_242)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_184),
.Y(n_286)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_187),
.Y(n_230)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx8_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_201),
.B(n_202),
.Y(n_194)
);

INVx8_ASAP7_75t_L g369 ( 
.A(n_196),
.Y(n_369)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx6_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_200),
.Y(n_377)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_200),
.Y(n_410)
);

BUFx24_ASAP7_75t_SL g462 ( 
.A(n_204),
.Y(n_462)
);

FAx1_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.CI(n_223),
.CON(n_204),
.SN(n_204)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_216),
.B(n_222),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_207),
.B(n_216),
.Y(n_222)
);

OAI21xp33_ASAP7_75t_SL g384 ( 
.A1(n_210),
.A2(n_302),
.B(n_374),
.Y(n_384)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

BUFx2_ASAP7_75t_L g386 ( 
.A(n_212),
.Y(n_386)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_213),
.Y(n_215)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_221),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g422 ( 
.A(n_217),
.Y(n_422)
);

BUFx3_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_226),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_287),
.B(n_458),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_237),
.B(n_240),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_237),
.B(n_240),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_243),
.C(n_245),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_241),
.B(n_243),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_SL g444 ( 
.A(n_245),
.B(n_445),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_253),
.C(n_280),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_246),
.B(n_280),
.Y(n_448)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_247),
.Y(n_434)
);

INVx1_ASAP7_75t_SL g249 ( 
.A(n_250),
.Y(n_249)
);

INVx6_ASAP7_75t_SL g250 ( 
.A(n_251),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_251),
.B(n_266),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_253),
.B(n_448),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_273),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_254),
.B(n_273),
.Y(n_430)
);

OAI32xp33_ASAP7_75t_L g254 ( 
.A1(n_255),
.A2(n_258),
.A3(n_261),
.B1(n_265),
.B2(n_268),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

BUFx12f_ASAP7_75t_L g388 ( 
.A(n_257),
.Y(n_388)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_259),
.Y(n_258)
);

INVx8_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_260),
.Y(n_439)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx8_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVxp33_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx2_ASAP7_75t_SL g270 ( 
.A(n_271),
.Y(n_270)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_272),
.Y(n_284)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx6_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_SL g336 ( 
.A(n_278),
.Y(n_336)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_281),
.Y(n_440)
);

INVx4_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx5_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_288),
.A2(n_442),
.B(n_455),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_290),
.A2(n_426),
.B(n_441),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_291),
.A2(n_399),
.B(n_425),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_292),
.A2(n_363),
.B(n_398),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_293),
.A2(n_331),
.B(n_362),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_314),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_294),
.B(n_314),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_300),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_295),
.B(n_300),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_302),
.B(n_356),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_302),
.B(n_375),
.Y(n_374)
);

INVx3_ASAP7_75t_SL g303 ( 
.A(n_304),
.Y(n_303)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_304),
.Y(n_397)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

BUFx3_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_307),
.Y(n_321)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

BUFx2_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_323),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_316),
.A2(n_317),
.B1(n_318),
.B2(n_322),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_316),
.B(n_322),
.C(n_323),
.Y(n_364)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_SL g322 ( 
.A(n_318),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_321),
.B(n_379),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_324),
.Y(n_338)
);

INVx3_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx6_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_332),
.A2(n_342),
.B(n_361),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_341),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_333),
.B(n_341),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_334),
.A2(n_337),
.B1(n_338),
.B2(n_339),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g342 ( 
.A1(n_343),
.A2(n_352),
.B(n_360),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_345),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_344),
.B(n_345),
.Y(n_360)
);

INVx4_ASAP7_75t_SL g347 ( 
.A(n_348),
.Y(n_347)
);

INVx5_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_353),
.B(n_354),
.Y(n_352)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_356),
.Y(n_414)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx8_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_365),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_364),
.B(n_365),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_382),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_366),
.B(n_383),
.C(n_389),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_SL g366 ( 
.A(n_367),
.B(n_381),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_367),
.B(n_381),
.Y(n_419)
);

OAI32xp33_ASAP7_75t_L g367 ( 
.A1(n_368),
.A2(n_370),
.A3(n_373),
.B1(n_374),
.B2(n_378),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx3_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx6_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_389),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_385),
.Y(n_405)
);

INVx3_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVxp67_ASAP7_75t_L g421 ( 
.A(n_390),
.Y(n_421)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_401),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_400),
.B(n_401),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_402),
.A2(n_403),
.B1(n_417),
.B2(n_418),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_402),
.B(n_420),
.C(n_423),
.Y(n_427)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_SL g403 ( 
.A(n_404),
.B(n_411),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_404),
.B(n_412),
.C(n_416),
.Y(n_431)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_412),
.A2(n_413),
.B1(n_415),
.B2(n_416),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_415),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_419),
.A2(n_420),
.B1(n_423),
.B2(n_424),
.Y(n_418)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_419),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_420),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_428),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_427),
.B(n_428),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_429),
.B(n_432),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_431),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_430),
.B(n_431),
.C(n_432),
.Y(n_452)
);

BUFx24_ASAP7_75t_SL g460 ( 
.A(n_432),
.Y(n_460)
);

FAx1_ASAP7_75t_L g432 ( 
.A(n_433),
.B(n_435),
.CI(n_436),
.CON(n_432),
.SN(n_432)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_433),
.B(n_435),
.C(n_436),
.Y(n_449)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_SL g442 ( 
.A(n_443),
.B(n_451),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_L g455 ( 
.A1(n_443),
.A2(n_456),
.B(n_457),
.Y(n_455)
);

NOR2xp67_ASAP7_75t_SL g443 ( 
.A(n_444),
.B(n_446),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_444),
.B(n_446),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_447),
.B(n_449),
.C(n_450),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_447),
.B(n_454),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_449),
.B(n_450),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_452),
.B(n_453),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_452),
.B(n_453),
.Y(n_456)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);


endmodule