module real_jpeg_29382_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_0),
.B(n_48),
.Y(n_47)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

HB1xp67_ASAP7_75t_L g154 ( 
.A(n_0),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g24 ( 
.A1(n_1),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

OAI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_1),
.A2(n_28),
.B1(n_85),
.B2(n_86),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_1),
.A2(n_28),
.B1(n_35),
.B2(n_36),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_1),
.A2(n_28),
.B1(n_48),
.B2(n_51),
.Y(n_147)
);

OAI22xp33_ASAP7_75t_L g38 ( 
.A1(n_2),
.A2(n_25),
.B1(n_26),
.B2(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_2),
.A2(n_35),
.B1(n_36),
.B2(n_39),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_2),
.A2(n_39),
.B1(n_48),
.B2(n_51),
.Y(n_141)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

BUFx8_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

INVx13_ASAP7_75t_L g86 ( 
.A(n_5),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_6),
.A2(n_35),
.B1(n_36),
.B2(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_6),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_6),
.A2(n_25),
.B1(n_26),
.B2(n_65),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_6),
.A2(n_48),
.B1(n_51),
.B2(n_65),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_7),
.A2(n_35),
.B1(n_36),
.B2(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_7),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_7),
.A2(n_48),
.B1(n_51),
.B2(n_67),
.Y(n_77)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_8),
.Y(n_61)
);

OAI32xp33_ASAP7_75t_L g124 ( 
.A1(n_8),
.A2(n_35),
.A3(n_51),
.B1(n_125),
.B2(n_126),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_9),
.A2(n_48),
.B1(n_51),
.B2(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_10),
.A2(n_48),
.B1(n_51),
.B2(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_10),
.Y(n_90)
);

BUFx24_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

A2O1A1Ixp33_ASAP7_75t_L g30 ( 
.A1(n_12),
.A2(n_25),
.B(n_31),
.C(n_34),
.Y(n_30)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_12),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_34)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_13),
.A2(n_48),
.B1(n_51),
.B2(n_52),
.Y(n_50)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_L g104 ( 
.A1(n_13),
.A2(n_35),
.B1(n_36),
.B2(n_52),
.Y(n_104)
);

INVx11_ASAP7_75t_SL g49 ( 
.A(n_14),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_15),
.B(n_43),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_15),
.Y(n_72)
);

AOI21xp33_ASAP7_75t_SL g84 ( 
.A1(n_15),
.A2(n_26),
.B(n_44),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_15),
.A2(n_72),
.B1(n_85),
.B2(n_86),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_15),
.A2(n_35),
.B(n_121),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_15),
.B(n_35),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_15),
.B(n_40),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_15),
.A2(n_54),
.B1(n_76),
.B2(n_147),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_15),
.A2(n_25),
.B(n_164),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_113),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_111),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_80),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_19),
.B(n_80),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_57),
.C(n_68),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_20),
.A2(n_21),
.B1(n_176),
.B2(n_177),
.Y(n_175)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_41),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_22),
.B(n_42),
.C(n_46),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_29),
.B1(n_38),
.B2(n_40),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_24),
.A2(n_30),
.B1(n_34),
.B2(n_163),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_32),
.Y(n_31)
);

AO22x1_ASAP7_75t_L g43 ( 
.A1(n_25),
.A2(n_26),
.B1(n_44),
.B2(n_45),
.Y(n_43)
);

OAI32xp33_ASAP7_75t_L g70 ( 
.A1(n_25),
.A2(n_32),
.A3(n_36),
.B1(n_71),
.B2(n_73),
.Y(n_70)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_26),
.B(n_72),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_30),
.A2(n_34),
.B1(n_98),
.B2(n_99),
.Y(n_97)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_32),
.Y(n_74)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

OAI22xp33_ASAP7_75t_L g62 ( 
.A1(n_35),
.A2(n_36),
.B1(n_60),
.B2(n_61),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_35),
.B(n_74),
.Y(n_73)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_38),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_46),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_43),
.A2(n_107),
.B1(n_109),
.B2(n_110),
.Y(n_106)
);

O2A1O1Ixp33_ASAP7_75t_L g107 ( 
.A1(n_43),
.A2(n_44),
.B(n_86),
.C(n_108),
.Y(n_107)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_44),
.Y(n_45)
);

NAND2xp33_ASAP7_75t_SL g108 ( 
.A(n_44),
.B(n_86),
.Y(n_108)
);

A2O1A1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_45),
.A2(n_72),
.B(n_84),
.C(n_85),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_50),
.B1(n_53),
.B2(n_55),
.Y(n_46)
);

CKINVDCx14_ASAP7_75t_R g76 ( 
.A(n_47),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_47),
.A2(n_55),
.B1(n_88),
.B2(n_89),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_47),
.A2(n_88),
.B1(n_140),
.B2(n_142),
.Y(n_139)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_48),
.A2(n_51),
.B1(n_60),
.B2(n_61),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_48),
.B(n_61),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_48),
.B(n_152),
.Y(n_151)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_50),
.Y(n_79)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

INVx5_ASAP7_75t_SL g136 ( 
.A(n_53),
.Y(n_136)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_57),
.A2(n_68),
.B1(n_69),
.B2(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_57),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_59),
.B1(n_63),
.B2(n_66),
.Y(n_57)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_58),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_58),
.A2(n_59),
.B1(n_120),
.B2(n_122),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_58),
.A2(n_59),
.B1(n_122),
.B2(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_59),
.B(n_62),
.Y(n_58)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_59),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_59),
.B(n_72),
.Y(n_148)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_64),
.A2(n_103),
.B1(n_105),
.B2(n_166),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_66),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_75),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_70),
.B(n_75),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_71),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_72),
.B(n_153),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_77),
.B1(n_78),
.B2(n_79),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_76),
.A2(n_77),
.B1(n_135),
.B2(n_136),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_76),
.A2(n_78),
.B1(n_141),
.B2(n_147),
.Y(n_146)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_94),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_91),
.B1(n_92),
.B2(n_93),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_82),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_87),
.Y(n_82)
);

CKINVDCx5p33_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_91),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_106),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_97),
.B1(n_100),
.B2(n_101),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_103),
.B1(n_104),
.B2(n_105),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_114),
.A2(n_173),
.B(n_179),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_158),
.B(n_172),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_137),
.B(n_157),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_127),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_117),
.B(n_127),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_118),
.B(n_123),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_118),
.A2(n_119),
.B1(n_123),
.B2(n_124),
.Y(n_143)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_121),
.Y(n_125)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_134),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_130),
.B1(n_131),
.B2(n_132),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_129),
.B(n_132),
.C(n_134),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_133),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_135),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_144),
.B(n_156),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_143),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_139),
.B(n_143),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_145),
.A2(n_149),
.B(n_155),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_148),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_146),
.B(n_148),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_150),
.B(n_151),
.Y(n_149)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_159),
.B(n_160),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_161),
.A2(n_169),
.B1(n_170),
.B2(n_171),
.Y(n_160)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_161),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_165),
.B1(n_167),
.B2(n_168),
.Y(n_161)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_162),
.Y(n_168)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_165),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_165),
.B(n_168),
.C(n_171),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_169),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_174),
.B(n_175),
.Y(n_179)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);


endmodule