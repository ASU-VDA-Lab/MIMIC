module real_jpeg_23646_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_215;
wire n_221;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_139;
wire n_33;
wire n_188;
wire n_65;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_193;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_15;
wire n_130;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_128;
wire n_202;
wire n_179;
wire n_167;
wire n_213;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

OAI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_2),
.A2(n_33),
.B1(n_35),
.B2(n_36),
.Y(n_32)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_2),
.A2(n_35),
.B1(n_51),
.B2(n_53),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_2),
.A2(n_35),
.B1(n_61),
.B2(n_62),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_2),
.A2(n_21),
.B1(n_24),
.B2(n_35),
.Y(n_146)
);

BUFx8_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g67 ( 
.A(n_4),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_6),
.A2(n_21),
.B1(n_24),
.B2(n_25),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_6),
.A2(n_25),
.B1(n_33),
.B2(n_36),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g28 ( 
.A1(n_7),
.A2(n_21),
.B1(n_24),
.B2(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_7),
.A2(n_29),
.B1(n_33),
.B2(n_36),
.Y(n_115)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_8),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_8),
.A2(n_9),
.B1(n_44),
.B2(n_70),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_9),
.A2(n_33),
.B1(n_36),
.B2(n_44),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_9),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_9),
.A2(n_44),
.B1(n_51),
.B2(n_53),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_9),
.A2(n_21),
.B1(n_24),
.B2(n_44),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_9),
.B(n_53),
.C(n_67),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_9),
.B(n_68),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_9),
.B(n_33),
.C(n_49),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_9),
.B(n_21),
.C(n_39),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_9),
.B(n_11),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_9),
.B(n_42),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_9),
.B(n_118),
.Y(n_203)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_11),
.Y(n_80)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_11),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_11),
.A2(n_145),
.B1(n_146),
.B2(n_147),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_122),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_121),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_102),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_16),
.B(n_102),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_74),
.C(n_86),
.Y(n_16)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_17),
.B(n_74),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_45),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_SL g120 ( 
.A(n_18),
.B(n_58),
.C(n_72),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_30),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_19),
.A2(n_30),
.B1(n_31),
.B2(n_232),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_19),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_23),
.B1(n_26),
.B2(n_28),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_20),
.B(n_78),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_20),
.B(n_93),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_20),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_22),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_21),
.Y(n_24)
);

OA22x2_ASAP7_75t_L g41 ( 
.A1(n_21),
.A2(n_24),
.B1(n_39),
.B2(n_40),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_21),
.B(n_193),
.Y(n_192)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_23),
.A2(n_90),
.B(n_91),
.Y(n_89)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_28),
.B(n_76),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_30),
.A2(n_31),
.B1(n_203),
.B2(n_204),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_30),
.A2(n_31),
.B1(n_172),
.B2(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_31),
.B(n_166),
.C(n_172),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_31),
.B(n_144),
.C(n_203),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_37),
.B1(n_42),
.B2(n_43),
.Y(n_31)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_32),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_33),
.Y(n_36)
);

OAI22xp33_ASAP7_75t_L g38 ( 
.A1(n_33),
.A2(n_36),
.B1(n_39),
.B2(n_40),
.Y(n_38)
);

OA22x2_ASAP7_75t_SL g47 ( 
.A1(n_33),
.A2(n_36),
.B1(n_48),
.B2(n_49),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_33),
.B(n_188),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_37),
.B(n_43),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_37),
.A2(n_42),
.B1(n_113),
.B2(n_114),
.Y(n_112)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_37),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_41),
.Y(n_37)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_39),
.Y(n_40)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_41),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_41),
.A2(n_83),
.B(n_84),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_41),
.A2(n_84),
.B(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_41),
.B(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_43),
.B(n_134),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_46),
.A2(n_58),
.B1(n_72),
.B2(n_73),
.Y(n_45)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_46),
.A2(n_72),
.B1(n_133),
.B2(n_156),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_46),
.A2(n_72),
.B1(n_94),
.B2(n_129),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_46),
.B(n_94),
.C(n_210),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_50),
.B(n_54),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_56),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_47),
.A2(n_97),
.B(n_98),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_47),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_48),
.A2(n_49),
.B1(n_51),
.B2(n_53),
.Y(n_56)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_50),
.Y(n_117)
);

INVx3_ASAP7_75t_SL g53 ( 
.A(n_51),
.Y(n_53)
);

AO22x1_ASAP7_75t_SL g68 ( 
.A1(n_51),
.A2(n_53),
.B1(n_66),
.B2(n_67),
.Y(n_68)
);

CKINVDCx6p67_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_53),
.B(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_55),
.B(n_57),
.Y(n_54)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_55),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_55),
.A2(n_57),
.B1(n_117),
.B2(n_118),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_57),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_58),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_58),
.A2(n_73),
.B1(n_116),
.B2(n_149),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_58),
.B(n_116),
.C(n_139),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_63),
.B1(n_68),
.B2(n_69),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_60),
.A2(n_100),
.B(n_101),
.Y(n_99)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_61),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_61),
.A2(n_65),
.B1(n_66),
.B2(n_67),
.Y(n_64)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_63),
.B(n_69),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_63),
.B(n_68),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_68),
.Y(n_63)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_68),
.Y(n_100)
);

INVxp33_ASAP7_75t_L g109 ( 
.A(n_69),
.Y(n_109)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_71),
.B(n_142),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_72),
.B(n_132),
.C(n_133),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_81),
.B1(n_82),
.B2(n_85),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_75),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_75),
.A2(n_85),
.B1(n_106),
.B2(n_107),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_75),
.B(n_82),
.Y(n_110)
);

INVxp33_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_77),
.B(n_147),
.Y(n_177)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_83),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_86),
.B(n_238),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_96),
.C(n_99),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_87),
.A2(n_88),
.B1(n_227),
.B2(n_228),
.Y(n_226)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_94),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_89),
.A2(n_94),
.B1(n_129),
.B2(n_130),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_89),
.Y(n_130)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_90),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_92),
.A2(n_146),
.B(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_93),
.Y(n_147)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_94),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_94),
.A2(n_129),
.B1(n_187),
.B2(n_189),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_94),
.B(n_189),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_96),
.A2(n_99),
.B1(n_132),
.B2(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_96),
.Y(n_229)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_99),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_99),
.A2(n_132),
.B1(n_154),
.B2(n_155),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_120),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_111),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_SL g104 ( 
.A(n_105),
.B(n_110),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_108),
.B(n_109),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_116),
.B(n_119),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_112),
.B(n_116),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_116),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_116),
.B(n_159),
.C(n_161),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_116),
.A2(n_149),
.B1(n_168),
.B2(n_169),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_235),
.B(n_239),
.Y(n_122)
);

A2O1A1Ixp33_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_162),
.B(n_221),
.C(n_234),
.Y(n_123)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_151),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_125),
.B(n_151),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_127),
.B1(n_138),
.B2(n_150),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_131),
.B1(n_136),
.B2(n_137),
.Y(n_127)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_128),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_128),
.B(n_137),
.C(n_150),
.Y(n_222)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_131),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_133),
.Y(n_156)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_138),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_148),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_143),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_140),
.A2(n_141),
.B1(n_143),
.B2(n_144),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_143),
.A2(n_144),
.B1(n_201),
.B2(n_202),
.Y(n_200)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_144),
.B(n_195),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_144),
.B(n_195),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_157),
.C(n_158),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_152),
.A2(n_153),
.B1(n_179),
.B2(n_180),
.Y(n_178)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_157),
.B(n_158),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_159),
.A2(n_161),
.B1(n_170),
.B2(n_171),
.Y(n_169)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_159),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_159),
.B(n_192),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_161),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_163),
.B(n_220),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_181),
.B(n_219),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_178),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_165),
.B(n_178),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_166),
.A2(n_167),
.B1(n_215),
.B2(n_217),
.Y(n_214)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_171),
.B(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_171),
.B(n_186),
.Y(n_197)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_172),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_176),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_173),
.A2(n_174),
.B1(n_176),
.B2(n_177),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_212),
.B(n_218),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_183),
.A2(n_206),
.B(n_211),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_198),
.B(n_205),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_185),
.A2(n_190),
.B(n_197),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_187),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_194),
.B(n_196),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_199),
.B(n_200),
.Y(n_205)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_203),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_207),
.B(n_208),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_213),
.B(n_214),
.Y(n_218)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_215),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_222),
.B(n_223),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_233),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_225),
.A2(n_226),
.B1(n_230),
.B2(n_231),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_225),
.B(n_231),
.C(n_233),
.Y(n_236)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

CKINVDCx14_ASAP7_75t_R g230 ( 
.A(n_231),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_236),
.B(n_237),
.Y(n_239)
);


endmodule