module fake_jpeg_23969_n_346 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_346);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_346;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_16),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_1),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_37),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_43),
.Y(n_53)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_23),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_41),
.A2(n_22),
.B1(n_28),
.B2(n_20),
.Y(n_61)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_45),
.Y(n_68)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_46),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_20),
.B(n_7),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_47),
.B(n_28),
.Y(n_66)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_49),
.Y(n_60)
);

AOI21xp33_ASAP7_75t_SL g51 ( 
.A1(n_40),
.A2(n_18),
.B(n_35),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_33),
.C(n_28),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_54),
.B(n_63),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_45),
.A2(n_23),
.B1(n_27),
.B2(n_33),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_55),
.A2(n_26),
.B1(n_36),
.B2(n_24),
.Y(n_99)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_45),
.A2(n_23),
.B1(n_27),
.B2(n_33),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_57),
.A2(n_48),
.B1(n_44),
.B2(n_22),
.Y(n_96)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_61),
.A2(n_64),
.B1(n_29),
.B2(n_32),
.Y(n_75)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_39),
.A2(n_27),
.B1(n_20),
.B2(n_29),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_66),
.B(n_32),
.Y(n_84)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_51),
.A2(n_39),
.B1(n_40),
.B2(n_43),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_71),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_72),
.B(n_98),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_67),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_74),
.B(n_79),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_75),
.A2(n_78),
.B1(n_99),
.B2(n_101),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_76),
.B(n_83),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_69),
.A2(n_32),
.B1(n_22),
.B2(n_29),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_67),
.Y(n_79)
);

OR2x2_ASAP7_75t_SL g80 ( 
.A(n_66),
.B(n_47),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_80),
.A2(n_34),
.B(n_24),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_SL g82 ( 
.A(n_53),
.B(n_42),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_82),
.B(n_35),
.C(n_31),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_67),
.Y(n_83)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_84),
.Y(n_114)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_86),
.Y(n_134)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_88),
.Y(n_106)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_52),
.B(n_18),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_90),
.B(n_93),
.Y(n_124)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_69),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g119 ( 
.A(n_91),
.Y(n_119)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_69),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_92),
.Y(n_133)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_57),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_52),
.B(n_17),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_94),
.B(n_105),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_58),
.Y(n_95)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_96),
.A2(n_25),
.B1(n_35),
.B2(n_31),
.Y(n_111)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_62),
.Y(n_97)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_97),
.Y(n_125)
);

AND2x4_ASAP7_75t_L g98 ( 
.A(n_62),
.B(n_37),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_56),
.A2(n_36),
.B(n_26),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_100),
.A2(n_105),
.B(n_98),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_50),
.A2(n_43),
.B1(n_26),
.B2(n_25),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_63),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_102),
.B(n_3),
.Y(n_135)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_50),
.Y(n_103)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_103),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_65),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_104),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_70),
.B(n_17),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_108),
.A2(n_102),
.B(n_81),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_88),
.A2(n_60),
.B1(n_59),
.B2(n_36),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_109),
.A2(n_110),
.B1(n_111),
.B2(n_120),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_71),
.A2(n_60),
.B1(n_59),
.B2(n_34),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_115),
.B(n_74),
.C(n_79),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_82),
.B(n_37),
.C(n_35),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_117),
.B(n_99),
.C(n_87),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_93),
.A2(n_31),
.B1(n_19),
.B2(n_2),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_122),
.A2(n_132),
.B(n_80),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_90),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_123),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_72),
.A2(n_31),
.B1(n_1),
.B2(n_2),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_127),
.A2(n_130),
.B1(n_73),
.B2(n_91),
.Y(n_156)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_98),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_128),
.B(n_92),
.Y(n_139)
);

OA22x2_ASAP7_75t_L g130 ( 
.A1(n_98),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_130)
);

O2A1O1Ixp33_ASAP7_75t_L g132 ( 
.A1(n_96),
.A2(n_0),
.B(n_3),
.C(n_4),
.Y(n_132)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_135),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_123),
.B(n_76),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_136),
.B(n_137),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_106),
.B(n_86),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_139),
.A2(n_142),
.B(n_133),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_140),
.B(n_144),
.C(n_154),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_106),
.B(n_100),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_141),
.A2(n_152),
.B(n_155),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_113),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_143),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_134),
.B(n_85),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g194 ( 
.A(n_146),
.Y(n_194)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_129),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_147),
.B(n_149),
.Y(n_197)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_124),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_119),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_150),
.B(n_151),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_131),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_124),
.B(n_89),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_109),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_153),
.B(n_157),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_117),
.B(n_104),
.C(n_77),
.Y(n_154)
);

OAI21xp33_ASAP7_75t_L g155 ( 
.A1(n_122),
.A2(n_16),
.B(n_4),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_156),
.A2(n_159),
.B1(n_73),
.B2(n_97),
.Y(n_193)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_135),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_110),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_158),
.B(n_163),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_121),
.A2(n_128),
.B1(n_115),
.B2(n_111),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_113),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_160),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_112),
.B(n_94),
.Y(n_161)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_161),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_134),
.B(n_85),
.Y(n_162)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_162),
.Y(n_176)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_120),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_130),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_164),
.B(n_166),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_107),
.B(n_103),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_165),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_163),
.A2(n_121),
.B1(n_118),
.B2(n_112),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_168),
.A2(n_159),
.B1(n_148),
.B2(n_156),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_140),
.B(n_112),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_169),
.B(n_174),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_161),
.B(n_127),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_170),
.B(n_173),
.C(n_145),
.Y(n_203)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_146),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_171),
.B(n_180),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_140),
.B(n_108),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_154),
.B(n_144),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_153),
.A2(n_114),
.B1(n_130),
.B2(n_132),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_177),
.A2(n_190),
.B1(n_193),
.B2(n_201),
.Y(n_215)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_162),
.Y(n_180)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_136),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_183),
.B(n_184),
.Y(n_213)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_137),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_143),
.B(n_133),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_185),
.B(n_126),
.Y(n_207)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_160),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_187),
.B(n_188),
.Y(n_216)
);

INVxp33_ASAP7_75t_L g188 ( 
.A(n_139),
.Y(n_188)
);

AOI22x1_ASAP7_75t_SL g190 ( 
.A1(n_142),
.A2(n_130),
.B1(n_107),
.B2(n_114),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_165),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_191),
.B(n_199),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_192),
.A2(n_166),
.B(n_157),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_147),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_195),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_152),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_141),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_200),
.B(n_148),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_138),
.A2(n_126),
.B1(n_116),
.B2(n_125),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_202),
.A2(n_167),
.B1(n_182),
.B2(n_190),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_203),
.B(n_227),
.C(n_170),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_181),
.A2(n_138),
.B(n_149),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_204),
.A2(n_209),
.B(n_220),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_196),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_206),
.Y(n_246)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_207),
.Y(n_238)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_201),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_208),
.B(n_219),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_189),
.B(n_145),
.Y(n_211)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_211),
.Y(n_243)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_212),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_198),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_214),
.B(n_218),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_197),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_172),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_192),
.A2(n_164),
.B(n_125),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_186),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_221),
.B(n_228),
.Y(n_234)
);

NOR2x1_ASAP7_75t_L g222 ( 
.A(n_195),
.B(n_164),
.Y(n_222)
);

OR2x2_ASAP7_75t_L g257 ( 
.A(n_222),
.B(n_218),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_193),
.A2(n_183),
.B1(n_179),
.B2(n_178),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_223),
.A2(n_226),
.B1(n_168),
.B2(n_200),
.Y(n_233)
);

O2A1O1Ixp33_ASAP7_75t_L g224 ( 
.A1(n_191),
.A2(n_95),
.B(n_116),
.C(n_81),
.Y(n_224)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_224),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_186),
.B(n_3),
.Y(n_225)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_225),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_177),
.A2(n_77),
.B1(n_95),
.B2(n_7),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_182),
.B(n_5),
.C(n_6),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_184),
.B(n_5),
.Y(n_228)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_187),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_230),
.B(n_180),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g231 ( 
.A(n_188),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_231),
.Y(n_251)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_233),
.Y(n_278)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_235),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_236),
.B(n_254),
.C(n_8),
.Y(n_276)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_237),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_208),
.A2(n_176),
.B1(n_194),
.B2(n_171),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_240),
.A2(n_205),
.B(n_219),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_203),
.B(n_169),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_241),
.B(n_249),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_216),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_242),
.B(n_255),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_202),
.A2(n_167),
.B1(n_174),
.B2(n_173),
.Y(n_247)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_247),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_210),
.B(n_175),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_210),
.B(n_175),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_250),
.B(n_223),
.Y(n_267)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_224),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_252),
.B(n_222),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_221),
.B(n_13),
.C(n_7),
.Y(n_254)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_229),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_212),
.A2(n_6),
.B1(n_8),
.B2(n_10),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_256),
.A2(n_228),
.B1(n_209),
.B2(n_220),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_257),
.B(n_211),
.Y(n_259)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_258),
.Y(n_292)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_259),
.Y(n_296)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_251),
.Y(n_260)
);

CKINVDCx11_ASAP7_75t_R g288 ( 
.A(n_260),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_253),
.A2(n_204),
.B(n_213),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_261),
.A2(n_266),
.B(n_271),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_234),
.B(n_225),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_262),
.B(n_265),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_263),
.B(n_268),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_234),
.B(n_243),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_253),
.A2(n_217),
.B(n_215),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_267),
.B(n_10),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_246),
.B(n_206),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_251),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_269),
.B(n_11),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_232),
.A2(n_230),
.B(n_214),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_273),
.A2(n_232),
.B1(n_237),
.B2(n_252),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_239),
.A2(n_205),
.B1(n_227),
.B2(n_225),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_274),
.A2(n_244),
.B1(n_256),
.B2(n_233),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_276),
.B(n_254),
.C(n_245),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_279),
.A2(n_289),
.B1(n_271),
.B2(n_284),
.Y(n_305)
);

BUFx2_ASAP7_75t_L g280 ( 
.A(n_260),
.Y(n_280)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_280),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_267),
.B(n_241),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_281),
.B(n_286),
.Y(n_297)
);

A2O1A1O1Ixp25_ASAP7_75t_L g282 ( 
.A1(n_266),
.A2(n_250),
.B(n_249),
.C(n_247),
.D(n_257),
.Y(n_282)
);

MAJx2_ASAP7_75t_L g301 ( 
.A(n_282),
.B(n_293),
.C(n_263),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_285),
.B(n_276),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_277),
.B(n_236),
.Y(n_286)
);

OA21x2_ASAP7_75t_SL g290 ( 
.A1(n_261),
.A2(n_248),
.B(n_238),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_290),
.A2(n_265),
.B(n_262),
.Y(n_300)
);

NOR3xp33_ASAP7_75t_SL g291 ( 
.A(n_259),
.B(n_10),
.C(n_11),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_291),
.B(n_12),
.Y(n_311)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_294),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_270),
.B(n_11),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_295),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_283),
.B(n_273),
.C(n_272),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_298),
.B(n_303),
.Y(n_313)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_299),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_300),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_301),
.A2(n_289),
.B1(n_296),
.B2(n_285),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_288),
.Y(n_303)
);

MAJx2_ASAP7_75t_L g304 ( 
.A(n_282),
.B(n_277),
.C(n_275),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_304),
.B(n_279),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_305),
.A2(n_280),
.B1(n_291),
.B2(n_13),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_287),
.B(n_269),
.C(n_264),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_306),
.B(n_309),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_292),
.B(n_274),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_293),
.B(n_278),
.C(n_12),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_310),
.B(n_311),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_306),
.B(n_281),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_312),
.B(n_315),
.Y(n_325)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_314),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_297),
.B(n_286),
.Y(n_315)
);

INVx11_ASAP7_75t_L g316 ( 
.A(n_303),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_316),
.B(n_321),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_320),
.B(n_323),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_308),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_313),
.B(n_298),
.C(n_302),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_326),
.B(n_329),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_318),
.A2(n_301),
.B(n_310),
.Y(n_327)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_327),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_319),
.B(n_297),
.C(n_304),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_323),
.B(n_307),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_330),
.B(n_322),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_315),
.B(n_312),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_331),
.B(n_314),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_326),
.B(n_316),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_334),
.B(n_335),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_324),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_337),
.B(n_338),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_336),
.B(n_317),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_341),
.A2(n_334),
.B(n_328),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_342),
.B(n_325),
.C(n_329),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_343),
.B(n_325),
.C(n_339),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_344),
.A2(n_340),
.B1(n_333),
.B2(n_332),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_345),
.B(n_332),
.Y(n_346)
);


endmodule