module real_aes_8973_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_504;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_527;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_617;
wire n_552;
wire n_602;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_713;
wire n_288;
wire n_404;
wire n_598;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_717;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_175;
wire n_168;
wire n_241;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g260 ( .A1(n_0), .A2(n_261), .B(n_262), .C(n_265), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_1), .B(n_202), .Y(n_266) );
INVx1_ASAP7_75t_L g111 ( .A(n_2), .Y(n_111) );
NAND2xp5_ASAP7_75t_SL g238 ( .A(n_3), .B(n_172), .Y(n_238) );
A2O1A1Ixp33_ASAP7_75t_L g449 ( .A1(n_4), .A2(n_142), .B(n_145), .C(n_450), .Y(n_449) );
AOI21xp5_ASAP7_75t_L g489 ( .A1(n_5), .A2(n_162), .B(n_490), .Y(n_489) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_6), .A2(n_102), .B1(n_113), .B2(n_739), .Y(n_101) );
AOI21xp5_ASAP7_75t_L g192 ( .A1(n_7), .A2(n_162), .B(n_193), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_8), .B(n_202), .Y(n_496) );
AO21x2_ASAP7_75t_L g181 ( .A1(n_9), .A2(n_129), .B(n_182), .Y(n_181) );
AND2x6_ASAP7_75t_L g142 ( .A(n_10), .B(n_143), .Y(n_142) );
A2O1A1Ixp33_ASAP7_75t_L g144 ( .A1(n_11), .A2(n_142), .B(n_145), .C(n_148), .Y(n_144) );
OAI22xp5_ASAP7_75t_L g115 ( .A1(n_12), .A2(n_45), .B1(n_116), .B2(n_117), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_12), .Y(n_116) );
NOR2xp33_ASAP7_75t_L g112 ( .A(n_13), .B(n_41), .Y(n_112) );
INVx1_ASAP7_75t_L g466 ( .A(n_14), .Y(n_466) );
NAND2xp5_ASAP7_75t_SL g452 ( .A(n_15), .B(n_152), .Y(n_452) );
INVx1_ASAP7_75t_L g134 ( .A(n_16), .Y(n_134) );
NAND2xp5_ASAP7_75t_SL g188 ( .A(n_17), .B(n_172), .Y(n_188) );
A2O1A1Ixp33_ASAP7_75t_L g473 ( .A1(n_18), .A2(n_150), .B(n_474), .C(n_476), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_19), .B(n_202), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_20), .B(n_226), .Y(n_509) );
A2O1A1Ixp33_ASAP7_75t_L g221 ( .A1(n_21), .A2(n_145), .B(n_189), .C(n_222), .Y(n_221) );
A2O1A1Ixp33_ASAP7_75t_L g482 ( .A1(n_22), .A2(n_154), .B(n_264), .C(n_483), .Y(n_482) );
NAND2xp5_ASAP7_75t_SL g528 ( .A(n_23), .B(n_152), .Y(n_528) );
CKINVDCx20_ASAP7_75t_R g736 ( .A(n_24), .Y(n_736) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_25), .B(n_152), .Y(n_517) );
CKINVDCx16_ASAP7_75t_R g524 ( .A(n_26), .Y(n_524) );
INVx1_ASAP7_75t_L g516 ( .A(n_27), .Y(n_516) );
A2O1A1Ixp33_ASAP7_75t_L g184 ( .A1(n_28), .A2(n_145), .B(n_185), .C(n_189), .Y(n_184) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_29), .Y(n_141) );
CKINVDCx20_ASAP7_75t_R g448 ( .A(n_30), .Y(n_448) );
INVx1_ASAP7_75t_L g507 ( .A(n_31), .Y(n_507) );
AOI21xp5_ASAP7_75t_L g257 ( .A1(n_32), .A2(n_162), .B(n_258), .Y(n_257) );
INVx2_ASAP7_75t_L g140 ( .A(n_33), .Y(n_140) );
A2O1A1Ixp33_ASAP7_75t_L g209 ( .A1(n_34), .A2(n_164), .B(n_175), .C(n_210), .Y(n_209) );
CKINVDCx20_ASAP7_75t_R g455 ( .A(n_35), .Y(n_455) );
A2O1A1Ixp33_ASAP7_75t_L g492 ( .A1(n_36), .A2(n_264), .B(n_493), .C(n_495), .Y(n_492) );
INVxp67_ASAP7_75t_L g508 ( .A(n_37), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_38), .B(n_187), .Y(n_186) );
CKINVDCx14_ASAP7_75t_R g491 ( .A(n_39), .Y(n_491) );
A2O1A1Ixp33_ASAP7_75t_L g514 ( .A1(n_40), .A2(n_145), .B(n_189), .C(n_515), .Y(n_514) );
A2O1A1Ixp33_ASAP7_75t_L g463 ( .A1(n_42), .A2(n_265), .B(n_464), .C(n_465), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_43), .B(n_220), .Y(n_219) );
CKINVDCx20_ASAP7_75t_R g157 ( .A(n_44), .Y(n_157) );
INVx1_ASAP7_75t_L g117 ( .A(n_45), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_46), .B(n_172), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_47), .B(n_162), .Y(n_183) );
CKINVDCx20_ASAP7_75t_R g519 ( .A(n_48), .Y(n_519) );
CKINVDCx20_ASAP7_75t_R g504 ( .A(n_49), .Y(n_504) );
A2O1A1Ixp33_ASAP7_75t_L g163 ( .A1(n_50), .A2(n_164), .B(n_166), .C(n_175), .Y(n_163) );
INVx1_ASAP7_75t_L g263 ( .A(n_51), .Y(n_263) );
INVx1_ASAP7_75t_L g167 ( .A(n_52), .Y(n_167) );
INVx1_ASAP7_75t_L g481 ( .A(n_53), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_54), .B(n_162), .Y(n_161) );
OAI22xp5_ASAP7_75t_SL g728 ( .A1(n_55), .A2(n_59), .B1(n_729), .B2(n_730), .Y(n_728) );
CKINVDCx20_ASAP7_75t_R g730 ( .A(n_55), .Y(n_730) );
CKINVDCx20_ASAP7_75t_R g716 ( .A(n_56), .Y(n_716) );
CKINVDCx20_ASAP7_75t_R g229 ( .A(n_57), .Y(n_229) );
CKINVDCx14_ASAP7_75t_R g462 ( .A(n_58), .Y(n_462) );
CKINVDCx20_ASAP7_75t_R g729 ( .A(n_59), .Y(n_729) );
INVx1_ASAP7_75t_L g143 ( .A(n_60), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_61), .B(n_162), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_62), .B(n_202), .Y(n_201) );
A2O1A1Ixp33_ASAP7_75t_L g195 ( .A1(n_63), .A2(n_196), .B(n_198), .C(n_200), .Y(n_195) );
INVx1_ASAP7_75t_L g133 ( .A(n_64), .Y(n_133) );
INVx1_ASAP7_75t_SL g494 ( .A(n_65), .Y(n_494) );
CKINVDCx20_ASAP7_75t_R g723 ( .A(n_66), .Y(n_723) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_67), .B(n_172), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_68), .B(n_202), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_69), .B(n_150), .Y(n_149) );
INVx1_ASAP7_75t_L g527 ( .A(n_70), .Y(n_527) );
CKINVDCx16_ASAP7_75t_R g259 ( .A(n_71), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_72), .B(n_169), .Y(n_223) );
A2O1A1Ixp33_ASAP7_75t_L g235 ( .A1(n_73), .A2(n_145), .B(n_175), .C(n_236), .Y(n_235) );
CKINVDCx16_ASAP7_75t_R g194 ( .A(n_74), .Y(n_194) );
INVx1_ASAP7_75t_L g106 ( .A(n_75), .Y(n_106) );
AOI21xp5_ASAP7_75t_L g460 ( .A1(n_76), .A2(n_162), .B(n_461), .Y(n_460) );
CKINVDCx20_ASAP7_75t_R g530 ( .A(n_77), .Y(n_530) );
AOI21xp5_ASAP7_75t_L g470 ( .A1(n_78), .A2(n_162), .B(n_471), .Y(n_470) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_79), .A2(n_220), .B(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g472 ( .A(n_80), .Y(n_472) );
CKINVDCx16_ASAP7_75t_R g513 ( .A(n_81), .Y(n_513) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_82), .B(n_168), .Y(n_224) );
CKINVDCx20_ASAP7_75t_R g214 ( .A(n_83), .Y(n_214) );
AOI21xp5_ASAP7_75t_L g479 ( .A1(n_84), .A2(n_162), .B(n_480), .Y(n_479) );
INVx1_ASAP7_75t_L g475 ( .A(n_85), .Y(n_475) );
INVx2_ASAP7_75t_L g131 ( .A(n_86), .Y(n_131) );
INVx1_ASAP7_75t_L g451 ( .A(n_87), .Y(n_451) );
CKINVDCx20_ASAP7_75t_R g243 ( .A(n_88), .Y(n_243) );
NAND2xp5_ASAP7_75t_SL g151 ( .A(n_89), .B(n_152), .Y(n_151) );
OR2x2_ASAP7_75t_L g108 ( .A(n_90), .B(n_109), .Y(n_108) );
OR2x2_ASAP7_75t_L g438 ( .A(n_90), .B(n_110), .Y(n_438) );
INVx2_ASAP7_75t_L g708 ( .A(n_90), .Y(n_708) );
A2O1A1Ixp33_ASAP7_75t_L g525 ( .A1(n_91), .A2(n_145), .B(n_175), .C(n_526), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_92), .B(n_162), .Y(n_208) );
INVx1_ASAP7_75t_L g211 ( .A(n_93), .Y(n_211) );
INVxp67_ASAP7_75t_L g199 ( .A(n_94), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_95), .B(n_129), .Y(n_467) );
INVx2_ASAP7_75t_L g484 ( .A(n_96), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_97), .B(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g136 ( .A(n_98), .Y(n_136) );
INVx1_ASAP7_75t_L g237 ( .A(n_99), .Y(n_237) );
AND2x2_ASAP7_75t_L g178 ( .A(n_100), .B(n_177), .Y(n_178) );
CKINVDCx6p67_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
INVx1_ASAP7_75t_L g740 ( .A(n_103), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g103 ( .A(n_104), .B(n_107), .Y(n_103) );
INVx1_ASAP7_75t_SL g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_SL g107 ( .A(n_108), .Y(n_107) );
INVx1_ASAP7_75t_SL g732 ( .A(n_108), .Y(n_732) );
INVx1_ASAP7_75t_SL g738 ( .A(n_108), .Y(n_738) );
NOR2x2_ASAP7_75t_L g720 ( .A(n_109), .B(n_708), .Y(n_720) );
INVx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
OR2x2_ASAP7_75t_L g707 ( .A(n_110), .B(n_708), .Y(n_707) );
AND2x2_ASAP7_75t_L g110 ( .A(n_111), .B(n_112), .Y(n_110) );
AO221x1_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_721), .B1(n_724), .B2(n_733), .C(n_735), .Y(n_113) );
OAI222xp33_ASAP7_75t_SL g114 ( .A1(n_115), .A2(n_118), .B1(n_709), .B2(n_710), .C1(n_716), .C2(n_717), .Y(n_114) );
INVx1_ASAP7_75t_L g709 ( .A(n_115), .Y(n_709) );
INVxp67_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
OAI22xp5_ASAP7_75t_SL g119 ( .A1(n_120), .A2(n_436), .B1(n_439), .B2(n_705), .Y(n_119) );
INVx2_ASAP7_75t_L g713 ( .A(n_120), .Y(n_713) );
AOI22xp5_ASAP7_75t_L g726 ( .A1(n_120), .A2(n_713), .B1(n_727), .B2(n_728), .Y(n_726) );
OR3x1_ASAP7_75t_L g120 ( .A(n_121), .B(n_334), .C(n_399), .Y(n_120) );
NAND4xp25_ASAP7_75t_SL g121 ( .A(n_122), .B(n_275), .C(n_301), .D(n_324), .Y(n_121) );
AOI221xp5_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_203), .B1(n_244), .B2(n_251), .C(n_267), .Y(n_122) );
CKINVDCx14_ASAP7_75t_R g123 ( .A(n_124), .Y(n_123) );
OAI22xp5_ASAP7_75t_L g422 ( .A1(n_124), .A2(n_268), .B1(n_292), .B2(n_423), .Y(n_422) );
OR2x2_ASAP7_75t_L g124 ( .A(n_125), .B(n_179), .Y(n_124) );
INVx1_ASAP7_75t_SL g328 ( .A(n_125), .Y(n_328) );
OR2x2_ASAP7_75t_L g125 ( .A(n_126), .B(n_159), .Y(n_125) );
OR2x2_ASAP7_75t_L g249 ( .A(n_126), .B(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g270 ( .A(n_126), .B(n_180), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_126), .B(n_190), .Y(n_283) );
AND2x2_ASAP7_75t_L g300 ( .A(n_126), .B(n_159), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_126), .B(n_247), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_126), .B(n_299), .Y(n_411) );
NOR2xp33_ASAP7_75t_L g421 ( .A(n_126), .B(n_179), .Y(n_421) );
AOI211xp5_ASAP7_75t_SL g432 ( .A1(n_126), .A2(n_338), .B(n_433), .C(n_434), .Y(n_432) );
INVx5_ASAP7_75t_SL g126 ( .A(n_127), .Y(n_126) );
NAND2xp5_ASAP7_75t_SL g304 ( .A(n_127), .B(n_180), .Y(n_304) );
AND2x2_ASAP7_75t_L g307 ( .A(n_127), .B(n_181), .Y(n_307) );
OR2x2_ASAP7_75t_L g352 ( .A(n_127), .B(n_180), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_127), .B(n_190), .Y(n_361) );
AO21x2_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_135), .B(n_156), .Y(n_127) );
INVx3_ASAP7_75t_L g202 ( .A(n_128), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g213 ( .A(n_128), .B(n_214), .Y(n_213) );
AO21x2_ASAP7_75t_L g233 ( .A1(n_128), .A2(n_234), .B(n_242), .Y(n_233) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_128), .B(n_243), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g454 ( .A(n_128), .B(n_455), .Y(n_454) );
NOR2xp33_ASAP7_75t_L g518 ( .A(n_128), .B(n_519), .Y(n_518) );
AO21x2_ASAP7_75t_L g522 ( .A1(n_128), .A2(n_523), .B(n_529), .Y(n_522) );
INVx4_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
AOI21xp5_ASAP7_75t_L g182 ( .A1(n_129), .A2(n_183), .B(n_184), .Y(n_182) );
HB1xp67_ASAP7_75t_L g191 ( .A(n_129), .Y(n_191) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx1_ASAP7_75t_L g158 ( .A(n_130), .Y(n_158) );
AND2x2_ASAP7_75t_L g130 ( .A(n_131), .B(n_132), .Y(n_130) );
AND2x2_ASAP7_75t_SL g177 ( .A(n_131), .B(n_132), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_133), .B(n_134), .Y(n_132) );
OAI21xp5_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_137), .B(n_144), .Y(n_135) );
OAI21xp5_ASAP7_75t_L g447 ( .A1(n_137), .A2(n_448), .B(n_449), .Y(n_447) );
O2A1O1Ixp33_ASAP7_75t_L g512 ( .A1(n_137), .A2(n_177), .B(n_513), .C(n_514), .Y(n_512) );
OAI21xp5_ASAP7_75t_L g523 ( .A1(n_137), .A2(n_524), .B(n_525), .Y(n_523) );
NAND2x1p5_ASAP7_75t_L g137 ( .A(n_138), .B(n_142), .Y(n_137) );
AND2x4_ASAP7_75t_L g162 ( .A(n_138), .B(n_142), .Y(n_162) );
AND2x2_ASAP7_75t_L g138 ( .A(n_139), .B(n_141), .Y(n_138) );
INVx1_ASAP7_75t_L g200 ( .A(n_139), .Y(n_200) );
INVx1_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx2_ASAP7_75t_L g146 ( .A(n_140), .Y(n_146) );
INVx1_ASAP7_75t_L g155 ( .A(n_140), .Y(n_155) );
INVx1_ASAP7_75t_L g147 ( .A(n_141), .Y(n_147) );
INVx3_ASAP7_75t_L g150 ( .A(n_141), .Y(n_150) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_141), .Y(n_152) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_141), .Y(n_170) );
INVx1_ASAP7_75t_L g187 ( .A(n_141), .Y(n_187) );
INVx4_ASAP7_75t_SL g176 ( .A(n_142), .Y(n_176) );
BUFx3_ASAP7_75t_L g189 ( .A(n_142), .Y(n_189) );
INVx5_ASAP7_75t_L g165 ( .A(n_145), .Y(n_165) );
AND2x6_ASAP7_75t_L g145 ( .A(n_146), .B(n_147), .Y(n_145) );
BUFx3_ASAP7_75t_L g174 ( .A(n_146), .Y(n_174) );
BUFx6f_ASAP7_75t_L g240 ( .A(n_146), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_151), .B(n_153), .Y(n_148) );
INVx5_ASAP7_75t_L g172 ( .A(n_150), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g465 ( .A(n_150), .B(n_466), .Y(n_465) );
INVx4_ASAP7_75t_L g264 ( .A(n_152), .Y(n_264) );
INVx2_ASAP7_75t_L g464 ( .A(n_152), .Y(n_464) );
AOI21xp5_ASAP7_75t_L g185 ( .A1(n_153), .A2(n_186), .B(n_188), .Y(n_185) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx3_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
NOR2xp33_ASAP7_75t_L g156 ( .A(n_157), .B(n_158), .Y(n_156) );
INVx2_ASAP7_75t_L g501 ( .A(n_158), .Y(n_501) );
INVx5_ASAP7_75t_SL g250 ( .A(n_159), .Y(n_250) );
AND2x2_ASAP7_75t_L g269 ( .A(n_159), .B(n_270), .Y(n_269) );
NOR2xp33_ASAP7_75t_L g351 ( .A(n_159), .B(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g355 ( .A(n_159), .B(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g387 ( .A(n_159), .B(n_190), .Y(n_387) );
OR2x2_ASAP7_75t_L g393 ( .A(n_159), .B(n_283), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_159), .B(n_343), .Y(n_402) );
OR2x6_ASAP7_75t_L g159 ( .A(n_160), .B(n_178), .Y(n_159) );
AOI21xp5_ASAP7_75t_L g160 ( .A1(n_161), .A2(n_163), .B(n_177), .Y(n_160) );
BUFx2_ASAP7_75t_L g220 ( .A(n_162), .Y(n_220) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
O2A1O1Ixp33_ASAP7_75t_L g193 ( .A1(n_165), .A2(n_176), .B(n_194), .C(n_195), .Y(n_193) );
O2A1O1Ixp33_ASAP7_75t_SL g258 ( .A1(n_165), .A2(n_176), .B(n_259), .C(n_260), .Y(n_258) );
O2A1O1Ixp33_ASAP7_75t_SL g461 ( .A1(n_165), .A2(n_176), .B(n_462), .C(n_463), .Y(n_461) );
O2A1O1Ixp33_ASAP7_75t_SL g471 ( .A1(n_165), .A2(n_176), .B(n_472), .C(n_473), .Y(n_471) );
O2A1O1Ixp33_ASAP7_75t_SL g480 ( .A1(n_165), .A2(n_176), .B(n_481), .C(n_482), .Y(n_480) );
O2A1O1Ixp33_ASAP7_75t_L g490 ( .A1(n_165), .A2(n_176), .B(n_491), .C(n_492), .Y(n_490) );
O2A1O1Ixp33_ASAP7_75t_SL g503 ( .A1(n_165), .A2(n_176), .B(n_504), .C(n_505), .Y(n_503) );
O2A1O1Ixp33_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_168), .B(n_171), .C(n_173), .Y(n_166) );
O2A1O1Ixp33_ASAP7_75t_L g210 ( .A1(n_168), .A2(n_173), .B(n_211), .C(n_212), .Y(n_210) );
O2A1O1Ixp5_ASAP7_75t_L g450 ( .A1(n_168), .A2(n_451), .B(n_452), .C(n_453), .Y(n_450) );
O2A1O1Ixp33_ASAP7_75t_L g526 ( .A1(n_168), .A2(n_453), .B(n_527), .C(n_528), .Y(n_526) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx4_ASAP7_75t_L g197 ( .A(n_170), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g198 ( .A(n_172), .B(n_199), .Y(n_198) );
INVx2_ASAP7_75t_L g261 ( .A(n_172), .Y(n_261) );
OAI22xp33_ASAP7_75t_L g506 ( .A1(n_172), .A2(n_197), .B1(n_507), .B2(n_508), .Y(n_506) );
O2A1O1Ixp33_ASAP7_75t_L g515 ( .A1(n_172), .A2(n_225), .B(n_516), .C(n_517), .Y(n_515) );
HB1xp67_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx2_ASAP7_75t_L g265 ( .A(n_174), .Y(n_265) );
INVx1_ASAP7_75t_L g476 ( .A(n_174), .Y(n_476) );
INVx1_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_177), .A2(n_208), .B(n_209), .Y(n_207) );
INVx2_ASAP7_75t_L g227 ( .A(n_177), .Y(n_227) );
INVx1_ASAP7_75t_L g230 ( .A(n_177), .Y(n_230) );
OA21x2_ASAP7_75t_L g459 ( .A1(n_177), .A2(n_460), .B(n_467), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_180), .B(n_190), .Y(n_179) );
AND2x2_ASAP7_75t_L g284 ( .A(n_180), .B(n_250), .Y(n_284) );
INVx1_ASAP7_75t_SL g297 ( .A(n_180), .Y(n_297) );
OR2x2_ASAP7_75t_L g332 ( .A(n_180), .B(n_333), .Y(n_332) );
OR2x2_ASAP7_75t_L g338 ( .A(n_180), .B(n_190), .Y(n_338) );
AND2x2_ASAP7_75t_L g396 ( .A(n_180), .B(n_247), .Y(n_396) );
INVx2_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_181), .B(n_250), .Y(n_323) );
INVx3_ASAP7_75t_L g247 ( .A(n_190), .Y(n_247) );
OR2x2_ASAP7_75t_L g289 ( .A(n_190), .B(n_250), .Y(n_289) );
AND2x2_ASAP7_75t_L g299 ( .A(n_190), .B(n_297), .Y(n_299) );
HB1xp67_ASAP7_75t_L g347 ( .A(n_190), .Y(n_347) );
AND2x2_ASAP7_75t_L g356 ( .A(n_190), .B(n_270), .Y(n_356) );
OA21x2_ASAP7_75t_L g190 ( .A1(n_191), .A2(n_192), .B(n_201), .Y(n_190) );
OA21x2_ASAP7_75t_L g469 ( .A1(n_191), .A2(n_470), .B(n_477), .Y(n_469) );
OA21x2_ASAP7_75t_L g478 ( .A1(n_191), .A2(n_479), .B(n_485), .Y(n_478) );
OA21x2_ASAP7_75t_L g488 ( .A1(n_191), .A2(n_489), .B(n_496), .Y(n_488) );
O2A1O1Ixp33_ASAP7_75t_L g236 ( .A1(n_196), .A2(n_237), .B(n_238), .C(n_239), .Y(n_236) );
INVx1_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g474 ( .A(n_197), .B(n_475), .Y(n_474) );
NOR2xp33_ASAP7_75t_L g483 ( .A(n_197), .B(n_484), .Y(n_483) );
INVx2_ASAP7_75t_L g225 ( .A(n_200), .Y(n_225) );
NAND2xp5_ASAP7_75t_SL g505 ( .A(n_200), .B(n_506), .Y(n_505) );
OA21x2_ASAP7_75t_L g256 ( .A1(n_202), .A2(n_257), .B(n_266), .Y(n_256) );
AOI221xp5_ASAP7_75t_L g372 ( .A1(n_203), .A2(n_373), .B1(n_375), .B2(n_377), .C(n_380), .Y(n_372) );
INVx2_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
OR2x2_ASAP7_75t_L g204 ( .A(n_205), .B(n_215), .Y(n_204) );
AND2x2_ASAP7_75t_L g346 ( .A(n_205), .B(n_327), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_205), .B(n_405), .Y(n_409) );
OR2x2_ASAP7_75t_L g430 ( .A(n_205), .B(n_431), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_205), .B(n_435), .Y(n_434) );
BUFx2_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
INVx5_ASAP7_75t_L g277 ( .A(n_206), .Y(n_277) );
AND2x2_ASAP7_75t_L g354 ( .A(n_206), .B(n_217), .Y(n_354) );
AND2x2_ASAP7_75t_L g415 ( .A(n_206), .B(n_294), .Y(n_415) );
AND2x2_ASAP7_75t_L g428 ( .A(n_206), .B(n_247), .Y(n_428) );
OR2x6_ASAP7_75t_L g206 ( .A(n_207), .B(n_213), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_216), .B(n_231), .Y(n_215) );
AND2x4_ASAP7_75t_L g254 ( .A(n_216), .B(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g273 ( .A(n_216), .B(n_274), .Y(n_273) );
INVx2_ASAP7_75t_L g280 ( .A(n_216), .Y(n_280) );
AND2x2_ASAP7_75t_L g349 ( .A(n_216), .B(n_327), .Y(n_349) );
AND2x2_ASAP7_75t_L g359 ( .A(n_216), .B(n_277), .Y(n_359) );
HB1xp67_ASAP7_75t_L g367 ( .A(n_216), .Y(n_367) );
AND2x2_ASAP7_75t_L g379 ( .A(n_216), .B(n_256), .Y(n_379) );
NOR2xp33_ASAP7_75t_L g383 ( .A(n_216), .B(n_311), .Y(n_383) );
AND2x2_ASAP7_75t_L g420 ( .A(n_216), .B(n_415), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_216), .B(n_294), .Y(n_431) );
OR2x2_ASAP7_75t_L g433 ( .A(n_216), .B(n_369), .Y(n_433) );
INVx5_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
AND2x2_ASAP7_75t_L g319 ( .A(n_217), .B(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g329 ( .A(n_217), .B(n_274), .Y(n_329) );
AND2x2_ASAP7_75t_L g341 ( .A(n_217), .B(n_256), .Y(n_341) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_217), .Y(n_371) );
AND2x4_ASAP7_75t_L g405 ( .A(n_217), .B(n_255), .Y(n_405) );
OR2x6_ASAP7_75t_L g217 ( .A(n_218), .B(n_228), .Y(n_217) );
AOI21xp5_ASAP7_75t_SL g218 ( .A1(n_219), .A2(n_221), .B(n_226), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_223), .A2(n_224), .B(n_225), .Y(n_222) );
INVx1_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g529 ( .A(n_227), .B(n_530), .Y(n_529) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_229), .B(n_230), .Y(n_228) );
AO21x2_ASAP7_75t_L g446 ( .A1(n_230), .A2(n_447), .B(n_454), .Y(n_446) );
BUFx2_ASAP7_75t_L g253 ( .A(n_231), .Y(n_253) );
HB1xp67_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
INVx2_ASAP7_75t_L g294 ( .A(n_232), .Y(n_294) );
AND2x2_ASAP7_75t_L g327 ( .A(n_232), .B(n_256), .Y(n_327) );
INVx2_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
AND2x2_ASAP7_75t_L g274 ( .A(n_233), .B(n_256), .Y(n_274) );
BUFx2_ASAP7_75t_L g320 ( .A(n_233), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_235), .B(n_241), .Y(n_234) );
HB1xp67_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
INVx3_ASAP7_75t_L g495 ( .A(n_240), .Y(n_495) );
INVx1_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_246), .B(n_248), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_246), .B(n_328), .Y(n_407) );
INVx1_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_247), .B(n_270), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_247), .B(n_250), .Y(n_309) );
AND2x2_ASAP7_75t_L g364 ( .A(n_247), .B(n_300), .Y(n_364) );
AOI221xp5_ASAP7_75t_SL g301 ( .A1(n_248), .A2(n_302), .B1(n_310), .B2(n_312), .C(n_316), .Y(n_301) );
INVx2_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
OR2x2_ASAP7_75t_L g296 ( .A(n_249), .B(n_297), .Y(n_296) );
OR2x2_ASAP7_75t_L g337 ( .A(n_249), .B(n_338), .Y(n_337) );
OAI321xp33_ASAP7_75t_L g344 ( .A1(n_249), .A2(n_303), .A3(n_345), .B1(n_347), .B2(n_348), .C(n_350), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_250), .B(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_253), .B(n_254), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_253), .B(n_405), .Y(n_423) );
AND2x2_ASAP7_75t_L g310 ( .A(n_254), .B(n_311), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_254), .B(n_314), .Y(n_313) );
HB1xp67_ASAP7_75t_L g286 ( .A(n_255), .Y(n_286) );
AND2x2_ASAP7_75t_L g293 ( .A(n_255), .B(n_294), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_255), .B(n_368), .Y(n_398) );
INVx1_ASAP7_75t_L g435 ( .A(n_255), .Y(n_435) );
INVx2_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
NOR2xp33_ASAP7_75t_L g262 ( .A(n_263), .B(n_264), .Y(n_262) );
NOR2xp33_ASAP7_75t_L g493 ( .A(n_264), .B(n_494), .Y(n_493) );
INVx2_ASAP7_75t_L g453 ( .A(n_265), .Y(n_453) );
AOI21xp5_ASAP7_75t_L g267 ( .A1(n_268), .A2(n_271), .B(n_272), .Y(n_267) );
INVx1_ASAP7_75t_SL g268 ( .A(n_269), .Y(n_268) );
A2O1A1Ixp33_ASAP7_75t_L g427 ( .A1(n_269), .A2(n_379), .B(n_428), .C(n_429), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_270), .B(n_288), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_270), .B(n_308), .Y(n_374) );
INVx1_ASAP7_75t_SL g272 ( .A(n_273), .Y(n_272) );
INVx1_ASAP7_75t_L g317 ( .A(n_274), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_274), .B(n_277), .Y(n_331) );
NOR2xp33_ASAP7_75t_L g340 ( .A(n_274), .B(n_341), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_274), .B(n_359), .Y(n_358) );
AOI22xp33_ASAP7_75t_L g275 ( .A1(n_276), .A2(n_278), .B1(n_290), .B2(n_295), .Y(n_275) );
HB1xp67_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
OR2x2_ASAP7_75t_L g291 ( .A(n_277), .B(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g314 ( .A(n_277), .B(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g326 ( .A(n_277), .B(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_277), .B(n_320), .Y(n_362) );
OR2x2_ASAP7_75t_L g369 ( .A(n_277), .B(n_294), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_277), .B(n_379), .Y(n_378) );
AND2x2_ASAP7_75t_L g419 ( .A(n_277), .B(n_405), .Y(n_419) );
OAI22xp33_ASAP7_75t_L g278 ( .A1(n_279), .A2(n_281), .B1(n_285), .B2(n_287), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g325 ( .A(n_280), .B(n_326), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_282), .B(n_284), .Y(n_281) );
INVx1_ASAP7_75t_SL g282 ( .A(n_283), .Y(n_282) );
OAI22xp33_ASAP7_75t_L g365 ( .A1(n_283), .A2(n_298), .B1(n_366), .B2(n_370), .Y(n_365) );
INVx1_ASAP7_75t_L g413 ( .A(n_284), .Y(n_413) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AOI221xp5_ASAP7_75t_L g324 ( .A1(n_288), .A2(n_325), .B1(n_328), .B2(n_329), .C(n_330), .Y(n_324) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
OR2x2_ASAP7_75t_L g303 ( .A(n_289), .B(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_293), .B(n_359), .Y(n_391) );
HB1xp67_ASAP7_75t_L g311 ( .A(n_294), .Y(n_311) );
INVx1_ASAP7_75t_L g315 ( .A(n_294), .Y(n_315) );
NAND2xp33_ASAP7_75t_L g295 ( .A(n_296), .B(n_298), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_299), .B(n_300), .Y(n_298) );
INVx1_ASAP7_75t_L g333 ( .A(n_300), .Y(n_333) );
AND2x2_ASAP7_75t_L g342 ( .A(n_300), .B(n_343), .Y(n_342) );
NAND2xp33_ASAP7_75t_L g302 ( .A(n_303), .B(n_305), .Y(n_302) );
INVx2_ASAP7_75t_SL g305 ( .A(n_306), .Y(n_305) );
AND2x4_ASAP7_75t_L g306 ( .A(n_307), .B(n_308), .Y(n_306) );
AND2x2_ASAP7_75t_L g386 ( .A(n_307), .B(n_387), .Y(n_386) );
INVx2_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
AOI221xp5_ASAP7_75t_L g335 ( .A1(n_310), .A2(n_336), .B1(n_339), .B2(n_342), .C(n_344), .Y(n_335) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_314), .B(n_371), .Y(n_370) );
AOI21xp33_ASAP7_75t_SL g316 ( .A1(n_317), .A2(n_318), .B(n_321), .Y(n_316) );
INVx2_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
CKINVDCx16_ASAP7_75t_R g418 ( .A(n_321), .Y(n_418) );
OR2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
OR2x2_ASAP7_75t_L g360 ( .A(n_323), .B(n_361), .Y(n_360) );
INVx1_ASAP7_75t_SL g381 ( .A(n_326), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_326), .B(n_386), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_329), .B(n_351), .Y(n_350) );
NOR2xp33_ASAP7_75t_L g330 ( .A(n_331), .B(n_332), .Y(n_330) );
NAND4xp25_ASAP7_75t_L g334 ( .A(n_335), .B(n_353), .C(n_372), .D(n_385), .Y(n_334) );
INVx1_ASAP7_75t_SL g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_SL g343 ( .A(n_338), .Y(n_343) );
INVxp67_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
OR2x2_ASAP7_75t_L g376 ( .A(n_347), .B(n_352), .Y(n_376) );
INVxp67_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
AOI211xp5_ASAP7_75t_L g353 ( .A1(n_354), .A2(n_355), .B(n_357), .C(n_365), .Y(n_353) );
AOI211xp5_ASAP7_75t_L g424 ( .A1(n_355), .A2(n_397), .B(n_425), .C(n_432), .Y(n_424) );
INVx1_ASAP7_75t_SL g384 ( .A(n_356), .Y(n_384) );
OAI22xp5_ASAP7_75t_L g357 ( .A1(n_358), .A2(n_360), .B1(n_362), .B2(n_363), .Y(n_357) );
INVx1_ASAP7_75t_L g388 ( .A(n_362), .Y(n_388) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_367), .B(n_368), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_368), .B(n_405), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_368), .B(n_379), .Y(n_412) );
INVx2_ASAP7_75t_SL g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_SL g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g389 ( .A(n_379), .Y(n_389) );
AOI21xp33_ASAP7_75t_L g380 ( .A1(n_381), .A2(n_382), .B(n_384), .Y(n_380) );
INVxp33_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
AOI322xp5_ASAP7_75t_L g385 ( .A1(n_386), .A2(n_388), .A3(n_389), .B1(n_390), .B2(n_392), .C1(n_394), .C2(n_397), .Y(n_385) );
INVxp67_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
NAND3xp33_ASAP7_75t_SL g399 ( .A(n_400), .B(n_417), .C(n_424), .Y(n_399) );
AOI221xp5_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_403), .B1(n_406), .B2(n_408), .C(n_410), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_SL g416 ( .A(n_405), .Y(n_416) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVxp67_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
OAI22xp33_ASAP7_75t_L g410 ( .A1(n_411), .A2(n_412), .B1(n_413), .B2(n_414), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_415), .B(n_416), .Y(n_414) );
AOI221xp5_ASAP7_75t_L g417 ( .A1(n_418), .A2(n_419), .B1(n_420), .B2(n_421), .C(n_422), .Y(n_417) );
NAND2xp33_ASAP7_75t_L g425 ( .A(n_426), .B(n_427), .Y(n_425) );
INVxp67_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx2_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx2_ASAP7_75t_L g712 ( .A(n_437), .Y(n_712) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx2_ASAP7_75t_L g714 ( .A(n_439), .Y(n_714) );
OR2x2_ASAP7_75t_SL g439 ( .A(n_440), .B(n_660), .Y(n_439) );
NAND5xp2_ASAP7_75t_L g440 ( .A(n_441), .B(n_572), .C(n_610), .D(n_631), .E(n_648), .Y(n_440) );
NOR3xp33_ASAP7_75t_L g441 ( .A(n_442), .B(n_544), .C(n_565), .Y(n_441) );
OAI221xp5_ASAP7_75t_SL g442 ( .A1(n_443), .A2(n_486), .B1(n_510), .B2(n_531), .C(n_535), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_444), .B(n_456), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_445), .B(n_533), .Y(n_552) );
OR2x2_ASAP7_75t_L g579 ( .A(n_445), .B(n_469), .Y(n_579) );
AND2x2_ASAP7_75t_L g593 ( .A(n_445), .B(n_469), .Y(n_593) );
NOR2xp33_ASAP7_75t_L g607 ( .A(n_445), .B(n_459), .Y(n_607) );
AND2x2_ASAP7_75t_L g645 ( .A(n_445), .B(n_609), .Y(n_645) );
AND2x2_ASAP7_75t_L g674 ( .A(n_445), .B(n_584), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_445), .B(n_556), .Y(n_691) );
INVx4_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
AND2x2_ASAP7_75t_L g571 ( .A(n_446), .B(n_468), .Y(n_571) );
BUFx3_ASAP7_75t_L g596 ( .A(n_446), .Y(n_596) );
AND2x2_ASAP7_75t_L g625 ( .A(n_446), .B(n_469), .Y(n_625) );
AND3x2_ASAP7_75t_L g638 ( .A(n_446), .B(n_639), .C(n_640), .Y(n_638) );
INVx1_ASAP7_75t_L g561 ( .A(n_456), .Y(n_561) );
AND2x2_ASAP7_75t_L g456 ( .A(n_457), .B(n_468), .Y(n_456) );
AOI32xp33_ASAP7_75t_L g616 ( .A1(n_457), .A2(n_568), .A3(n_617), .B1(n_620), .B2(n_621), .Y(n_616) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
AND2x2_ASAP7_75t_L g543 ( .A(n_458), .B(n_468), .Y(n_543) );
NAND2xp5_ASAP7_75t_SL g614 ( .A(n_458), .B(n_571), .Y(n_614) );
AND2x2_ASAP7_75t_L g621 ( .A(n_458), .B(n_593), .Y(n_621) );
OR2x2_ASAP7_75t_L g627 ( .A(n_458), .B(n_628), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_458), .B(n_582), .Y(n_652) );
OR2x2_ASAP7_75t_L g670 ( .A(n_458), .B(n_498), .Y(n_670) );
BUFx3_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
AND2x2_ASAP7_75t_L g534 ( .A(n_459), .B(n_478), .Y(n_534) );
INVx2_ASAP7_75t_L g556 ( .A(n_459), .Y(n_556) );
OR2x2_ASAP7_75t_L g578 ( .A(n_459), .B(n_478), .Y(n_578) );
AND2x2_ASAP7_75t_L g583 ( .A(n_459), .B(n_584), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_459), .B(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_L g639 ( .A(n_459), .B(n_533), .Y(n_639) );
INVx1_ASAP7_75t_SL g690 ( .A(n_468), .Y(n_690) );
AND2x2_ASAP7_75t_L g468 ( .A(n_469), .B(n_478), .Y(n_468) );
INVx1_ASAP7_75t_SL g533 ( .A(n_469), .Y(n_533) );
HB1xp67_ASAP7_75t_L g582 ( .A(n_469), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_469), .B(n_619), .Y(n_618) );
NAND3xp33_ASAP7_75t_L g685 ( .A(n_469), .B(n_556), .C(n_674), .Y(n_685) );
INVx2_ASAP7_75t_L g584 ( .A(n_478), .Y(n_584) );
HB1xp67_ASAP7_75t_L g598 ( .A(n_478), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_487), .B(n_497), .Y(n_486) );
INVx1_ASAP7_75t_L g620 ( .A(n_487), .Y(n_620) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
AND2x2_ASAP7_75t_L g538 ( .A(n_488), .B(n_521), .Y(n_538) );
INVx2_ASAP7_75t_L g555 ( .A(n_488), .Y(n_555) );
AND2x2_ASAP7_75t_L g560 ( .A(n_488), .B(n_522), .Y(n_560) );
AND2x2_ASAP7_75t_L g575 ( .A(n_488), .B(n_511), .Y(n_575) );
AND2x2_ASAP7_75t_L g587 ( .A(n_488), .B(n_559), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_497), .B(n_603), .Y(n_602) );
NAND2x1p5_ASAP7_75t_L g659 ( .A(n_497), .B(n_560), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_497), .B(n_679), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_497), .B(n_554), .Y(n_682) );
BUFx3_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
OR2x2_ASAP7_75t_L g520 ( .A(n_498), .B(n_521), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_498), .B(n_538), .Y(n_537) );
AND2x2_ASAP7_75t_L g564 ( .A(n_498), .B(n_511), .Y(n_564) );
AND2x2_ASAP7_75t_L g590 ( .A(n_498), .B(n_521), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_498), .B(n_630), .Y(n_629) );
OA21x2_ASAP7_75t_L g498 ( .A1(n_499), .A2(n_502), .B(n_509), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
AO21x2_ASAP7_75t_L g548 ( .A1(n_500), .A2(n_549), .B(n_550), .Y(n_548) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g549 ( .A(n_502), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_509), .Y(n_550) );
OR2x2_ASAP7_75t_L g510 ( .A(n_511), .B(n_520), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_511), .B(n_541), .Y(n_540) );
AND2x4_ASAP7_75t_L g554 ( .A(n_511), .B(n_555), .Y(n_554) );
INVx3_ASAP7_75t_SL g559 ( .A(n_511), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_511), .B(n_546), .Y(n_612) );
OR2x2_ASAP7_75t_L g622 ( .A(n_511), .B(n_548), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_511), .B(n_590), .Y(n_650) );
OR2x2_ASAP7_75t_L g680 ( .A(n_511), .B(n_521), .Y(n_680) );
AND2x2_ASAP7_75t_L g684 ( .A(n_511), .B(n_522), .Y(n_684) );
NAND2xp5_ASAP7_75t_SL g697 ( .A(n_511), .B(n_560), .Y(n_697) );
AND2x2_ASAP7_75t_L g704 ( .A(n_511), .B(n_586), .Y(n_704) );
OR2x6_ASAP7_75t_L g511 ( .A(n_512), .B(n_518), .Y(n_511) );
INVx1_ASAP7_75t_SL g647 ( .A(n_520), .Y(n_647) );
AND2x2_ASAP7_75t_L g586 ( .A(n_521), .B(n_548), .Y(n_586) );
AND2x2_ASAP7_75t_L g600 ( .A(n_521), .B(n_555), .Y(n_600) );
AND2x2_ASAP7_75t_L g603 ( .A(n_521), .B(n_559), .Y(n_603) );
INVx1_ASAP7_75t_L g630 ( .A(n_521), .Y(n_630) );
INVx2_ASAP7_75t_SL g521 ( .A(n_522), .Y(n_521) );
BUFx2_ASAP7_75t_L g542 ( .A(n_522), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_532), .B(n_534), .Y(n_531) );
A2O1A1Ixp33_ASAP7_75t_L g701 ( .A1(n_532), .A2(n_578), .B(n_702), .C(n_703), .Y(n_701) );
HB1xp67_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
AND2x2_ASAP7_75t_L g608 ( .A(n_533), .B(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_534), .B(n_551), .Y(n_566) );
AND2x2_ASAP7_75t_L g592 ( .A(n_534), .B(n_593), .Y(n_592) );
OAI21xp5_ASAP7_75t_SL g535 ( .A1(n_536), .A2(n_539), .B(n_543), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
NOR2xp33_ASAP7_75t_L g636 ( .A(n_537), .B(n_637), .Y(n_636) );
AND2x2_ASAP7_75t_L g563 ( .A(n_538), .B(n_564), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_538), .B(n_559), .Y(n_604) );
AND2x2_ASAP7_75t_L g695 ( .A(n_538), .B(n_546), .Y(n_695) );
INVxp67_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
AND2x2_ASAP7_75t_L g568 ( .A(n_542), .B(n_555), .Y(n_568) );
OR2x2_ASAP7_75t_L g569 ( .A(n_542), .B(n_553), .Y(n_569) );
OAI322xp33_ASAP7_75t_L g544 ( .A1(n_545), .A2(n_552), .A3(n_553), .B1(n_556), .B2(n_557), .C1(n_561), .C2(n_562), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_546), .B(n_551), .Y(n_545) );
AND2x2_ASAP7_75t_L g656 ( .A(n_546), .B(n_568), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_546), .B(n_620), .Y(n_702) );
INVx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx1_ASAP7_75t_SL g547 ( .A(n_548), .Y(n_547) );
AND2x2_ASAP7_75t_L g599 ( .A(n_548), .B(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
OR2x2_ASAP7_75t_L g665 ( .A(n_552), .B(n_578), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_553), .B(n_647), .Y(n_646) );
INVx3_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_554), .B(n_586), .Y(n_643) );
AND2x2_ASAP7_75t_L g589 ( .A(n_555), .B(n_559), .Y(n_589) );
AND2x2_ASAP7_75t_L g597 ( .A(n_556), .B(n_598), .Y(n_597) );
A2O1A1Ixp33_ASAP7_75t_L g694 ( .A1(n_556), .A2(n_635), .B(n_695), .C(n_696), .Y(n_694) );
AOI21xp33_ASAP7_75t_L g667 ( .A1(n_557), .A2(n_570), .B(n_668), .Y(n_667) );
INVx1_ASAP7_75t_SL g557 ( .A(n_558), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_559), .B(n_560), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_559), .B(n_586), .Y(n_626) );
AND2x2_ASAP7_75t_L g632 ( .A(n_559), .B(n_600), .Y(n_632) );
AND2x2_ASAP7_75t_L g666 ( .A(n_559), .B(n_568), .Y(n_666) );
NOR2xp33_ASAP7_75t_L g574 ( .A(n_560), .B(n_575), .Y(n_574) );
INVx2_ASAP7_75t_SL g676 ( .A(n_560), .Y(n_676) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
AOI22xp5_ASAP7_75t_L g591 ( .A1(n_564), .A2(n_592), .B1(n_594), .B2(n_599), .Y(n_591) );
OAI22xp5_ASAP7_75t_SL g565 ( .A1(n_566), .A2(n_567), .B1(n_569), .B2(n_570), .Y(n_565) );
OAI22xp33_ASAP7_75t_L g601 ( .A1(n_566), .A2(n_602), .B1(n_604), .B2(n_605), .Y(n_601) );
INVxp67_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx1_ASAP7_75t_SL g570 ( .A(n_571), .Y(n_570) );
AOI221xp5_ASAP7_75t_L g672 ( .A1(n_571), .A2(n_673), .B1(n_675), .B2(n_677), .C(n_681), .Y(n_672) );
AOI211xp5_ASAP7_75t_L g572 ( .A1(n_573), .A2(n_576), .B(n_580), .C(n_601), .Y(n_572) );
INVxp67_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
OR2x2_ASAP7_75t_L g577 ( .A(n_578), .B(n_579), .Y(n_577) );
OR2x2_ASAP7_75t_L g642 ( .A(n_578), .B(n_595), .Y(n_642) );
INVx1_ASAP7_75t_L g693 ( .A(n_578), .Y(n_693) );
OAI221xp5_ASAP7_75t_L g580 ( .A1(n_579), .A2(n_581), .B1(n_585), .B2(n_588), .C(n_591), .Y(n_580) );
INVx2_ASAP7_75t_SL g635 ( .A(n_579), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_582), .B(n_583), .Y(n_581) );
INVx1_ASAP7_75t_L g700 ( .A(n_582), .Y(n_700) );
AND2x2_ASAP7_75t_L g624 ( .A(n_583), .B(n_625), .Y(n_624) );
INVx2_ASAP7_75t_L g609 ( .A(n_584), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_586), .B(n_587), .Y(n_585) );
INVx1_ASAP7_75t_L g671 ( .A(n_587), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .Y(n_588) );
AND2x2_ASAP7_75t_L g594 ( .A(n_595), .B(n_597), .Y(n_594) );
NOR2xp33_ASAP7_75t_L g696 ( .A(n_595), .B(n_697), .Y(n_696) );
CKINVDCx16_ASAP7_75t_R g595 ( .A(n_596), .Y(n_595) );
INVxp67_ASAP7_75t_L g640 ( .A(n_598), .Y(n_640) );
O2A1O1Ixp33_ASAP7_75t_L g610 ( .A1(n_599), .A2(n_611), .B(n_613), .C(n_615), .Y(n_610) );
INVx1_ASAP7_75t_L g688 ( .A(n_602), .Y(n_688) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
NOR2xp33_ASAP7_75t_L g663 ( .A(n_606), .B(n_664), .Y(n_663) );
AND2x2_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .Y(n_606) );
INVx2_ASAP7_75t_L g619 ( .A(n_609), .Y(n_619) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
OAI222xp33_ASAP7_75t_L g615 ( .A1(n_616), .A2(n_622), .B1(n_623), .B2(n_626), .C1(n_627), .C2(n_629), .Y(n_615) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_SL g655 ( .A(n_619), .Y(n_655) );
NOR2xp33_ASAP7_75t_L g675 ( .A(n_622), .B(n_676), .Y(n_675) );
NAND2xp33_ASAP7_75t_SL g653 ( .A(n_623), .B(n_654), .Y(n_653) );
INVx1_ASAP7_75t_SL g623 ( .A(n_624), .Y(n_623) );
INVx1_ASAP7_75t_SL g628 ( .A(n_625), .Y(n_628) );
AND2x2_ASAP7_75t_L g692 ( .A(n_625), .B(n_693), .Y(n_692) );
OR2x2_ASAP7_75t_L g658 ( .A(n_628), .B(n_655), .Y(n_658) );
INVx1_ASAP7_75t_L g687 ( .A(n_629), .Y(n_687) );
AOI211xp5_ASAP7_75t_L g631 ( .A1(n_632), .A2(n_633), .B(n_636), .C(n_641), .Y(n_631) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_635), .B(n_655), .Y(n_654) );
INVx2_ASAP7_75t_SL g637 ( .A(n_638), .Y(n_637) );
AOI322xp5_ASAP7_75t_L g686 ( .A1(n_638), .A2(n_666), .A3(n_671), .B1(n_687), .B2(n_688), .C1(n_689), .C2(n_692), .Y(n_686) );
AND2x2_ASAP7_75t_L g673 ( .A(n_639), .B(n_674), .Y(n_673) );
OAI22xp33_ASAP7_75t_L g641 ( .A1(n_642), .A2(n_643), .B1(n_644), .B2(n_646), .Y(n_641) );
INVxp33_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
AOI221xp5_ASAP7_75t_L g648 ( .A1(n_649), .A2(n_651), .B1(n_653), .B2(n_656), .C(n_657), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
NOR2xp33_ASAP7_75t_L g657 ( .A(n_658), .B(n_659), .Y(n_657) );
NAND5xp2_ASAP7_75t_L g660 ( .A(n_661), .B(n_672), .C(n_686), .D(n_694), .E(n_698), .Y(n_660) );
AOI21xp5_ASAP7_75t_L g661 ( .A1(n_662), .A2(n_666), .B(n_667), .Y(n_661) );
INVxp67_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx2_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVxp33_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
NOR2xp33_ASAP7_75t_L g669 ( .A(n_670), .B(n_671), .Y(n_669) );
A2O1A1Ixp33_ASAP7_75t_L g698 ( .A1(n_674), .A2(n_699), .B(n_700), .C(n_701), .Y(n_698) );
AOI31xp33_ASAP7_75t_L g681 ( .A1(n_676), .A2(n_682), .A3(n_683), .B(n_685), .Y(n_681) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
NOR2xp33_ASAP7_75t_L g689 ( .A(n_690), .B(n_691), .Y(n_689) );
INVx1_ASAP7_75t_L g699 ( .A(n_697), .Y(n_699) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx2_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx2_ASAP7_75t_L g715 ( .A(n_706), .Y(n_715) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVxp67_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
OAI22x1_ASAP7_75t_SL g711 ( .A1(n_712), .A2(n_713), .B1(n_714), .B2(n_715), .Y(n_711) );
INVx1_ASAP7_75t_SL g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx2_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
BUFx2_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx2_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g734 ( .A(n_723), .Y(n_734) );
INVxp67_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
NAND2xp5_ASAP7_75t_SL g725 ( .A(n_726), .B(n_731), .Y(n_725) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_SL g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
NOR2xp33_ASAP7_75t_L g735 ( .A(n_736), .B(n_737), .Y(n_735) );
INVx1_ASAP7_75t_SL g737 ( .A(n_738), .Y(n_737) );
INVx2_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
endmodule