module fake_jpeg_14107_n_59 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_59);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_59;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_51;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_15;

INVx8_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_8),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_SL g13 ( 
.A(n_7),
.B(n_5),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_13),
.B(n_0),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_18),
.B(n_19),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_13),
.B(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_20),
.B(n_21),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_15),
.B(n_3),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_24),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_23),
.Y(n_30)
);

INVx2_ASAP7_75t_SL g24 ( 
.A(n_10),
.Y(n_24)
);

OA22x2_ASAP7_75t_L g28 ( 
.A1(n_21),
.A2(n_11),
.B1(n_9),
.B2(n_12),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_28),
.A2(n_29),
.B1(n_14),
.B2(n_17),
.Y(n_37)
);

A2O1A1Ixp33_ASAP7_75t_SL g29 ( 
.A1(n_21),
.A2(n_11),
.B(n_0),
.C(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_24),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_16),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_25),
.A2(n_23),
.B1(n_24),
.B2(n_20),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_32),
.A2(n_34),
.B1(n_30),
.B2(n_14),
.Y(n_41)
);

AND2x2_ASAP7_75t_SL g33 ( 
.A(n_28),
.B(n_23),
.Y(n_33)
);

XOR2xp5_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_29),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_30),
.A2(n_14),
.B1(n_17),
.B2(n_16),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_15),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_36),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_37),
.A2(n_4),
.B(n_6),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_26),
.A2(n_18),
.B(n_5),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_4),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_41),
.Y(n_47)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_44),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_43),
.B(n_35),
.C(n_33),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_45),
.B(n_39),
.C(n_42),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_41),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_48),
.B(n_33),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_50),
.B(n_51),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_46),
.B(n_6),
.Y(n_52)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_52),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_53),
.A2(n_47),
.B(n_49),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_55),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_54),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_57),
.A2(n_47),
.B1(n_56),
.B2(n_37),
.Y(n_58)
);

BUFx24_ASAP7_75t_SL g59 ( 
.A(n_58),
.Y(n_59)
);


endmodule