module real_aes_3117_n_105 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_104, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_105);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_104;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_105;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_980;
wire n_618;
wire n_800;
wire n_778;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_977;
wire n_943;
wire n_287;
wire n_635;
wire n_357;
wire n_503;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_905;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_979;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_852;
wire n_766;
wire n_974;
wire n_132;
wire n_919;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_923;
wire n_894;
wire n_952;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_937;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_963;
wire n_865;
wire n_666;
wire n_320;
wire n_537;
wire n_551;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_983;
wire n_767;
wire n_138;
wire n_696;
wire n_889;
wire n_955;
wire n_975;
wire n_704;
wire n_941;
wire n_379;
wire n_453;
wire n_374;
wire n_647;
wire n_235;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_958;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_961;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_953;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_966;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_356;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_892;
wire n_495;
wire n_370;
wire n_938;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_935;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_951;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_981;
wire n_976;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_906;
wire n_477;
wire n_515;
wire n_230;
wire n_984;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_962;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_298;
wire n_523;
wire n_909;
wire n_439;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_960;
wire n_164;
wire n_671;
wire n_973;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_950;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_236;
wire n_278;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_936;
wire n_610;
wire n_581;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_940;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_142;
wire n_947;
wire n_970;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_964;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_913;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_917;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_985;
wire n_777;
wire n_488;
wire n_501;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_957;
wire n_296;
wire n_702;
wire n_954;
wire n_969;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_945;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_649;
wire n_193;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_397;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_915;
wire n_851;
wire n_133;
wire n_934;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_927;
wire n_965;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_972;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_291;
wire n_978;
wire n_907;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_939;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_155;
wire n_928;
wire n_243;
wire n_899;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_926;
wire n_922;
wire n_149;
wire n_942;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_134;
wire n_946;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_982;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_836;
wire n_888;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_929;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_949;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_967;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_921;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_968;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
INVx1_ASAP7_75t_L g640 ( .A(n_0), .Y(n_640) );
INVx1_ASAP7_75t_L g292 ( .A(n_1), .Y(n_292) );
AOI22xp5_ASAP7_75t_L g200 ( .A1(n_2), .A2(n_19), .B1(n_184), .B2(n_191), .Y(n_200) );
OAI22xp5_ASAP7_75t_SL g938 ( .A1(n_3), .A2(n_101), .B1(n_939), .B2(n_940), .Y(n_938) );
INVx1_ASAP7_75t_L g939 ( .A(n_3), .Y(n_939) );
AOI22xp5_ASAP7_75t_L g935 ( .A1(n_4), .A2(n_936), .B1(n_937), .B2(n_938), .Y(n_935) );
CKINVDCx5p33_ASAP7_75t_R g936 ( .A(n_4), .Y(n_936) );
INVx2_ASAP7_75t_L g169 ( .A(n_5), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_6), .B(n_563), .Y(n_580) );
INVx1_ASAP7_75t_SL g249 ( .A(n_7), .Y(n_249) );
BUFx2_ASAP7_75t_L g112 ( .A(n_8), .Y(n_112) );
INVx1_ASAP7_75t_L g124 ( .A(n_8), .Y(n_124) );
INVx1_ASAP7_75t_L g548 ( .A(n_8), .Y(n_548) );
INVxp67_ASAP7_75t_L g953 ( .A(n_8), .Y(n_953) );
NAND2xp5_ASAP7_75t_SL g581 ( .A(n_9), .B(n_264), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g678 ( .A1(n_10), .A2(n_40), .B1(n_594), .B2(n_679), .Y(n_678) );
AOI22xp5_ASAP7_75t_L g662 ( .A1(n_11), .A2(n_47), .B1(n_189), .B2(n_607), .Y(n_662) );
AOI22xp5_ASAP7_75t_L g654 ( .A1(n_12), .A2(n_71), .B1(n_648), .B2(n_649), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_13), .B(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_14), .B(n_268), .Y(n_267) );
INVx1_ASAP7_75t_L g635 ( .A(n_15), .Y(n_635) );
AOI22xp33_ASAP7_75t_L g262 ( .A1(n_16), .A2(n_58), .B1(n_263), .B2(n_264), .Y(n_262) );
INVx1_ASAP7_75t_L g638 ( .A(n_17), .Y(n_638) );
OA21x2_ASAP7_75t_L g148 ( .A1(n_18), .A2(n_75), .B(n_149), .Y(n_148) );
OA21x2_ASAP7_75t_L g209 ( .A1(n_18), .A2(n_75), .B(n_149), .Y(n_209) );
AOI22xp5_ASAP7_75t_L g647 ( .A1(n_20), .A2(n_73), .B1(n_648), .B2(n_649), .Y(n_647) );
NOR2xp33_ASAP7_75t_L g316 ( .A(n_21), .B(n_165), .Y(n_316) );
AOI22xp5_ASAP7_75t_L g151 ( .A1(n_22), .A2(n_85), .B1(n_152), .B2(n_155), .Y(n_151) );
INVx2_ASAP7_75t_L g196 ( .A(n_23), .Y(n_196) );
INVx1_ASAP7_75t_L g632 ( .A(n_24), .Y(n_632) );
AOI22xp5_ASAP7_75t_L g201 ( .A1(n_25), .A2(n_29), .B1(n_202), .B2(n_204), .Y(n_201) );
BUFx3_ASAP7_75t_L g957 ( .A(n_26), .Y(n_957) );
O2A1O1Ixp5_ASAP7_75t_L g188 ( .A1(n_27), .A2(n_189), .B(n_190), .C(n_193), .Y(n_188) );
AOI22xp33_ASAP7_75t_L g161 ( .A1(n_28), .A2(n_67), .B1(n_162), .B2(n_164), .Y(n_161) );
CKINVDCx5p33_ASAP7_75t_R g235 ( .A(n_30), .Y(n_235) );
AO22x1_ASAP7_75t_L g577 ( .A1(n_31), .A2(n_83), .B1(n_254), .B2(n_578), .Y(n_577) );
CKINVDCx5p33_ASAP7_75t_R g597 ( .A(n_32), .Y(n_597) );
AND2x2_ASAP7_75t_L g606 ( .A(n_33), .B(n_607), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_34), .B(n_254), .Y(n_601) );
AOI22xp5_ASAP7_75t_L g270 ( .A1(n_35), .A2(n_86), .B1(n_271), .B2(n_273), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_36), .B(n_84), .Y(n_115) );
INVx1_ASAP7_75t_L g128 ( .A(n_36), .Y(n_128) );
INVx1_ASAP7_75t_L g181 ( .A(n_37), .Y(n_181) );
AOI22x1_ASAP7_75t_L g664 ( .A1(n_38), .A2(n_102), .B1(n_648), .B2(n_665), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_39), .B(n_667), .Y(n_680) );
AND2x2_ASAP7_75t_L g113 ( .A(n_41), .B(n_114), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_42), .B(n_177), .Y(n_287) );
INVx2_ASAP7_75t_L g192 ( .A(n_43), .Y(n_192) );
CKINVDCx5p33_ASAP7_75t_R g237 ( .A(n_44), .Y(n_237) );
XNOR2x1_ASAP7_75t_L g974 ( .A(n_45), .B(n_975), .Y(n_974) );
NAND2xp5_ASAP7_75t_SL g615 ( .A(n_46), .B(n_561), .Y(n_615) );
INVx2_ASAP7_75t_L g315 ( .A(n_48), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g949 ( .A(n_49), .B(n_950), .Y(n_949) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_50), .B(n_285), .Y(n_284) );
INVx1_ASAP7_75t_SL g253 ( .A(n_51), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_52), .B(n_204), .Y(n_565) );
INVx1_ASAP7_75t_L g230 ( .A(n_53), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_54), .B(n_183), .Y(n_600) );
OAI22xp5_ASAP7_75t_L g978 ( .A1(n_55), .A2(n_642), .B1(n_979), .B2(n_980), .Y(n_978) );
INVx1_ASAP7_75t_L g979 ( .A(n_55), .Y(n_979) );
INVx1_ASAP7_75t_L g149 ( .A(n_56), .Y(n_149) );
AND2x2_ASAP7_75t_L g985 ( .A(n_57), .B(n_986), .Y(n_985) );
AND2x4_ASAP7_75t_L g143 ( .A(n_59), .B(n_144), .Y(n_143) );
AND2x4_ASAP7_75t_L g186 ( .A(n_59), .B(n_144), .Y(n_186) );
INVx1_ASAP7_75t_L g258 ( .A(n_60), .Y(n_258) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_61), .Y(n_160) );
INVx2_ASAP7_75t_L g651 ( .A(n_62), .Y(n_651) );
AOI22xp33_ASAP7_75t_L g675 ( .A1(n_63), .A2(n_78), .B1(n_594), .B2(n_665), .Y(n_675) );
CKINVDCx5p33_ASAP7_75t_R g945 ( .A(n_64), .Y(n_945) );
CKINVDCx14_ASAP7_75t_R g584 ( .A(n_65), .Y(n_584) );
AND2x2_ASAP7_75t_L g613 ( .A(n_66), .B(n_254), .Y(n_613) );
NOR2xp33_ASAP7_75t_L g319 ( .A(n_68), .B(n_251), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_69), .B(n_285), .Y(n_566) );
OAI22x1_ASAP7_75t_SL g976 ( .A1(n_70), .A2(n_93), .B1(n_130), .B2(n_977), .Y(n_976) );
INVx1_ASAP7_75t_L g977 ( .A(n_70), .Y(n_977) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_72), .B(n_279), .Y(n_557) );
NAND2x1p5_ASAP7_75t_L g616 ( .A(n_74), .B(n_575), .Y(n_616) );
CKINVDCx14_ASAP7_75t_R g669 ( .A(n_76), .Y(n_669) );
CKINVDCx5p33_ASAP7_75t_R g223 ( .A(n_77), .Y(n_223) );
CKINVDCx5p33_ASAP7_75t_R g179 ( .A(n_79), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_80), .B(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g110 ( .A(n_81), .Y(n_110) );
OR2x6_ASAP7_75t_L g125 ( .A(n_81), .B(n_126), .Y(n_125) );
NOR2xp33_ASAP7_75t_L g255 ( .A(n_82), .B(n_156), .Y(n_255) );
INVx1_ASAP7_75t_L g127 ( .A(n_84), .Y(n_127) );
OAI22xp5_ASAP7_75t_L g933 ( .A1(n_87), .A2(n_934), .B1(n_935), .B2(n_941), .Y(n_933) );
CKINVDCx5p33_ASAP7_75t_R g941 ( .A(n_87), .Y(n_941) );
INVx1_ASAP7_75t_L g114 ( .A(n_88), .Y(n_114) );
INVx1_ASAP7_75t_L g154 ( .A(n_89), .Y(n_154) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_89), .Y(n_157) );
BUFx5_ASAP7_75t_L g203 ( .A(n_89), .Y(n_203) );
INVx2_ASAP7_75t_L g642 ( .A(n_90), .Y(n_642) );
NOR2xp33_ASAP7_75t_L g250 ( .A(n_91), .B(n_251), .Y(n_250) );
INVx2_ASAP7_75t_L g318 ( .A(n_92), .Y(n_318) );
INVx2_ASAP7_75t_L g130 ( .A(n_93), .Y(n_130) );
INVx1_ASAP7_75t_L g322 ( .A(n_94), .Y(n_322) );
NAND2xp33_ASAP7_75t_L g609 ( .A(n_95), .B(n_610), .Y(n_609) );
INVx2_ASAP7_75t_L g241 ( .A(n_96), .Y(n_241) );
INVx2_ASAP7_75t_SL g144 ( .A(n_97), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_98), .B(n_561), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_99), .B(n_227), .Y(n_598) );
NAND2xp5_ASAP7_75t_SL g278 ( .A(n_100), .B(n_279), .Y(n_278) );
INVx1_ASAP7_75t_L g940 ( .A(n_101), .Y(n_940) );
AO32x2_ASAP7_75t_L g198 ( .A1(n_103), .A2(n_194), .A3(n_199), .B1(n_206), .B2(n_207), .Y(n_198) );
AO22x2_ASAP7_75t_L g341 ( .A1(n_103), .A2(n_199), .B1(n_342), .B2(n_344), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_104), .B(n_573), .Y(n_603) );
AOI21xp5_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_116), .B(n_985), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
BUFx2_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
BUFx24_ASAP7_75t_L g986 ( .A(n_108), .Y(n_986) );
OR2x2_ASAP7_75t_SL g108 ( .A(n_109), .B(n_115), .Y(n_108) );
NAND3xp33_ASAP7_75t_L g109 ( .A(n_110), .B(n_111), .C(n_113), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_112), .Y(n_111) );
AND2x4_ASAP7_75t_L g116 ( .A(n_117), .B(n_966), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g117 ( .A(n_118), .B(n_958), .Y(n_117) );
AOI21xp33_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_933), .B(n_942), .Y(n_118) );
OAI21x1_ASAP7_75t_SL g119 ( .A1(n_120), .A2(n_129), .B(n_545), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
BUFx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
HB1xp67_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx1_ASAP7_75t_L g962 ( .A(n_123), .Y(n_962) );
AND2x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_125), .Y(n_123) );
OR2x6_ASAP7_75t_L g948 ( .A(n_124), .B(n_125), .Y(n_948) );
INVx8_ASAP7_75t_L g549 ( .A(n_125), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g126 ( .A(n_127), .B(n_128), .Y(n_126) );
INVx2_ASAP7_75t_L g960 ( .A(n_129), .Y(n_960) );
XNOR2x1_ASAP7_75t_L g129 ( .A(n_130), .B(n_131), .Y(n_129) );
INVx2_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
XNOR2x1_ASAP7_75t_L g975 ( .A(n_132), .B(n_976), .Y(n_975) );
OR2x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_439), .Y(n_132) );
NAND3xp33_ASAP7_75t_L g133 ( .A(n_134), .B(n_336), .C(n_391), .Y(n_133) );
AOI211xp5_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_214), .B(n_304), .C(n_334), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_136), .B(n_210), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
AND2x2_ASAP7_75t_L g137 ( .A(n_138), .B(n_197), .Y(n_137) );
AND2x4_ASAP7_75t_L g397 ( .A(n_138), .B(n_361), .Y(n_397) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx1_ASAP7_75t_L g339 ( .A(n_139), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_140), .B(n_171), .Y(n_139) );
OR2x2_ASAP7_75t_L g212 ( .A(n_140), .B(n_171), .Y(n_212) );
AND2x2_ASAP7_75t_L g390 ( .A(n_140), .B(n_341), .Y(n_390) );
INVx1_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx1_ASAP7_75t_L g309 ( .A(n_141), .Y(n_309) );
INVx1_ASAP7_75t_L g366 ( .A(n_141), .Y(n_366) );
AOI21x1_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_150), .B(n_168), .Y(n_141) );
AND2x2_ASAP7_75t_L g142 ( .A(n_143), .B(n_145), .Y(n_142) );
BUFx6f_ASAP7_75t_L g206 ( .A(n_143), .Y(n_206) );
INVx3_ASAP7_75t_L g246 ( .A(n_143), .Y(n_246) );
AND2x2_ASAP7_75t_L g342 ( .A(n_143), .B(n_343), .Y(n_342) );
INVx3_ASAP7_75t_L g569 ( .A(n_143), .Y(n_569) );
INVx1_ASAP7_75t_L g572 ( .A(n_143), .Y(n_572) );
AOI21xp33_ASAP7_75t_SL g618 ( .A1(n_145), .A2(n_619), .B(n_620), .Y(n_618) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_146), .B(n_246), .Y(n_245) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx3_ASAP7_75t_L g575 ( .A(n_147), .Y(n_575) );
INVx4_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g170 ( .A(n_148), .Y(n_170) );
BUFx3_ASAP7_75t_L g239 ( .A(n_148), .Y(n_239) );
OAI22xp5_ASAP7_75t_L g150 ( .A1(n_151), .A2(n_158), .B1(n_161), .B2(n_166), .Y(n_150) );
INVx2_ASAP7_75t_L g578 ( .A(n_152), .Y(n_578) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx2_ASAP7_75t_L g224 ( .A(n_153), .Y(n_224) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g163 ( .A(n_154), .Y(n_163) );
INVx1_ASAP7_75t_L g649 ( .A(n_155), .Y(n_649) );
INVx1_ASAP7_75t_L g679 ( .A(n_155), .Y(n_679) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx2_ASAP7_75t_L g204 ( .A(n_156), .Y(n_204) );
INVx1_ASAP7_75t_L g264 ( .A(n_156), .Y(n_264) );
INVx1_ASAP7_75t_L g283 ( .A(n_156), .Y(n_283) );
INVx3_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx6_ASAP7_75t_L g165 ( .A(n_157), .Y(n_165) );
INVx2_ASAP7_75t_L g184 ( .A(n_157), .Y(n_184) );
INVx2_ASAP7_75t_L g228 ( .A(n_157), .Y(n_228) );
AOI21x1_ASAP7_75t_L g576 ( .A1(n_158), .A2(n_577), .B(n_579), .Y(n_576) );
INVx1_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx1_ASAP7_75t_L g205 ( .A(n_159), .Y(n_205) );
A2O1A1Ixp33_ASAP7_75t_L g247 ( .A1(n_159), .A2(n_248), .B(n_249), .C(n_250), .Y(n_247) );
NAND2xp5_ASAP7_75t_SL g265 ( .A(n_159), .B(n_266), .Y(n_265) );
A2O1A1Ixp33_ASAP7_75t_L g317 ( .A1(n_159), .A2(n_224), .B(n_318), .C(n_319), .Y(n_317) );
INVx1_ASAP7_75t_L g567 ( .A(n_159), .Y(n_567) );
INVx2_ASAP7_75t_SL g582 ( .A(n_159), .Y(n_582) );
INVxp67_ASAP7_75t_L g602 ( .A(n_159), .Y(n_602) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx3_ASAP7_75t_L g167 ( .A(n_160), .Y(n_167) );
INVx4_ASAP7_75t_L g178 ( .A(n_160), .Y(n_178) );
BUFx6f_ASAP7_75t_L g193 ( .A(n_160), .Y(n_193) );
INVx1_ASAP7_75t_L g275 ( .A(n_160), .Y(n_275) );
INVxp67_ASAP7_75t_L g611 ( .A(n_160), .Y(n_611) );
NOR2xp33_ASAP7_75t_L g631 ( .A(n_160), .B(n_632), .Y(n_631) );
NOR2xp33_ASAP7_75t_L g634 ( .A(n_160), .B(n_635), .Y(n_634) );
INVx3_ASAP7_75t_L g189 ( .A(n_162), .Y(n_189) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx1_ASAP7_75t_L g251 ( .A(n_163), .Y(n_251) );
INVx1_ASAP7_75t_L g314 ( .A(n_164), .Y(n_314) );
INVx1_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx2_ASAP7_75t_L g175 ( .A(n_165), .Y(n_175) );
INVx2_ASAP7_75t_SL g191 ( .A(n_165), .Y(n_191) );
INVx2_ASAP7_75t_L g236 ( .A(n_165), .Y(n_236) );
INVx1_ASAP7_75t_L g561 ( .A(n_165), .Y(n_561) );
INVx1_ASAP7_75t_L g610 ( .A(n_165), .Y(n_610) );
NOR2xp33_ASAP7_75t_L g225 ( .A(n_166), .B(n_185), .Y(n_225) );
NOR3xp33_ASAP7_75t_L g229 ( .A(n_166), .B(n_185), .C(n_230), .Y(n_229) );
NAND3xp33_ASAP7_75t_L g653 ( .A(n_166), .B(n_619), .C(n_628), .Y(n_653) );
INVx3_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
A2O1A1Ixp33_ASAP7_75t_L g252 ( .A1(n_167), .A2(n_253), .B(n_254), .C(n_255), .Y(n_252) );
A2O1A1Ixp33_ASAP7_75t_L g313 ( .A1(n_167), .A2(n_314), .B(n_315), .C(n_316), .Y(n_313) );
NOR2xp33_ASAP7_75t_L g168 ( .A(n_169), .B(n_170), .Y(n_168) );
BUFx3_ASAP7_75t_L g194 ( .A(n_170), .Y(n_194) );
NOR2xp33_ASAP7_75t_L g195 ( .A(n_170), .B(n_196), .Y(n_195) );
INVx3_ASAP7_75t_L g279 ( .A(n_170), .Y(n_279) );
NOR2xp33_ASAP7_75t_L g641 ( .A(n_170), .B(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g323 ( .A(n_171), .Y(n_323) );
INVx2_ASAP7_75t_L g329 ( .A(n_171), .Y(n_329) );
AND2x2_ASAP7_75t_L g351 ( .A(n_171), .B(n_345), .Y(n_351) );
AND2x2_ASAP7_75t_L g360 ( .A(n_171), .B(n_311), .Y(n_360) );
AO31x2_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_187), .A3(n_194), .B(n_195), .Y(n_171) );
AOI221x1_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_176), .B1(n_180), .B2(n_182), .C(n_185), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
AND2x2_ASAP7_75t_L g176 ( .A(n_177), .B(n_179), .Y(n_176) );
AND2x2_ASAP7_75t_L g180 ( .A(n_177), .B(n_181), .Y(n_180) );
INVx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g291 ( .A(n_178), .B(n_292), .Y(n_291) );
NOR2xp33_ASAP7_75t_SL g637 ( .A(n_178), .B(n_638), .Y(n_637) );
NOR2xp33_ASAP7_75t_L g639 ( .A(n_178), .B(n_640), .Y(n_639) );
NAND3xp33_ASAP7_75t_SL g646 ( .A(n_178), .B(n_619), .C(n_628), .Y(n_646) );
INVx1_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_183), .B(n_634), .Y(n_633) );
AOI22xp5_ASAP7_75t_L g636 ( .A1(n_183), .A2(n_254), .B1(n_637), .B2(n_639), .Y(n_636) );
INVx2_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVxp67_ASAP7_75t_SL g273 ( .A(n_184), .Y(n_273) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_185), .B(n_233), .Y(n_232) );
INVx4_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
INVx1_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_191), .B(n_192), .Y(n_190) );
OAI22xp5_ASAP7_75t_L g199 ( .A1(n_193), .A2(n_200), .B1(n_201), .B2(n_205), .Y(n_199) );
INVx4_ASAP7_75t_L g233 ( .A(n_193), .Y(n_233) );
AOI21xp5_ASAP7_75t_L g281 ( .A1(n_193), .A2(n_282), .B(n_284), .Y(n_281) );
AOI21xp5_ASAP7_75t_L g559 ( .A1(n_193), .A2(n_560), .B(n_562), .Y(n_559) );
OAI22xp5_ASAP7_75t_L g593 ( .A1(n_193), .A2(n_594), .B1(n_595), .B2(n_598), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_193), .B(n_674), .Y(n_673) );
INVx2_ASAP7_75t_L g344 ( .A(n_194), .Y(n_344) );
INVx2_ASAP7_75t_L g213 ( .A(n_197), .Y(n_213) );
AND2x2_ASAP7_75t_L g350 ( .A(n_197), .B(n_351), .Y(n_350) );
OR2x2_ASAP7_75t_L g384 ( .A(n_197), .B(n_385), .Y(n_384) );
AND2x4_ASAP7_75t_L g462 ( .A(n_197), .B(n_365), .Y(n_462) );
AND2x2_ASAP7_75t_L g515 ( .A(n_197), .B(n_360), .Y(n_515) );
AND2x2_ASAP7_75t_SL g531 ( .A(n_197), .B(n_310), .Y(n_531) );
BUFx3_ASAP7_75t_L g541 ( .A(n_197), .Y(n_541) );
BUFx8_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
INVx2_ASAP7_75t_L g327 ( .A(n_198), .Y(n_327) );
AND2x2_ASAP7_75t_L g431 ( .A(n_198), .B(n_432), .Y(n_431) );
OAI22xp33_ASAP7_75t_L g234 ( .A1(n_202), .A2(n_235), .B1(n_236), .B2(n_237), .Y(n_234) );
INVx2_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
INVx2_ASAP7_75t_L g254 ( .A(n_203), .Y(n_254) );
INVx2_ASAP7_75t_L g263 ( .A(n_203), .Y(n_263) );
INVx2_ASAP7_75t_L g285 ( .A(n_203), .Y(n_285) );
INVx1_ASAP7_75t_L g289 ( .A(n_203), .Y(n_289) );
INVx2_ASAP7_75t_L g563 ( .A(n_203), .Y(n_563) );
INVx1_ASAP7_75t_L g248 ( .A(n_204), .Y(n_248) );
OAI21x1_ASAP7_75t_L g592 ( .A1(n_206), .A2(n_593), .B(n_599), .Y(n_592) );
AO31x2_ASAP7_75t_L g660 ( .A1(n_206), .A2(n_661), .A3(n_666), .B(n_668), .Y(n_660) );
AO31x2_ASAP7_75t_L g689 ( .A1(n_206), .A2(n_661), .A3(n_666), .B(n_668), .Y(n_689) );
INVxp67_ASAP7_75t_L g303 ( .A(n_207), .Y(n_303) );
INVx1_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_208), .B(n_241), .Y(n_240) );
INVx1_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx1_ASAP7_75t_L g257 ( .A(n_209), .Y(n_257) );
NOR2xp67_ASAP7_75t_L g266 ( .A(n_209), .B(n_246), .Y(n_266) );
BUFx3_ASAP7_75t_L g268 ( .A(n_209), .Y(n_268) );
NOR2xp33_ASAP7_75t_L g293 ( .A(n_209), .B(n_246), .Y(n_293) );
NOR2xp33_ASAP7_75t_L g320 ( .A(n_209), .B(n_246), .Y(n_320) );
INVx1_ASAP7_75t_L g343 ( .A(n_209), .Y(n_343) );
INVx2_ASAP7_75t_L g628 ( .A(n_209), .Y(n_628) );
NOR2xp33_ASAP7_75t_L g674 ( .A(n_209), .B(n_246), .Y(n_674) );
HB1xp67_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
NAND3xp33_ASAP7_75t_SL g526 ( .A(n_211), .B(n_527), .C(n_530), .Y(n_526) );
OR2x2_ASAP7_75t_L g211 ( .A(n_212), .B(n_213), .Y(n_211) );
INVx2_ASAP7_75t_L g405 ( .A(n_212), .Y(n_405) );
NAND2x1_ASAP7_75t_L g214 ( .A(n_215), .B(n_294), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g334 ( .A(n_215), .B(n_335), .Y(n_334) );
INVx2_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
AND2x2_ASAP7_75t_L g216 ( .A(n_217), .B(n_259), .Y(n_216) );
INVx1_ASAP7_75t_L g352 ( .A(n_217), .Y(n_352) );
AND2x2_ASAP7_75t_L g482 ( .A(n_217), .B(n_483), .Y(n_482) );
AND2x2_ASAP7_75t_L g520 ( .A(n_217), .B(n_373), .Y(n_520) );
AND2x4_ASAP7_75t_L g217 ( .A(n_218), .B(n_242), .Y(n_217) );
OR2x2_ASAP7_75t_L g387 ( .A(n_218), .B(n_301), .Y(n_387) );
AND2x2_ASAP7_75t_L g474 ( .A(n_218), .B(n_348), .Y(n_474) );
INVx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
AND2x2_ASAP7_75t_L g375 ( .A(n_219), .B(n_333), .Y(n_375) );
BUFx2_ASAP7_75t_L g379 ( .A(n_219), .Y(n_379) );
OR2x2_ASAP7_75t_L g396 ( .A(n_219), .B(n_244), .Y(n_396) );
AO21x2_ASAP7_75t_L g219 ( .A1(n_220), .A2(n_238), .B(n_240), .Y(n_219) );
AO21x2_ASAP7_75t_L g302 ( .A1(n_220), .A2(n_240), .B(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_221), .B(n_231), .Y(n_220) );
AOI22xp5_ASAP7_75t_L g221 ( .A1(n_222), .A2(n_225), .B1(n_226), .B2(n_229), .Y(n_221) );
NOR2xp67_ASAP7_75t_L g222 ( .A(n_223), .B(n_224), .Y(n_222) );
INVx1_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
INVx2_ASAP7_75t_L g272 ( .A(n_228), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_232), .B(n_234), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_233), .B(n_596), .Y(n_595) );
OAI22x1_ASAP7_75t_L g661 ( .A1(n_233), .A2(n_662), .B1(n_663), .B2(n_664), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_236), .B(n_291), .Y(n_290) );
INVx2_ASAP7_75t_L g607 ( .A(n_236), .Y(n_607) );
OR2x2_ASAP7_75t_L g583 ( .A(n_238), .B(n_584), .Y(n_583) );
NOR2xp67_ASAP7_75t_SL g668 ( .A(n_238), .B(n_669), .Y(n_668) );
INVx3_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
OA21x2_ASAP7_75t_L g591 ( .A1(n_239), .A2(n_592), .B(n_603), .Y(n_591) );
OA21x2_ASAP7_75t_L g695 ( .A1(n_239), .A2(n_592), .B(n_603), .Y(n_695) );
INVx1_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
AND2x2_ASAP7_75t_L g426 ( .A(n_243), .B(n_277), .Y(n_426) );
INVx2_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
INVx1_ASAP7_75t_L g299 ( .A(n_244), .Y(n_299) );
INVx2_ASAP7_75t_L g333 ( .A(n_244), .Y(n_333) );
AND2x2_ASAP7_75t_L g407 ( .A(n_244), .B(n_302), .Y(n_407) );
INVx1_ASAP7_75t_L g459 ( .A(n_244), .Y(n_459) );
HB1xp67_ASAP7_75t_L g493 ( .A(n_244), .Y(n_493) );
AO31x2_ASAP7_75t_L g244 ( .A1(n_245), .A2(n_247), .A3(n_252), .B(n_256), .Y(n_244) );
NOR2xp33_ASAP7_75t_SL g256 ( .A(n_257), .B(n_258), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g321 ( .A(n_257), .B(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g667 ( .A(n_257), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_259), .B(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g411 ( .A(n_259), .B(n_407), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_259), .B(n_379), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_259), .B(n_378), .Y(n_542) );
NAND2xp67_ASAP7_75t_L g543 ( .A(n_259), .B(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_L g259 ( .A(n_260), .B(n_276), .Y(n_259) );
INVx1_ASAP7_75t_L g297 ( .A(n_260), .Y(n_297) );
INVx2_ASAP7_75t_L g348 ( .A(n_260), .Y(n_348) );
INVx1_ASAP7_75t_L g356 ( .A(n_260), .Y(n_356) );
AND2x2_ASAP7_75t_L g418 ( .A(n_260), .B(n_277), .Y(n_418) );
NAND2x1p5_ASAP7_75t_L g260 ( .A(n_261), .B(n_269), .Y(n_260) );
AND2x2_ASAP7_75t_SL g455 ( .A(n_261), .B(n_269), .Y(n_455) );
OA21x2_ASAP7_75t_L g261 ( .A1(n_262), .A2(n_265), .B(n_267), .Y(n_261) );
INVx2_ASAP7_75t_L g648 ( .A(n_263), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_266), .B(n_275), .Y(n_274) );
OR2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_274), .Y(n_269) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
INVx1_ASAP7_75t_L g663 ( .A(n_275), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_275), .B(n_674), .Y(n_677) );
OR2x2_ASAP7_75t_L g358 ( .A(n_276), .B(n_302), .Y(n_358) );
INVx2_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
INVx1_ASAP7_75t_L g301 ( .A(n_277), .Y(n_301) );
INVx1_ASAP7_75t_L g382 ( .A(n_277), .Y(n_382) );
HB1xp67_ASAP7_75t_L g450 ( .A(n_277), .Y(n_450) );
AND2x4_ASAP7_75t_L g277 ( .A(n_278), .B(n_280), .Y(n_277) );
NOR2x1_ASAP7_75t_L g568 ( .A(n_279), .B(n_569), .Y(n_568) );
OAI21xp5_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_286), .B(n_293), .Y(n_280) );
OAI21xp5_ASAP7_75t_L g286 ( .A1(n_287), .A2(n_288), .B(n_290), .Y(n_286) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx2_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
AOI22xp5_ASAP7_75t_L g487 ( .A1(n_295), .A2(n_488), .B1(n_490), .B2(n_492), .Y(n_487) );
AND2x4_ASAP7_75t_L g295 ( .A(n_296), .B(n_300), .Y(n_295) );
AND2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
BUFx3_ASAP7_75t_L g402 ( .A(n_297), .Y(n_402) );
AND2x2_ASAP7_75t_L g449 ( .A(n_298), .B(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
AND2x2_ASAP7_75t_L g458 ( .A(n_301), .B(n_459), .Y(n_458) );
AND2x2_ASAP7_75t_L g347 ( .A(n_302), .B(n_348), .Y(n_347) );
AOI21xp33_ASAP7_75t_L g304 ( .A1(n_305), .A2(n_324), .B(n_330), .Y(n_304) );
OAI21xp5_ASAP7_75t_L g427 ( .A1(n_305), .A2(n_428), .B(n_429), .Y(n_427) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g306 ( .A(n_307), .B(n_310), .Y(n_306) );
AND2x4_ASAP7_75t_L g325 ( .A(n_307), .B(n_326), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_307), .B(n_340), .Y(n_460) );
INVx4_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g416 ( .A(n_308), .B(n_310), .Y(n_416) );
INVx2_ASAP7_75t_L g467 ( .A(n_308), .Y(n_467) );
NAND2xp5_ASAP7_75t_SL g521 ( .A(n_308), .B(n_351), .Y(n_521) );
BUFx3_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g432 ( .A(n_309), .Y(n_432) );
INVx2_ASAP7_75t_L g335 ( .A(n_310), .Y(n_335) );
INVx2_ASAP7_75t_L g385 ( .A(n_310), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_310), .B(n_390), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_310), .B(n_375), .Y(n_478) );
AND2x4_ASAP7_75t_L g310 ( .A(n_311), .B(n_323), .Y(n_310) );
INVx2_ASAP7_75t_L g345 ( .A(n_311), .Y(n_345) );
INVx1_ASAP7_75t_L g368 ( .A(n_311), .Y(n_368) );
BUFx3_ASAP7_75t_L g399 ( .A(n_311), .Y(n_399) );
AND2x4_ASAP7_75t_L g469 ( .A(n_311), .B(n_327), .Y(n_469) );
INVx3_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
AO31x2_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_317), .A3(n_320), .B(n_321), .Y(n_312) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g415 ( .A(n_326), .Y(n_415) );
AND2x2_ASAP7_75t_L g326 ( .A(n_327), .B(n_328), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_327), .B(n_432), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_328), .B(n_424), .Y(n_423) );
INVx2_ASAP7_75t_SL g328 ( .A(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g365 ( .A(n_329), .B(n_366), .Y(n_365) );
BUFx3_ASAP7_75t_L g409 ( .A(n_329), .Y(n_409) );
INVx1_ASAP7_75t_L g491 ( .A(n_329), .Y(n_491) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
NOR2xp67_ASAP7_75t_L g421 ( .A(n_332), .B(n_387), .Y(n_421) );
HB1xp67_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
OR2x2_ASAP7_75t_L g437 ( .A(n_333), .B(n_424), .Y(n_437) );
INVxp67_ASAP7_75t_SL g537 ( .A(n_333), .Y(n_537) );
NOR3xp33_ASAP7_75t_L g336 ( .A(n_337), .B(n_353), .C(n_362), .Y(n_336) );
OAI22xp33_ASAP7_75t_SL g337 ( .A1(n_338), .A2(n_346), .B1(n_349), .B2(n_352), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_339), .B(n_340), .Y(n_338) );
INVx2_ASAP7_75t_L g512 ( .A(n_339), .Y(n_512) );
AND2x4_ASAP7_75t_L g404 ( .A(n_340), .B(n_405), .Y(n_404) );
INVx4_ASAP7_75t_L g420 ( .A(n_340), .Y(n_420) );
AND2x4_ASAP7_75t_L g340 ( .A(n_341), .B(n_345), .Y(n_340) );
INVx1_ASAP7_75t_L g361 ( .A(n_341), .Y(n_361) );
INVx1_ASAP7_75t_L g369 ( .A(n_341), .Y(n_369) );
AND2x4_ASAP7_75t_L g398 ( .A(n_341), .B(n_399), .Y(n_398) );
AND2x2_ASAP7_75t_L g410 ( .A(n_345), .B(n_366), .Y(n_410) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_SL g457 ( .A(n_347), .B(n_458), .Y(n_457) );
AND2x2_ASAP7_75t_L g510 ( .A(n_347), .B(n_426), .Y(n_510) );
BUFx2_ASAP7_75t_L g373 ( .A(n_348), .Y(n_373) );
HB1xp67_ASAP7_75t_L g499 ( .A(n_348), .Y(n_499) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
NOR2x1_ASAP7_75t_L g363 ( .A(n_350), .B(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g430 ( .A(n_351), .B(n_431), .Y(n_430) );
AND2x2_ASAP7_75t_L g470 ( .A(n_351), .B(n_471), .Y(n_470) );
AND2x2_ASAP7_75t_L g505 ( .A(n_351), .B(n_424), .Y(n_505) );
AND2x2_ASAP7_75t_L g353 ( .A(n_354), .B(n_359), .Y(n_353) );
INVx3_ASAP7_75t_L g428 ( .A(n_354), .Y(n_428) );
AND2x4_ASAP7_75t_L g354 ( .A(n_355), .B(n_357), .Y(n_354) );
AND2x2_ASAP7_75t_L g452 ( .A(n_355), .B(n_407), .Y(n_452) );
INVx1_ASAP7_75t_L g534 ( .A(n_355), .Y(n_534) );
INVx2_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g425 ( .A(n_356), .B(n_426), .Y(n_425) );
INVxp67_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g435 ( .A(n_358), .Y(n_435) );
INVxp67_ASAP7_75t_SL g500 ( .A(n_358), .Y(n_500) );
OR2x6_ASAP7_75t_L g536 ( .A(n_358), .B(n_537), .Y(n_536) );
OAI31xp33_ASAP7_75t_L g451 ( .A1(n_359), .A2(n_371), .A3(n_452), .B(n_453), .Y(n_451) );
AND2x2_ASAP7_75t_L g359 ( .A(n_360), .B(n_361), .Y(n_359) );
INVx2_ASAP7_75t_L g446 ( .A(n_360), .Y(n_446) );
INVx2_ASAP7_75t_L g529 ( .A(n_360), .Y(n_529) );
OAI21xp5_ASAP7_75t_SL g362 ( .A1(n_363), .A2(n_370), .B(n_376), .Y(n_362) );
AND2x2_ASAP7_75t_L g364 ( .A(n_365), .B(n_367), .Y(n_364) );
INVxp67_ASAP7_75t_SL g539 ( .A(n_365), .Y(n_539) );
HB1xp67_ASAP7_75t_L g401 ( .A(n_366), .Y(n_401) );
INVx2_ASAP7_75t_L g424 ( .A(n_366), .Y(n_424) );
AOI33xp33_ASAP7_75t_L g419 ( .A1(n_367), .A2(n_420), .A3(n_421), .B1(n_422), .B2(n_423), .B3(n_425), .Y(n_419) );
AND2x2_ASAP7_75t_L g486 ( .A(n_367), .B(n_424), .Y(n_486) );
AND2x2_ASAP7_75t_L g488 ( .A(n_367), .B(n_489), .Y(n_488) );
AND2x4_ASAP7_75t_SL g367 ( .A(n_368), .B(n_369), .Y(n_367) );
INVxp67_ASAP7_75t_SL g370 ( .A(n_371), .Y(n_370) );
NOR2x1p5_ASAP7_75t_L g371 ( .A(n_372), .B(n_374), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g406 ( .A(n_373), .B(n_407), .Y(n_406) );
INVx2_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AND2x4_ASAP7_75t_L g400 ( .A(n_375), .B(n_401), .Y(n_400) );
NAND2x1p5_ASAP7_75t_L g463 ( .A(n_375), .B(n_464), .Y(n_463) );
AND2x2_ASAP7_75t_L g524 ( .A(n_375), .B(n_418), .Y(n_524) );
AOI22xp5_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_383), .B1(n_386), .B2(n_388), .Y(n_376) );
AND2x2_ASAP7_75t_L g377 ( .A(n_378), .B(n_380), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
AND2x2_ASAP7_75t_L g444 ( .A(n_379), .B(n_418), .Y(n_444) );
INVx2_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_381), .B(n_402), .Y(n_476) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_L g483 ( .A(n_382), .B(n_455), .Y(n_483) );
AND2x2_ASAP7_75t_L g517 ( .A(n_382), .B(n_455), .Y(n_517) );
INVx2_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
NOR2xp67_ASAP7_75t_SL g453 ( .A(n_387), .B(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVxp67_ASAP7_75t_L g477 ( .A(n_390), .Y(n_477) );
NOR3xp33_ASAP7_75t_L g391 ( .A(n_392), .B(n_412), .C(n_427), .Y(n_391) );
OAI21xp5_ASAP7_75t_SL g392 ( .A1(n_393), .A2(n_402), .B(n_403), .Y(n_392) );
AOI22xp5_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_397), .B1(n_398), .B2(n_400), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
HB1xp67_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx2_ASAP7_75t_L g544 ( .A(n_396), .Y(n_544) );
INVx2_ASAP7_75t_L g495 ( .A(n_398), .Y(n_495) );
INVx1_ASAP7_75t_L g528 ( .A(n_401), .Y(n_528) );
AOI22xp5_ASAP7_75t_L g403 ( .A1(n_404), .A2(n_406), .B1(n_408), .B2(n_411), .Y(n_403) );
AND2x2_ASAP7_75t_L g417 ( .A(n_407), .B(n_418), .Y(n_417) );
OAI21xp5_ASAP7_75t_L g522 ( .A1(n_408), .A2(n_523), .B(n_524), .Y(n_522) );
AND2x2_ASAP7_75t_L g408 ( .A(n_409), .B(n_410), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_413), .B(n_419), .Y(n_412) );
OAI21xp33_ASAP7_75t_L g413 ( .A1(n_414), .A2(n_416), .B(n_417), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g438 ( .A(n_418), .Y(n_438) );
AND2x2_ASAP7_75t_L g492 ( .A(n_418), .B(n_493), .Y(n_492) );
NOR3xp33_ASAP7_75t_L g436 ( .A(n_420), .B(n_437), .C(n_438), .Y(n_436) );
OAI221xp5_ASAP7_75t_L g480 ( .A1(n_420), .A2(n_481), .B1(n_484), .B2(n_485), .C(n_487), .Y(n_480) );
INVx2_ASAP7_75t_L g442 ( .A(n_422), .Y(n_442) );
INVx2_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g489 ( .A(n_424), .Y(n_489) );
BUFx3_ASAP7_75t_L g514 ( .A(n_424), .Y(n_514) );
AND2x2_ASAP7_75t_L g523 ( .A(n_426), .B(n_474), .Y(n_523) );
AOI21xp5_ASAP7_75t_L g429 ( .A1(n_430), .A2(n_433), .B(n_436), .Y(n_429) );
AND2x4_ASAP7_75t_SL g490 ( .A(n_431), .B(n_491), .Y(n_490) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx2_ASAP7_75t_L g497 ( .A(n_437), .Y(n_497) );
NAND4xp25_ASAP7_75t_L g439 ( .A(n_440), .B(n_479), .C(n_507), .D(n_525), .Y(n_439) );
NOR2xp33_ASAP7_75t_L g440 ( .A(n_441), .B(n_456), .Y(n_440) );
OAI221xp5_ASAP7_75t_SL g441 ( .A1(n_442), .A2(n_443), .B1(n_445), .B2(n_448), .C(n_451), .Y(n_441) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
OR2x2_ASAP7_75t_L g445 ( .A(n_446), .B(n_447), .Y(n_445) );
INVx1_ASAP7_75t_L g471 ( .A(n_447), .Y(n_471) );
INVx1_ASAP7_75t_L g502 ( .A(n_447), .Y(n_502) );
INVxp67_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g473 ( .A(n_450), .Y(n_473) );
INVx1_ASAP7_75t_SL g484 ( .A(n_452), .Y(n_484) );
INVx2_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g464 ( .A(n_455), .Y(n_464) );
OAI221xp5_ASAP7_75t_L g456 ( .A1(n_457), .A2(n_460), .B1(n_461), .B2(n_463), .C(n_465), .Y(n_456) );
AND2x2_ASAP7_75t_L g516 ( .A(n_459), .B(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx2_ASAP7_75t_L g506 ( .A(n_463), .Y(n_506) );
O2A1O1Ixp5_ASAP7_75t_L g465 ( .A1(n_466), .A2(n_470), .B(n_472), .C(n_475), .Y(n_465) );
NOR2x1_ASAP7_75t_L g466 ( .A(n_467), .B(n_468), .Y(n_466) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
AND2x4_ASAP7_75t_L g472 ( .A(n_473), .B(n_474), .Y(n_472) );
AOI21xp5_ASAP7_75t_L g475 ( .A1(n_476), .A2(n_477), .B(n_478), .Y(n_475) );
NOR2xp33_ASAP7_75t_L g479 ( .A(n_480), .B(n_494), .Y(n_479) );
INVx2_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVxp67_ASAP7_75t_SL g485 ( .A(n_486), .Y(n_485) );
OAI21xp33_ASAP7_75t_L g494 ( .A1(n_495), .A2(n_496), .B(n_501), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_497), .B(n_498), .Y(n_496) );
AND2x4_ASAP7_75t_L g498 ( .A(n_499), .B(n_500), .Y(n_498) );
AOI22xp5_ASAP7_75t_L g501 ( .A1(n_502), .A2(n_503), .B1(n_505), .B2(n_506), .Y(n_501) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
AOI221xp5_ASAP7_75t_L g507 ( .A1(n_508), .A2(n_511), .B1(n_513), .B2(n_516), .C(n_518), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
CKINVDCx5p33_ASAP7_75t_R g511 ( .A(n_512), .Y(n_511) );
AND2x2_ASAP7_75t_L g513 ( .A(n_514), .B(n_515), .Y(n_513) );
OAI21xp5_ASAP7_75t_L g518 ( .A1(n_519), .A2(n_521), .B(n_522), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
AOI22xp5_ASAP7_75t_L g525 ( .A1(n_526), .A2(n_532), .B1(n_538), .B2(n_540), .Y(n_525) );
OR2x2_ASAP7_75t_L g527 ( .A(n_528), .B(n_529), .Y(n_527) );
INVx2_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
AND2x4_ASAP7_75t_L g532 ( .A(n_533), .B(n_535), .Y(n_532) );
INVxp67_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVxp67_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
OAI21xp33_ASAP7_75t_L g540 ( .A1(n_541), .A2(n_542), .B(n_543), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_546), .B(n_550), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g963 ( .A(n_546), .B(n_964), .Y(n_963) );
CKINVDCx5p33_ASAP7_75t_R g546 ( .A(n_547), .Y(n_546) );
OR2x6_ASAP7_75t_L g547 ( .A(n_548), .B(n_549), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g952 ( .A(n_549), .B(n_953), .Y(n_952) );
INVx2_ASAP7_75t_L g964 ( .A(n_550), .Y(n_964) );
OR2x2_ASAP7_75t_L g550 ( .A(n_551), .B(n_837), .Y(n_550) );
NAND4xp25_ASAP7_75t_L g551 ( .A(n_552), .B(n_732), .C(n_773), .D(n_808), .Y(n_551) );
AOI211xp5_ASAP7_75t_L g552 ( .A1(n_553), .A2(n_585), .B(n_681), .C(n_703), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
OR2x2_ASAP7_75t_L g801 ( .A(n_554), .B(n_710), .Y(n_801) );
OR2x2_ASAP7_75t_L g822 ( .A(n_554), .B(n_701), .Y(n_822) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g683 ( .A(n_555), .B(n_684), .Y(n_683) );
AND2x2_ASAP7_75t_L g870 ( .A(n_555), .B(n_701), .Y(n_870) );
AND2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_570), .Y(n_555) );
AND2x2_ASAP7_75t_L g698 ( .A(n_556), .B(n_699), .Y(n_698) );
INVx3_ASAP7_75t_L g718 ( .A(n_556), .Y(n_718) );
INVx2_ASAP7_75t_L g722 ( .A(n_556), .Y(n_722) );
AND2x4_ASAP7_75t_L g556 ( .A(n_557), .B(n_558), .Y(n_556) );
OAI21x1_ASAP7_75t_L g558 ( .A1(n_559), .A2(n_564), .B(n_568), .Y(n_558) );
INVx2_ASAP7_75t_L g594 ( .A(n_563), .Y(n_594) );
AOI21xp5_ASAP7_75t_L g564 ( .A1(n_565), .A2(n_566), .B(n_567), .Y(n_564) );
INVx2_ASAP7_75t_L g619 ( .A(n_569), .Y(n_619) );
INVx2_ASAP7_75t_SL g699 ( .A(n_570), .Y(n_699) );
AND2x2_ASAP7_75t_L g825 ( .A(n_570), .B(n_718), .Y(n_825) );
OAI21x1_ASAP7_75t_L g570 ( .A1(n_571), .A2(n_576), .B(n_583), .Y(n_570) );
OAI21xp5_ASAP7_75t_L g771 ( .A1(n_571), .A2(n_576), .B(n_583), .Y(n_771) );
OR2x2_ASAP7_75t_L g571 ( .A(n_572), .B(n_573), .Y(n_571) );
NOR2xp33_ASAP7_75t_L g626 ( .A(n_572), .B(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
OR2x2_ASAP7_75t_L g650 ( .A(n_574), .B(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
AOI21x1_ASAP7_75t_L g579 ( .A1(n_580), .A2(n_581), .B(n_582), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_582), .B(n_616), .Y(n_617) );
AO21x1_ASAP7_75t_L g585 ( .A1(n_586), .A2(n_621), .B(n_655), .Y(n_585) );
AOI22xp5_ASAP7_75t_L g844 ( .A1(n_586), .A2(n_845), .B1(n_850), .B2(n_853), .Y(n_844) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g656 ( .A(n_589), .Y(n_656) );
INVx1_ASAP7_75t_L g799 ( .A(n_589), .Y(n_799) );
OR2x2_ASAP7_75t_L g883 ( .A(n_589), .B(n_884), .Y(n_883) );
INVx2_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g757 ( .A(n_590), .B(n_692), .Y(n_757) );
AND2x2_ASAP7_75t_L g899 ( .A(n_590), .B(n_884), .Y(n_899) );
AND2x2_ASAP7_75t_L g590 ( .A(n_591), .B(n_604), .Y(n_590) );
AND2x2_ASAP7_75t_L g793 ( .A(n_591), .B(n_671), .Y(n_793) );
AND2x2_ASAP7_75t_L g807 ( .A(n_591), .B(n_686), .Y(n_807) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
AOI21xp5_ASAP7_75t_L g599 ( .A1(n_600), .A2(n_601), .B(n_602), .Y(n_599) );
AND2x2_ASAP7_75t_L g688 ( .A(n_604), .B(n_689), .Y(n_688) );
AND2x4_ASAP7_75t_L g746 ( .A(n_604), .B(n_747), .Y(n_746) );
OR2x2_ASAP7_75t_L g753 ( .A(n_604), .B(n_689), .Y(n_753) );
AO21x2_ASAP7_75t_L g604 ( .A1(n_605), .A2(n_612), .B(n_618), .Y(n_604) );
AO21x2_ASAP7_75t_L g708 ( .A1(n_605), .A2(n_612), .B(n_618), .Y(n_708) );
OAI21x1_ASAP7_75t_L g605 ( .A1(n_606), .A2(n_608), .B(n_611), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_607), .B(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx2_ASAP7_75t_L g665 ( .A(n_610), .Y(n_665) );
OAI21x1_ASAP7_75t_SL g612 ( .A1(n_613), .A2(n_614), .B(n_617), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
INVx1_ASAP7_75t_L g620 ( .A(n_616), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
OR2x2_ASAP7_75t_L g819 ( .A(n_622), .B(n_820), .Y(n_819) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
AND2x2_ASAP7_75t_L g750 ( .A(n_623), .B(n_735), .Y(n_750) );
AND2x2_ASAP7_75t_L g803 ( .A(n_623), .B(n_698), .Y(n_803) );
AND2x2_ASAP7_75t_L g623 ( .A(n_624), .B(n_643), .Y(n_623) );
AND2x2_ASAP7_75t_L g711 ( .A(n_624), .B(n_644), .Y(n_711) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g724 ( .A(n_625), .Y(n_724) );
INVx1_ASAP7_75t_L g739 ( .A(n_625), .Y(n_739) );
AND2x2_ASAP7_75t_L g760 ( .A(n_625), .B(n_699), .Y(n_760) );
AND2x2_ASAP7_75t_L g772 ( .A(n_625), .B(n_644), .Y(n_772) );
OR2x2_ASAP7_75t_L g782 ( .A(n_625), .B(n_771), .Y(n_782) );
INVxp67_ASAP7_75t_L g930 ( .A(n_625), .Y(n_930) );
AO21x2_ASAP7_75t_L g625 ( .A1(n_626), .A2(n_629), .B(n_641), .Y(n_625) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
NAND3xp33_ASAP7_75t_SL g629 ( .A(n_630), .B(n_633), .C(n_636), .Y(n_629) );
CKINVDCx5p33_ASAP7_75t_R g980 ( .A(n_642), .Y(n_980) );
INVx2_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g702 ( .A(n_644), .Y(n_702) );
NOR2x1_ASAP7_75t_L g738 ( .A(n_644), .B(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g764 ( .A(n_644), .Y(n_764) );
HB1xp67_ASAP7_75t_L g788 ( .A(n_644), .Y(n_788) );
INVx1_ASAP7_75t_L g836 ( .A(n_644), .Y(n_836) );
AND2x2_ASAP7_75t_L g854 ( .A(n_644), .B(n_718), .Y(n_854) );
OR2x6_ASAP7_75t_L g644 ( .A(n_645), .B(n_652), .Y(n_644) );
OAI21x1_ASAP7_75t_L g645 ( .A1(n_646), .A2(n_647), .B(n_650), .Y(n_645) );
NOR2xp67_ASAP7_75t_L g652 ( .A(n_653), .B(n_654), .Y(n_652) );
INVx1_ASAP7_75t_L g889 ( .A(n_655), .Y(n_889) );
AND2x4_ASAP7_75t_L g655 ( .A(n_656), .B(n_657), .Y(n_655) );
AND2x2_ASAP7_75t_L g657 ( .A(n_658), .B(n_670), .Y(n_657) );
INVx2_ASAP7_75t_L g692 ( .A(n_658), .Y(n_692) );
INVx1_ASAP7_75t_L g791 ( .A(n_658), .Y(n_791) );
INVx2_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g745 ( .A(n_659), .Y(n_745) );
AND2x2_ASAP7_75t_L g766 ( .A(n_659), .B(n_729), .Y(n_766) );
AND2x2_ASAP7_75t_L g831 ( .A(n_659), .B(n_708), .Y(n_831) );
INVx3_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
AND2x2_ASAP7_75t_L g780 ( .A(n_660), .B(n_694), .Y(n_780) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx2_ASAP7_75t_L g884 ( .A(n_670), .Y(n_884) );
INVx2_ASAP7_75t_L g907 ( .A(n_670), .Y(n_907) );
INVx2_ASAP7_75t_SL g670 ( .A(n_671), .Y(n_670) );
AND2x2_ASAP7_75t_L g671 ( .A(n_672), .B(n_676), .Y(n_671) );
NAND2x1p5_ASAP7_75t_L g686 ( .A(n_672), .B(n_676), .Y(n_686) );
OR2x2_ASAP7_75t_L g672 ( .A(n_673), .B(n_675), .Y(n_672) );
OA21x2_ASAP7_75t_L g676 ( .A1(n_677), .A2(n_678), .B(n_680), .Y(n_676) );
O2A1O1Ixp33_ASAP7_75t_SL g681 ( .A1(n_682), .A2(n_687), .B(n_690), .C(n_700), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
OR2x2_ASAP7_75t_L g901 ( .A(n_684), .B(n_886), .Y(n_901) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g743 ( .A(n_685), .Y(n_743) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
AND2x2_ASAP7_75t_L g693 ( .A(n_686), .B(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g715 ( .A(n_686), .Y(n_715) );
INVx2_ASAP7_75t_L g729 ( .A(n_686), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g848 ( .A(n_686), .B(n_849), .Y(n_848) );
OAI21xp33_ASAP7_75t_L g839 ( .A1(n_687), .A2(n_840), .B(n_844), .Y(n_839) );
INVx2_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
AND2x4_ASAP7_75t_L g706 ( .A(n_689), .B(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g814 ( .A(n_689), .Y(n_814) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_691), .B(n_696), .Y(n_690) );
AND2x2_ASAP7_75t_L g691 ( .A(n_692), .B(n_693), .Y(n_691) );
INVx1_ASAP7_75t_L g798 ( .A(n_692), .Y(n_798) );
AND2x2_ASAP7_75t_L g827 ( .A(n_692), .B(n_746), .Y(n_827) );
INVx1_ASAP7_75t_L g861 ( .A(n_693), .Y(n_861) );
INVx2_ASAP7_75t_L g920 ( .A(n_693), .Y(n_920) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_694), .B(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g847 ( .A(n_694), .Y(n_847) );
INVx2_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx2_ASAP7_75t_L g747 ( .A(n_695), .Y(n_747) );
HB1xp67_ASAP7_75t_L g834 ( .A(n_695), .Y(n_834) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx2_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
NAND2x1_ASAP7_75t_SL g877 ( .A(n_698), .B(n_772), .Y(n_877) );
INVx1_ASAP7_75t_L g725 ( .A(n_699), .Y(n_725) );
INVx1_ASAP7_75t_L g821 ( .A(n_699), .Y(n_821) );
INVx2_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
OR2x2_ASAP7_75t_L g851 ( .A(n_701), .B(n_852), .Y(n_851) );
OR2x2_ASAP7_75t_SL g922 ( .A(n_701), .B(n_824), .Y(n_922) );
INVx2_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
AND2x2_ASAP7_75t_L g842 ( .A(n_702), .B(n_843), .Y(n_842) );
OAI32xp33_ASAP7_75t_L g703 ( .A1(n_704), .A2(n_709), .A3(n_712), .B1(n_719), .B2(n_730), .Y(n_703) );
OAI22xp33_ASAP7_75t_SL g761 ( .A1(n_704), .A2(n_762), .B1(n_765), .B2(n_767), .Y(n_761) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
BUFx3_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx3_ASAP7_75t_L g731 ( .A(n_706), .Y(n_731) );
AND2x4_ASAP7_75t_L g924 ( .A(n_706), .B(n_793), .Y(n_924) );
AND2x2_ASAP7_75t_L g931 ( .A(n_706), .B(n_907), .Y(n_931) );
INVx1_ASAP7_75t_L g779 ( .A(n_707), .Y(n_779) );
INVx2_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVxp67_ASAP7_75t_L g806 ( .A(n_708), .Y(n_806) );
INVx1_ASAP7_75t_L g849 ( .A(n_708), .Y(n_849) );
HB1xp67_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx2_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g816 ( .A(n_711), .B(n_817), .Y(n_816) );
AND2x2_ASAP7_75t_L g887 ( .A(n_711), .B(n_825), .Y(n_887) );
NAND2xp5_ASAP7_75t_L g913 ( .A(n_711), .B(n_725), .Y(n_913) );
INVx2_ASAP7_75t_SL g712 ( .A(n_713), .Y(n_712) );
AND2x2_ASAP7_75t_L g841 ( .A(n_713), .B(n_842), .Y(n_841) );
AND2x2_ASAP7_75t_L g713 ( .A(n_714), .B(n_716), .Y(n_713) );
INVx2_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g903 ( .A(n_716), .Y(n_903) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
OR2x2_ASAP7_75t_L g852 ( .A(n_717), .B(n_821), .Y(n_852) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_720), .B(n_726), .Y(n_719) );
AND2x2_ASAP7_75t_L g720 ( .A(n_721), .B(n_723), .Y(n_720) );
HB1xp67_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx2_ASAP7_75t_L g735 ( .A(n_722), .Y(n_735) );
AND2x2_ASAP7_75t_L g763 ( .A(n_722), .B(n_764), .Y(n_763) );
OR2x2_ASAP7_75t_L g785 ( .A(n_722), .B(n_782), .Y(n_785) );
NOR2xp33_ASAP7_75t_L g929 ( .A(n_722), .B(n_930), .Y(n_929) );
INVx1_ASAP7_75t_L g890 ( .A(n_723), .Y(n_890) );
AND2x2_ASAP7_75t_L g723 ( .A(n_724), .B(n_725), .Y(n_723) );
INVx2_ASAP7_75t_L g896 ( .A(n_724), .Y(n_896) );
AND2x2_ASAP7_75t_L g918 ( .A(n_724), .B(n_735), .Y(n_918) );
HB1xp67_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g755 ( .A(n_727), .Y(n_755) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVxp67_ASAP7_75t_L g812 ( .A(n_728), .Y(n_812) );
OR2x2_ASAP7_75t_L g868 ( .A(n_728), .B(n_869), .Y(n_868) );
INVx1_ASAP7_75t_L g830 ( .A(n_729), .Y(n_830) );
A2O1A1Ixp33_ASAP7_75t_L g914 ( .A1(n_730), .A2(n_915), .B(n_917), .C(n_919), .Y(n_914) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
AOI211xp5_ASAP7_75t_L g732 ( .A1(n_733), .A2(n_740), .B(n_748), .C(n_761), .Y(n_732) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_735), .B(n_736), .Y(n_734) );
INVx1_ASAP7_75t_L g817 ( .A(n_735), .Y(n_817) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx2_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
AND2x4_ASAP7_75t_L g863 ( .A(n_738), .B(n_825), .Y(n_863) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
NAND2xp67_ASAP7_75t_L g741 ( .A(n_742), .B(n_744), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_742), .B(n_776), .Y(n_775) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_743), .B(n_795), .Y(n_794) );
AND2x2_ASAP7_75t_L g865 ( .A(n_743), .B(n_866), .Y(n_865) );
AND2x4_ASAP7_75t_SL g744 ( .A(n_745), .B(n_746), .Y(n_744) );
INVx1_ASAP7_75t_L g875 ( .A(n_745), .Y(n_875) );
AND2x2_ASAP7_75t_L g932 ( .A(n_745), .B(n_807), .Y(n_932) );
BUFx3_ASAP7_75t_L g795 ( .A(n_746), .Y(n_795) );
NAND2xp5_ASAP7_75t_L g897 ( .A(n_746), .B(n_766), .Y(n_897) );
NAND2xp5_ASAP7_75t_L g886 ( .A(n_747), .B(n_814), .Y(n_886) );
OAI32xp33_ASAP7_75t_L g748 ( .A1(n_749), .A2(n_751), .A3(n_754), .B1(n_756), .B2(n_758), .Y(n_748) );
INVx2_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
NAND2x1_ASAP7_75t_L g906 ( .A(n_752), .B(n_907), .Y(n_906) );
INVx2_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx2_ASAP7_75t_L g866 ( .A(n_753), .Y(n_866) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVx1_ASAP7_75t_L g911 ( .A(n_755), .Y(n_911) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
INVxp67_ASAP7_75t_SL g758 ( .A(n_759), .Y(n_758) );
NAND2x2_ASAP7_75t_L g762 ( .A(n_759), .B(n_763), .Y(n_762) );
BUFx3_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g835 ( .A(n_760), .B(n_836), .Y(n_835) );
AND2x4_ASAP7_75t_L g853 ( .A(n_760), .B(n_854), .Y(n_853) );
OR2x2_ASAP7_75t_L g823 ( .A(n_764), .B(n_824), .Y(n_823) );
INVx2_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g832 ( .A(n_766), .B(n_833), .Y(n_832) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_768), .B(n_772), .Y(n_767) );
INVxp67_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
INVx1_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
AND2x2_ASAP7_75t_L g916 ( .A(n_770), .B(n_836), .Y(n_916) );
BUFx2_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
AND2x2_ASAP7_75t_L g874 ( .A(n_772), .B(n_820), .Y(n_874) );
INVx1_ASAP7_75t_L g880 ( .A(n_772), .Y(n_880) );
HB1xp67_ASAP7_75t_L g902 ( .A(n_772), .Y(n_902) );
AOI221xp5_ASAP7_75t_L g773 ( .A1(n_774), .A2(n_781), .B1(n_783), .B2(n_789), .C(n_800), .Y(n_773) );
INVx1_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
INVx1_ASAP7_75t_L g891 ( .A(n_776), .Y(n_891) );
INVx2_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
AND2x2_ASAP7_75t_L g925 ( .A(n_777), .B(n_926), .Y(n_925) );
NAND2x1p5_ASAP7_75t_L g777 ( .A(n_778), .B(n_780), .Y(n_777) );
INVx1_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
NOR2xp33_ASAP7_75t_L g833 ( .A(n_779), .B(n_834), .Y(n_833) );
INVx1_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
INVx2_ASAP7_75t_L g843 ( .A(n_782), .Y(n_843) );
INVx1_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
OR2x2_ASAP7_75t_L g784 ( .A(n_785), .B(n_786), .Y(n_784) );
INVx1_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
HB1xp67_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
AND2x2_ASAP7_75t_L g894 ( .A(n_788), .B(n_843), .Y(n_894) );
NAND3xp33_ASAP7_75t_SL g789 ( .A(n_790), .B(n_794), .C(n_796), .Y(n_789) );
INVx2_ASAP7_75t_L g857 ( .A(n_790), .Y(n_857) );
OR2x2_ASAP7_75t_L g790 ( .A(n_791), .B(n_792), .Y(n_790) );
OR2x2_ASAP7_75t_L g860 ( .A(n_791), .B(n_861), .Y(n_860) );
INVx1_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
INVx1_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
AND2x2_ASAP7_75t_L g797 ( .A(n_798), .B(n_799), .Y(n_797) );
AOI21xp33_ASAP7_75t_L g800 ( .A1(n_801), .A2(n_802), .B(n_804), .Y(n_800) );
INVx2_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
OAI221xp5_ASAP7_75t_L g872 ( .A1(n_804), .A2(n_873), .B1(n_878), .B2(n_879), .C(n_881), .Y(n_872) );
INVx2_ASAP7_75t_SL g804 ( .A(n_805), .Y(n_804) );
AND2x2_ASAP7_75t_L g805 ( .A(n_806), .B(n_807), .Y(n_805) );
INVx1_ASAP7_75t_L g878 ( .A(n_807), .Y(n_878) );
NAND2xp5_ASAP7_75t_L g926 ( .A(n_807), .B(n_866), .Y(n_926) );
AOI221xp5_ASAP7_75t_L g808 ( .A1(n_809), .A2(n_815), .B1(n_818), .B2(n_826), .C(n_828), .Y(n_808) );
HB1xp67_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
INVx2_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
NAND2xp5_ASAP7_75t_L g811 ( .A(n_812), .B(n_813), .Y(n_811) );
INVx1_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
INVx1_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
NAND3xp33_ASAP7_75t_L g818 ( .A(n_819), .B(n_822), .C(n_823), .Y(n_818) );
INVxp67_ASAP7_75t_SL g820 ( .A(n_821), .Y(n_820) );
OAI221xp5_ASAP7_75t_SL g921 ( .A1(n_822), .A2(n_922), .B1(n_923), .B2(n_925), .C(n_927), .Y(n_921) );
OAI211xp5_ASAP7_75t_L g905 ( .A1(n_823), .A2(n_906), .B(n_908), .C(n_914), .Y(n_905) );
OR2x2_ASAP7_75t_L g879 ( .A(n_824), .B(n_880), .Y(n_879) );
INVx2_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
HB1xp67_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
NAND2xp5_ASAP7_75t_L g893 ( .A(n_827), .B(n_894), .Y(n_893) );
AOI21xp33_ASAP7_75t_L g828 ( .A1(n_829), .A2(n_832), .B(n_835), .Y(n_828) );
NAND2xp5_ASAP7_75t_L g829 ( .A(n_830), .B(n_831), .Y(n_829) );
NAND3xp33_ASAP7_75t_L g837 ( .A(n_838), .B(n_871), .C(n_904), .Y(n_837) );
NOR2xp33_ASAP7_75t_L g838 ( .A(n_839), .B(n_855), .Y(n_838) );
INVxp67_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
INVx1_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
OR2x2_ASAP7_75t_L g846 ( .A(n_847), .B(n_848), .Y(n_846) );
INVx1_ASAP7_75t_L g869 ( .A(n_849), .Y(n_869) );
INVxp67_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
HB1xp67_ASAP7_75t_L g892 ( .A(n_852), .Y(n_892) );
NOR2xp33_ASAP7_75t_L g862 ( .A(n_853), .B(n_863), .Y(n_862) );
A2O1A1Ixp33_ASAP7_75t_L g855 ( .A1(n_856), .A2(n_858), .B(n_862), .C(n_864), .Y(n_855) );
INVx1_ASAP7_75t_L g856 ( .A(n_857), .Y(n_856) );
INVx1_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
INVx1_ASAP7_75t_L g859 ( .A(n_860), .Y(n_859) );
AOI22xp5_ASAP7_75t_L g864 ( .A1(n_863), .A2(n_865), .B1(n_867), .B2(n_870), .Y(n_864) );
INVx1_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
AOI22xp33_ASAP7_75t_L g927 ( .A1(n_870), .A2(n_928), .B1(n_931), .B2(n_932), .Y(n_927) );
NOR3xp33_ASAP7_75t_L g871 ( .A(n_872), .B(n_888), .C(n_895), .Y(n_871) );
AOI21xp33_ASAP7_75t_L g873 ( .A1(n_874), .A2(n_875), .B(n_876), .Y(n_873) );
INVxp67_ASAP7_75t_SL g876 ( .A(n_877), .Y(n_876) );
OAI21xp5_ASAP7_75t_L g881 ( .A1(n_882), .A2(n_885), .B(n_887), .Y(n_881) );
INVx2_ASAP7_75t_L g882 ( .A(n_883), .Y(n_882) );
INVx2_ASAP7_75t_SL g885 ( .A(n_886), .Y(n_885) );
OAI221xp5_ASAP7_75t_L g888 ( .A1(n_889), .A2(n_890), .B1(n_891), .B2(n_892), .C(n_893), .Y(n_888) );
INVx2_ASAP7_75t_L g910 ( .A(n_894), .Y(n_910) );
O2A1O1Ixp33_ASAP7_75t_L g895 ( .A1(n_896), .A2(n_897), .B(n_898), .C(n_903), .Y(n_895) );
OAI21xp5_ASAP7_75t_L g898 ( .A1(n_899), .A2(n_900), .B(n_902), .Y(n_898) );
AOI22xp33_ASAP7_75t_L g908 ( .A1(n_899), .A2(n_909), .B1(n_911), .B2(n_912), .Y(n_908) );
INVxp67_ASAP7_75t_L g900 ( .A(n_901), .Y(n_900) );
NOR2xp33_ASAP7_75t_L g904 ( .A(n_905), .B(n_921), .Y(n_904) );
INVx1_ASAP7_75t_L g909 ( .A(n_910), .Y(n_909) );
INVx1_ASAP7_75t_L g912 ( .A(n_913), .Y(n_912) );
HB1xp67_ASAP7_75t_L g915 ( .A(n_916), .Y(n_915) );
AND2x2_ASAP7_75t_L g917 ( .A(n_916), .B(n_918), .Y(n_917) );
AND2x2_ASAP7_75t_L g928 ( .A(n_916), .B(n_929), .Y(n_928) );
INVx2_ASAP7_75t_L g919 ( .A(n_920), .Y(n_919) );
INVx1_ASAP7_75t_L g923 ( .A(n_924), .Y(n_923) );
INVx1_ASAP7_75t_L g965 ( .A(n_933), .Y(n_965) );
INVx1_ASAP7_75t_L g934 ( .A(n_935), .Y(n_934) );
INVx1_ASAP7_75t_L g937 ( .A(n_938), .Y(n_937) );
NAND3xp33_ASAP7_75t_L g942 ( .A(n_943), .B(n_949), .C(n_954), .Y(n_942) );
INVx1_ASAP7_75t_L g943 ( .A(n_944), .Y(n_943) );
NOR2xp33_ASAP7_75t_L g944 ( .A(n_945), .B(n_946), .Y(n_944) );
BUFx3_ASAP7_75t_L g946 ( .A(n_947), .Y(n_946) );
HB1xp67_ASAP7_75t_L g947 ( .A(n_948), .Y(n_947) );
INVx1_ASAP7_75t_L g984 ( .A(n_949), .Y(n_984) );
INVx3_ASAP7_75t_L g950 ( .A(n_951), .Y(n_950) );
BUFx6f_ASAP7_75t_L g971 ( .A(n_951), .Y(n_971) );
BUFx6f_ASAP7_75t_L g951 ( .A(n_952), .Y(n_951) );
CKINVDCx5p33_ASAP7_75t_R g954 ( .A(n_955), .Y(n_954) );
CKINVDCx5p33_ASAP7_75t_R g955 ( .A(n_956), .Y(n_955) );
BUFx3_ASAP7_75t_L g956 ( .A(n_957), .Y(n_956) );
CKINVDCx20_ASAP7_75t_R g983 ( .A(n_957), .Y(n_983) );
NAND2xp5_ASAP7_75t_SL g958 ( .A(n_959), .B(n_965), .Y(n_958) );
OAI21xp5_ASAP7_75t_L g959 ( .A1(n_960), .A2(n_961), .B(n_963), .Y(n_959) );
BUFx4_ASAP7_75t_SL g961 ( .A(n_962), .Y(n_961) );
OAI21x1_ASAP7_75t_L g966 ( .A1(n_967), .A2(n_972), .B(n_981), .Y(n_966) );
HB1xp67_ASAP7_75t_SL g967 ( .A(n_968), .Y(n_967) );
INVx1_ASAP7_75t_L g968 ( .A(n_969), .Y(n_968) );
INVx2_ASAP7_75t_L g969 ( .A(n_970), .Y(n_969) );
INVx5_ASAP7_75t_SL g970 ( .A(n_971), .Y(n_970) );
XOR2x1_ASAP7_75t_L g972 ( .A(n_973), .B(n_978), .Y(n_972) );
INVx2_ASAP7_75t_L g973 ( .A(n_974), .Y(n_973) );
NOR2xp33_ASAP7_75t_L g981 ( .A(n_982), .B(n_984), .Y(n_981) );
CKINVDCx20_ASAP7_75t_R g982 ( .A(n_983), .Y(n_982) );
endmodule