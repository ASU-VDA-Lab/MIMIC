module fake_jpeg_20431_n_135 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_135);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_135;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_93;
wire n_91;
wire n_54;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_42),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_18),
.B(n_16),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_21),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_20),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_9),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_38),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

BUFx16f_ASAP7_75t_L g57 ( 
.A(n_0),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_3),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_24),
.Y(n_60)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

BUFx24_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_7),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_63),
.Y(n_67)
);

CKINVDCx6p67_ASAP7_75t_R g82 ( 
.A(n_67),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_63),
.Y(n_68)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

O2A1O1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_69),
.A2(n_59),
.B(n_65),
.C(n_47),
.Y(n_75)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_62),
.Y(n_71)
);

AOI21xp33_ASAP7_75t_L g78 ( 
.A1(n_71),
.A2(n_66),
.B(n_53),
.Y(n_78)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

BUFx10_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_75),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_73),
.A2(n_46),
.B1(n_64),
.B2(n_66),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_76),
.B(n_80),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_78),
.A2(n_48),
.B(n_60),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_71),
.B(n_45),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_72),
.A2(n_61),
.B1(n_51),
.B2(n_52),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_81),
.B(n_74),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_86),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_80),
.B(n_79),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_88),
.B(n_93),
.Y(n_99)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_89),
.B(n_55),
.Y(n_97)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_84),
.Y(n_90)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_82),
.Y(n_91)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_49),
.Y(n_93)
);

INVx2_ASAP7_75t_R g94 ( 
.A(n_83),
.Y(n_94)
);

OA21x2_ASAP7_75t_L g107 ( 
.A1(n_94),
.A2(n_6),
.B(n_8),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_83),
.B(n_54),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_95),
.B(n_58),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_87),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_96),
.B(n_100),
.Y(n_111)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_97),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_56),
.Y(n_98)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_92),
.B(n_0),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_1),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_102),
.B(n_103),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_94),
.B(n_1),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_104),
.B(n_13),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_105),
.A2(n_107),
.B1(n_106),
.B2(n_101),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_107),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_108),
.B(n_109),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_99),
.B(n_14),
.Y(n_109)
);

OA21x2_ASAP7_75t_L g117 ( 
.A1(n_110),
.A2(n_17),
.B(n_23),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_99),
.B(n_15),
.Y(n_114)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_114),
.Y(n_120)
);

O2A1O1Ixp33_ASAP7_75t_L g124 ( 
.A1(n_117),
.A2(n_118),
.B(n_122),
.C(n_112),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_115),
.Y(n_118)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_116),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_121),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_111),
.Y(n_122)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_124),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_125),
.A2(n_123),
.B(n_121),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_126),
.B(n_113),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_127),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_128),
.A2(n_120),
.B1(n_108),
.B2(n_119),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_129),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_26),
.Y(n_131)
);

OAI321xp33_ASAP7_75t_L g132 ( 
.A1(n_131),
.A2(n_27),
.A3(n_28),
.B1(n_30),
.B2(n_31),
.C(n_35),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_132),
.A2(n_36),
.B(n_40),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_133),
.B(n_41),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_43),
.Y(n_135)
);


endmodule