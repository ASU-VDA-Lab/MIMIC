module fake_jpeg_21825_n_43 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_43);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_43;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_40;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_32;

INVx3_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_20),
.B(n_15),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_23),
.B(n_0),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_27),
.B(n_4),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_23),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_28),
.A2(n_1),
.B1(n_2),
.B2(n_25),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_22),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_29),
.B(n_24),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_30),
.B(n_33),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_32),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_5),
.Y(n_34)
);

HAxp5_ASAP7_75t_SL g36 ( 
.A(n_34),
.B(n_35),
.CON(n_36),
.SN(n_36)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_27),
.B(n_6),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_37),
.B(n_31),
.C(n_12),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_39),
.A2(n_31),
.B1(n_38),
.B2(n_36),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_40),
.B(n_36),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_41),
.A2(n_11),
.B1(n_13),
.B2(n_16),
.Y(n_42)
);

AO21x1_ASAP7_75t_L g43 ( 
.A1(n_42),
.A2(n_19),
.B(n_17),
.Y(n_43)
);


endmodule