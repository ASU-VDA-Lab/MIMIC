module fake_jpeg_18525_n_55 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_55);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_55;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_51;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

NOR2xp33_ASAP7_75t_L g8 ( 
.A(n_3),
.B(n_7),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

INVx3_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

INVx3_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

INVx8_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_2),
.B(n_3),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_5),
.B(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_15),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_17),
.B(n_22),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g18 ( 
.A1(n_13),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_18)
);

OAI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_18),
.A2(n_10),
.B1(n_13),
.B2(n_1),
.Y(n_26)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_20),
.B(n_21),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_16),
.B(n_0),
.Y(n_21)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

OA22x2_ASAP7_75t_L g34 ( 
.A1(n_26),
.A2(n_22),
.B1(n_18),
.B2(n_19),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_17),
.B(n_16),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_23),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_33),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_SL g33 ( 
.A1(n_24),
.A2(n_21),
.B(n_17),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_34),
.A2(n_23),
.B1(n_20),
.B2(n_28),
.Y(n_37)
);

AO22x1_ASAP7_75t_L g35 ( 
.A1(n_24),
.A2(n_21),
.B1(n_20),
.B2(n_22),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_35),
.B(n_30),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_37),
.A2(n_38),
.B1(n_14),
.B2(n_2),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_34),
.A2(n_10),
.B1(n_13),
.B2(n_19),
.Y(n_38)
);

OAI21xp33_ASAP7_75t_L g45 ( 
.A1(n_39),
.A2(n_40),
.B(n_1),
.Y(n_45)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_39),
.A2(n_35),
.B1(n_14),
.B2(n_9),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_43),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_41),
.B(n_9),
.C(n_12),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_44),
.B(n_38),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_45),
.B(n_6),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_48),
.B(n_8),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_50),
.B(n_36),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_51),
.A2(n_52),
.B1(n_47),
.B2(n_44),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_49),
.B(n_43),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_53),
.B(n_37),
.C(n_12),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g55 ( 
.A(n_54),
.B(n_12),
.Y(n_55)
);


endmodule