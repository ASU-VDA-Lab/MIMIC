module fake_jpeg_20723_n_154 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_154);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_154;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_149;
wire n_87;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_4),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_41),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_9),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_24),
.B(n_8),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_46),
.Y(n_56)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_7),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_14),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_13),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_6),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_8),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_39),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_15),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_10),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_34),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_31),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

HB1xp67_ASAP7_75t_L g77 ( 
.A(n_20),
.Y(n_77)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_62),
.B(n_19),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_79),
.B(n_80),
.Y(n_92)
);

AOI21xp33_ASAP7_75t_L g80 ( 
.A1(n_55),
.A2(n_51),
.B(n_64),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_81),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_82),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_49),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_83),
.A2(n_57),
.B1(n_52),
.B2(n_50),
.Y(n_86)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_84),
.Y(n_88)
);

INVx3_ASAP7_75t_SL g85 ( 
.A(n_69),
.Y(n_85)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

NAND3xp33_ASAP7_75t_L g99 ( 
.A(n_86),
.B(n_66),
.C(n_77),
.Y(n_99)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_89),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_85),
.A2(n_81),
.B1(n_78),
.B2(n_84),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_90),
.A2(n_96),
.B1(n_61),
.B2(n_63),
.Y(n_109)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_85),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_79),
.A2(n_76),
.B1(n_71),
.B2(n_58),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_92),
.B(n_72),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_98),
.B(n_100),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_99),
.A2(n_26),
.B(n_47),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_96),
.B(n_53),
.Y(n_100)
);

INVx4_ASAP7_75t_SL g101 ( 
.A(n_95),
.Y(n_101)
);

INVx13_ASAP7_75t_L g117 ( 
.A(n_101),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_94),
.B(n_54),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_103),
.B(n_108),
.Y(n_114)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_94),
.Y(n_104)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_104),
.Y(n_111)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_93),
.Y(n_105)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_105),
.Y(n_120)
);

CKINVDCx5p33_ASAP7_75t_R g106 ( 
.A(n_93),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g110 ( 
.A(n_106),
.Y(n_110)
);

BUFx16f_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_107),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_87),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_109),
.A2(n_71),
.B1(n_63),
.B2(n_61),
.Y(n_121)
);

AND2x6_ASAP7_75t_L g112 ( 
.A(n_109),
.B(n_77),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_112),
.B(n_121),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_103),
.B(n_75),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_113),
.B(n_0),
.C(n_1),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_97),
.A2(n_68),
.B1(n_70),
.B2(n_74),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_116),
.B(n_119),
.Y(n_126)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_102),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_118),
.B(n_123),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_107),
.B(n_73),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_122),
.A2(n_124),
.B(n_56),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_100),
.A2(n_59),
.B1(n_60),
.B2(n_65),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_100),
.B(n_0),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_111),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_127),
.B(n_128),
.Y(n_137)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_120),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_114),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_129),
.A2(n_130),
.B(n_131),
.Y(n_138)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_114),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_133),
.B(n_125),
.Y(n_139)
);

OAI22xp33_ASAP7_75t_L g135 ( 
.A1(n_110),
.A2(n_18),
.B1(n_42),
.B2(n_38),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_135),
.A2(n_136),
.B1(n_117),
.B2(n_2),
.Y(n_141)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_119),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_139),
.B(n_133),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_132),
.A2(n_110),
.B1(n_124),
.B2(n_115),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_140),
.A2(n_141),
.B1(n_135),
.B2(n_134),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_142),
.A2(n_143),
.B1(n_126),
.B2(n_139),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_144),
.A2(n_138),
.B(n_137),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_145),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_16),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_17),
.C(n_37),
.Y(n_148)
);

OR2x2_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_11),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_43),
.Y(n_150)
);

AOI322xp5_ASAP7_75t_L g151 ( 
.A1(n_150),
.A2(n_36),
.A3(n_32),
.B1(n_28),
.B2(n_27),
.C1(n_22),
.C2(n_6),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_1),
.Y(n_152)
);

OAI221xp5_ASAP7_75t_L g153 ( 
.A1(n_152),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.C(n_5),
.Y(n_153)
);

BUFx24_ASAP7_75t_SL g154 ( 
.A(n_153),
.Y(n_154)
);


endmodule