module fake_jpeg_9268_n_204 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_204);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_204;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx4f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx11_ASAP7_75t_SL g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_33),
.Y(n_34)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_38),
.Y(n_50)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_46),
.Y(n_51)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_40),
.A2(n_36),
.B1(n_37),
.B2(n_28),
.Y(n_70)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_43),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_24),
.B(n_0),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_1),
.Y(n_58)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_32),
.Y(n_60)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_39),
.A2(n_20),
.B1(n_24),
.B2(n_28),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_47),
.A2(n_19),
.B1(n_16),
.B2(n_32),
.Y(n_83)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_49),
.B(n_52),
.Y(n_71)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_53),
.B(n_57),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_25),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_55),
.B(n_58),
.Y(n_72)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_59),
.B(n_67),
.Y(n_79)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_35),
.B(n_25),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_64),
.B(n_1),
.Y(n_94)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_37),
.B(n_19),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_69),
.B(n_31),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_70),
.A2(n_31),
.B1(n_30),
.B2(n_21),
.Y(n_95)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_75),
.B(n_78),
.Y(n_103)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_80),
.B(n_82),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_51),
.B(n_40),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_83),
.A2(n_84),
.B1(n_95),
.B2(n_48),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_70),
.A2(n_40),
.B1(n_16),
.B2(n_18),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_85),
.B(n_86),
.Y(n_115)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_66),
.A2(n_17),
.B1(n_21),
.B2(n_30),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_87),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_58),
.B(n_26),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_89),
.B(n_2),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_68),
.A2(n_17),
.B(n_34),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_90),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_91),
.B(n_93),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_92),
.Y(n_101)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_62),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_94),
.B(n_97),
.Y(n_104)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_62),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_96),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_66),
.B(n_1),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_76),
.A2(n_48),
.B1(n_67),
.B2(n_59),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_98),
.A2(n_102),
.B1(n_87),
.B2(n_96),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_99),
.B(n_3),
.Y(n_138)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_100),
.B(n_108),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_82),
.B(n_63),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_106),
.B(n_111),
.Y(n_125)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_79),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_71),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_109),
.B(n_110),
.Y(n_139)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_97),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g111 ( 
.A(n_83),
.B(n_52),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_89),
.B(n_2),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_113),
.B(n_116),
.Y(n_130)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_114),
.B(n_118),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_94),
.B(n_3),
.Y(n_116)
);

BUFx24_ASAP7_75t_SL g118 ( 
.A(n_78),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_115),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_120),
.B(n_121),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_103),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g122 ( 
.A(n_101),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_122),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_109),
.B(n_72),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_123),
.B(n_133),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_124),
.A2(n_129),
.B1(n_107),
.B2(n_114),
.Y(n_140)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_106),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_126),
.B(n_132),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_105),
.A2(n_84),
.B1(n_76),
.B2(n_73),
.Y(n_129)
);

A2O1A1O1Ixp25_ASAP7_75t_L g131 ( 
.A1(n_112),
.A2(n_94),
.B(n_90),
.C(n_86),
.D(n_81),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_131),
.A2(n_137),
.B(n_125),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_99),
.B(n_81),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_100),
.B(n_74),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_113),
.B(n_88),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_134),
.B(n_137),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_117),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_135),
.B(n_111),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_119),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_136),
.A2(n_119),
.B(n_101),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_111),
.B(n_88),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_138),
.B(n_15),
.Y(n_155)
);

AOI221xp5_ASAP7_75t_L g166 ( 
.A1(n_140),
.A2(n_148),
.B1(n_12),
.B2(n_10),
.C(n_7),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_132),
.B(n_110),
.C(n_108),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_142),
.B(n_154),
.C(n_130),
.Y(n_157)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_143),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_126),
.A2(n_107),
.B1(n_104),
.B2(n_116),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_145),
.A2(n_153),
.B1(n_4),
.B2(n_5),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_149),
.A2(n_139),
.B(n_136),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_128),
.B(n_104),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_150),
.B(n_151),
.Y(n_160)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_127),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_125),
.A2(n_104),
.B1(n_74),
.B2(n_119),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_92),
.C(n_41),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_155),
.B(n_15),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_134),
.B(n_4),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_156),
.B(n_122),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_157),
.B(n_159),
.C(n_161),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_158),
.B(n_162),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_144),
.B(n_138),
.C(n_120),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_144),
.B(n_131),
.C(n_121),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_148),
.A2(n_52),
.B(n_41),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_163),
.B(n_146),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_164),
.B(n_166),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_147),
.A2(n_122),
.B1(n_5),
.B2(n_6),
.Y(n_165)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_165),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_142),
.B(n_122),
.C(n_12),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_167),
.B(n_168),
.Y(n_179)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_160),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_173),
.B(n_174),
.Y(n_185)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_168),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_161),
.A2(n_147),
.B1(n_153),
.B2(n_154),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_176),
.A2(n_145),
.B1(n_169),
.B2(n_159),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_167),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_177),
.A2(n_178),
.B(n_156),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_171),
.B(n_157),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_180),
.B(n_187),
.C(n_175),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_181),
.B(n_183),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_176),
.A2(n_172),
.B1(n_170),
.B2(n_146),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_182),
.A2(n_186),
.B1(n_9),
.B2(n_180),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_170),
.A2(n_151),
.B1(n_152),
.B2(n_171),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_184),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_179),
.A2(n_149),
.B1(n_141),
.B2(n_164),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_179),
.B(n_155),
.C(n_8),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_188),
.B(n_192),
.C(n_193),
.Y(n_196)
);

INVx6_ASAP7_75t_L g190 ( 
.A(n_185),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_190),
.B(n_9),
.Y(n_197)
);

NOR2xp67_ASAP7_75t_L g191 ( 
.A(n_181),
.B(n_175),
.Y(n_191)
);

OR2x2_ASAP7_75t_L g195 ( 
.A(n_191),
.B(n_186),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_193),
.A2(n_182),
.B(n_187),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_194),
.B(n_196),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_195),
.B(n_197),
.Y(n_198)
);

NOR2xp67_ASAP7_75t_SL g200 ( 
.A(n_195),
.B(n_192),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_200),
.B(n_189),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_201),
.A2(n_202),
.B(n_190),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_198),
.B(n_188),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_203),
.B(n_199),
.Y(n_204)
);


endmodule