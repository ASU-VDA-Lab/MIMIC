module fake_netlist_6_2543_n_985 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_985);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_985;

wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_881;
wire n_875;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_828;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_933;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_978;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_969;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_628;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_845;
wire n_255;
wire n_807;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_955;
wire n_865;
wire n_893;
wire n_214;
wire n_925;
wire n_485;
wire n_443;
wire n_246;
wire n_892;
wire n_768;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_669;
wire n_200;
wire n_447;
wire n_872;
wire n_198;
wire n_300;
wire n_222;
wire n_248;
wire n_517;
wire n_718;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_901;
wire n_504;
wire n_923;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_945;
wire n_977;
wire n_603;
wire n_957;
wire n_235;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_658;
wire n_616;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_822;
wire n_693;
wire n_631;
wire n_516;
wire n_720;
wire n_525;
wire n_758;
wire n_842;
wire n_611;
wire n_943;
wire n_491;
wire n_878;
wire n_656;
wire n_772;
wire n_843;
wire n_797;
wire n_666;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_844;
wire n_448;
wire n_886;
wire n_953;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_236;
wire n_653;
wire n_887;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_224;
wire n_926;
wire n_927;
wire n_839;
wire n_734;
wire n_708;
wire n_196;
wire n_919;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_800;
wire n_779;
wire n_929;
wire n_460;
wire n_907;
wire n_854;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_594;
wire n_565;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_619;
wire n_885;
wire n_216;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_527;
wire n_474;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_981;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_821;
wire n_325;
wire n_938;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_964;
wire n_982;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_707;
wire n_322;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_692;
wire n_733;
wire n_754;
wire n_941;
wire n_975;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_811;
wire n_882;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_257;
wire n_920;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_816;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_205;
wire n_604;
wire n_848;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_438;
wire n_267;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_983;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_961;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_457;
wire n_391;
wire n_697;
wire n_687;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_897;
wire n_900;
wire n_846;
wire n_501;
wire n_841;
wire n_956;
wire n_960;
wire n_531;
wire n_827;
wire n_508;
wire n_361;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_332;
wire n_891;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_664;
wire n_949;
wire n_678;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_185),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_117),
.Y(n_196)
);

BUFx10_ASAP7_75t_L g197 ( 
.A(n_157),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_139),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_28),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_5),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_61),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_22),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_188),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_125),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_27),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_192),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_20),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_6),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_87),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_6),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_112),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_114),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_91),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_7),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_155),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_86),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_44),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_133),
.Y(n_218)
);

INVxp67_ASAP7_75t_SL g219 ( 
.A(n_50),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_4),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_17),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g222 ( 
.A(n_145),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_177),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_137),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_52),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_180),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_22),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_25),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_150),
.Y(n_229)
);

CKINVDCx14_ASAP7_75t_R g230 ( 
.A(n_42),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_41),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_80),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_166),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_73),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_161),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_144),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_165),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_126),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_168),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_13),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_14),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_107),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_1),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_57),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_111),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_158),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_51),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_53),
.Y(n_248)
);

CKINVDCx14_ASAP7_75t_R g249 ( 
.A(n_123),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_56),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_189),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_116),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_35),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_58),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_21),
.Y(n_255)
);

BUFx10_ASAP7_75t_L g256 ( 
.A(n_10),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_93),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_59),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_43),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_67),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_17),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_12),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_74),
.Y(n_263)
);

BUFx2_ASAP7_75t_SL g264 ( 
.A(n_190),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_69),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_138),
.Y(n_266)
);

BUFx10_ASAP7_75t_L g267 ( 
.A(n_159),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_115),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_9),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_178),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_31),
.Y(n_271)
);

INVx2_ASAP7_75t_SL g272 ( 
.A(n_68),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_129),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_164),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_240),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_220),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_256),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_195),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_204),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_220),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_220),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_211),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_212),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_220),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_202),
.Y(n_285)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_222),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_215),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_207),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_210),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_216),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_223),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_214),
.Y(n_292)
);

INVxp67_ASAP7_75t_SL g293 ( 
.A(n_274),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_241),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_199),
.Y(n_295)
);

BUFx2_ASAP7_75t_L g296 ( 
.A(n_200),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_255),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_225),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_232),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_272),
.B(n_0),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_261),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_252),
.B(n_258),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_258),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_218),
.Y(n_304)
);

BUFx2_ASAP7_75t_SL g305 ( 
.A(n_201),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_209),
.B(n_233),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_234),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_235),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_226),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_196),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_198),
.Y(n_311)
);

HB1xp67_ASAP7_75t_L g312 ( 
.A(n_205),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_203),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_238),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_239),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_213),
.Y(n_316)
);

INVxp33_ASAP7_75t_SL g317 ( 
.A(n_208),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_201),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_206),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_217),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_206),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_257),
.Y(n_322)
);

INVxp33_ASAP7_75t_L g323 ( 
.A(n_224),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_227),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_245),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_229),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_276),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_306),
.B(n_230),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g329 ( 
.A(n_295),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_280),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_305),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_280),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_281),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_305),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_281),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_284),
.Y(n_336)
);

OA21x2_ASAP7_75t_L g337 ( 
.A1(n_304),
.A2(n_237),
.B(n_231),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_304),
.Y(n_338)
);

OR2x6_ASAP7_75t_L g339 ( 
.A(n_277),
.B(n_264),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_278),
.B(n_249),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_279),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g342 ( 
.A(n_286),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_282),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_284),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_283),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_310),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_310),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_317),
.B(n_222),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_318),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_287),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_311),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_311),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_290),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_313),
.Y(n_354)
);

BUFx2_ASAP7_75t_L g355 ( 
.A(n_291),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_313),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_303),
.Y(n_357)
);

INVxp67_ASAP7_75t_SL g358 ( 
.A(n_286),
.Y(n_358)
);

INVx3_ASAP7_75t_L g359 ( 
.A(n_303),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_316),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_298),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_319),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_316),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_321),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_299),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_320),
.Y(n_366)
);

BUFx8_ASAP7_75t_L g367 ( 
.A(n_296),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_307),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_322),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_308),
.Y(n_370)
);

AND2x4_ASAP7_75t_L g371 ( 
.A(n_286),
.B(n_274),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_320),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_326),
.Y(n_373)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_294),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_312),
.B(n_236),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_326),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_314),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_285),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_315),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_325),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_285),
.Y(n_381)
);

NOR2xp67_ASAP7_75t_L g382 ( 
.A(n_324),
.B(n_242),
.Y(n_382)
);

INVx3_ASAP7_75t_L g383 ( 
.A(n_288),
.Y(n_383)
);

BUFx3_ASAP7_75t_L g384 ( 
.A(n_342),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_328),
.B(n_218),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_371),
.B(n_218),
.Y(n_386)
);

INVx4_ASAP7_75t_L g387 ( 
.A(n_378),
.Y(n_387)
);

INVx3_ASAP7_75t_L g388 ( 
.A(n_338),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_346),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_378),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_347),
.Y(n_391)
);

BUFx3_ASAP7_75t_L g392 ( 
.A(n_342),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_351),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_348),
.B(n_296),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_352),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_354),
.Y(n_396)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_338),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_359),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_371),
.B(n_218),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_356),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_360),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_358),
.B(n_293),
.Y(n_402)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_359),
.Y(n_403)
);

BUFx2_ASAP7_75t_L g404 ( 
.A(n_331),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_371),
.B(n_244),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_340),
.B(n_302),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_366),
.Y(n_407)
);

AND2x6_ASAP7_75t_L g408 ( 
.A(n_375),
.B(n_236),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_341),
.B(n_343),
.Y(n_409)
);

AND2x4_ASAP7_75t_L g410 ( 
.A(n_372),
.B(n_288),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_373),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_382),
.B(n_246),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_359),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_330),
.Y(n_414)
);

INVx3_ASAP7_75t_L g415 ( 
.A(n_337),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_376),
.Y(n_416)
);

INVx3_ASAP7_75t_L g417 ( 
.A(n_337),
.Y(n_417)
);

BUFx2_ASAP7_75t_L g418 ( 
.A(n_331),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_345),
.B(n_254),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_381),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_374),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_345),
.B(n_300),
.Y(n_422)
);

INVx4_ASAP7_75t_L g423 ( 
.A(n_378),
.Y(n_423)
);

INVx3_ASAP7_75t_L g424 ( 
.A(n_337),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_374),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_379),
.B(n_275),
.Y(n_426)
);

INVxp33_ASAP7_75t_L g427 ( 
.A(n_329),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_378),
.Y(n_428)
);

AND2x4_ASAP7_75t_L g429 ( 
.A(n_383),
.B(n_327),
.Y(n_429)
);

INVx1_ASAP7_75t_SL g430 ( 
.A(n_349),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_332),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_333),
.Y(n_432)
);

NOR2x1p5_ASAP7_75t_L g433 ( 
.A(n_380),
.B(n_228),
.Y(n_433)
);

BUFx4f_ASAP7_75t_L g434 ( 
.A(n_374),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_335),
.Y(n_435)
);

INVx4_ASAP7_75t_SL g436 ( 
.A(n_374),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_350),
.B(n_323),
.Y(n_437)
);

INVx2_ASAP7_75t_SL g438 ( 
.A(n_339),
.Y(n_438)
);

AND2x4_ASAP7_75t_L g439 ( 
.A(n_383),
.B(n_289),
.Y(n_439)
);

AND2x6_ASAP7_75t_L g440 ( 
.A(n_383),
.B(n_289),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_336),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_344),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_363),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_363),
.B(n_247),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_350),
.B(n_309),
.Y(n_445)
);

INVx5_ASAP7_75t_L g446 ( 
.A(n_357),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_357),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_339),
.B(n_248),
.Y(n_448)
);

AND2x2_ASAP7_75t_SL g449 ( 
.A(n_355),
.B(n_292),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_339),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_339),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_353),
.Y(n_452)
);

OAI22xp33_ASAP7_75t_SL g453 ( 
.A1(n_334),
.A2(n_262),
.B1(n_243),
.B2(n_271),
.Y(n_453)
);

INVx8_ASAP7_75t_L g454 ( 
.A(n_353),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_361),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_361),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_334),
.Y(n_457)
);

INVxp33_ASAP7_75t_L g458 ( 
.A(n_349),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_406),
.A2(n_377),
.B1(n_370),
.B2(n_365),
.Y(n_459)
);

AOI22xp33_ASAP7_75t_L g460 ( 
.A1(n_440),
.A2(n_417),
.B1(n_424),
.B2(n_415),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_394),
.A2(n_377),
.B1(n_370),
.B2(n_365),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_449),
.B(n_368),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_389),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_447),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_447),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_398),
.Y(n_466)
);

INVx8_ASAP7_75t_L g467 ( 
.A(n_454),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_437),
.B(n_368),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_402),
.B(n_257),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_419),
.B(n_263),
.Y(n_470)
);

INVxp67_ASAP7_75t_L g471 ( 
.A(n_426),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_398),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_449),
.B(n_457),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_391),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_393),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_403),
.B(n_219),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_413),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_403),
.B(n_250),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_457),
.B(n_367),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_403),
.B(n_251),
.Y(n_480)
);

BUFx3_ASAP7_75t_L g481 ( 
.A(n_384),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_429),
.B(n_259),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_419),
.B(n_263),
.Y(n_483)
);

OAI22xp33_ASAP7_75t_L g484 ( 
.A1(n_438),
.A2(n_266),
.B1(n_268),
.B2(n_270),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_429),
.B(n_260),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_457),
.B(n_429),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_395),
.B(n_265),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_422),
.B(n_266),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_413),
.Y(n_489)
);

INVx3_ASAP7_75t_L g490 ( 
.A(n_439),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_457),
.B(n_367),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_396),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_388),
.Y(n_493)
);

AND2x2_ASAP7_75t_SL g494 ( 
.A(n_457),
.B(n_292),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_422),
.B(n_268),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_438),
.B(n_367),
.Y(n_496)
);

AND2x4_ASAP7_75t_SL g497 ( 
.A(n_450),
.B(n_451),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_408),
.A2(n_270),
.B1(n_273),
.B2(n_269),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_450),
.B(n_451),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_453),
.B(n_197),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_448),
.B(n_197),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_400),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_401),
.B(n_297),
.Y(n_503)
);

AND2x6_ASAP7_75t_SL g504 ( 
.A(n_445),
.B(n_409),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_407),
.B(n_221),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_411),
.B(n_297),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_416),
.B(n_301),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_404),
.B(n_197),
.Y(n_508)
);

NOR2x1p5_ASAP7_75t_L g509 ( 
.A(n_452),
.B(n_301),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_418),
.B(n_267),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_388),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_420),
.B(n_415),
.Y(n_512)
);

AND2x2_ASAP7_75t_L g513 ( 
.A(n_427),
.B(n_256),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_415),
.B(n_267),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_388),
.Y(n_515)
);

AOI21xp5_ASAP7_75t_L g516 ( 
.A1(n_417),
.A2(n_267),
.B(n_40),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_417),
.B(n_39),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_397),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_384),
.B(n_256),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_397),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_397),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_444),
.B(n_0),
.Y(n_522)
);

INVx2_ASAP7_75t_SL g523 ( 
.A(n_410),
.Y(n_523)
);

BUFx12f_ASAP7_75t_L g524 ( 
.A(n_433),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_424),
.B(n_45),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_424),
.B(n_46),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_439),
.Y(n_527)
);

AOI22xp33_ASAP7_75t_L g528 ( 
.A1(n_440),
.A2(n_269),
.B1(n_253),
.B2(n_362),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_442),
.B(n_47),
.Y(n_529)
);

BUFx12f_ASAP7_75t_L g530 ( 
.A(n_410),
.Y(n_530)
);

O2A1O1Ixp5_ASAP7_75t_L g531 ( 
.A1(n_386),
.A2(n_98),
.B(n_194),
.C(n_193),
.Y(n_531)
);

AND2x4_ASAP7_75t_L g532 ( 
.A(n_392),
.B(n_48),
.Y(n_532)
);

AOI22xp33_ASAP7_75t_L g533 ( 
.A1(n_440),
.A2(n_253),
.B1(n_364),
.B2(n_362),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_385),
.B(n_49),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_439),
.Y(n_535)
);

BUFx5_ASAP7_75t_L g536 ( 
.A(n_440),
.Y(n_536)
);

OR2x6_ASAP7_75t_L g537 ( 
.A(n_454),
.B(n_455),
.Y(n_537)
);

INVx3_ASAP7_75t_L g538 ( 
.A(n_392),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_443),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_414),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_405),
.B(n_1),
.Y(n_541)
);

OR2x6_ASAP7_75t_L g542 ( 
.A(n_467),
.B(n_454),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_527),
.Y(n_543)
);

BUFx2_ASAP7_75t_L g544 ( 
.A(n_530),
.Y(n_544)
);

BUFx6f_ASAP7_75t_L g545 ( 
.A(n_481),
.Y(n_545)
);

NOR3xp33_ASAP7_75t_SL g546 ( 
.A(n_484),
.B(n_456),
.C(n_405),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_535),
.Y(n_547)
);

BUFx2_ASAP7_75t_L g548 ( 
.A(n_481),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_460),
.B(n_440),
.Y(n_549)
);

AO22x1_ASAP7_75t_L g550 ( 
.A1(n_470),
.A2(n_427),
.B1(n_408),
.B2(n_458),
.Y(n_550)
);

BUFx2_ASAP7_75t_L g551 ( 
.A(n_532),
.Y(n_551)
);

AND2x2_ASAP7_75t_L g552 ( 
.A(n_471),
.B(n_430),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_469),
.B(n_458),
.Y(n_553)
);

BUFx10_ASAP7_75t_L g554 ( 
.A(n_504),
.Y(n_554)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_467),
.Y(n_555)
);

INVx6_ASAP7_75t_L g556 ( 
.A(n_524),
.Y(n_556)
);

BUFx4f_ASAP7_75t_L g557 ( 
.A(n_467),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_540),
.Y(n_558)
);

BUFx8_ASAP7_75t_L g559 ( 
.A(n_468),
.Y(n_559)
);

INVx4_ASAP7_75t_L g560 ( 
.A(n_490),
.Y(n_560)
);

CKINVDCx8_ASAP7_75t_R g561 ( 
.A(n_537),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_469),
.B(n_364),
.Y(n_562)
);

BUFx2_ASAP7_75t_L g563 ( 
.A(n_532),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_540),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_494),
.B(n_408),
.Y(n_565)
);

HB1xp67_ASAP7_75t_L g566 ( 
.A(n_509),
.Y(n_566)
);

OR2x6_ASAP7_75t_L g567 ( 
.A(n_537),
.B(n_454),
.Y(n_567)
);

OAI22xp5_ASAP7_75t_L g568 ( 
.A1(n_470),
.A2(n_483),
.B1(n_495),
.B2(n_488),
.Y(n_568)
);

INVx1_ASAP7_75t_SL g569 ( 
.A(n_494),
.Y(n_569)
);

AND2x4_ASAP7_75t_L g570 ( 
.A(n_497),
.B(n_410),
.Y(n_570)
);

NAND2xp33_ASAP7_75t_R g571 ( 
.A(n_488),
.B(n_369),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_460),
.B(n_440),
.Y(n_572)
);

BUFx6f_ASAP7_75t_L g573 ( 
.A(n_538),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_473),
.B(n_434),
.Y(n_574)
);

NOR3xp33_ASAP7_75t_SL g575 ( 
.A(n_483),
.B(n_412),
.C(n_385),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_490),
.Y(n_576)
);

BUFx3_ASAP7_75t_L g577 ( 
.A(n_497),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_466),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_466),
.Y(n_579)
);

AOI22xp33_ASAP7_75t_L g580 ( 
.A1(n_541),
.A2(n_408),
.B1(n_386),
.B2(n_399),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_505),
.B(n_495),
.Y(n_581)
);

INVx3_ASAP7_75t_L g582 ( 
.A(n_538),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_472),
.Y(n_583)
);

NOR2xp67_ASAP7_75t_L g584 ( 
.A(n_459),
.B(n_399),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_523),
.B(n_461),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_512),
.B(n_414),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_463),
.B(n_408),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_472),
.Y(n_588)
);

INVx4_ASAP7_75t_L g589 ( 
.A(n_537),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_477),
.Y(n_590)
);

AND2x4_ASAP7_75t_L g591 ( 
.A(n_499),
.B(n_431),
.Y(n_591)
);

INVx4_ASAP7_75t_L g592 ( 
.A(n_536),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_462),
.B(n_508),
.Y(n_593)
);

A2O1A1Ixp33_ASAP7_75t_L g594 ( 
.A1(n_541),
.A2(n_432),
.B(n_441),
.C(n_435),
.Y(n_594)
);

INVxp67_ASAP7_75t_SL g595 ( 
.A(n_486),
.Y(n_595)
);

INVx1_ASAP7_75t_SL g596 ( 
.A(n_513),
.Y(n_596)
);

AND2x4_ASAP7_75t_L g597 ( 
.A(n_474),
.B(n_431),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_477),
.Y(n_598)
);

AOI21xp5_ASAP7_75t_L g599 ( 
.A1(n_517),
.A2(n_434),
.B(n_423),
.Y(n_599)
);

NOR3xp33_ASAP7_75t_SL g600 ( 
.A(n_500),
.B(n_412),
.C(n_369),
.Y(n_600)
);

BUFx6f_ASAP7_75t_L g601 ( 
.A(n_486),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_489),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_522),
.B(n_432),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_489),
.Y(n_604)
);

OAI21x1_ASAP7_75t_L g605 ( 
.A1(n_599),
.A2(n_526),
.B(n_525),
.Y(n_605)
);

BUFx6f_ASAP7_75t_L g606 ( 
.A(n_555),
.Y(n_606)
);

AO32x2_ASAP7_75t_L g607 ( 
.A1(n_568),
.A2(n_387),
.A3(n_423),
.B1(n_522),
.B2(n_408),
.Y(n_607)
);

AOI21xp33_ASAP7_75t_L g608 ( 
.A1(n_568),
.A2(n_528),
.B(n_498),
.Y(n_608)
);

BUFx4_ASAP7_75t_SL g609 ( 
.A(n_544),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_581),
.B(n_505),
.Y(n_610)
);

OAI21x1_ASAP7_75t_L g611 ( 
.A1(n_586),
.A2(n_511),
.B(n_493),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_569),
.B(n_533),
.Y(n_612)
);

OAI21x1_ASAP7_75t_L g613 ( 
.A1(n_586),
.A2(n_511),
.B(n_493),
.Y(n_613)
);

AO31x2_ASAP7_75t_L g614 ( 
.A1(n_594),
.A2(n_516),
.A3(n_534),
.B(n_529),
.Y(n_614)
);

AOI21xp5_ASAP7_75t_L g615 ( 
.A1(n_592),
.A2(n_434),
.B(n_514),
.Y(n_615)
);

AOI21xp5_ASAP7_75t_L g616 ( 
.A1(n_592),
.A2(n_476),
.B(n_423),
.Y(n_616)
);

AOI21xp5_ASAP7_75t_L g617 ( 
.A1(n_565),
.A2(n_387),
.B(n_482),
.Y(n_617)
);

INVxp67_ASAP7_75t_SL g618 ( 
.A(n_573),
.Y(n_618)
);

OAI22xp5_ASAP7_75t_L g619 ( 
.A1(n_569),
.A2(n_528),
.B1(n_533),
.B2(n_485),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_603),
.B(n_475),
.Y(n_620)
);

INVx5_ASAP7_75t_L g621 ( 
.A(n_542),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_559),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_558),
.Y(n_623)
);

OAI22xp5_ASAP7_75t_L g624 ( 
.A1(n_551),
.A2(n_563),
.B1(n_572),
.B2(n_549),
.Y(n_624)
);

OAI21xp5_ASAP7_75t_L g625 ( 
.A1(n_549),
.A2(n_465),
.B(n_464),
.Y(n_625)
);

OA21x2_ASAP7_75t_L g626 ( 
.A1(n_603),
.A2(n_465),
.B(n_464),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_596),
.B(n_492),
.Y(n_627)
);

AO31x2_ASAP7_75t_L g628 ( 
.A1(n_587),
.A2(n_572),
.A3(n_564),
.B(n_593),
.Y(n_628)
);

OAI21x1_ASAP7_75t_L g629 ( 
.A1(n_578),
.A2(n_518),
.B(n_515),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_596),
.B(n_502),
.Y(n_630)
);

AOI21xp5_ASAP7_75t_L g631 ( 
.A1(n_574),
.A2(n_387),
.B(n_478),
.Y(n_631)
);

OAI22x1_ASAP7_75t_L g632 ( 
.A1(n_562),
.A2(n_479),
.B1(n_491),
.B2(n_496),
.Y(n_632)
);

BUFx3_ASAP7_75t_L g633 ( 
.A(n_556),
.Y(n_633)
);

OAI21xp5_ASAP7_75t_L g634 ( 
.A1(n_595),
.A2(n_518),
.B(n_515),
.Y(n_634)
);

OAI21x1_ASAP7_75t_L g635 ( 
.A1(n_579),
.A2(n_521),
.B(n_520),
.Y(n_635)
);

AOI22xp5_ASAP7_75t_L g636 ( 
.A1(n_584),
.A2(n_539),
.B1(n_441),
.B2(n_435),
.Y(n_636)
);

OAI21x1_ASAP7_75t_L g637 ( 
.A1(n_583),
.A2(n_521),
.B(n_520),
.Y(n_637)
);

NAND3x1_ASAP7_75t_L g638 ( 
.A(n_553),
.B(n_506),
.C(n_503),
.Y(n_638)
);

BUFx6f_ASAP7_75t_L g639 ( 
.A(n_555),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_597),
.B(n_507),
.Y(n_640)
);

OA21x2_ASAP7_75t_L g641 ( 
.A1(n_588),
.A2(n_539),
.B(n_480),
.Y(n_641)
);

OAI21x1_ASAP7_75t_L g642 ( 
.A1(n_590),
.A2(n_531),
.B(n_425),
.Y(n_642)
);

NOR2x1_ASAP7_75t_L g643 ( 
.A(n_560),
.B(n_487),
.Y(n_643)
);

AOI21xp5_ASAP7_75t_L g644 ( 
.A1(n_580),
.A2(n_536),
.B(n_428),
.Y(n_644)
);

AOI21xp5_ASAP7_75t_L g645 ( 
.A1(n_560),
.A2(n_536),
.B(n_428),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_597),
.B(n_501),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_552),
.B(n_510),
.Y(n_647)
);

OAI21x1_ASAP7_75t_L g648 ( 
.A1(n_598),
.A2(n_604),
.B(n_602),
.Y(n_648)
);

OAI21xp5_ASAP7_75t_L g649 ( 
.A1(n_575),
.A2(n_421),
.B(n_519),
.Y(n_649)
);

AOI21xp5_ASAP7_75t_L g650 ( 
.A1(n_582),
.A2(n_536),
.B(n_428),
.Y(n_650)
);

AOI21xp5_ASAP7_75t_L g651 ( 
.A1(n_582),
.A2(n_536),
.B(n_428),
.Y(n_651)
);

A2O1A1Ixp33_ASAP7_75t_L g652 ( 
.A1(n_546),
.A2(n_390),
.B(n_536),
.C(n_446),
.Y(n_652)
);

OAI21x1_ASAP7_75t_L g653 ( 
.A1(n_576),
.A2(n_436),
.B(n_390),
.Y(n_653)
);

AOI22xp5_ASAP7_75t_L g654 ( 
.A1(n_543),
.A2(n_390),
.B1(n_436),
.B2(n_446),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_547),
.B(n_390),
.Y(n_655)
);

OAI21xp5_ASAP7_75t_L g656 ( 
.A1(n_591),
.A2(n_446),
.B(n_436),
.Y(n_656)
);

INVx2_ASAP7_75t_SL g657 ( 
.A(n_566),
.Y(n_657)
);

OAI21x1_ASAP7_75t_L g658 ( 
.A1(n_585),
.A2(n_436),
.B(n_390),
.Y(n_658)
);

AOI22xp5_ASAP7_75t_L g659 ( 
.A1(n_571),
.A2(n_446),
.B1(n_96),
.B2(n_97),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_573),
.B(n_446),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_623),
.Y(n_661)
);

OAI21xp5_ASAP7_75t_L g662 ( 
.A1(n_608),
.A2(n_591),
.B(n_600),
.Y(n_662)
);

OAI21x1_ASAP7_75t_L g663 ( 
.A1(n_611),
.A2(n_601),
.B(n_589),
.Y(n_663)
);

AOI22xp33_ASAP7_75t_L g664 ( 
.A1(n_619),
.A2(n_570),
.B1(n_601),
.B2(n_545),
.Y(n_664)
);

OAI21xp5_ASAP7_75t_L g665 ( 
.A1(n_610),
.A2(n_570),
.B(n_557),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_630),
.Y(n_666)
);

AO21x2_ASAP7_75t_L g667 ( 
.A1(n_605),
.A2(n_601),
.B(n_550),
.Y(n_667)
);

OAI22xp5_ASAP7_75t_L g668 ( 
.A1(n_620),
.A2(n_573),
.B1(n_557),
.B2(n_542),
.Y(n_668)
);

OAI22xp5_ASAP7_75t_L g669 ( 
.A1(n_612),
.A2(n_542),
.B1(n_545),
.B2(n_567),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_640),
.B(n_545),
.Y(n_670)
);

CKINVDCx6p67_ASAP7_75t_R g671 ( 
.A(n_633),
.Y(n_671)
);

A2O1A1Ixp33_ASAP7_75t_L g672 ( 
.A1(n_647),
.A2(n_577),
.B(n_548),
.C(n_555),
.Y(n_672)
);

OA21x2_ASAP7_75t_L g673 ( 
.A1(n_613),
.A2(n_561),
.B(n_589),
.Y(n_673)
);

NAND3xp33_ASAP7_75t_L g674 ( 
.A(n_649),
.B(n_559),
.C(n_567),
.Y(n_674)
);

AO21x2_ASAP7_75t_L g675 ( 
.A1(n_652),
.A2(n_567),
.B(n_99),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_627),
.Y(n_676)
);

OAI21x1_ASAP7_75t_L g677 ( 
.A1(n_629),
.A2(n_95),
.B(n_136),
.Y(n_677)
);

AOI22xp33_ASAP7_75t_SL g678 ( 
.A1(n_646),
.A2(n_554),
.B1(n_556),
.B2(n_4),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_648),
.Y(n_679)
);

NOR2x1_ASAP7_75t_SL g680 ( 
.A(n_624),
.B(n_54),
.Y(n_680)
);

OAI22xp5_ASAP7_75t_L g681 ( 
.A1(n_638),
.A2(n_636),
.B1(n_654),
.B2(n_621),
.Y(n_681)
);

OAI21x1_ASAP7_75t_L g682 ( 
.A1(n_635),
.A2(n_100),
.B(n_191),
.Y(n_682)
);

BUFx3_ASAP7_75t_L g683 ( 
.A(n_606),
.Y(n_683)
);

OAI21x1_ASAP7_75t_L g684 ( 
.A1(n_637),
.A2(n_94),
.B(n_187),
.Y(n_684)
);

BUFx2_ASAP7_75t_L g685 ( 
.A(n_657),
.Y(n_685)
);

BUFx6f_ASAP7_75t_L g686 ( 
.A(n_606),
.Y(n_686)
);

NAND2x1p5_ASAP7_75t_L g687 ( 
.A(n_621),
.B(n_658),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_626),
.Y(n_688)
);

OA21x2_ASAP7_75t_L g689 ( 
.A1(n_625),
.A2(n_2),
.B(n_3),
.Y(n_689)
);

OAI21x1_ASAP7_75t_SL g690 ( 
.A1(n_644),
.A2(n_92),
.B(n_186),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_655),
.Y(n_691)
);

BUFx3_ASAP7_75t_L g692 ( 
.A(n_606),
.Y(n_692)
);

BUFx6f_ASAP7_75t_SL g693 ( 
.A(n_639),
.Y(n_693)
);

A2O1A1Ixp33_ASAP7_75t_L g694 ( 
.A1(n_636),
.A2(n_554),
.B(n_3),
.C(n_5),
.Y(n_694)
);

OAI21x1_ASAP7_75t_L g695 ( 
.A1(n_642),
.A2(n_90),
.B(n_183),
.Y(n_695)
);

NOR2xp67_ASAP7_75t_SL g696 ( 
.A(n_621),
.B(n_55),
.Y(n_696)
);

OAI21x1_ASAP7_75t_L g697 ( 
.A1(n_653),
.A2(n_615),
.B(n_631),
.Y(n_697)
);

AOI221xp5_ASAP7_75t_L g698 ( 
.A1(n_632),
.A2(n_2),
.B1(n_7),
.B2(n_8),
.C(n_9),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_618),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_626),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_641),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_628),
.Y(n_702)
);

HB1xp67_ASAP7_75t_L g703 ( 
.A(n_609),
.Y(n_703)
);

OAI21xp33_ASAP7_75t_SL g704 ( 
.A1(n_654),
.A2(n_8),
.B(n_10),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_628),
.Y(n_705)
);

OAI21x1_ASAP7_75t_L g706 ( 
.A1(n_617),
.A2(n_634),
.B(n_645),
.Y(n_706)
);

CKINVDCx8_ASAP7_75t_R g707 ( 
.A(n_622),
.Y(n_707)
);

NAND2x1p5_ASAP7_75t_L g708 ( 
.A(n_643),
.B(n_60),
.Y(n_708)
);

AO21x2_ASAP7_75t_L g709 ( 
.A1(n_656),
.A2(n_104),
.B(n_182),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_641),
.Y(n_710)
);

AND2x4_ASAP7_75t_L g711 ( 
.A(n_683),
.B(n_692),
.Y(n_711)
);

AOI22xp33_ASAP7_75t_L g712 ( 
.A1(n_698),
.A2(n_659),
.B1(n_643),
.B2(n_639),
.Y(n_712)
);

OAI22xp5_ASAP7_75t_L g713 ( 
.A1(n_672),
.A2(n_659),
.B1(n_639),
.B2(n_660),
.Y(n_713)
);

AOI22xp5_ASAP7_75t_L g714 ( 
.A1(n_674),
.A2(n_616),
.B1(n_650),
.B2(n_651),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_661),
.Y(n_715)
);

BUFx12f_ASAP7_75t_L g716 ( 
.A(n_685),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_688),
.Y(n_717)
);

AND2x4_ASAP7_75t_L g718 ( 
.A(n_683),
.B(n_628),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_661),
.Y(n_719)
);

OAI21x1_ASAP7_75t_L g720 ( 
.A1(n_697),
.A2(n_614),
.B(n_607),
.Y(n_720)
);

AOI22xp33_ASAP7_75t_SL g721 ( 
.A1(n_689),
.A2(n_607),
.B1(n_12),
.B2(n_13),
.Y(n_721)
);

AND2x4_ASAP7_75t_L g722 ( 
.A(n_692),
.B(n_614),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_688),
.Y(n_723)
);

AOI21xp5_ASAP7_75t_L g724 ( 
.A1(n_706),
.A2(n_607),
.B(n_614),
.Y(n_724)
);

AOI22xp33_ASAP7_75t_SL g725 ( 
.A1(n_689),
.A2(n_11),
.B1(n_14),
.B2(n_15),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_666),
.B(n_11),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_676),
.B(n_15),
.Y(n_727)
);

OAI22xp33_ASAP7_75t_L g728 ( 
.A1(n_689),
.A2(n_16),
.B1(n_18),
.B2(n_19),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_701),
.Y(n_729)
);

AND2x2_ASAP7_75t_L g730 ( 
.A(n_670),
.B(n_16),
.Y(n_730)
);

NOR2x1_ASAP7_75t_SL g731 ( 
.A(n_675),
.B(n_62),
.Y(n_731)
);

A2O1A1Ixp33_ASAP7_75t_L g732 ( 
.A1(n_662),
.A2(n_18),
.B(n_19),
.C(n_20),
.Y(n_732)
);

NAND2xp33_ASAP7_75t_R g733 ( 
.A(n_673),
.B(n_63),
.Y(n_733)
);

INVx3_ASAP7_75t_L g734 ( 
.A(n_686),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_691),
.B(n_21),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_665),
.B(n_23),
.Y(n_736)
);

BUFx2_ASAP7_75t_L g737 ( 
.A(n_685),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_707),
.Y(n_738)
);

BUFx3_ASAP7_75t_L g739 ( 
.A(n_671),
.Y(n_739)
);

OAI22xp33_ASAP7_75t_L g740 ( 
.A1(n_681),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_740)
);

AOI22xp33_ASAP7_75t_L g741 ( 
.A1(n_678),
.A2(n_24),
.B1(n_26),
.B2(n_27),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_699),
.B(n_26),
.Y(n_742)
);

AOI22xp33_ASAP7_75t_L g743 ( 
.A1(n_696),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_702),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_664),
.B(n_29),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_705),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_694),
.B(n_30),
.Y(n_747)
);

NAND2x1p5_ASAP7_75t_L g748 ( 
.A(n_696),
.B(n_64),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_700),
.Y(n_749)
);

AND2x4_ASAP7_75t_L g750 ( 
.A(n_686),
.B(n_65),
.Y(n_750)
);

AND2x2_ASAP7_75t_L g751 ( 
.A(n_686),
.B(n_31),
.Y(n_751)
);

AOI22xp33_ASAP7_75t_L g752 ( 
.A1(n_704),
.A2(n_709),
.B1(n_669),
.B2(n_675),
.Y(n_752)
);

INVx4_ASAP7_75t_L g753 ( 
.A(n_693),
.Y(n_753)
);

OAI22xp33_ASAP7_75t_SL g754 ( 
.A1(n_708),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_754)
);

NAND2xp33_ASAP7_75t_SL g755 ( 
.A(n_693),
.B(n_32),
.Y(n_755)
);

CKINVDCx6p67_ASAP7_75t_R g756 ( 
.A(n_693),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_701),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_710),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_700),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_679),
.Y(n_760)
);

AOI22xp33_ASAP7_75t_L g761 ( 
.A1(n_709),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_761)
);

OAI22xp5_ASAP7_75t_L g762 ( 
.A1(n_668),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.Y(n_762)
);

CKINVDCx20_ASAP7_75t_R g763 ( 
.A(n_707),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_679),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_663),
.Y(n_765)
);

AND2x4_ASAP7_75t_L g766 ( 
.A(n_686),
.B(n_66),
.Y(n_766)
);

CKINVDCx20_ASAP7_75t_R g767 ( 
.A(n_671),
.Y(n_767)
);

OAI22xp5_ASAP7_75t_L g768 ( 
.A1(n_708),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.Y(n_768)
);

OAI21x1_ASAP7_75t_L g769 ( 
.A1(n_697),
.A2(n_695),
.B(n_706),
.Y(n_769)
);

OR2x2_ASAP7_75t_L g770 ( 
.A(n_686),
.B(n_70),
.Y(n_770)
);

AOI22xp5_ASAP7_75t_L g771 ( 
.A1(n_675),
.A2(n_71),
.B1(n_72),
.B2(n_75),
.Y(n_771)
);

OAI22xp33_ASAP7_75t_L g772 ( 
.A1(n_747),
.A2(n_708),
.B1(n_703),
.B2(n_687),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_716),
.B(n_680),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_730),
.B(n_680),
.Y(n_774)
);

OR2x6_ASAP7_75t_L g775 ( 
.A(n_748),
.B(n_663),
.Y(n_775)
);

OAI22xp5_ASAP7_75t_L g776 ( 
.A1(n_741),
.A2(n_687),
.B1(n_673),
.B2(n_710),
.Y(n_776)
);

OAI211xp5_ASAP7_75t_L g777 ( 
.A1(n_741),
.A2(n_673),
.B(n_695),
.C(n_684),
.Y(n_777)
);

OAI22xp33_ASAP7_75t_L g778 ( 
.A1(n_740),
.A2(n_771),
.B1(n_733),
.B2(n_736),
.Y(n_778)
);

OAI22xp5_ASAP7_75t_L g779 ( 
.A1(n_712),
.A2(n_687),
.B1(n_690),
.B2(n_709),
.Y(n_779)
);

OAI21x1_ASAP7_75t_L g780 ( 
.A1(n_769),
.A2(n_684),
.B(n_682),
.Y(n_780)
);

AOI22xp33_ASAP7_75t_SL g781 ( 
.A1(n_768),
.A2(n_690),
.B1(n_667),
.B2(n_677),
.Y(n_781)
);

AOI221xp5_ASAP7_75t_SL g782 ( 
.A1(n_740),
.A2(n_667),
.B1(n_682),
.B2(n_677),
.C(n_79),
.Y(n_782)
);

OAI22xp5_ASAP7_75t_L g783 ( 
.A1(n_712),
.A2(n_667),
.B1(n_77),
.B2(n_78),
.Y(n_783)
);

AOI22xp33_ASAP7_75t_L g784 ( 
.A1(n_743),
.A2(n_76),
.B1(n_81),
.B2(n_82),
.Y(n_784)
);

OAI221xp5_ASAP7_75t_L g785 ( 
.A1(n_732),
.A2(n_83),
.B1(n_84),
.B2(n_85),
.C(n_88),
.Y(n_785)
);

AOI222xp33_ASAP7_75t_L g786 ( 
.A1(n_743),
.A2(n_89),
.B1(n_101),
.B2(n_102),
.C1(n_103),
.C2(n_105),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_715),
.Y(n_787)
);

AND2x4_ASAP7_75t_L g788 ( 
.A(n_753),
.B(n_106),
.Y(n_788)
);

OAI221xp5_ASAP7_75t_L g789 ( 
.A1(n_732),
.A2(n_108),
.B1(n_109),
.B2(n_110),
.C(n_113),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_738),
.B(n_118),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_719),
.Y(n_791)
);

AOI22xp33_ASAP7_75t_L g792 ( 
.A1(n_761),
.A2(n_755),
.B1(n_762),
.B2(n_745),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_749),
.Y(n_793)
);

AOI22xp5_ASAP7_75t_L g794 ( 
.A1(n_755),
.A2(n_119),
.B1(n_120),
.B2(n_121),
.Y(n_794)
);

OAI221xp5_ASAP7_75t_SL g795 ( 
.A1(n_761),
.A2(n_122),
.B1(n_124),
.B2(n_127),
.C(n_128),
.Y(n_795)
);

INVx3_ASAP7_75t_L g796 ( 
.A(n_734),
.Y(n_796)
);

AOI22xp33_ASAP7_75t_L g797 ( 
.A1(n_725),
.A2(n_130),
.B1(n_131),
.B2(n_132),
.Y(n_797)
);

INVx3_ASAP7_75t_L g798 ( 
.A(n_734),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_759),
.Y(n_799)
);

BUFx6f_ASAP7_75t_L g800 ( 
.A(n_739),
.Y(n_800)
);

OAI22xp33_ASAP7_75t_L g801 ( 
.A1(n_733),
.A2(n_134),
.B1(n_135),
.B2(n_140),
.Y(n_801)
);

AOI22xp33_ASAP7_75t_SL g802 ( 
.A1(n_754),
.A2(n_141),
.B1(n_142),
.B2(n_143),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_763),
.B(n_146),
.Y(n_803)
);

AOI22xp5_ASAP7_75t_L g804 ( 
.A1(n_713),
.A2(n_147),
.B1(n_148),
.B2(n_149),
.Y(n_804)
);

NAND3xp33_ASAP7_75t_L g805 ( 
.A(n_725),
.B(n_151),
.C(n_152),
.Y(n_805)
);

AOI22xp33_ASAP7_75t_L g806 ( 
.A1(n_728),
.A2(n_153),
.B1(n_154),
.B2(n_156),
.Y(n_806)
);

OAI221xp5_ASAP7_75t_L g807 ( 
.A1(n_752),
.A2(n_160),
.B1(n_162),
.B2(n_163),
.C(n_167),
.Y(n_807)
);

OAI22xp5_ASAP7_75t_L g808 ( 
.A1(n_756),
.A2(n_169),
.B1(n_170),
.B2(n_171),
.Y(n_808)
);

NAND3xp33_ASAP7_75t_L g809 ( 
.A(n_752),
.B(n_172),
.C(n_173),
.Y(n_809)
);

INVx3_ASAP7_75t_L g810 ( 
.A(n_711),
.Y(n_810)
);

AOI22xp33_ASAP7_75t_SL g811 ( 
.A1(n_748),
.A2(n_174),
.B1(n_175),
.B2(n_176),
.Y(n_811)
);

OAI22xp33_ASAP7_75t_L g812 ( 
.A1(n_727),
.A2(n_179),
.B1(n_181),
.B2(n_184),
.Y(n_812)
);

OAI211xp5_ASAP7_75t_L g813 ( 
.A1(n_721),
.A2(n_735),
.B(n_726),
.C(n_742),
.Y(n_813)
);

CKINVDCx6p67_ASAP7_75t_R g814 ( 
.A(n_767),
.Y(n_814)
);

OAI22xp33_ASAP7_75t_L g815 ( 
.A1(n_728),
.A2(n_753),
.B1(n_739),
.B2(n_737),
.Y(n_815)
);

AOI21x1_ASAP7_75t_L g816 ( 
.A1(n_724),
.A2(n_765),
.B(n_722),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_711),
.Y(n_817)
);

AOI22xp33_ASAP7_75t_L g818 ( 
.A1(n_722),
.A2(n_721),
.B1(n_718),
.B2(n_751),
.Y(n_818)
);

OAI22xp5_ASAP7_75t_L g819 ( 
.A1(n_714),
.A2(n_718),
.B1(n_770),
.B2(n_766),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_744),
.Y(n_820)
);

OAI22xp5_ASAP7_75t_L g821 ( 
.A1(n_750),
.A2(n_766),
.B1(n_746),
.B2(n_764),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_760),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_750),
.B(n_717),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_L g824 ( 
.A(n_803),
.B(n_790),
.Y(n_824)
);

OA21x2_ASAP7_75t_L g825 ( 
.A1(n_782),
.A2(n_720),
.B(n_729),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_822),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_799),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_820),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_793),
.B(n_717),
.Y(n_829)
);

INVx1_ASAP7_75t_SL g830 ( 
.A(n_823),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_787),
.Y(n_831)
);

INVxp67_ASAP7_75t_L g832 ( 
.A(n_791),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_816),
.B(n_723),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_772),
.B(n_723),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_774),
.B(n_729),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_775),
.Y(n_836)
);

INVx2_ASAP7_75t_SL g837 ( 
.A(n_800),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_775),
.Y(n_838)
);

AND2x2_ASAP7_75t_L g839 ( 
.A(n_818),
.B(n_757),
.Y(n_839)
);

INVxp67_ASAP7_75t_L g840 ( 
.A(n_817),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_776),
.B(n_757),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_775),
.Y(n_842)
);

HB1xp67_ASAP7_75t_L g843 ( 
.A(n_819),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_780),
.Y(n_844)
);

OR2x2_ASAP7_75t_L g845 ( 
.A(n_779),
.B(n_758),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_796),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_796),
.B(n_758),
.Y(n_847)
);

INVxp67_ASAP7_75t_SL g848 ( 
.A(n_798),
.Y(n_848)
);

INVx2_ASAP7_75t_SL g849 ( 
.A(n_800),
.Y(n_849)
);

AND2x2_ASAP7_75t_L g850 ( 
.A(n_798),
.B(n_731),
.Y(n_850)
);

BUFx3_ASAP7_75t_L g851 ( 
.A(n_800),
.Y(n_851)
);

INVxp67_ASAP7_75t_SL g852 ( 
.A(n_810),
.Y(n_852)
);

AOI222xp33_ASAP7_75t_L g853 ( 
.A1(n_778),
.A2(n_792),
.B1(n_805),
.B2(n_789),
.C1(n_785),
.C2(n_784),
.Y(n_853)
);

NOR2x1p5_ASAP7_75t_L g854 ( 
.A(n_809),
.B(n_810),
.Y(n_854)
);

OA21x2_ASAP7_75t_L g855 ( 
.A1(n_777),
.A2(n_809),
.B(n_807),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_821),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_781),
.Y(n_857)
);

AOI21xp33_ASAP7_75t_L g858 ( 
.A1(n_815),
.A2(n_813),
.B(n_786),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_773),
.B(n_806),
.Y(n_859)
);

BUFx5_ASAP7_75t_L g860 ( 
.A(n_788),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_783),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_797),
.B(n_802),
.Y(n_862)
);

NAND2x1_ASAP7_75t_L g863 ( 
.A(n_788),
.B(n_804),
.Y(n_863)
);

INVx2_ASAP7_75t_SL g864 ( 
.A(n_851),
.Y(n_864)
);

OAI211xp5_ASAP7_75t_L g865 ( 
.A1(n_858),
.A2(n_795),
.B(n_794),
.C(n_811),
.Y(n_865)
);

AO21x2_ASAP7_75t_L g866 ( 
.A1(n_844),
.A2(n_801),
.B(n_812),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_827),
.Y(n_867)
);

AOI221xp5_ASAP7_75t_L g868 ( 
.A1(n_858),
.A2(n_808),
.B1(n_814),
.B2(n_857),
.C(n_843),
.Y(n_868)
);

NOR3xp33_ASAP7_75t_SL g869 ( 
.A(n_857),
.B(n_824),
.C(n_842),
.Y(n_869)
);

OAI221xp5_ASAP7_75t_L g870 ( 
.A1(n_853),
.A2(n_863),
.B1(n_862),
.B2(n_855),
.C(n_859),
.Y(n_870)
);

AOI22xp33_ASAP7_75t_L g871 ( 
.A1(n_853),
.A2(n_862),
.B1(n_854),
.B2(n_859),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_827),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_826),
.Y(n_873)
);

BUFx3_ASAP7_75t_L g874 ( 
.A(n_851),
.Y(n_874)
);

OAI211xp5_ASAP7_75t_L g875 ( 
.A1(n_855),
.A2(n_861),
.B(n_856),
.C(n_863),
.Y(n_875)
);

NAND3xp33_ASAP7_75t_L g876 ( 
.A(n_855),
.B(n_861),
.C(n_834),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_835),
.B(n_836),
.Y(n_877)
);

HB1xp67_ASAP7_75t_L g878 ( 
.A(n_830),
.Y(n_878)
);

NOR2xp33_ASAP7_75t_L g879 ( 
.A(n_840),
.B(n_851),
.Y(n_879)
);

AOI22xp33_ASAP7_75t_L g880 ( 
.A1(n_854),
.A2(n_855),
.B1(n_856),
.B2(n_839),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_L g881 ( 
.A(n_830),
.B(n_837),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_826),
.Y(n_882)
);

NOR4xp25_ASAP7_75t_SL g883 ( 
.A(n_836),
.B(n_838),
.C(n_842),
.D(n_848),
.Y(n_883)
);

AOI222xp33_ASAP7_75t_L g884 ( 
.A1(n_839),
.A2(n_834),
.B1(n_832),
.B2(n_841),
.C1(n_828),
.C2(n_831),
.Y(n_884)
);

OAI33xp33_ASAP7_75t_L g885 ( 
.A1(n_832),
.A2(n_828),
.A3(n_831),
.B1(n_838),
.B2(n_845),
.B3(n_827),
.Y(n_885)
);

OAI22xp33_ASAP7_75t_L g886 ( 
.A1(n_845),
.A2(n_837),
.B1(n_849),
.B2(n_852),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_829),
.Y(n_887)
);

NOR2x1_ASAP7_75t_L g888 ( 
.A(n_876),
.B(n_846),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_873),
.Y(n_889)
);

AND2x4_ASAP7_75t_SL g890 ( 
.A(n_878),
.B(n_850),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_867),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_877),
.B(n_835),
.Y(n_892)
);

AND2x2_ASAP7_75t_L g893 ( 
.A(n_877),
.B(n_841),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_873),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_884),
.B(n_846),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_887),
.B(n_833),
.Y(n_896)
);

BUFx3_ASAP7_75t_L g897 ( 
.A(n_874),
.Y(n_897)
);

NAND2x1_ASAP7_75t_L g898 ( 
.A(n_867),
.B(n_872),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_882),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_882),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_872),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_887),
.Y(n_902)
);

AND2x2_ASAP7_75t_L g903 ( 
.A(n_884),
.B(n_833),
.Y(n_903)
);

INVx4_ASAP7_75t_L g904 ( 
.A(n_874),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_903),
.B(n_876),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_889),
.Y(n_906)
);

AND2x2_ASAP7_75t_L g907 ( 
.A(n_903),
.B(n_883),
.Y(n_907)
);

INVx3_ASAP7_75t_L g908 ( 
.A(n_898),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_889),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_895),
.B(n_880),
.Y(n_910)
);

NOR2x1p5_ASAP7_75t_L g911 ( 
.A(n_897),
.B(n_874),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_890),
.B(n_883),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_896),
.B(n_875),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_890),
.B(n_864),
.Y(n_914)
);

AND2x2_ASAP7_75t_L g915 ( 
.A(n_893),
.B(n_864),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_894),
.Y(n_916)
);

AND2x2_ASAP7_75t_L g917 ( 
.A(n_893),
.B(n_896),
.Y(n_917)
);

OR2x2_ASAP7_75t_L g918 ( 
.A(n_905),
.B(n_892),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_917),
.B(n_892),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_906),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_R g921 ( 
.A(n_907),
.B(n_871),
.Y(n_921)
);

HB1xp67_ASAP7_75t_L g922 ( 
.A(n_906),
.Y(n_922)
);

OR2x2_ASAP7_75t_L g923 ( 
.A(n_913),
.B(n_902),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_916),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_916),
.Y(n_925)
);

AOI31xp67_ASAP7_75t_SL g926 ( 
.A1(n_910),
.A2(n_870),
.A3(n_869),
.B(n_888),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_917),
.B(n_897),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_911),
.B(n_904),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_927),
.B(n_915),
.Y(n_929)
);

AOI322xp5_ASAP7_75t_L g930 ( 
.A1(n_926),
.A2(n_907),
.A3(n_868),
.B1(n_912),
.B2(n_915),
.C1(n_886),
.C2(n_914),
.Y(n_930)
);

INVxp33_ASAP7_75t_L g931 ( 
.A(n_921),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_922),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_921),
.B(n_912),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_922),
.Y(n_934)
);

OAI22xp5_ASAP7_75t_L g935 ( 
.A1(n_933),
.A2(n_926),
.B1(n_918),
.B2(n_928),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_932),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_931),
.B(n_928),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_930),
.B(n_919),
.Y(n_938)
);

OAI21xp33_ASAP7_75t_L g939 ( 
.A1(n_938),
.A2(n_931),
.B(n_934),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_936),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_937),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_SL g942 ( 
.A(n_935),
.B(n_929),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_937),
.Y(n_943)
);

NOR3xp33_ASAP7_75t_L g944 ( 
.A(n_939),
.B(n_865),
.C(n_923),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_941),
.B(n_943),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_940),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_943),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_942),
.B(n_925),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_SL g949 ( 
.A(n_943),
.B(n_908),
.Y(n_949)
);

INVxp67_ASAP7_75t_SL g950 ( 
.A(n_941),
.Y(n_950)
);

NAND3xp33_ASAP7_75t_SL g951 ( 
.A(n_944),
.B(n_904),
.C(n_920),
.Y(n_951)
);

AOI221xp5_ASAP7_75t_L g952 ( 
.A1(n_950),
.A2(n_948),
.B1(n_947),
.B2(n_945),
.C(n_946),
.Y(n_952)
);

NOR2xp33_ASAP7_75t_L g953 ( 
.A(n_950),
.B(n_924),
.Y(n_953)
);

AOI221xp5_ASAP7_75t_L g954 ( 
.A1(n_949),
.A2(n_885),
.B1(n_879),
.B2(n_909),
.C(n_904),
.Y(n_954)
);

NAND2xp33_ASAP7_75t_R g955 ( 
.A(n_945),
.B(n_908),
.Y(n_955)
);

OAI21xp5_ASAP7_75t_L g956 ( 
.A1(n_944),
.A2(n_908),
.B(n_914),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_953),
.Y(n_957)
);

INVxp67_ASAP7_75t_L g958 ( 
.A(n_955),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_952),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_951),
.Y(n_960)
);

NOR2xp67_ASAP7_75t_L g961 ( 
.A(n_956),
.B(n_849),
.Y(n_961)
);

AOI22xp5_ASAP7_75t_SL g962 ( 
.A1(n_954),
.A2(n_881),
.B1(n_902),
.B2(n_899),
.Y(n_962)
);

OR2x2_ASAP7_75t_L g963 ( 
.A(n_957),
.B(n_901),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_959),
.A2(n_958),
.B(n_961),
.Y(n_964)
);

AO22x2_ASAP7_75t_L g965 ( 
.A1(n_960),
.A2(n_900),
.B1(n_894),
.B2(n_898),
.Y(n_965)
);

NOR3x2_ASAP7_75t_L g966 ( 
.A(n_962),
.B(n_860),
.C(n_866),
.Y(n_966)
);

AND2x4_ASAP7_75t_L g967 ( 
.A(n_958),
.B(n_891),
.Y(n_967)
);

INVxp67_ASAP7_75t_L g968 ( 
.A(n_964),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_963),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_967),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_965),
.B(n_900),
.Y(n_971)
);

HB1xp67_ASAP7_75t_L g972 ( 
.A(n_970),
.Y(n_972)
);

HB1xp67_ASAP7_75t_L g973 ( 
.A(n_969),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_972),
.Y(n_974)
);

OAI22xp5_ASAP7_75t_L g975 ( 
.A1(n_973),
.A2(n_968),
.B1(n_971),
.B2(n_966),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_975),
.A2(n_974),
.B(n_866),
.Y(n_976)
);

OAI22xp5_ASAP7_75t_SL g977 ( 
.A1(n_974),
.A2(n_891),
.B1(n_846),
.B2(n_860),
.Y(n_977)
);

OR2x2_ASAP7_75t_L g978 ( 
.A(n_976),
.B(n_866),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_977),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_979),
.A2(n_844),
.B(n_850),
.Y(n_980)
);

OAI21xp5_ASAP7_75t_L g981 ( 
.A1(n_978),
.A2(n_844),
.B(n_847),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_981),
.Y(n_982)
);

HB1xp67_ASAP7_75t_L g983 ( 
.A(n_982),
.Y(n_983)
);

OAI221xp5_ASAP7_75t_L g984 ( 
.A1(n_983),
.A2(n_980),
.B1(n_825),
.B2(n_829),
.C(n_847),
.Y(n_984)
);

AOI211xp5_ASAP7_75t_L g985 ( 
.A1(n_984),
.A2(n_825),
.B(n_860),
.C(n_968),
.Y(n_985)
);


endmodule