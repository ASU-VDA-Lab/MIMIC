module fake_jpeg_16563_n_58 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_58);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_58;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_27;
wire n_55;
wire n_47;
wire n_51;
wire n_40;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_44;
wire n_38;
wire n_26;
wire n_28;
wire n_36;
wire n_25;
wire n_31;
wire n_56;
wire n_37;
wire n_29;
wire n_43;
wire n_50;
wire n_32;

INVx1_ASAP7_75t_L g24 ( 
.A(n_23),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_7),
.B(n_18),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_24),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_34),
.Y(n_41)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_25),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_35),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_26),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_37),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_38),
.B(n_27),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_40),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_5),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_44),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_28),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_41),
.B(n_31),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_46),
.B(n_47),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_42),
.B(n_6),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_45),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_49),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_51),
.B(n_50),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_53),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_54),
.A2(n_52),
.B1(n_48),
.B2(n_10),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_55),
.B(n_8),
.Y(n_56)
);

AOI322xp5_ASAP7_75t_L g57 ( 
.A1(n_56),
.A2(n_9),
.A3(n_11),
.B1(n_12),
.B2(n_13),
.C1(n_14),
.C2(n_15),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_22),
.Y(n_58)
);


endmodule