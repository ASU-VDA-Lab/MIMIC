module fake_ariane_2064_n_1244 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_169, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1244);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1244;

wire n_913;
wire n_589;
wire n_1174;
wire n_691;
wire n_423;
wire n_603;
wire n_373;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_319;
wire n_690;
wire n_416;
wire n_1109;
wire n_525;
wire n_187;
wire n_1238;
wire n_817;
wire n_924;
wire n_781;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_524;
wire n_1214;
wire n_634;
wire n_1138;
wire n_214;
wire n_764;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_232;
wire n_568;
wire n_1088;
wire n_766;
wire n_377;
wire n_520;
wire n_870;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_672;
wire n_740;
wire n_1018;
wire n_259;
wire n_953;
wire n_1224;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_200;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1195;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_868;
wire n_884;
wire n_1034;
wire n_1085;
wire n_277;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_611;
wire n_238;
wire n_365;
wire n_1013;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_440;
wire n_273;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_579;
wire n_844;
wire n_1012;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_491;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_461;
wire n_1121;
wire n_490;
wire n_209;
wire n_225;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_676;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_851;
wire n_444;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_912;
wire n_460;
wire n_366;
wire n_762;
wire n_555;
wire n_804;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_514;
wire n_418;
wire n_513;
wire n_288;
wire n_179;
wire n_1178;
wire n_1026;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_746;
wire n_292;
wire n_1079;
wire n_615;
wire n_1139;
wire n_517;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1101;
wire n_563;
wire n_990;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_767;
wire n_964;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1220;
wire n_356;
wire n_698;
wire n_307;
wire n_1209;
wire n_1020;
wire n_646;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_299;
wire n_836;
wire n_564;
wire n_205;
wire n_1029;
wire n_760;
wire n_522;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_776;
wire n_424;
wire n_466;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_637;
wire n_327;
wire n_1177;
wire n_1231;
wire n_980;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_487;
wire n_855;
wire n_808;
wire n_553;
wire n_814;
wire n_578;
wire n_405;
wire n_320;
wire n_1134;
wire n_647;
wire n_481;
wire n_600;
wire n_1053;
wire n_529;
wire n_502;
wire n_218;
wire n_247;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_545;
wire n_1015;
wire n_1162;
wire n_536;
wire n_325;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_442;
wire n_777;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_887;
wire n_729;
wire n_1122;
wire n_1205;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_233;
wire n_957;
wire n_388;
wire n_1242;
wire n_1218;
wire n_321;
wire n_221;
wire n_861;
wire n_877;
wire n_1119;
wire n_616;
wire n_1055;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_888;
wire n_845;
wire n_178;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_742;
wire n_1081;
wire n_769;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1171;
wire n_1030;
wire n_785;
wire n_999;
wire n_456;
wire n_852;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1243;
wire n_342;
wire n_358;
wire n_608;
wire n_1037;
wire n_317;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_687;
wire n_797;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_595;
wire n_602;
wire n_592;
wire n_854;
wire n_393;
wire n_474;
wire n_805;
wire n_295;
wire n_190;
wire n_1072;
wire n_695;
wire n_180;
wire n_730;
wire n_386;
wire n_516;
wire n_1137;
wire n_197;
wire n_640;
wire n_463;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_878;
wire n_771;
wire n_752;
wire n_985;
wire n_421;
wire n_906;
wire n_1180;
wire n_283;
wire n_806;
wire n_649;
wire n_374;
wire n_643;
wire n_226;
wire n_682;
wire n_819;
wire n_586;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1130;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_979;
wire n_897;
wire n_949;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_818;
wire n_779;
wire n_594;
wire n_1052;
wire n_272;
wire n_833;
wire n_879;
wire n_1117;
wire n_422;
wire n_597;
wire n_1047;
wire n_1050;
wire n_566;
wire n_1201;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1192;
wire n_224;
wire n_894;
wire n_420;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_538;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1128;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1065;
wire n_453;
wire n_810;
wire n_181;
wire n_617;
wire n_543;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_743;
wire n_1194;
wire n_907;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_284;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_613;
wire n_1022;
wire n_1033;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_820;
wire n_872;
wire n_254;
wire n_1157;
wire n_234;
wire n_848;
wire n_280;
wire n_629;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_223;
wire n_750;
wire n_834;
wire n_800;
wire n_395;
wire n_621;
wire n_213;
wire n_1014;
wire n_724;
wire n_493;
wire n_1100;
wire n_585;
wire n_875;
wire n_827;
wire n_697;
wire n_622;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_739;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_580;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1124;
wire n_932;
wire n_1183;
wire n_981;
wire n_1110;
wire n_243;
wire n_185;
wire n_1204;
wire n_994;
wire n_973;
wire n_268;
wire n_972;
wire n_184;
wire n_856;
wire n_1176;
wire n_1054;
wire n_508;
wire n_353;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_828;
wire n_322;
wire n_558;
wire n_653;
wire n_783;
wire n_556;
wire n_1127;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1167;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_318;
wire n_244;
wire n_679;
wire n_220;
wire n_663;
wire n_443;
wire n_528;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_385;
wire n_917;
wire n_372;
wire n_631;
wire n_399;
wire n_1170;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1064;
wire n_633;
wire n_900;
wire n_1093;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_835;
wire n_446;
wire n_1076;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_309;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_291;
wire n_822;
wire n_1094;
wire n_840;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_188;
wire n_323;
wire n_550;
wire n_997;
wire n_635;
wire n_694;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1236;
wire n_228;
wire n_671;
wire n_1148;
wire n_654;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1144;
wire n_383;
wire n_838;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_658;
wire n_630;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_235;
wire n_881;
wire n_1019;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_902;
wire n_1031;
wire n_853;
wire n_716;
wire n_196;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1229;
wire n_415;
wire n_544;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1126;
wire n_195;
wire n_938;
wire n_895;
wire n_304;
wire n_583;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_946;
wire n_757;
wire n_375;
wire n_1146;
wire n_1203;
wire n_998;
wire n_472;
wire n_937;
wire n_265;
wire n_208;
wire n_174;
wire n_275;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_963;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1001;
wire n_1115;
wire n_1002;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_250;
wire n_773;
wire n_1010;
wire n_882;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_289;
wire n_548;
wire n_523;
wire n_457;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_447;
wire n_1233;
wire n_893;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_573;
wire n_796;
wire n_531;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_160),
.Y(n_172)
);

BUFx2_ASAP7_75t_SL g173 ( 
.A(n_105),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_23),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_23),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_7),
.Y(n_176)
);

BUFx5_ASAP7_75t_L g177 ( 
.A(n_94),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_149),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_167),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_158),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_98),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_40),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_143),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_163),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_161),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_110),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_113),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_138),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_169),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_44),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_60),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_20),
.Y(n_192)
);

INVx2_ASAP7_75t_SL g193 ( 
.A(n_170),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_76),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_122),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_47),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_164),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_168),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_32),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_171),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_117),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_32),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_140),
.Y(n_203)
);

INVx2_ASAP7_75t_SL g204 ( 
.A(n_97),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_107),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_111),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_46),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_130),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_99),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_96),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_24),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_103),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_100),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_89),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_135),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_12),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_119),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_120),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_157),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_137),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_166),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_132),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_114),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_112),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_80),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_30),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_155),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_109),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_68),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_174),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_192),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_202),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_213),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_179),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_179),
.Y(n_235)
);

BUFx10_ASAP7_75t_L g236 ( 
.A(n_193),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_205),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_175),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_211),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_172),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_186),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_187),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_219),
.Y(n_243)
);

BUFx10_ASAP7_75t_L g244 ( 
.A(n_193),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_189),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_190),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_176),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_182),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_219),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_216),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_195),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_213),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_196),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_197),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_199),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_226),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_199),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_184),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_198),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_243),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_238),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_257),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_238),
.Y(n_263)
);

NOR2xp67_ASAP7_75t_L g264 ( 
.A(n_240),
.B(n_204),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_247),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_241),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_247),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_248),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_248),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_252),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_242),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_245),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_252),
.Y(n_273)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_249),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_237),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_233),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_246),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_251),
.Y(n_278)
);

BUFx2_ASAP7_75t_SL g279 ( 
.A(n_236),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_234),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_255),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_230),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_237),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_234),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_237),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_231),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_235),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_235),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_253),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_254),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_259),
.Y(n_291)
);

NOR2xp67_ASAP7_75t_L g292 ( 
.A(n_232),
.B(n_204),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_239),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_236),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_233),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_233),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_250),
.Y(n_297)
);

INVxp33_ASAP7_75t_SL g298 ( 
.A(n_256),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_258),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_236),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_236),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_244),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_244),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_237),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_244),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_244),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_237),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_237),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_237),
.Y(n_309)
);

INVx1_ASAP7_75t_SL g310 ( 
.A(n_257),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_238),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_280),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_284),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_266),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_287),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_288),
.Y(n_316)
);

HB1xp67_ASAP7_75t_L g317 ( 
.A(n_310),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_282),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_270),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_273),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_275),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_261),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_263),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_286),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_265),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_267),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_268),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_269),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_311),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_295),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_296),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_260),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_266),
.Y(n_333)
);

BUFx3_ASAP7_75t_L g334 ( 
.A(n_276),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_271),
.Y(n_335)
);

INVxp33_ASAP7_75t_L g336 ( 
.A(n_262),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_271),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_272),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_281),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_275),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_276),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_299),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_283),
.Y(n_343)
);

INVxp67_ASAP7_75t_SL g344 ( 
.A(n_298),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_283),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_293),
.Y(n_346)
);

BUFx3_ASAP7_75t_L g347 ( 
.A(n_308),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_272),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_277),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_285),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_277),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_285),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_307),
.Y(n_353)
);

INVxp33_ASAP7_75t_SL g354 ( 
.A(n_293),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_274),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_278),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_307),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_304),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_304),
.Y(n_359)
);

HB1xp67_ASAP7_75t_L g360 ( 
.A(n_298),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_308),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_317),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_314),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_312),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_322),
.B(n_279),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_333),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_312),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_318),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_313),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_313),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_335),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_337),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_324),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_315),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_338),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_315),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_348),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_332),
.Y(n_378)
);

HB1xp67_ASAP7_75t_L g379 ( 
.A(n_360),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_339),
.Y(n_380)
);

INVxp67_ASAP7_75t_SL g381 ( 
.A(n_347),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_349),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_351),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_354),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_346),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_316),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_356),
.Y(n_387)
);

CKINVDCx16_ASAP7_75t_R g388 ( 
.A(n_334),
.Y(n_388)
);

INVxp67_ASAP7_75t_SL g389 ( 
.A(n_355),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_316),
.Y(n_390)
);

NOR2xp67_ASAP7_75t_L g391 ( 
.A(n_342),
.B(n_278),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_319),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_344),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_334),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_319),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_341),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_336),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_320),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_320),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_330),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_322),
.B(n_289),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_323),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_325),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_325),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_330),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_326),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_364),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_364),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_367),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_363),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_392),
.Y(n_411)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_367),
.Y(n_412)
);

AOI22x1_ASAP7_75t_SL g413 ( 
.A1(n_385),
.A2(n_290),
.B1(n_291),
.B2(n_289),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_369),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_369),
.B(n_326),
.Y(n_415)
);

INVx3_ASAP7_75t_L g416 ( 
.A(n_370),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_370),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_392),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_401),
.A2(n_291),
.B1(n_290),
.B2(n_303),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_395),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_374),
.Y(n_421)
);

AND2x4_ASAP7_75t_L g422 ( 
.A(n_394),
.B(n_327),
.Y(n_422)
);

INVx3_ASAP7_75t_L g423 ( 
.A(n_374),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_376),
.B(n_327),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_376),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_386),
.B(n_328),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_400),
.A2(n_264),
.B1(n_302),
.B2(n_306),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_386),
.Y(n_428)
);

INVxp33_ASAP7_75t_SL g429 ( 
.A(n_366),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_390),
.B(n_328),
.Y(n_430)
);

BUFx8_ASAP7_75t_L g431 ( 
.A(n_378),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_395),
.Y(n_432)
);

HB1xp67_ASAP7_75t_L g433 ( 
.A(n_379),
.Y(n_433)
);

AND2x2_ASAP7_75t_SL g434 ( 
.A(n_390),
.B(n_200),
.Y(n_434)
);

BUFx2_ASAP7_75t_L g435 ( 
.A(n_397),
.Y(n_435)
);

OAI21x1_ASAP7_75t_L g436 ( 
.A1(n_399),
.A2(n_358),
.B(n_359),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_403),
.Y(n_437)
);

INVx6_ASAP7_75t_L g438 ( 
.A(n_388),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_403),
.Y(n_439)
);

OR2x2_ASAP7_75t_L g440 ( 
.A(n_362),
.B(n_297),
.Y(n_440)
);

OA21x2_ASAP7_75t_L g441 ( 
.A1(n_404),
.A2(n_345),
.B(n_343),
.Y(n_441)
);

AND2x6_ASAP7_75t_L g442 ( 
.A(n_404),
.B(n_329),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_405),
.A2(n_301),
.B1(n_306),
.B2(n_294),
.Y(n_443)
);

AOI22x1_ASAP7_75t_SL g444 ( 
.A1(n_368),
.A2(n_294),
.B1(n_301),
.B2(n_227),
.Y(n_444)
);

HB1xp67_ASAP7_75t_L g445 ( 
.A(n_380),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_406),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_393),
.A2(n_292),
.B1(n_305),
.B2(n_361),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_399),
.B(n_329),
.Y(n_448)
);

OAI21x1_ASAP7_75t_L g449 ( 
.A1(n_365),
.A2(n_358),
.B(n_359),
.Y(n_449)
);

AND2x4_ASAP7_75t_L g450 ( 
.A(n_391),
.B(n_331),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_398),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_381),
.B(n_350),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_396),
.Y(n_453)
);

BUFx6f_ASAP7_75t_L g454 ( 
.A(n_371),
.Y(n_454)
);

BUFx6f_ASAP7_75t_L g455 ( 
.A(n_372),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_375),
.Y(n_456)
);

INVx3_ASAP7_75t_L g457 ( 
.A(n_377),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_387),
.B(n_300),
.Y(n_458)
);

OAI22x1_ASAP7_75t_R g459 ( 
.A1(n_373),
.A2(n_181),
.B1(n_227),
.B2(n_224),
.Y(n_459)
);

AND2x4_ASAP7_75t_L g460 ( 
.A(n_402),
.B(n_357),
.Y(n_460)
);

CKINVDCx6p67_ASAP7_75t_R g461 ( 
.A(n_382),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_383),
.A2(n_203),
.B1(n_181),
.B2(n_223),
.Y(n_462)
);

HB1xp67_ASAP7_75t_L g463 ( 
.A(n_384),
.Y(n_463)
);

BUFx2_ASAP7_75t_L g464 ( 
.A(n_389),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_392),
.Y(n_465)
);

BUFx8_ASAP7_75t_L g466 ( 
.A(n_378),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_L g467 ( 
.A1(n_364),
.A2(n_183),
.B1(n_228),
.B2(n_188),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_364),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_L g469 ( 
.A1(n_364),
.A2(n_214),
.B1(n_191),
.B2(n_194),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_364),
.B(n_352),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_392),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_364),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_364),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_392),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_364),
.B(n_352),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_364),
.Y(n_476)
);

BUFx12f_ASAP7_75t_L g477 ( 
.A(n_363),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_363),
.Y(n_478)
);

INVx3_ASAP7_75t_L g479 ( 
.A(n_364),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_362),
.B(n_353),
.Y(n_480)
);

AND2x4_ASAP7_75t_L g481 ( 
.A(n_394),
.B(n_357),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_401),
.B(n_353),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_401),
.A2(n_224),
.B1(n_203),
.B2(n_223),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_385),
.A2(n_173),
.B1(n_229),
.B2(n_178),
.Y(n_484)
);

AND2x4_ASAP7_75t_L g485 ( 
.A(n_394),
.B(n_321),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_L g486 ( 
.A1(n_364),
.A2(n_221),
.B1(n_218),
.B2(n_225),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_364),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_364),
.B(n_340),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_363),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_364),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_364),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_401),
.B(n_180),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_392),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_488),
.Y(n_494)
);

AND2x2_ASAP7_75t_SL g495 ( 
.A(n_434),
.B(n_205),
.Y(n_495)
);

INVx4_ASAP7_75t_L g496 ( 
.A(n_442),
.Y(n_496)
);

OR2x2_ASAP7_75t_L g497 ( 
.A(n_415),
.B(n_0),
.Y(n_497)
);

INVx3_ASAP7_75t_L g498 ( 
.A(n_442),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_492),
.B(n_185),
.Y(n_499)
);

BUFx6f_ASAP7_75t_L g500 ( 
.A(n_408),
.Y(n_500)
);

AND2x4_ASAP7_75t_L g501 ( 
.A(n_412),
.B(n_201),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_488),
.Y(n_502)
);

HB1xp67_ASAP7_75t_L g503 ( 
.A(n_433),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_408),
.Y(n_504)
);

HB1xp67_ASAP7_75t_L g505 ( 
.A(n_433),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_412),
.B(n_217),
.Y(n_506)
);

OA21x2_ASAP7_75t_L g507 ( 
.A1(n_449),
.A2(n_229),
.B(n_207),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_416),
.Y(n_508)
);

INVx3_ASAP7_75t_L g509 ( 
.A(n_442),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_470),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_423),
.B(n_0),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_470),
.Y(n_512)
);

AND2x4_ASAP7_75t_SL g513 ( 
.A(n_408),
.B(n_205),
.Y(n_513)
);

HB1xp67_ASAP7_75t_L g514 ( 
.A(n_414),
.Y(n_514)
);

BUFx3_ASAP7_75t_L g515 ( 
.A(n_442),
.Y(n_515)
);

HB1xp67_ASAP7_75t_L g516 ( 
.A(n_414),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_451),
.B(n_206),
.Y(n_517)
);

HB1xp67_ASAP7_75t_L g518 ( 
.A(n_414),
.Y(n_518)
);

AND2x4_ASAP7_75t_L g519 ( 
.A(n_479),
.B(n_41),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_411),
.B(n_1),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_436),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_407),
.B(n_177),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_475),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_475),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_441),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_442),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_418),
.B(n_1),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_409),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_417),
.B(n_177),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_420),
.B(n_432),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_425),
.B(n_177),
.Y(n_531)
);

INVx3_ASAP7_75t_L g532 ( 
.A(n_421),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_468),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_472),
.Y(n_534)
);

NAND2xp33_ASAP7_75t_L g535 ( 
.A(n_421),
.B(n_177),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_473),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_441),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_476),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_487),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_490),
.Y(n_540)
);

AND2x4_ASAP7_75t_L g541 ( 
.A(n_421),
.B(n_42),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_L g542 ( 
.A1(n_415),
.A2(n_212),
.B1(n_208),
.B2(n_209),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_465),
.Y(n_543)
);

BUFx3_ASAP7_75t_L g544 ( 
.A(n_438),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_471),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_491),
.B(n_177),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_474),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_493),
.Y(n_548)
);

AND2x4_ASAP7_75t_L g549 ( 
.A(n_428),
.B(n_43),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_424),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_528),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_543),
.Y(n_552)
);

OAI22xp5_ASAP7_75t_SL g553 ( 
.A1(n_495),
.A2(n_419),
.B1(n_434),
.B2(n_492),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_544),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_499),
.B(n_464),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_503),
.B(n_422),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_495),
.B(n_437),
.Y(n_557)
);

OAI22xp33_ASAP7_75t_SL g558 ( 
.A1(n_499),
.A2(n_486),
.B1(n_469),
.B2(n_467),
.Y(n_558)
);

OAI22xp33_ASAP7_75t_L g559 ( 
.A1(n_497),
.A2(n_483),
.B1(n_443),
.B2(n_427),
.Y(n_559)
);

AOI22xp5_ASAP7_75t_L g560 ( 
.A1(n_495),
.A2(n_422),
.B1(n_462),
.B2(n_478),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_543),
.Y(n_561)
);

INVxp67_ASAP7_75t_L g562 ( 
.A(n_503),
.Y(n_562)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_530),
.B(n_437),
.Y(n_563)
);

AOI22xp5_ASAP7_75t_L g564 ( 
.A1(n_550),
.A2(n_489),
.B1(n_478),
.B2(n_410),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_543),
.Y(n_565)
);

AND2x2_ASAP7_75t_L g566 ( 
.A(n_530),
.B(n_437),
.Y(n_566)
);

AND2x2_ASAP7_75t_SL g567 ( 
.A(n_496),
.B(n_439),
.Y(n_567)
);

AND2x4_ASAP7_75t_L g568 ( 
.A(n_515),
.B(n_439),
.Y(n_568)
);

NAND3x1_ASAP7_75t_L g569 ( 
.A(n_528),
.B(n_457),
.C(n_447),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_530),
.B(n_439),
.Y(n_570)
);

OAI22xp5_ASAP7_75t_L g571 ( 
.A1(n_550),
.A2(n_482),
.B1(n_424),
.B2(n_426),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_545),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_533),
.Y(n_573)
);

AO22x2_ASAP7_75t_L g574 ( 
.A1(n_525),
.A2(n_486),
.B1(n_469),
.B2(n_467),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_520),
.B(n_446),
.Y(n_575)
);

OAI22xp33_ASAP7_75t_L g576 ( 
.A1(n_497),
.A2(n_453),
.B1(n_440),
.B2(n_445),
.Y(n_576)
);

OAI22xp33_ASAP7_75t_L g577 ( 
.A1(n_497),
.A2(n_453),
.B1(n_445),
.B2(n_454),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_545),
.Y(n_578)
);

OA22x2_ASAP7_75t_L g579 ( 
.A1(n_505),
.A2(n_460),
.B1(n_481),
.B2(n_450),
.Y(n_579)
);

OAI22xp5_ASAP7_75t_L g580 ( 
.A1(n_510),
.A2(n_482),
.B1(n_523),
.B2(n_512),
.Y(n_580)
);

OAI22xp33_ASAP7_75t_SL g581 ( 
.A1(n_542),
.A2(n_460),
.B1(n_450),
.B2(n_458),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_520),
.B(n_446),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_533),
.Y(n_583)
);

OAI22xp33_ASAP7_75t_L g584 ( 
.A1(n_496),
.A2(n_453),
.B1(n_454),
.B2(n_455),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_534),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_545),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_544),
.Y(n_587)
);

OAI22xp33_ASAP7_75t_SL g588 ( 
.A1(n_542),
.A2(n_458),
.B1(n_430),
.B2(n_448),
.Y(n_588)
);

OAI22xp33_ASAP7_75t_SL g589 ( 
.A1(n_510),
.A2(n_448),
.B1(n_426),
.B2(n_430),
.Y(n_589)
);

AO22x2_ASAP7_75t_L g590 ( 
.A1(n_525),
.A2(n_481),
.B1(n_485),
.B2(n_452),
.Y(n_590)
);

AO22x2_ASAP7_75t_L g591 ( 
.A1(n_525),
.A2(n_537),
.B1(n_523),
.B2(n_524),
.Y(n_591)
);

INVx3_ASAP7_75t_L g592 ( 
.A(n_567),
.Y(n_592)
);

BUFx3_ASAP7_75t_L g593 ( 
.A(n_554),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_555),
.B(n_505),
.Y(n_594)
);

HB1xp67_ASAP7_75t_L g595 ( 
.A(n_562),
.Y(n_595)
);

AOI22xp5_ASAP7_75t_L g596 ( 
.A1(n_553),
.A2(n_527),
.B1(n_520),
.B2(n_524),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_591),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_552),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_564),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_552),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_554),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_561),
.Y(n_602)
);

INVx1_ASAP7_75t_SL g603 ( 
.A(n_587),
.Y(n_603)
);

BUFx10_ASAP7_75t_L g604 ( 
.A(n_568),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_580),
.B(n_500),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_561),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_591),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_591),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_565),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_565),
.Y(n_610)
);

INVx3_ASAP7_75t_L g611 ( 
.A(n_567),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_572),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_572),
.Y(n_613)
);

BUFx6f_ASAP7_75t_SL g614 ( 
.A(n_568),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_577),
.B(n_500),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_578),
.Y(n_616)
);

BUFx2_ASAP7_75t_L g617 ( 
.A(n_590),
.Y(n_617)
);

CKINVDCx20_ASAP7_75t_R g618 ( 
.A(n_587),
.Y(n_618)
);

INVxp67_ASAP7_75t_SL g619 ( 
.A(n_571),
.Y(n_619)
);

BUFx6f_ASAP7_75t_L g620 ( 
.A(n_568),
.Y(n_620)
);

AOI21x1_ASAP7_75t_L g621 ( 
.A1(n_574),
.A2(n_521),
.B(n_507),
.Y(n_621)
);

BUFx6f_ASAP7_75t_L g622 ( 
.A(n_575),
.Y(n_622)
);

OAI21xp33_ASAP7_75t_SL g623 ( 
.A1(n_551),
.A2(n_512),
.B(n_496),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_586),
.Y(n_624)
);

OAI22xp5_ASAP7_75t_L g625 ( 
.A1(n_559),
.A2(n_560),
.B1(n_576),
.B2(n_496),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_573),
.Y(n_626)
);

BUFx6f_ASAP7_75t_L g627 ( 
.A(n_575),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_583),
.Y(n_628)
);

AOI22xp33_ASAP7_75t_L g629 ( 
.A1(n_558),
.A2(n_485),
.B1(n_502),
.B2(n_494),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_585),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_590),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_563),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_590),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_563),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_589),
.Y(n_635)
);

INVxp33_ASAP7_75t_SL g636 ( 
.A(n_556),
.Y(n_636)
);

INVx3_ASAP7_75t_L g637 ( 
.A(n_582),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_566),
.Y(n_638)
);

NAND2xp33_ASAP7_75t_L g639 ( 
.A(n_569),
.B(n_454),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_566),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_570),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_570),
.Y(n_642)
);

INVx2_ASAP7_75t_SL g643 ( 
.A(n_582),
.Y(n_643)
);

AND2x2_ASAP7_75t_SL g644 ( 
.A(n_557),
.B(n_496),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_574),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_584),
.B(n_527),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_557),
.B(n_527),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_581),
.B(n_588),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_574),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_579),
.B(n_500),
.Y(n_650)
);

INVx3_ASAP7_75t_L g651 ( 
.A(n_569),
.Y(n_651)
);

BUFx3_ASAP7_75t_L g652 ( 
.A(n_579),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_591),
.Y(n_653)
);

NAND2xp33_ASAP7_75t_L g654 ( 
.A(n_553),
.B(n_455),
.Y(n_654)
);

BUFx4f_ASAP7_75t_L g655 ( 
.A(n_567),
.Y(n_655)
);

INVxp67_ASAP7_75t_L g656 ( 
.A(n_556),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_580),
.B(n_500),
.Y(n_657)
);

INVx2_ASAP7_75t_SL g658 ( 
.A(n_563),
.Y(n_658)
);

INVx3_ASAP7_75t_L g659 ( 
.A(n_567),
.Y(n_659)
);

NAND2xp33_ASAP7_75t_SL g660 ( 
.A(n_571),
.B(n_410),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_591),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_580),
.B(n_500),
.Y(n_662)
);

INVx2_ASAP7_75t_SL g663 ( 
.A(n_563),
.Y(n_663)
);

BUFx6f_ASAP7_75t_L g664 ( 
.A(n_567),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_552),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_552),
.Y(n_666)
);

INVxp67_ASAP7_75t_L g667 ( 
.A(n_556),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_564),
.B(n_429),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_552),
.Y(n_669)
);

BUFx10_ASAP7_75t_L g670 ( 
.A(n_568),
.Y(n_670)
);

INVx3_ASAP7_75t_L g671 ( 
.A(n_567),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_552),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_594),
.B(n_534),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_598),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_626),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_619),
.B(n_536),
.Y(n_676)
);

INVx3_ASAP7_75t_L g677 ( 
.A(n_622),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_598),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_626),
.Y(n_679)
);

INVx5_ASAP7_75t_L g680 ( 
.A(n_664),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_601),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_638),
.B(n_544),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_660),
.B(n_500),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_595),
.B(n_536),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_600),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_628),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_628),
.Y(n_687)
);

BUFx3_ASAP7_75t_L g688 ( 
.A(n_593),
.Y(n_688)
);

INVx3_ASAP7_75t_L g689 ( 
.A(n_622),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_625),
.B(n_500),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_630),
.Y(n_691)
);

AND2x6_ASAP7_75t_L g692 ( 
.A(n_664),
.B(n_515),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_638),
.B(n_514),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_655),
.B(n_596),
.Y(n_694)
);

BUFx3_ASAP7_75t_L g695 ( 
.A(n_593),
.Y(n_695)
);

INVx2_ASAP7_75t_SL g696 ( 
.A(n_601),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_656),
.B(n_538),
.Y(n_697)
);

INVx5_ASAP7_75t_L g698 ( 
.A(n_664),
.Y(n_698)
);

INVxp67_ASAP7_75t_L g699 ( 
.A(n_635),
.Y(n_699)
);

OR2x6_ASAP7_75t_L g700 ( 
.A(n_651),
.B(n_515),
.Y(n_700)
);

BUFx2_ASAP7_75t_L g701 ( 
.A(n_618),
.Y(n_701)
);

AND2x4_ASAP7_75t_L g702 ( 
.A(n_637),
.B(n_541),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_637),
.B(n_514),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_599),
.B(n_532),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_599),
.B(n_636),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_636),
.B(n_654),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_655),
.B(n_504),
.Y(n_707)
);

XOR2xp5_ASAP7_75t_L g708 ( 
.A(n_632),
.B(n_413),
.Y(n_708)
);

BUFx3_ASAP7_75t_L g709 ( 
.A(n_622),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_637),
.B(n_516),
.Y(n_710)
);

AO21x2_ASAP7_75t_L g711 ( 
.A1(n_621),
.A2(n_650),
.B(n_648),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_667),
.B(n_538),
.Y(n_712)
);

INVx5_ASAP7_75t_L g713 ( 
.A(n_664),
.Y(n_713)
);

AND2x2_ASAP7_75t_SL g714 ( 
.A(n_617),
.B(n_513),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_630),
.Y(n_715)
);

INVx2_ASAP7_75t_SL g716 ( 
.A(n_603),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_609),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_639),
.B(n_532),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_655),
.B(n_596),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_622),
.B(n_516),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_609),
.Y(n_721)
);

CKINVDCx20_ASAP7_75t_R g722 ( 
.A(n_668),
.Y(n_722)
);

INVx3_ASAP7_75t_L g723 ( 
.A(n_622),
.Y(n_723)
);

INVx4_ASAP7_75t_L g724 ( 
.A(n_620),
.Y(n_724)
);

INVx2_ASAP7_75t_SL g725 ( 
.A(n_627),
.Y(n_725)
);

OAI22xp5_ASAP7_75t_L g726 ( 
.A1(n_629),
.A2(n_498),
.B1(n_526),
.B2(n_509),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_613),
.Y(n_727)
);

BUFx6f_ASAP7_75t_L g728 ( 
.A(n_620),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_600),
.Y(n_729)
);

AND2x4_ASAP7_75t_L g730 ( 
.A(n_632),
.B(n_541),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_651),
.B(n_504),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_L g732 ( 
.A(n_635),
.B(n_532),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_613),
.Y(n_733)
);

INVx5_ASAP7_75t_L g734 ( 
.A(n_664),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_616),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_602),
.Y(n_736)
);

AND2x4_ASAP7_75t_L g737 ( 
.A(n_634),
.B(n_541),
.Y(n_737)
);

INVx3_ASAP7_75t_L g738 ( 
.A(n_627),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_616),
.Y(n_739)
);

INVx2_ASAP7_75t_SL g740 ( 
.A(n_627),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_634),
.B(n_539),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_624),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_651),
.B(n_504),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_640),
.B(n_539),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_640),
.B(n_540),
.Y(n_745)
);

INVx3_ASAP7_75t_L g746 ( 
.A(n_627),
.Y(n_746)
);

CKINVDCx16_ASAP7_75t_R g747 ( 
.A(n_614),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_624),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_602),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_606),
.Y(n_750)
);

INVx2_ASAP7_75t_SL g751 ( 
.A(n_627),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_641),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_606),
.Y(n_753)
);

INVx4_ASAP7_75t_L g754 ( 
.A(n_620),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_610),
.Y(n_755)
);

AND2x4_ASAP7_75t_L g756 ( 
.A(n_643),
.B(n_549),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_641),
.B(n_540),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_706),
.B(n_489),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_722),
.B(n_429),
.Y(n_759)
);

AOI21xp5_ASAP7_75t_L g760 ( 
.A1(n_683),
.A2(n_623),
.B(n_605),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_673),
.B(n_645),
.Y(n_761)
);

INVx3_ASAP7_75t_L g762 ( 
.A(n_688),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_676),
.B(n_645),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_693),
.B(n_643),
.Y(n_764)
);

AND2x4_ASAP7_75t_L g765 ( 
.A(n_709),
.B(n_700),
.Y(n_765)
);

NOR2xp67_ASAP7_75t_L g766 ( 
.A(n_716),
.B(n_623),
.Y(n_766)
);

BUFx6f_ASAP7_75t_L g767 ( 
.A(n_728),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_699),
.B(n_649),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_691),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_706),
.B(n_455),
.Y(n_770)
);

INVxp67_ASAP7_75t_L g771 ( 
.A(n_705),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_675),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_679),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_686),
.Y(n_774)
);

NOR2xp67_ASAP7_75t_L g775 ( 
.A(n_699),
.B(n_457),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_687),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_684),
.B(n_649),
.Y(n_777)
);

NAND2xp33_ASAP7_75t_L g778 ( 
.A(n_681),
.B(n_456),
.Y(n_778)
);

INVx2_ASAP7_75t_SL g779 ( 
.A(n_688),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_715),
.Y(n_780)
);

INVxp67_ASAP7_75t_L g781 ( 
.A(n_705),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_722),
.B(n_456),
.Y(n_782)
);

NOR3xp33_ASAP7_75t_L g783 ( 
.A(n_683),
.B(n_517),
.C(n_657),
.Y(n_783)
);

BUFx3_ASAP7_75t_L g784 ( 
.A(n_701),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_752),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_674),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_704),
.B(n_456),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_704),
.B(n_695),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_674),
.Y(n_789)
);

INVxp67_ASAP7_75t_SL g790 ( 
.A(n_731),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_741),
.B(n_744),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_717),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_745),
.B(n_597),
.Y(n_793)
);

INVxp67_ASAP7_75t_L g794 ( 
.A(n_695),
.Y(n_794)
);

XOR2xp5_ASAP7_75t_L g795 ( 
.A(n_708),
.B(n_444),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_721),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_697),
.B(n_712),
.Y(n_797)
);

BUFx6f_ASAP7_75t_L g798 ( 
.A(n_728),
.Y(n_798)
);

HB1xp67_ASAP7_75t_L g799 ( 
.A(n_711),
.Y(n_799)
);

NOR3xp33_ASAP7_75t_L g800 ( 
.A(n_732),
.B(n_662),
.C(n_615),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_732),
.B(n_642),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_727),
.Y(n_802)
);

NAND3xp33_ASAP7_75t_L g803 ( 
.A(n_690),
.B(n_484),
.C(n_646),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_757),
.B(n_597),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_SL g805 ( 
.A(n_747),
.B(n_477),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_696),
.B(n_620),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_703),
.B(n_642),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_718),
.B(n_620),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_718),
.B(n_658),
.Y(n_809)
);

INVx2_ASAP7_75t_SL g810 ( 
.A(n_682),
.Y(n_810)
);

AND2x2_ASAP7_75t_L g811 ( 
.A(n_709),
.B(n_658),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_681),
.B(n_461),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_733),
.B(n_607),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_735),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_739),
.Y(n_815)
);

BUFx6f_ASAP7_75t_L g816 ( 
.A(n_728),
.Y(n_816)
);

INVx3_ASAP7_75t_L g817 ( 
.A(n_677),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_678),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_742),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_724),
.B(n_463),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_748),
.B(n_607),
.Y(n_821)
);

BUFx6f_ASAP7_75t_L g822 ( 
.A(n_728),
.Y(n_822)
);

NOR2xp67_ASAP7_75t_L g823 ( 
.A(n_680),
.B(n_608),
.Y(n_823)
);

INVx4_ASAP7_75t_L g824 ( 
.A(n_724),
.Y(n_824)
);

NOR2xp67_ASAP7_75t_L g825 ( 
.A(n_680),
.B(n_608),
.Y(n_825)
);

AOI22xp33_ASAP7_75t_L g826 ( 
.A1(n_694),
.A2(n_652),
.B1(n_617),
.B2(n_633),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_694),
.B(n_663),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_711),
.B(n_653),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_719),
.B(n_663),
.Y(n_829)
);

INVx3_ASAP7_75t_L g830 ( 
.A(n_677),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_731),
.B(n_653),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_719),
.B(n_644),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_775),
.B(n_754),
.Y(n_833)
);

INVx3_ASAP7_75t_L g834 ( 
.A(n_762),
.Y(n_834)
);

A2O1A1Ixp33_ASAP7_75t_L g835 ( 
.A1(n_803),
.A2(n_652),
.B(n_690),
.C(n_714),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_786),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_797),
.B(n_791),
.Y(n_837)
);

AOI22xp33_ASAP7_75t_L g838 ( 
.A1(n_800),
.A2(n_647),
.B1(n_633),
.B2(n_631),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_791),
.B(n_710),
.Y(n_839)
);

AND2x4_ASAP7_75t_SL g840 ( 
.A(n_765),
.B(n_720),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_771),
.B(n_743),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_L g842 ( 
.A(n_759),
.B(n_463),
.Y(n_842)
);

AOI22xp33_ASAP7_75t_L g843 ( 
.A1(n_826),
.A2(n_631),
.B1(n_547),
.B2(n_548),
.Y(n_843)
);

NOR2xp33_ASAP7_75t_L g844 ( 
.A(n_781),
.B(n_743),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_766),
.B(n_754),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_784),
.Y(n_846)
);

AND2x6_ASAP7_75t_SL g847 ( 
.A(n_812),
.B(n_431),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_772),
.Y(n_848)
);

A2O1A1Ixp33_ASAP7_75t_L g849 ( 
.A1(n_760),
.A2(n_714),
.B(n_661),
.C(n_541),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_789),
.Y(n_850)
);

INVxp67_ASAP7_75t_L g851 ( 
.A(n_782),
.Y(n_851)
);

AOI22xp33_ASAP7_75t_L g852 ( 
.A1(n_832),
.A2(n_547),
.B1(n_548),
.B2(n_501),
.Y(n_852)
);

AOI22xp5_ASAP7_75t_L g853 ( 
.A1(n_783),
.A2(n_700),
.B1(n_756),
.B2(n_692),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_763),
.B(n_689),
.Y(n_854)
);

AOI22xp33_ASAP7_75t_L g855 ( 
.A1(n_795),
.A2(n_501),
.B1(n_737),
.B2(n_730),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_L g856 ( 
.A(n_778),
.B(n_431),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_805),
.B(n_466),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_SL g858 ( 
.A(n_762),
.B(n_779),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_818),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_763),
.B(n_764),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_794),
.B(n_689),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_758),
.B(n_466),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_SL g863 ( 
.A(n_820),
.B(n_725),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_769),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_773),
.B(n_723),
.Y(n_865)
);

INVx1_ASAP7_75t_SL g866 ( 
.A(n_810),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_774),
.B(n_723),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_780),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_776),
.B(n_738),
.Y(n_869)
);

NAND3xp33_ASAP7_75t_L g870 ( 
.A(n_799),
.B(n_707),
.C(n_740),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_777),
.B(n_738),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_785),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_L g873 ( 
.A(n_788),
.B(n_746),
.Y(n_873)
);

AND2x4_ASAP7_75t_SL g874 ( 
.A(n_765),
.B(n_746),
.Y(n_874)
);

NAND3xp33_ASAP7_75t_L g875 ( 
.A(n_828),
.B(n_831),
.C(n_790),
.Y(n_875)
);

AND2x2_ASAP7_75t_L g876 ( 
.A(n_811),
.B(n_751),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_792),
.Y(n_877)
);

BUFx8_ASAP7_75t_L g878 ( 
.A(n_767),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_777),
.B(n_707),
.Y(n_879)
);

INVxp67_ASAP7_75t_SL g880 ( 
.A(n_828),
.Y(n_880)
);

AOI22xp33_ASAP7_75t_L g881 ( 
.A1(n_768),
.A2(n_501),
.B1(n_737),
.B2(n_730),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_817),
.B(n_680),
.Y(n_882)
);

O2A1O1Ixp33_ASAP7_75t_L g883 ( 
.A1(n_787),
.A2(n_459),
.B(n_726),
.C(n_506),
.Y(n_883)
);

AND2x6_ASAP7_75t_SL g884 ( 
.A(n_801),
.B(n_435),
.Y(n_884)
);

BUFx3_ASAP7_75t_L g885 ( 
.A(n_807),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_SL g886 ( 
.A(n_770),
.B(n_680),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_796),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_802),
.B(n_661),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_806),
.B(n_592),
.Y(n_889)
);

OAI22xp5_ASAP7_75t_L g890 ( 
.A1(n_827),
.A2(n_700),
.B1(n_611),
.B2(n_659),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_767),
.Y(n_891)
);

NOR2xp33_ASAP7_75t_L g892 ( 
.A(n_809),
.B(n_592),
.Y(n_892)
);

OAI22xp33_ASAP7_75t_L g893 ( 
.A1(n_829),
.A2(n_592),
.B1(n_659),
.B2(n_611),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_814),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_824),
.B(n_698),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_815),
.B(n_702),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_L g897 ( 
.A(n_819),
.B(n_611),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_761),
.B(n_702),
.Y(n_898)
);

OAI22xp5_ASAP7_75t_L g899 ( 
.A1(n_808),
.A2(n_659),
.B1(n_671),
.B2(n_644),
.Y(n_899)
);

BUFx3_ASAP7_75t_L g900 ( 
.A(n_767),
.Y(n_900)
);

NOR3xp33_ASAP7_75t_L g901 ( 
.A(n_817),
.B(n_621),
.C(n_506),
.Y(n_901)
);

NOR2xp33_ASAP7_75t_L g902 ( 
.A(n_830),
.B(n_671),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_SL g903 ( 
.A(n_824),
.B(n_698),
.Y(n_903)
);

NOR2xp33_ASAP7_75t_L g904 ( 
.A(n_798),
.B(n_438),
.Y(n_904)
);

NOR2xp33_ASAP7_75t_L g905 ( 
.A(n_798),
.B(n_438),
.Y(n_905)
);

BUFx2_ASAP7_75t_SL g906 ( 
.A(n_798),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_SL g907 ( 
.A(n_816),
.B(n_698),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_813),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_761),
.B(n_831),
.Y(n_909)
);

O2A1O1Ixp33_ASAP7_75t_L g910 ( 
.A1(n_813),
.A2(n_511),
.B(n_518),
.C(n_501),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_816),
.B(n_698),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_793),
.B(n_730),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_821),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_908),
.Y(n_914)
);

AO22x2_ASAP7_75t_L g915 ( 
.A1(n_875),
.A2(n_768),
.B1(n_804),
.B2(n_793),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_837),
.B(n_804),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_913),
.Y(n_917)
);

BUFx2_ASAP7_75t_L g918 ( 
.A(n_834),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_877),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_848),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_841),
.B(n_830),
.Y(n_921)
);

OAI221xp5_ASAP7_75t_L g922 ( 
.A1(n_849),
.A2(n_821),
.B1(n_823),
.B2(n_825),
.C(n_671),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_887),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_894),
.Y(n_924)
);

INVx4_ASAP7_75t_L g925 ( 
.A(n_846),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_836),
.Y(n_926)
);

AOI22xp5_ASAP7_75t_L g927 ( 
.A1(n_835),
.A2(n_838),
.B1(n_893),
.B2(n_853),
.Y(n_927)
);

HB1xp67_ASAP7_75t_L g928 ( 
.A(n_854),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_872),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_909),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_888),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_L g932 ( 
.A(n_851),
.B(n_822),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_864),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_SL g934 ( 
.A(n_863),
.B(n_822),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_SL g935 ( 
.A(n_844),
.B(n_822),
.Y(n_935)
);

BUFx8_ASAP7_75t_L g936 ( 
.A(n_847),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_844),
.B(n_737),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_SL g938 ( 
.A(n_891),
.B(n_713),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_868),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_860),
.B(n_756),
.Y(n_940)
);

AO22x2_ASAP7_75t_L g941 ( 
.A1(n_880),
.A2(n_859),
.B1(n_850),
.B2(n_870),
.Y(n_941)
);

AO22x2_ASAP7_75t_L g942 ( 
.A1(n_866),
.A2(n_685),
.B1(n_729),
.B2(n_678),
.Y(n_942)
);

AND2x4_ASAP7_75t_L g943 ( 
.A(n_840),
.B(n_713),
.Y(n_943)
);

BUFx2_ASAP7_75t_L g944 ( 
.A(n_834),
.Y(n_944)
);

OAI221xp5_ASAP7_75t_L g945 ( 
.A1(n_883),
.A2(n_529),
.B1(n_522),
.B2(n_531),
.C(n_546),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_871),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_865),
.Y(n_947)
);

AND2x4_ASAP7_75t_L g948 ( 
.A(n_874),
.B(n_713),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_867),
.Y(n_949)
);

INVxp67_ASAP7_75t_L g950 ( 
.A(n_842),
.Y(n_950)
);

NAND2xp33_ASAP7_75t_L g951 ( 
.A(n_845),
.B(n_692),
.Y(n_951)
);

OAI221xp5_ASAP7_75t_L g952 ( 
.A1(n_879),
.A2(n_535),
.B1(n_518),
.B2(n_507),
.C(n_713),
.Y(n_952)
);

AO22x2_ASAP7_75t_L g953 ( 
.A1(n_890),
.A2(n_755),
.B1(n_753),
.B2(n_750),
.Y(n_953)
);

OAI221xp5_ASAP7_75t_L g954 ( 
.A1(n_855),
.A2(n_507),
.B1(n_734),
.B2(n_750),
.C(n_749),
.Y(n_954)
);

INVxp67_ASAP7_75t_L g955 ( 
.A(n_858),
.Y(n_955)
);

AO21x1_ASAP7_75t_L g956 ( 
.A1(n_893),
.A2(n_519),
.B(n_541),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_885),
.Y(n_957)
);

AO22x2_ASAP7_75t_L g958 ( 
.A1(n_899),
.A2(n_755),
.B1(n_753),
.B2(n_749),
.Y(n_958)
);

CKINVDCx20_ASAP7_75t_R g959 ( 
.A(n_878),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_869),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_839),
.Y(n_961)
);

NAND2x1p5_ASAP7_75t_L g962 ( 
.A(n_900),
.B(n_734),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_898),
.B(n_734),
.Y(n_963)
);

AO22x2_ASAP7_75t_L g964 ( 
.A1(n_896),
.A2(n_736),
.B1(n_685),
.B2(n_729),
.Y(n_964)
);

AO22x2_ASAP7_75t_L g965 ( 
.A1(n_912),
.A2(n_736),
.B1(n_669),
.B2(n_666),
.Y(n_965)
);

AOI22xp5_ASAP7_75t_L g966 ( 
.A1(n_892),
.A2(n_692),
.B1(n_644),
.B2(n_614),
.Y(n_966)
);

AO22x2_ASAP7_75t_L g967 ( 
.A1(n_861),
.A2(n_665),
.B1(n_612),
.B2(n_672),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_876),
.Y(n_968)
);

AND2x6_ASAP7_75t_SL g969 ( 
.A(n_936),
.B(n_857),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_930),
.B(n_950),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_951),
.A2(n_833),
.B(n_886),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_931),
.B(n_884),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_SL g973 ( 
.A(n_956),
.B(n_873),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_947),
.B(n_897),
.Y(n_974)
);

AND2x6_ASAP7_75t_L g975 ( 
.A(n_927),
.B(n_856),
.Y(n_975)
);

CKINVDCx11_ASAP7_75t_R g976 ( 
.A(n_959),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_949),
.B(n_960),
.Y(n_977)
);

OAI21xp33_ASAP7_75t_L g978 ( 
.A1(n_941),
.A2(n_897),
.B(n_873),
.Y(n_978)
);

BUFx6f_ASAP7_75t_L g979 ( 
.A(n_925),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_915),
.A2(n_903),
.B(n_895),
.Y(n_980)
);

AOI21x1_ASAP7_75t_L g981 ( 
.A1(n_941),
.A2(n_911),
.B(n_907),
.Y(n_981)
);

AOI22xp5_ASAP7_75t_L g982 ( 
.A1(n_915),
.A2(n_958),
.B1(n_961),
.B2(n_945),
.Y(n_982)
);

AND2x2_ASAP7_75t_L g983 ( 
.A(n_955),
.B(n_882),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_914),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_934),
.A2(n_910),
.B(n_892),
.Y(n_985)
);

NOR3xp33_ASAP7_75t_L g986 ( 
.A(n_952),
.B(n_862),
.C(n_901),
.Y(n_986)
);

BUFx6f_ASAP7_75t_L g987 ( 
.A(n_962),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_916),
.B(n_943),
.Y(n_988)
);

CKINVDCx20_ASAP7_75t_R g989 ( 
.A(n_932),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_L g990 ( 
.A(n_921),
.B(n_904),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_942),
.Y(n_991)
);

AO21x1_ASAP7_75t_L g992 ( 
.A1(n_920),
.A2(n_889),
.B(n_905),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_942),
.Y(n_993)
);

OAI22xp5_ASAP7_75t_L g994 ( 
.A1(n_966),
.A2(n_889),
.B1(n_855),
.B2(n_902),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_935),
.A2(n_902),
.B(n_852),
.Y(n_995)
);

INVx4_ASAP7_75t_L g996 ( 
.A(n_918),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_938),
.A2(n_852),
.B(n_881),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_946),
.B(n_881),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_922),
.A2(n_843),
.B(n_734),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_SL g1000 ( 
.A(n_943),
.B(n_928),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_917),
.B(n_878),
.Y(n_1001)
);

CKINVDCx10_ASAP7_75t_R g1002 ( 
.A(n_957),
.Y(n_1002)
);

NAND2x1p5_ASAP7_75t_L g1003 ( 
.A(n_948),
.B(n_549),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_923),
.B(n_906),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_964),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_924),
.B(n_919),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_929),
.B(n_843),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_937),
.B(n_507),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_963),
.A2(n_958),
.B(n_954),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_953),
.A2(n_507),
.B(n_549),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_940),
.B(n_692),
.Y(n_1011)
);

OR2x2_ASAP7_75t_L g1012 ( 
.A(n_968),
.B(n_944),
.Y(n_1012)
);

AOI21x1_ASAP7_75t_L g1013 ( 
.A1(n_953),
.A2(n_521),
.B(n_537),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_933),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_964),
.B(n_692),
.Y(n_1015)
);

AOI22xp5_ASAP7_75t_L g1016 ( 
.A1(n_967),
.A2(n_614),
.B1(n_549),
.B2(n_501),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_965),
.B(n_511),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_965),
.B(n_177),
.Y(n_1018)
);

AOI22xp5_ASAP7_75t_L g1019 ( 
.A1(n_967),
.A2(n_604),
.B1(n_670),
.B2(n_513),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_926),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_939),
.B(n_2),
.Y(n_1021)
);

O2A1O1Ixp33_ASAP7_75t_L g1022 ( 
.A1(n_950),
.A2(n_519),
.B(n_526),
.C(n_498),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_914),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_930),
.B(n_2),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_SL g1025 ( 
.A(n_950),
.B(n_604),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_936),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_SL g1027 ( 
.A(n_950),
.B(n_604),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_930),
.B(n_3),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_SL g1029 ( 
.A(n_936),
.B(n_604),
.Y(n_1029)
);

A2O1A1Ixp33_ASAP7_75t_L g1030 ( 
.A1(n_927),
.A2(n_509),
.B(n_498),
.C(n_526),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_1013),
.Y(n_1031)
);

BUFx3_ASAP7_75t_L g1032 ( 
.A(n_1026),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_SL g1033 ( 
.A(n_992),
.B(n_981),
.Y(n_1033)
);

BUFx6f_ASAP7_75t_L g1034 ( 
.A(n_976),
.Y(n_1034)
);

INVx5_ASAP7_75t_L g1035 ( 
.A(n_969),
.Y(n_1035)
);

INVx5_ASAP7_75t_L g1036 ( 
.A(n_975),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_1006),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_985),
.B(n_3),
.Y(n_1038)
);

CKINVDCx8_ASAP7_75t_R g1039 ( 
.A(n_979),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_1005),
.Y(n_1040)
);

OR2x2_ASAP7_75t_SL g1041 ( 
.A(n_972),
.B(n_508),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_991),
.Y(n_1042)
);

BUFx6f_ASAP7_75t_L g1043 ( 
.A(n_979),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_L g1044 ( 
.A(n_979),
.B(n_4),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_975),
.B(n_4),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_977),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_984),
.Y(n_1047)
);

AND2x2_ASAP7_75t_L g1048 ( 
.A(n_996),
.B(n_983),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_975),
.B(n_5),
.Y(n_1049)
);

BUFx6f_ASAP7_75t_L g1050 ( 
.A(n_1018),
.Y(n_1050)
);

NAND2x1p5_ASAP7_75t_L g1051 ( 
.A(n_996),
.B(n_509),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_L g1052 ( 
.A(n_1034),
.B(n_989),
.Y(n_1052)
);

NOR2xp33_ASAP7_75t_L g1053 ( 
.A(n_1034),
.B(n_1002),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_1041),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_1046),
.B(n_1037),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_1047),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_1041),
.Y(n_1057)
);

INVxp67_ASAP7_75t_L g1058 ( 
.A(n_1034),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_1040),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_L g1060 ( 
.A(n_1034),
.B(n_973),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_1033),
.A2(n_978),
.B(n_1009),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_1045),
.B(n_975),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_SL g1063 ( 
.A(n_1036),
.B(n_980),
.Y(n_1063)
);

CKINVDCx10_ASAP7_75t_R g1064 ( 
.A(n_1032),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_1033),
.A2(n_982),
.B(n_998),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_1049),
.B(n_986),
.Y(n_1066)
);

AND2x4_ASAP7_75t_L g1067 ( 
.A(n_1048),
.B(n_1000),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_1036),
.A2(n_970),
.B(n_1024),
.Y(n_1068)
);

CKINVDCx20_ASAP7_75t_R g1069 ( 
.A(n_1034),
.Y(n_1069)
);

NOR2xp33_ASAP7_75t_L g1070 ( 
.A(n_1032),
.B(n_1028),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_1040),
.Y(n_1071)
);

AOI22xp5_ASAP7_75t_L g1072 ( 
.A1(n_1038),
.A2(n_1017),
.B1(n_1007),
.B2(n_1016),
.Y(n_1072)
);

AOI22xp5_ASAP7_75t_L g1073 ( 
.A1(n_1036),
.A2(n_1008),
.B1(n_1015),
.B2(n_994),
.Y(n_1073)
);

BUFx2_ASAP7_75t_L g1074 ( 
.A(n_1043),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_1036),
.B(n_1023),
.Y(n_1075)
);

OAI22xp5_ASAP7_75t_L g1076 ( 
.A1(n_1036),
.A2(n_1030),
.B1(n_997),
.B2(n_995),
.Y(n_1076)
);

BUFx12f_ASAP7_75t_L g1077 ( 
.A(n_1064),
.Y(n_1077)
);

A2O1A1Ixp33_ASAP7_75t_L g1078 ( 
.A1(n_1061),
.A2(n_1035),
.B(n_1050),
.C(n_1031),
.Y(n_1078)
);

OAI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_1076),
.A2(n_1044),
.B(n_1035),
.Y(n_1079)
);

AOI21xp33_ASAP7_75t_L g1080 ( 
.A1(n_1076),
.A2(n_1050),
.B(n_1042),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_SL g1081 ( 
.A(n_1067),
.B(n_1035),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_1065),
.A2(n_1035),
.B(n_1048),
.Y(n_1082)
);

OAI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_1063),
.A2(n_1035),
.B(n_1051),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_1081),
.Y(n_1084)
);

OR2x2_ASAP7_75t_L g1085 ( 
.A(n_1082),
.B(n_1055),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_1084),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_1085),
.A2(n_1078),
.B(n_1079),
.Y(n_1087)
);

OR2x2_ASAP7_75t_L g1088 ( 
.A(n_1085),
.B(n_1058),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_1088),
.B(n_1066),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_1086),
.Y(n_1090)
);

INVx4_ASAP7_75t_L g1091 ( 
.A(n_1087),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_1091),
.Y(n_1092)
);

INVx6_ASAP7_75t_L g1093 ( 
.A(n_1091),
.Y(n_1093)
);

BUFx2_ASAP7_75t_SL g1094 ( 
.A(n_1092),
.Y(n_1094)
);

CKINVDCx6p67_ASAP7_75t_R g1095 ( 
.A(n_1093),
.Y(n_1095)
);

OA21x2_ASAP7_75t_L g1096 ( 
.A1(n_1095),
.A2(n_1089),
.B(n_1090),
.Y(n_1096)
);

OAI22xp5_ASAP7_75t_L g1097 ( 
.A1(n_1094),
.A2(n_1069),
.B1(n_1060),
.B2(n_1052),
.Y(n_1097)
);

AOI22xp33_ASAP7_75t_SL g1098 ( 
.A1(n_1096),
.A2(n_1077),
.B1(n_1050),
.B2(n_1070),
.Y(n_1098)
);

AOI22xp33_ASAP7_75t_L g1099 ( 
.A1(n_1097),
.A2(n_1080),
.B1(n_1050),
.B2(n_1042),
.Y(n_1099)
);

BUFx2_ASAP7_75t_L g1100 ( 
.A(n_1098),
.Y(n_1100)
);

BUFx6f_ASAP7_75t_L g1101 ( 
.A(n_1099),
.Y(n_1101)
);

OAI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_1100),
.A2(n_1068),
.B(n_1083),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_1101),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_1103),
.Y(n_1104)
);

AND2x2_ASAP7_75t_L g1105 ( 
.A(n_1102),
.B(n_1101),
.Y(n_1105)
);

BUFx3_ASAP7_75t_L g1106 ( 
.A(n_1103),
.Y(n_1106)
);

AND2x2_ASAP7_75t_L g1107 ( 
.A(n_1106),
.B(n_1053),
.Y(n_1107)
);

OR2x2_ASAP7_75t_L g1108 ( 
.A(n_1106),
.B(n_1074),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_1104),
.Y(n_1109)
);

HB1xp67_ASAP7_75t_L g1110 ( 
.A(n_1107),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_1108),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_1110),
.Y(n_1112)
);

BUFx2_ASAP7_75t_L g1113 ( 
.A(n_1111),
.Y(n_1113)
);

OR2x2_ASAP7_75t_L g1114 ( 
.A(n_1113),
.B(n_1109),
.Y(n_1114)
);

INVx3_ASAP7_75t_L g1115 ( 
.A(n_1112),
.Y(n_1115)
);

NOR3xp33_ASAP7_75t_L g1116 ( 
.A(n_1115),
.B(n_1105),
.C(n_1062),
.Y(n_1116)
);

OR2x2_ASAP7_75t_L g1117 ( 
.A(n_1114),
.B(n_1105),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_1117),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_1116),
.B(n_1059),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_1118),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1119),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_1120),
.Y(n_1122)
);

OA21x2_ASAP7_75t_L g1123 ( 
.A1(n_1121),
.A2(n_1067),
.B(n_1056),
.Y(n_1123)
);

OA21x2_ASAP7_75t_L g1124 ( 
.A1(n_1120),
.A2(n_1075),
.B(n_1071),
.Y(n_1124)
);

OAI22xp5_ASAP7_75t_L g1125 ( 
.A1(n_1122),
.A2(n_1039),
.B1(n_1043),
.B2(n_1075),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_1124),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1123),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1126),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1127),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_1129),
.B(n_1125),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1128),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_1131),
.B(n_1043),
.Y(n_1132)
);

HB1xp67_ASAP7_75t_L g1133 ( 
.A(n_1130),
.Y(n_1133)
);

NOR2xp67_ASAP7_75t_L g1134 ( 
.A(n_1133),
.B(n_5),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1132),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1135),
.Y(n_1136)
);

AOI22xp5_ASAP7_75t_L g1137 ( 
.A1(n_1134),
.A2(n_1043),
.B1(n_1050),
.B2(n_1072),
.Y(n_1137)
);

NOR3x1_ASAP7_75t_L g1138 ( 
.A(n_1136),
.B(n_1137),
.C(n_1039),
.Y(n_1138)
);

AOI22xp33_ASAP7_75t_L g1139 ( 
.A1(n_1136),
.A2(n_1054),
.B1(n_1057),
.B2(n_205),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1138),
.Y(n_1140)
);

OAI22xp5_ASAP7_75t_L g1141 ( 
.A1(n_1139),
.A2(n_1073),
.B1(n_210),
.B2(n_222),
.Y(n_1141)
);

OAI21xp5_ASAP7_75t_SL g1142 ( 
.A1(n_1138),
.A2(n_480),
.B(n_6),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_1140),
.B(n_6),
.Y(n_1143)
);

AND2x2_ASAP7_75t_L g1144 ( 
.A(n_1142),
.B(n_7),
.Y(n_1144)
);

OR2x2_ASAP7_75t_L g1145 ( 
.A(n_1141),
.B(n_8),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1143),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_1144),
.B(n_8),
.Y(n_1147)
);

NOR2xp33_ASAP7_75t_L g1148 ( 
.A(n_1147),
.B(n_1145),
.Y(n_1148)
);

NOR3xp33_ASAP7_75t_L g1149 ( 
.A(n_1146),
.B(n_220),
.C(n_215),
.Y(n_1149)
);

OAI22x1_ASAP7_75t_L g1150 ( 
.A1(n_1148),
.A2(n_993),
.B1(n_1021),
.B2(n_1001),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1149),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1151),
.Y(n_1152)
);

NOR2xp33_ASAP7_75t_L g1153 ( 
.A(n_1150),
.B(n_304),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_1152),
.A2(n_309),
.B(n_304),
.Y(n_1154)
);

XNOR2xp5_ASAP7_75t_L g1155 ( 
.A(n_1153),
.B(n_9),
.Y(n_1155)
);

NOR3xp33_ASAP7_75t_L g1156 ( 
.A(n_1154),
.B(n_9),
.C(n_10),
.Y(n_1156)
);

NAND4xp75_ASAP7_75t_L g1157 ( 
.A(n_1155),
.B(n_10),
.C(n_11),
.D(n_12),
.Y(n_1157)
);

NOR4xp25_ASAP7_75t_L g1158 ( 
.A(n_1157),
.B(n_1031),
.C(n_1004),
.D(n_990),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1156),
.Y(n_1159)
);

AOI22xp5_ASAP7_75t_L g1160 ( 
.A1(n_1156),
.A2(n_1029),
.B1(n_304),
.B2(n_309),
.Y(n_1160)
);

AOI211x1_ASAP7_75t_SL g1161 ( 
.A1(n_1159),
.A2(n_971),
.B(n_974),
.C(n_1027),
.Y(n_1161)
);

AOI221xp5_ASAP7_75t_L g1162 ( 
.A1(n_1158),
.A2(n_309),
.B1(n_987),
.B2(n_14),
.C(n_15),
.Y(n_1162)
);

AOI311xp33_ASAP7_75t_L g1163 ( 
.A1(n_1160),
.A2(n_1014),
.A3(n_13),
.B(n_14),
.C(n_15),
.Y(n_1163)
);

AOI22x1_ASAP7_75t_L g1164 ( 
.A1(n_1163),
.A2(n_309),
.B1(n_987),
.B2(n_16),
.Y(n_1164)
);

XNOR2xp5_ASAP7_75t_L g1165 ( 
.A(n_1162),
.B(n_11),
.Y(n_1165)
);

AOI211xp5_ASAP7_75t_L g1166 ( 
.A1(n_1165),
.A2(n_1161),
.B(n_16),
.C(n_17),
.Y(n_1166)
);

AOI221xp5_ASAP7_75t_L g1167 ( 
.A1(n_1164),
.A2(n_13),
.B1(n_17),
.B2(n_18),
.C(n_19),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1166),
.Y(n_1168)
);

XNOR2xp5_ASAP7_75t_L g1169 ( 
.A(n_1167),
.B(n_18),
.Y(n_1169)
);

NOR2x1_ASAP7_75t_L g1170 ( 
.A(n_1168),
.B(n_987),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1169),
.B(n_19),
.Y(n_1171)
);

NOR3xp33_ASAP7_75t_L g1172 ( 
.A(n_1171),
.B(n_20),
.C(n_21),
.Y(n_1172)
);

NOR2x1_ASAP7_75t_L g1173 ( 
.A(n_1170),
.B(n_21),
.Y(n_1173)
);

OAI321xp33_ASAP7_75t_L g1174 ( 
.A1(n_1172),
.A2(n_22),
.A3(n_24),
.B1(n_25),
.B2(n_26),
.C(n_27),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1173),
.Y(n_1175)
);

INVx1_ASAP7_75t_SL g1176 ( 
.A(n_1175),
.Y(n_1176)
);

BUFx6f_ASAP7_75t_L g1177 ( 
.A(n_1174),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1175),
.Y(n_1178)
);

AOI221xp5_ASAP7_75t_L g1179 ( 
.A1(n_1176),
.A2(n_22),
.B1(n_25),
.B2(n_26),
.C(n_27),
.Y(n_1179)
);

NOR3xp33_ASAP7_75t_L g1180 ( 
.A(n_1178),
.B(n_28),
.C(n_29),
.Y(n_1180)
);

BUFx4f_ASAP7_75t_SL g1181 ( 
.A(n_1177),
.Y(n_1181)
);

AOI22x1_ASAP7_75t_L g1182 ( 
.A1(n_1181),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_1182)
);

AOI22x1_ASAP7_75t_L g1183 ( 
.A1(n_1180),
.A2(n_31),
.B1(n_33),
.B2(n_34),
.Y(n_1183)
);

INVxp67_ASAP7_75t_SL g1184 ( 
.A(n_1183),
.Y(n_1184)
);

AOI22xp5_ASAP7_75t_L g1185 ( 
.A1(n_1182),
.A2(n_1179),
.B1(n_33),
.B2(n_34),
.Y(n_1185)
);

OAI22xp5_ASAP7_75t_L g1186 ( 
.A1(n_1184),
.A2(n_1051),
.B1(n_35),
.B2(n_36),
.Y(n_1186)
);

AND2x2_ASAP7_75t_L g1187 ( 
.A(n_1185),
.B(n_31),
.Y(n_1187)
);

OAI22xp5_ASAP7_75t_L g1188 ( 
.A1(n_1187),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_1188)
);

XNOR2x1_ASAP7_75t_L g1189 ( 
.A(n_1186),
.B(n_37),
.Y(n_1189)
);

OAI221xp5_ASAP7_75t_L g1190 ( 
.A1(n_1189),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.C(n_1012),
.Y(n_1190)
);

HB1xp67_ASAP7_75t_L g1191 ( 
.A(n_1188),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1191),
.Y(n_1192)
);

OAI21xp5_ASAP7_75t_SL g1193 ( 
.A1(n_1190),
.A2(n_38),
.B(n_39),
.Y(n_1193)
);

INVx2_ASAP7_75t_SL g1194 ( 
.A(n_1191),
.Y(n_1194)
);

OAI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_1192),
.A2(n_988),
.B(n_1025),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1194),
.Y(n_1196)
);

OR2x6_ASAP7_75t_L g1197 ( 
.A(n_1193),
.B(n_999),
.Y(n_1197)
);

AOI22x1_ASAP7_75t_L g1198 ( 
.A1(n_1192),
.A2(n_1003),
.B1(n_48),
.B2(n_49),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1196),
.Y(n_1199)
);

CKINVDCx20_ASAP7_75t_R g1200 ( 
.A(n_1197),
.Y(n_1200)
);

INVx1_ASAP7_75t_SL g1201 ( 
.A(n_1195),
.Y(n_1201)
);

AOI22xp33_ASAP7_75t_R g1202 ( 
.A1(n_1198),
.A2(n_45),
.B1(n_50),
.B2(n_51),
.Y(n_1202)
);

OAI22xp33_ASAP7_75t_L g1203 ( 
.A1(n_1199),
.A2(n_1011),
.B1(n_53),
.B2(n_54),
.Y(n_1203)
);

NAND2xp33_ASAP7_75t_L g1204 ( 
.A(n_1201),
.B(n_1200),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1202),
.B(n_52),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1199),
.Y(n_1206)
);

AOI221xp5_ASAP7_75t_L g1207 ( 
.A1(n_1199),
.A2(n_55),
.B1(n_56),
.B2(n_57),
.C(n_58),
.Y(n_1207)
);

AOI21xp33_ASAP7_75t_SL g1208 ( 
.A1(n_1199),
.A2(n_59),
.B(n_61),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1199),
.B(n_62),
.Y(n_1209)
);

OAI22xp5_ASAP7_75t_L g1210 ( 
.A1(n_1199),
.A2(n_63),
.B1(n_64),
.B2(n_65),
.Y(n_1210)
);

AOI22xp33_ASAP7_75t_SL g1211 ( 
.A1(n_1199),
.A2(n_66),
.B1(n_67),
.B2(n_69),
.Y(n_1211)
);

OAI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1199),
.A2(n_70),
.B(n_71),
.Y(n_1212)
);

AOI22xp5_ASAP7_75t_L g1213 ( 
.A1(n_1199),
.A2(n_72),
.B1(n_73),
.B2(n_74),
.Y(n_1213)
);

OAI22xp5_ASAP7_75t_SL g1214 ( 
.A1(n_1199),
.A2(n_75),
.B1(n_77),
.B2(n_78),
.Y(n_1214)
);

XNOR2x1_ASAP7_75t_L g1215 ( 
.A(n_1204),
.B(n_79),
.Y(n_1215)
);

O2A1O1Ixp33_ASAP7_75t_L g1216 ( 
.A1(n_1206),
.A2(n_81),
.B(n_82),
.C(n_83),
.Y(n_1216)
);

HB1xp67_ASAP7_75t_L g1217 ( 
.A(n_1212),
.Y(n_1217)
);

OR3x1_ASAP7_75t_L g1218 ( 
.A(n_1208),
.B(n_84),
.C(n_85),
.Y(n_1218)
);

AOI22xp33_ASAP7_75t_L g1219 ( 
.A1(n_1205),
.A2(n_86),
.B1(n_87),
.B2(n_88),
.Y(n_1219)
);

AOI211xp5_ASAP7_75t_L g1220 ( 
.A1(n_1207),
.A2(n_90),
.B(n_91),
.C(n_92),
.Y(n_1220)
);

OAI322xp33_ASAP7_75t_L g1221 ( 
.A1(n_1213),
.A2(n_1211),
.A3(n_1209),
.B1(n_1214),
.B2(n_1210),
.C1(n_1203),
.C2(n_106),
.Y(n_1221)
);

OAI22xp5_ASAP7_75t_L g1222 ( 
.A1(n_1204),
.A2(n_93),
.B1(n_95),
.B2(n_101),
.Y(n_1222)
);

AOI211xp5_ASAP7_75t_L g1223 ( 
.A1(n_1204),
.A2(n_102),
.B(n_104),
.C(n_108),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1217),
.B(n_115),
.Y(n_1224)
);

AOI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1223),
.A2(n_1010),
.B(n_118),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1220),
.A2(n_116),
.B(n_121),
.Y(n_1226)
);

AOI221x1_ASAP7_75t_L g1227 ( 
.A1(n_1218),
.A2(n_123),
.B1(n_124),
.B2(n_125),
.C(n_126),
.Y(n_1227)
);

NOR2xp67_ASAP7_75t_L g1228 ( 
.A(n_1219),
.B(n_127),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1216),
.B(n_128),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1215),
.A2(n_129),
.B(n_131),
.Y(n_1230)
);

OAI22xp5_ASAP7_75t_L g1231 ( 
.A1(n_1221),
.A2(n_1019),
.B1(n_134),
.B2(n_136),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1228),
.B(n_1222),
.Y(n_1232)
);

OA22x2_ASAP7_75t_L g1233 ( 
.A1(n_1224),
.A2(n_133),
.B1(n_139),
.B2(n_141),
.Y(n_1233)
);

OAI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1226),
.A2(n_1229),
.B(n_1227),
.Y(n_1234)
);

OAI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1232),
.A2(n_1230),
.B(n_1225),
.Y(n_1235)
);

AOI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1235),
.A2(n_1234),
.B(n_1233),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1236),
.Y(n_1237)
);

AND2x2_ASAP7_75t_SL g1238 ( 
.A(n_1237),
.B(n_1231),
.Y(n_1238)
);

AO21x2_ASAP7_75t_L g1239 ( 
.A1(n_1238),
.A2(n_142),
.B(n_144),
.Y(n_1239)
);

OAI221xp5_ASAP7_75t_R g1240 ( 
.A1(n_1239),
.A2(n_145),
.B1(n_146),
.B2(n_147),
.C(n_148),
.Y(n_1240)
);

AND4x1_ASAP7_75t_L g1241 ( 
.A(n_1240),
.B(n_150),
.C(n_151),
.D(n_152),
.Y(n_1241)
);

AOI22xp5_ASAP7_75t_L g1242 ( 
.A1(n_1241),
.A2(n_670),
.B1(n_1020),
.B2(n_156),
.Y(n_1242)
);

AOI211xp5_ASAP7_75t_L g1243 ( 
.A1(n_1242),
.A2(n_1022),
.B(n_154),
.C(n_159),
.Y(n_1243)
);

AOI211xp5_ASAP7_75t_L g1244 ( 
.A1(n_1243),
.A2(n_153),
.B(n_162),
.C(n_165),
.Y(n_1244)
);


endmodule