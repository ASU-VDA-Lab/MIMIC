module fake_jpeg_17224_n_82 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_82);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_82;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

INVx1_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

BUFx5_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

CKINVDCx16_ASAP7_75t_R g13 ( 
.A(n_0),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_10),
.B(n_14),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_20),
.B(n_21),
.Y(n_29)
);

OR2x2_ASAP7_75t_L g21 ( 
.A(n_13),
.B(n_0),
.Y(n_21)
);

NAND3xp33_ASAP7_75t_L g22 ( 
.A(n_14),
.B(n_1),
.C(n_2),
.Y(n_22)
);

NOR3xp33_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_13),
.C(n_10),
.Y(n_27)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_26),
.Y(n_28)
);

OR2x2_ASAP7_75t_L g43 ( 
.A(n_27),
.B(n_31),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_25),
.A2(n_19),
.B1(n_1),
.B2(n_11),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_21),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_SL g31 ( 
.A1(n_20),
.A2(n_19),
.B(n_11),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_21),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_42),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_36),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_16),
.Y(n_37)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_39),
.Y(n_48)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_32),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_41),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_22),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_28),
.B(n_16),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_15),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_18),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_26),
.C(n_12),
.Y(n_49)
);

XOR2xp5_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_53),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_50),
.B(n_51),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_12),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_43),
.Y(n_52)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_52),
.Y(n_57)
);

BUFx12f_ASAP7_75t_SL g55 ( 
.A(n_51),
.Y(n_55)
);

NAND3xp33_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_53),
.C(n_49),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_58),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_46),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_43),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_60),
.B(n_47),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_45),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_61),
.B(n_15),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_62),
.B(n_65),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_64),
.A2(n_67),
.B(n_5),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_57),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_66),
.Y(n_70)
);

NOR3xp33_ASAP7_75t_L g67 ( 
.A(n_60),
.B(n_15),
.C(n_6),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_63),
.A2(n_55),
.B1(n_54),
.B2(n_59),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_68),
.A2(n_69),
.B1(n_59),
.B2(n_70),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_71),
.B(n_7),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_72),
.B(n_26),
.C(n_8),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_69),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_73),
.B(n_74),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g75 ( 
.A(n_72),
.B(n_62),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_75),
.B(n_76),
.C(n_17),
.Y(n_79)
);

AOI21xp33_ASAP7_75t_L g78 ( 
.A1(n_75),
.A2(n_7),
.B(n_9),
.Y(n_78)
);

AOI322xp5_ASAP7_75t_L g80 ( 
.A1(n_78),
.A2(n_79),
.A3(n_77),
.B1(n_18),
.B2(n_24),
.C1(n_23),
.C2(n_34),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_80),
.B(n_23),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_81),
.B(n_24),
.Y(n_82)
);


endmodule