module fake_netlist_6_3096_n_1174 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_235, n_256, n_298, n_18, n_21, n_193, n_147, n_269, n_258, n_281, n_154, n_191, n_88, n_3, n_209, n_98, n_277, n_260, n_265, n_283, n_113, n_39, n_63, n_223, n_278, n_270, n_73, n_279, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_226, n_228, n_252, n_266, n_296, n_166, n_28, n_184, n_212, n_268, n_271, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_299, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_297, n_178, n_247, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_227, n_132, n_188, n_102, n_186, n_204, n_245, n_0, n_87, n_195, n_285, n_261, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_257, n_100, n_292, n_129, n_13, n_121, n_294, n_197, n_11, n_137, n_17, n_23, n_203, n_254, n_142, n_286, n_20, n_143, n_207, n_2, n_242, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_291, n_75, n_109, n_150, n_233, n_263, n_122, n_264, n_45, n_255, n_284, n_205, n_34, n_140, n_218, n_70, n_120, n_234, n_251, n_301, n_214, n_274, n_37, n_15, n_67, n_33, n_82, n_27, n_236, n_246, n_38, n_110, n_151, n_289, n_61, n_112, n_172, n_237, n_81, n_59, n_244, n_181, n_76, n_36, n_182, n_26, n_124, n_238, n_239, n_55, n_126, n_202, n_94, n_97, n_108, n_267, n_282, n_58, n_116, n_280, n_211, n_287, n_64, n_220, n_288, n_290, n_117, n_118, n_175, n_224, n_48, n_231, n_65, n_230, n_25, n_40, n_93, n_80, n_141, n_240, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_259, n_177, n_176, n_273, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_243, n_9, n_248, n_300, n_107, n_10, n_295, n_71, n_74, n_229, n_253, n_6, n_190, n_14, n_123, n_262, n_136, n_72, n_187, n_89, n_249, n_173, n_201, n_250, n_103, n_111, n_60, n_159, n_272, n_157, n_162, n_170, n_185, n_35, n_183, n_232, n_115, n_12, n_69, n_128, n_241, n_30, n_79, n_275, n_43, n_194, n_171, n_293, n_31, n_192, n_57, n_169, n_53, n_276, n_51, n_44, n_56, n_221, n_1174);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_235;
input n_256;
input n_298;
input n_18;
input n_21;
input n_193;
input n_147;
input n_269;
input n_258;
input n_281;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_277;
input n_260;
input n_265;
input n_283;
input n_113;
input n_39;
input n_63;
input n_223;
input n_278;
input n_270;
input n_73;
input n_279;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_226;
input n_228;
input n_252;
input n_266;
input n_296;
input n_166;
input n_28;
input n_184;
input n_212;
input n_268;
input n_271;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_299;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_297;
input n_178;
input n_247;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_227;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_245;
input n_0;
input n_87;
input n_195;
input n_285;
input n_261;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_257;
input n_100;
input n_292;
input n_129;
input n_13;
input n_121;
input n_294;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_254;
input n_142;
input n_286;
input n_20;
input n_143;
input n_207;
input n_2;
input n_242;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_291;
input n_75;
input n_109;
input n_150;
input n_233;
input n_263;
input n_122;
input n_264;
input n_45;
input n_255;
input n_284;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_234;
input n_251;
input n_301;
input n_214;
input n_274;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_236;
input n_246;
input n_38;
input n_110;
input n_151;
input n_289;
input n_61;
input n_112;
input n_172;
input n_237;
input n_81;
input n_59;
input n_244;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_238;
input n_239;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_267;
input n_282;
input n_58;
input n_116;
input n_280;
input n_211;
input n_287;
input n_64;
input n_220;
input n_288;
input n_290;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_231;
input n_65;
input n_230;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_240;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_259;
input n_177;
input n_176;
input n_273;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_243;
input n_9;
input n_248;
input n_300;
input n_107;
input n_10;
input n_295;
input n_71;
input n_74;
input n_229;
input n_253;
input n_6;
input n_190;
input n_14;
input n_123;
input n_262;
input n_136;
input n_72;
input n_187;
input n_89;
input n_249;
input n_173;
input n_201;
input n_250;
input n_103;
input n_111;
input n_60;
input n_159;
input n_272;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_232;
input n_115;
input n_12;
input n_69;
input n_128;
input n_241;
input n_30;
input n_79;
input n_275;
input n_43;
input n_194;
input n_171;
input n_293;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_276;
input n_51;
input n_44;
input n_56;
input n_221;

output n_1174;

wire n_992;
wire n_591;
wire n_435;
wire n_1115;
wire n_793;
wire n_326;
wire n_801;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_881;
wire n_875;
wire n_465;
wire n_367;
wire n_760;
wire n_680;
wire n_741;
wire n_1008;
wire n_1027;
wire n_590;
wire n_625;
wire n_661;
wire n_1079;
wire n_341;
wire n_362;
wire n_828;
wire n_462;
wire n_1033;
wire n_607;
wire n_671;
wire n_726;
wire n_1052;
wire n_316;
wire n_419;
wire n_304;
wire n_700;
wire n_694;
wire n_1103;
wire n_933;
wire n_740;
wire n_1038;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_1061;
wire n_384;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_1044;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_1164;
wire n_310;
wire n_509;
wire n_368;
wire n_575;
wire n_994;
wire n_1072;
wire n_677;
wire n_969;
wire n_988;
wire n_805;
wire n_1151;
wire n_396;
wire n_495;
wire n_1065;
wire n_815;
wire n_350;
wire n_1100;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_1128;
wire n_382;
wire n_673;
wire n_1020;
wire n_1009;
wire n_1042;
wire n_1071;
wire n_628;
wire n_1067;
wire n_1160;
wire n_883;
wire n_557;
wire n_823;
wire n_1132;
wire n_349;
wire n_643;
wire n_898;
wire n_617;
wire n_698;
wire n_1074;
wire n_1032;
wire n_845;
wire n_807;
wire n_1036;
wire n_739;
wire n_400;
wire n_337;
wire n_955;
wire n_865;
wire n_1138;
wire n_893;
wire n_925;
wire n_485;
wire n_1101;
wire n_1026;
wire n_443;
wire n_1099;
wire n_892;
wire n_768;
wire n_1097;
wire n_471;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_1130;
wire n_1127;
wire n_1095;
wire n_573;
wire n_769;
wire n_320;
wire n_639;
wire n_963;
wire n_676;
wire n_327;
wire n_794;
wire n_727;
wire n_894;
wire n_369;
wire n_1120;
wire n_597;
wire n_685;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_447;
wire n_872;
wire n_1139;
wire n_718;
wire n_517;
wire n_1018;
wire n_1172;
wire n_747;
wire n_852;
wire n_667;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_1105;
wire n_621;
wire n_305;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_691;
wire n_535;
wire n_544;
wire n_372;
wire n_468;
wire n_901;
wire n_1078;
wire n_504;
wire n_923;
wire n_314;
wire n_1140;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1057;
wire n_1147;
wire n_360;
wire n_945;
wire n_977;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_1143;
wire n_536;
wire n_895;
wire n_1126;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_1108;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_1119;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_631;
wire n_516;
wire n_720;
wire n_758;
wire n_525;
wire n_842;
wire n_1163;
wire n_1173;
wire n_1116;
wire n_611;
wire n_943;
wire n_1168;
wire n_491;
wire n_878;
wire n_656;
wire n_843;
wire n_989;
wire n_772;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_538;
wire n_1035;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_844;
wire n_343;
wire n_886;
wire n_448;
wire n_953;
wire n_1017;
wire n_1004;
wire n_1094;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_1083;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_1112;
wire n_454;
wire n_638;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_653;
wire n_887;
wire n_1117;
wire n_1087;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_1049;
wire n_576;
wire n_1028;
wire n_472;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_809;
wire n_1043;
wire n_1011;
wire n_926;
wire n_927;
wire n_986;
wire n_839;
wire n_734;
wire n_1088;
wire n_708;
wire n_919;
wire n_1081;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_779;
wire n_800;
wire n_929;
wire n_460;
wire n_1084;
wire n_1171;
wire n_1104;
wire n_907;
wire n_854;
wire n_1058;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_1122;
wire n_374;
wire n_659;
wire n_709;
wire n_904;
wire n_366;
wire n_870;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_526;
wire n_1109;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_1148;
wire n_1054;
wire n_334;
wire n_559;
wire n_370;
wire n_1161;
wire n_458;
wire n_1070;
wire n_1085;
wire n_650;
wire n_998;
wire n_1046;
wire n_717;
wire n_1145;
wire n_330;
wire n_771;
wire n_1121;
wire n_1152;
wire n_470;
wire n_475;
wire n_924;
wire n_1102;
wire n_492;
wire n_972;
wire n_551;
wire n_699;
wire n_456;
wire n_1149;
wire n_564;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_1073;
wire n_1000;
wire n_686;
wire n_796;
wire n_1041;
wire n_757;
wire n_594;
wire n_565;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_1062;
wire n_619;
wire n_885;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_1090;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_1156;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_1142;
wire n_503;
wire n_716;
wire n_623;
wire n_1048;
wire n_1123;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_868;
wire n_731;
wire n_859;
wire n_570;
wire n_406;
wire n_483;
wire n_735;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_307;
wire n_469;
wire n_1137;
wire n_433;
wire n_500;
wire n_942;
wire n_880;
wire n_981;
wire n_476;
wire n_792;
wire n_714;
wire n_543;
wire n_1144;
wire n_889;
wire n_357;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_1162;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_1068;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_982;
wire n_964;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_1075;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_584;
wire n_1110;
wire n_399;
wire n_979;
wire n_548;
wire n_905;
wire n_436;
wire n_833;
wire n_523;
wire n_707;
wire n_322;
wire n_993;
wire n_345;
wire n_409;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_1155;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_558;
wire n_810;
wire n_1133;
wire n_635;
wire n_787;
wire n_311;
wire n_1064;
wire n_403;
wire n_1080;
wire n_723;
wire n_1051;
wire n_634;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_1146;
wire n_1141;
wire n_386;
wire n_764;
wire n_1039;
wire n_556;
wire n_1034;
wire n_1086;
wire n_1066;
wire n_692;
wire n_733;
wire n_1158;
wire n_754;
wire n_1136;
wire n_941;
wire n_975;
wire n_1031;
wire n_487;
wire n_550;
wire n_1125;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_1107;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_1159;
wire n_569;
wire n_1092;
wire n_441;
wire n_882;
wire n_811;
wire n_1060;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_1111;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_1053;
wire n_530;
wire n_520;
wire n_1029;
wire n_418;
wire n_1093;
wire n_618;
wire n_1055;
wire n_790;
wire n_1106;
wire n_582;
wire n_1167;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_404;
wire n_651;
wire n_439;
wire n_1153;
wire n_518;
wire n_679;
wire n_1069;
wire n_453;
wire n_612;
wire n_633;
wire n_1170;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1047;
wire n_1010;
wire n_355;
wire n_1165;
wire n_426;
wire n_317;
wire n_1040;
wire n_915;
wire n_632;
wire n_702;
wire n_1166;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_1131;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_920;
wire n_730;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_670;
wire n_834;
wire n_928;
wire n_835;
wire n_690;
wire n_850;
wire n_1089;
wire n_1135;
wire n_1169;
wire n_401;
wire n_324;
wire n_743;
wire n_816;
wire n_766;
wire n_1157;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_604;
wire n_848;
wire n_1019;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_1096;
wire n_1063;
wire n_729;
wire n_1091;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_438;
wire n_1124;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_515;
wire n_983;
wire n_427;
wire n_1059;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_1077;
wire n_961;
wire n_862;
wire n_869;
wire n_351;
wire n_437;
wire n_1082;
wire n_1154;
wire n_1113;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_1098;
wire n_697;
wire n_687;
wire n_364;
wire n_890;
wire n_637;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_484;
wire n_613;
wire n_736;
wire n_897;
wire n_900;
wire n_846;
wire n_501;
wire n_956;
wire n_841;
wire n_960;
wire n_531;
wire n_827;
wire n_1001;
wire n_361;
wire n_508;
wire n_663;
wire n_856;
wire n_1050;
wire n_379;
wire n_778;
wire n_1025;
wire n_1134;
wire n_332;
wire n_891;
wire n_336;
wire n_1150;
wire n_410;
wire n_398;
wire n_1129;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_664;
wire n_949;
wire n_678;
wire n_1007;
wire n_649;

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_277),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_16),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_173),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_136),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_78),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_123),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_204),
.Y(n_308)
);

BUFx3_ASAP7_75t_L g309 ( 
.A(n_20),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_167),
.Y(n_310)
);

INVx1_ASAP7_75t_SL g311 ( 
.A(n_29),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_60),
.Y(n_312)
);

BUFx3_ASAP7_75t_L g313 ( 
.A(n_13),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_10),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_35),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_255),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_181),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_129),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_26),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_73),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_125),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_205),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_290),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_139),
.Y(n_324)
);

BUFx10_ASAP7_75t_L g325 ( 
.A(n_234),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_111),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_94),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_53),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_212),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_145),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_287),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_135),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_177),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_27),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_288),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_113),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_301),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_201),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_251),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_10),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_146),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_295),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_175),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_95),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_68),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_99),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_160),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_46),
.Y(n_348)
);

BUFx5_ASAP7_75t_L g349 ( 
.A(n_223),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_198),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_231),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_278),
.Y(n_352)
);

INVx1_ASAP7_75t_SL g353 ( 
.A(n_32),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_81),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_259),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_196),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_153),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_104),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_11),
.Y(n_359)
);

BUFx2_ASAP7_75t_L g360 ( 
.A(n_276),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_239),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_202),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_130),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_245),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_216),
.Y(n_365)
);

CKINVDCx14_ASAP7_75t_R g366 ( 
.A(n_106),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_291),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_211),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_241),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_103),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_191),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_89),
.Y(n_372)
);

BUFx2_ASAP7_75t_L g373 ( 
.A(n_17),
.Y(n_373)
);

BUFx3_ASAP7_75t_L g374 ( 
.A(n_186),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_266),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_215),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g377 ( 
.A(n_187),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_300),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_154),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_8),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_230),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_206),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_262),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_76),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_183),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_268),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_272),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_269),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_69),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_298),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_87),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_264),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_178),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_42),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_34),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_101),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_263),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_199),
.Y(n_398)
);

INVx2_ASAP7_75t_SL g399 ( 
.A(n_40),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_296),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_220),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_214),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_270),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_240),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_292),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_67),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_284),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_261),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_275),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_116),
.Y(n_410)
);

CKINVDCx14_ASAP7_75t_R g411 ( 
.A(n_274),
.Y(n_411)
);

BUFx3_ASAP7_75t_L g412 ( 
.A(n_51),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_289),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_297),
.Y(n_414)
);

INVxp67_ASAP7_75t_L g415 ( 
.A(n_57),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_19),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_27),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_294),
.Y(n_418)
);

BUFx10_ASAP7_75t_L g419 ( 
.A(n_128),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_279),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g421 ( 
.A(n_260),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_28),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_258),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_127),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_70),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_6),
.Y(n_426)
);

BUFx2_ASAP7_75t_SL g427 ( 
.A(n_7),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_184),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_5),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_33),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_31),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_242),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_120),
.Y(n_433)
);

BUFx5_ASAP7_75t_L g434 ( 
.A(n_16),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_133),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_150),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_32),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_63),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_98),
.Y(n_439)
);

BUFx3_ASAP7_75t_L g440 ( 
.A(n_72),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_85),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_18),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_203),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_140),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_58),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_96),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_155),
.Y(n_447)
);

HB1xp67_ASAP7_75t_L g448 ( 
.A(n_256),
.Y(n_448)
);

CKINVDCx16_ASAP7_75t_R g449 ( 
.A(n_197),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_267),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_143),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_189),
.Y(n_452)
);

BUFx3_ASAP7_75t_L g453 ( 
.A(n_282),
.Y(n_453)
);

BUFx3_ASAP7_75t_L g454 ( 
.A(n_185),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_97),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_84),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_163),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_2),
.Y(n_458)
);

INVx2_ASAP7_75t_SL g459 ( 
.A(n_281),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_23),
.Y(n_460)
);

INVx1_ASAP7_75t_SL g461 ( 
.A(n_52),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_176),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_192),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_29),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_280),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_115),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_221),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_218),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_285),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_194),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_252),
.Y(n_471)
);

BUFx5_ASAP7_75t_L g472 ( 
.A(n_157),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_293),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_151),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_148),
.Y(n_475)
);

INVx3_ASAP7_75t_L g476 ( 
.A(n_132),
.Y(n_476)
);

INVx1_ASAP7_75t_SL g477 ( 
.A(n_208),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_19),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_14),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_92),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_265),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_118),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_168),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_182),
.Y(n_484)
);

BUFx8_ASAP7_75t_SL g485 ( 
.A(n_74),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_273),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_271),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_105),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_54),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_377),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_434),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_373),
.B(n_0),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_360),
.B(n_0),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_309),
.B(n_1),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_313),
.B(n_1),
.Y(n_495)
);

AND2x4_ASAP7_75t_L g496 ( 
.A(n_374),
.B(n_412),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_434),
.Y(n_497)
);

BUFx3_ASAP7_75t_L g498 ( 
.A(n_325),
.Y(n_498)
);

INVx5_ASAP7_75t_L g499 ( 
.A(n_377),
.Y(n_499)
);

AND2x4_ASAP7_75t_L g500 ( 
.A(n_440),
.B(n_453),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_476),
.B(n_399),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_377),
.Y(n_502)
);

BUFx12f_ASAP7_75t_L g503 ( 
.A(n_325),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_434),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_485),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_366),
.B(n_2),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g507 ( 
.A(n_377),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_454),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_448),
.B(n_3),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_434),
.Y(n_510)
);

INVx5_ASAP7_75t_L g511 ( 
.A(n_476),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_372),
.Y(n_512)
);

AND2x4_ASAP7_75t_L g513 ( 
.A(n_459),
.B(n_3),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_434),
.Y(n_514)
);

INVx3_ASAP7_75t_L g515 ( 
.A(n_340),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_411),
.B(n_302),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_434),
.B(n_4),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_349),
.Y(n_518)
);

BUFx3_ASAP7_75t_L g519 ( 
.A(n_419),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_484),
.B(n_4),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_306),
.B(n_5),
.Y(n_521)
);

AND2x4_ASAP7_75t_L g522 ( 
.A(n_305),
.B(n_6),
.Y(n_522)
);

AND2x4_ASAP7_75t_L g523 ( 
.A(n_308),
.B(n_7),
.Y(n_523)
);

INVx5_ASAP7_75t_L g524 ( 
.A(n_419),
.Y(n_524)
);

AND2x4_ASAP7_75t_L g525 ( 
.A(n_310),
.B(n_8),
.Y(n_525)
);

AND2x6_ASAP7_75t_L g526 ( 
.A(n_316),
.B(n_318),
.Y(n_526)
);

BUFx12f_ASAP7_75t_L g527 ( 
.A(n_314),
.Y(n_527)
);

AND2x4_ASAP7_75t_L g528 ( 
.A(n_321),
.B(n_9),
.Y(n_528)
);

HB1xp67_ASAP7_75t_L g529 ( 
.A(n_319),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_426),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_449),
.B(n_9),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_304),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g533 ( 
.A(n_328),
.Y(n_533)
);

BUFx6f_ASAP7_75t_L g534 ( 
.A(n_329),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_338),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_341),
.Y(n_536)
);

AND2x4_ASAP7_75t_L g537 ( 
.A(n_345),
.B(n_11),
.Y(n_537)
);

BUFx6f_ASAP7_75t_L g538 ( 
.A(n_347),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_334),
.B(n_12),
.Y(n_539)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_303),
.Y(n_540)
);

BUFx3_ASAP7_75t_L g541 ( 
.A(n_307),
.Y(n_541)
);

INVx4_ASAP7_75t_L g542 ( 
.A(n_317),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_349),
.Y(n_543)
);

BUFx12f_ASAP7_75t_L g544 ( 
.A(n_359),
.Y(n_544)
);

BUFx6f_ASAP7_75t_L g545 ( 
.A(n_350),
.Y(n_545)
);

BUFx8_ASAP7_75t_L g546 ( 
.A(n_315),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_320),
.Y(n_547)
);

BUFx6f_ASAP7_75t_L g548 ( 
.A(n_354),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_430),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_349),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_323),
.B(n_12),
.Y(n_551)
);

BUFx6f_ASAP7_75t_L g552 ( 
.A(n_355),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_479),
.Y(n_553)
);

HB1xp67_ASAP7_75t_L g554 ( 
.A(n_380),
.Y(n_554)
);

AND2x6_ASAP7_75t_L g555 ( 
.A(n_357),
.B(n_37),
.Y(n_555)
);

INVx5_ASAP7_75t_L g556 ( 
.A(n_349),
.Y(n_556)
);

INVx4_ASAP7_75t_L g557 ( 
.A(n_322),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_323),
.B(n_13),
.Y(n_558)
);

AND2x4_ASAP7_75t_L g559 ( 
.A(n_358),
.B(n_14),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_361),
.Y(n_560)
);

INVxp67_ASAP7_75t_L g561 ( 
.A(n_427),
.Y(n_561)
);

HB1xp67_ASAP7_75t_L g562 ( 
.A(n_395),
.Y(n_562)
);

INVx3_ASAP7_75t_L g563 ( 
.A(n_416),
.Y(n_563)
);

AND2x4_ASAP7_75t_L g564 ( 
.A(n_363),
.B(n_15),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_349),
.Y(n_565)
);

INVx2_ASAP7_75t_SL g566 ( 
.A(n_417),
.Y(n_566)
);

AND2x2_ASAP7_75t_L g567 ( 
.A(n_311),
.B(n_15),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_349),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_353),
.B(n_429),
.Y(n_569)
);

BUFx6f_ASAP7_75t_L g570 ( 
.A(n_371),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_375),
.Y(n_571)
);

AND2x4_ASAP7_75t_L g572 ( 
.A(n_388),
.B(n_17),
.Y(n_572)
);

BUFx6f_ASAP7_75t_L g573 ( 
.A(n_391),
.Y(n_573)
);

HB1xp67_ASAP7_75t_L g574 ( 
.A(n_431),
.Y(n_574)
);

AND2x4_ASAP7_75t_L g575 ( 
.A(n_396),
.B(n_401),
.Y(n_575)
);

INVx2_ASAP7_75t_SL g576 ( 
.A(n_458),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_356),
.B(n_18),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_SL g578 ( 
.A(n_356),
.B(n_20),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_415),
.B(n_21),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_403),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_415),
.B(n_21),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_SL g582 ( 
.A(n_421),
.B(n_22),
.Y(n_582)
);

AND2x4_ASAP7_75t_L g583 ( 
.A(n_404),
.B(n_22),
.Y(n_583)
);

AND2x4_ASAP7_75t_L g584 ( 
.A(n_406),
.B(n_23),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_472),
.Y(n_585)
);

BUFx6f_ASAP7_75t_L g586 ( 
.A(n_407),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_421),
.B(n_24),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_472),
.B(n_24),
.Y(n_588)
);

HB1xp67_ASAP7_75t_L g589 ( 
.A(n_460),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_472),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_472),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_472),
.B(n_25),
.Y(n_592)
);

INVx5_ASAP7_75t_L g593 ( 
.A(n_472),
.Y(n_593)
);

AO22x2_ASAP7_75t_L g594 ( 
.A1(n_492),
.A2(n_410),
.B1(n_414),
.B2(n_408),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_516),
.B(n_461),
.Y(n_595)
);

AO22x2_ASAP7_75t_L g596 ( 
.A1(n_513),
.A2(n_423),
.B1(n_425),
.B2(n_420),
.Y(n_596)
);

AOI22xp5_ASAP7_75t_L g597 ( 
.A1(n_521),
.A2(n_327),
.B1(n_344),
.B2(n_312),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_542),
.B(n_477),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_532),
.B(n_433),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_490),
.Y(n_600)
);

OAI22xp33_ASAP7_75t_L g601 ( 
.A1(n_578),
.A2(n_478),
.B1(n_437),
.B2(n_442),
.Y(n_601)
);

INVx8_ASAP7_75t_L g602 ( 
.A(n_505),
.Y(n_602)
);

AO22x2_ASAP7_75t_L g603 ( 
.A1(n_513),
.A2(n_531),
.B1(n_522),
.B2(n_525),
.Y(n_603)
);

AOI22xp5_ASAP7_75t_L g604 ( 
.A1(n_506),
.A2(n_368),
.B1(n_397),
.B2(n_364),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_571),
.Y(n_605)
);

AOI22xp5_ASAP7_75t_L g606 ( 
.A1(n_493),
.A2(n_457),
.B1(n_480),
.B2(n_418),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_547),
.B(n_438),
.Y(n_607)
);

AOI22xp5_ASAP7_75t_L g608 ( 
.A1(n_509),
.A2(n_464),
.B1(n_422),
.B2(n_326),
.Y(n_608)
);

AO22x2_ASAP7_75t_L g609 ( 
.A1(n_522),
.A2(n_445),
.B1(n_451),
.B2(n_439),
.Y(n_609)
);

AOI22xp5_ASAP7_75t_L g610 ( 
.A1(n_582),
.A2(n_330),
.B1(n_331),
.B2(n_324),
.Y(n_610)
);

OAI22xp5_ASAP7_75t_SL g611 ( 
.A1(n_587),
.A2(n_455),
.B1(n_456),
.B2(n_487),
.Y(n_611)
);

OAI22xp33_ASAP7_75t_SL g612 ( 
.A1(n_579),
.A2(n_462),
.B1(n_463),
.B2(n_466),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_580),
.Y(n_613)
);

OR2x6_ASAP7_75t_L g614 ( 
.A(n_527),
.B(n_544),
.Y(n_614)
);

AOI22xp5_ASAP7_75t_L g615 ( 
.A1(n_569),
.A2(n_398),
.B1(n_488),
.B2(n_486),
.Y(n_615)
);

OR2x2_ASAP7_75t_L g616 ( 
.A(n_529),
.B(n_25),
.Y(n_616)
);

AOI22xp5_ASAP7_75t_L g617 ( 
.A1(n_567),
.A2(n_393),
.B1(n_333),
.B2(n_482),
.Y(n_617)
);

OAI22xp33_ASAP7_75t_SL g618 ( 
.A1(n_551),
.A2(n_467),
.B1(n_483),
.B2(n_469),
.Y(n_618)
);

AO22x2_ASAP7_75t_L g619 ( 
.A1(n_523),
.A2(n_471),
.B1(n_473),
.B2(n_475),
.Y(n_619)
);

INVx1_ASAP7_75t_SL g620 ( 
.A(n_524),
.Y(n_620)
);

AO22x2_ASAP7_75t_L g621 ( 
.A1(n_523),
.A2(n_26),
.B1(n_28),
.B2(n_30),
.Y(n_621)
);

INVx3_ASAP7_75t_L g622 ( 
.A(n_508),
.Y(n_622)
);

OAI22xp5_ASAP7_75t_L g623 ( 
.A1(n_558),
.A2(n_489),
.B1(n_481),
.B2(n_474),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_490),
.Y(n_624)
);

BUFx2_ASAP7_75t_L g625 ( 
.A(n_498),
.Y(n_625)
);

AOI22xp5_ASAP7_75t_L g626 ( 
.A1(n_554),
.A2(n_386),
.B1(n_468),
.B2(n_465),
.Y(n_626)
);

OA22x2_ASAP7_75t_L g627 ( 
.A1(n_562),
.A2(n_470),
.B1(n_452),
.B2(n_450),
.Y(n_627)
);

AOI22xp5_ASAP7_75t_L g628 ( 
.A1(n_574),
.A2(n_383),
.B1(n_446),
.B2(n_444),
.Y(n_628)
);

AOI22xp5_ASAP7_75t_L g629 ( 
.A1(n_589),
.A2(n_576),
.B1(n_566),
.B2(n_539),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_490),
.Y(n_630)
);

AO22x2_ASAP7_75t_L g631 ( 
.A1(n_525),
.A2(n_30),
.B1(n_31),
.B2(n_33),
.Y(n_631)
);

OR2x2_ASAP7_75t_L g632 ( 
.A(n_561),
.B(n_34),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_502),
.Y(n_633)
);

OAI22xp33_ASAP7_75t_SL g634 ( 
.A1(n_577),
.A2(n_447),
.B1(n_443),
.B2(n_441),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_563),
.B(n_332),
.Y(n_635)
);

AO22x2_ASAP7_75t_L g636 ( 
.A1(n_528),
.A2(n_35),
.B1(n_36),
.B2(n_436),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_563),
.B(n_335),
.Y(n_637)
);

AO22x2_ASAP7_75t_L g638 ( 
.A1(n_528),
.A2(n_36),
.B1(n_435),
.B2(n_432),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_524),
.B(n_336),
.Y(n_639)
);

AND2x2_ASAP7_75t_SL g640 ( 
.A(n_494),
.B(n_337),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_512),
.Y(n_641)
);

AND2x2_ASAP7_75t_L g642 ( 
.A(n_524),
.B(n_496),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_512),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_496),
.B(n_339),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_542),
.B(n_342),
.Y(n_645)
);

OAI22xp33_ASAP7_75t_SL g646 ( 
.A1(n_581),
.A2(n_428),
.B1(n_424),
.B2(n_413),
.Y(n_646)
);

OAI22xp33_ASAP7_75t_SL g647 ( 
.A1(n_501),
.A2(n_592),
.B1(n_588),
.B2(n_517),
.Y(n_647)
);

XNOR2xp5_ASAP7_75t_L g648 ( 
.A(n_495),
.B(n_343),
.Y(n_648)
);

OAI22xp5_ASAP7_75t_SL g649 ( 
.A1(n_519),
.A2(n_409),
.B1(n_405),
.B2(n_402),
.Y(n_649)
);

AO22x2_ASAP7_75t_L g650 ( 
.A1(n_537),
.A2(n_400),
.B1(n_394),
.B2(n_392),
.Y(n_650)
);

OAI22xp33_ASAP7_75t_L g651 ( 
.A1(n_520),
.A2(n_390),
.B1(n_389),
.B2(n_387),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_500),
.B(n_541),
.Y(n_652)
);

AOI22xp5_ASAP7_75t_L g653 ( 
.A1(n_503),
.A2(n_369),
.B1(n_384),
.B2(n_382),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_500),
.B(n_346),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_502),
.Y(n_655)
);

OAI22xp5_ASAP7_75t_SL g656 ( 
.A1(n_537),
.A2(n_385),
.B1(n_381),
.B2(n_379),
.Y(n_656)
);

OAI22xp5_ASAP7_75t_L g657 ( 
.A1(n_559),
.A2(n_378),
.B1(n_376),
.B2(n_370),
.Y(n_657)
);

OAI22xp5_ASAP7_75t_SL g658 ( 
.A1(n_559),
.A2(n_367),
.B1(n_365),
.B2(n_362),
.Y(n_658)
);

AOI22xp5_ASAP7_75t_L g659 ( 
.A1(n_564),
.A2(n_352),
.B1(n_351),
.B2(n_348),
.Y(n_659)
);

AO22x2_ASAP7_75t_L g660 ( 
.A1(n_564),
.A2(n_38),
.B1(n_39),
.B2(n_41),
.Y(n_660)
);

OAI22xp33_ASAP7_75t_SL g661 ( 
.A1(n_572),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_661)
);

INVx3_ASAP7_75t_L g662 ( 
.A(n_508),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_512),
.Y(n_663)
);

OA22x2_ASAP7_75t_L g664 ( 
.A1(n_549),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_502),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_507),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_508),
.Y(n_667)
);

OAI22xp5_ASAP7_75t_L g668 ( 
.A1(n_572),
.A2(n_50),
.B1(n_55),
.B2(n_56),
.Y(n_668)
);

OA22x2_ASAP7_75t_L g669 ( 
.A1(n_553),
.A2(n_59),
.B1(n_61),
.B2(n_62),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_507),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_557),
.B(n_64),
.Y(n_671)
);

INVx3_ASAP7_75t_L g672 ( 
.A(n_533),
.Y(n_672)
);

AO22x2_ASAP7_75t_L g673 ( 
.A1(n_583),
.A2(n_65),
.B1(n_66),
.B2(n_71),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_557),
.B(n_75),
.Y(n_674)
);

AND2x2_ASAP7_75t_SL g675 ( 
.A(n_583),
.B(n_77),
.Y(n_675)
);

INVxp67_ASAP7_75t_L g676 ( 
.A(n_595),
.Y(n_676)
);

AND2x4_ASAP7_75t_L g677 ( 
.A(n_652),
.B(n_575),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_605),
.Y(n_678)
);

BUFx3_ASAP7_75t_L g679 ( 
.A(n_622),
.Y(n_679)
);

XOR2xp5_ASAP7_75t_L g680 ( 
.A(n_606),
.B(n_79),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_599),
.B(n_575),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_613),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_641),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_643),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_663),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_607),
.B(n_584),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_600),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_624),
.Y(n_688)
);

CKINVDCx14_ASAP7_75t_R g689 ( 
.A(n_597),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_630),
.Y(n_690)
);

BUFx3_ASAP7_75t_L g691 ( 
.A(n_662),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_633),
.Y(n_692)
);

INVxp33_ASAP7_75t_SL g693 ( 
.A(n_648),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_640),
.B(n_598),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_655),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_665),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_635),
.B(n_533),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_666),
.Y(n_698)
);

HB1xp67_ASAP7_75t_L g699 ( 
.A(n_642),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_670),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_647),
.B(n_491),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_672),
.Y(n_702)
);

INVx2_ASAP7_75t_SL g703 ( 
.A(n_639),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_667),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_602),
.Y(n_705)
);

BUFx2_ASAP7_75t_R g706 ( 
.A(n_625),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_615),
.B(n_584),
.Y(n_707)
);

OAI21xp5_ASAP7_75t_L g708 ( 
.A1(n_669),
.A2(n_555),
.B(n_526),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_603),
.B(n_497),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_644),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_654),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_664),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_637),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_603),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_632),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_616),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_596),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_609),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_609),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_620),
.B(n_604),
.Y(n_720)
);

OR2x2_ASAP7_75t_L g721 ( 
.A(n_608),
.B(n_657),
.Y(n_721)
);

XNOR2x2_ASAP7_75t_L g722 ( 
.A(n_621),
.B(n_553),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_602),
.Y(n_723)
);

XOR2xp5_ASAP7_75t_L g724 ( 
.A(n_653),
.B(n_80),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_619),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_619),
.Y(n_726)
);

BUFx6f_ASAP7_75t_L g727 ( 
.A(n_675),
.Y(n_727)
);

AND2x2_ASAP7_75t_L g728 ( 
.A(n_626),
.B(n_511),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_610),
.B(n_560),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_671),
.B(n_504),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_596),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_668),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_594),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_594),
.Y(n_734)
);

INVx4_ASAP7_75t_L g735 ( 
.A(n_674),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_645),
.B(n_560),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_627),
.Y(n_737)
);

BUFx6f_ASAP7_75t_L g738 ( 
.A(n_614),
.Y(n_738)
);

INVxp67_ASAP7_75t_L g739 ( 
.A(n_649),
.Y(n_739)
);

INVx2_ASAP7_75t_SL g740 ( 
.A(n_650),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_628),
.B(n_511),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_617),
.B(n_659),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_621),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_612),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_611),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_660),
.Y(n_746)
);

AND2x2_ASAP7_75t_L g747 ( 
.A(n_629),
.B(n_511),
.Y(n_747)
);

INVx1_ASAP7_75t_SL g748 ( 
.A(n_636),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_660),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_673),
.Y(n_750)
);

XOR2xp5_ASAP7_75t_L g751 ( 
.A(n_634),
.B(n_82),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_673),
.Y(n_752)
);

AOI21xp5_ASAP7_75t_L g753 ( 
.A1(n_618),
.A2(n_514),
.B(n_510),
.Y(n_753)
);

XNOR2x2_ASAP7_75t_L g754 ( 
.A(n_631),
.B(n_530),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_661),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_631),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_636),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_651),
.B(n_510),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_656),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_658),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_650),
.Y(n_761)
);

XOR2x2_ASAP7_75t_L g762 ( 
.A(n_646),
.B(n_546),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_678),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_686),
.B(n_623),
.Y(n_764)
);

INVx2_ASAP7_75t_SL g765 ( 
.A(n_677),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_736),
.B(n_526),
.Y(n_766)
);

HB1xp67_ASAP7_75t_L g767 ( 
.A(n_676),
.Y(n_767)
);

AND2x2_ASAP7_75t_L g768 ( 
.A(n_676),
.B(n_638),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_692),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_713),
.B(n_638),
.Y(n_770)
);

OAI21xp5_ASAP7_75t_L g771 ( 
.A1(n_701),
.A2(n_555),
.B(n_526),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_697),
.B(n_526),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_697),
.B(n_555),
.Y(n_773)
);

AND2x4_ASAP7_75t_L g774 ( 
.A(n_714),
.B(n_555),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_700),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_681),
.B(n_533),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_682),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_712),
.B(n_540),
.Y(n_778)
);

AND2x2_ASAP7_75t_L g779 ( 
.A(n_677),
.B(n_540),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_701),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_730),
.B(n_534),
.Y(n_781)
);

INVx3_ASAP7_75t_L g782 ( 
.A(n_687),
.Y(n_782)
);

AND2x2_ASAP7_75t_L g783 ( 
.A(n_729),
.B(n_530),
.Y(n_783)
);

AND2x4_ASAP7_75t_L g784 ( 
.A(n_703),
.B(n_717),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_688),
.Y(n_785)
);

HB1xp67_ASAP7_75t_L g786 ( 
.A(n_699),
.Y(n_786)
);

BUFx4f_ASAP7_75t_L g787 ( 
.A(n_727),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_699),
.B(n_707),
.Y(n_788)
);

BUFx3_ASAP7_75t_L g789 ( 
.A(n_679),
.Y(n_789)
);

BUFx3_ASAP7_75t_L g790 ( 
.A(n_691),
.Y(n_790)
);

AND2x2_ASAP7_75t_L g791 ( 
.A(n_710),
.B(n_518),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_690),
.Y(n_792)
);

BUFx6f_ASAP7_75t_L g793 ( 
.A(n_709),
.Y(n_793)
);

AND2x4_ASAP7_75t_L g794 ( 
.A(n_711),
.B(n_83),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_727),
.B(n_708),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_695),
.Y(n_796)
);

AND2x2_ASAP7_75t_SL g797 ( 
.A(n_727),
.B(n_543),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_708),
.B(n_755),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_715),
.B(n_550),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_744),
.B(n_565),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_696),
.Y(n_801)
);

AND2x2_ASAP7_75t_L g802 ( 
.A(n_732),
.B(n_568),
.Y(n_802)
);

HB1xp67_ASAP7_75t_L g803 ( 
.A(n_737),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_716),
.B(n_614),
.Y(n_804)
);

INVx4_ASAP7_75t_L g805 ( 
.A(n_735),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_730),
.B(n_534),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_720),
.B(n_515),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_735),
.B(n_534),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_698),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_704),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_683),
.Y(n_811)
);

HB1xp67_ASAP7_75t_L g812 ( 
.A(n_731),
.Y(n_812)
);

INVx4_ASAP7_75t_L g813 ( 
.A(n_684),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_685),
.Y(n_814)
);

BUFx6f_ASAP7_75t_L g815 ( 
.A(n_709),
.Y(n_815)
);

AND2x2_ASAP7_75t_L g816 ( 
.A(n_758),
.B(n_585),
.Y(n_816)
);

OR2x2_ASAP7_75t_L g817 ( 
.A(n_721),
.B(n_601),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_758),
.B(n_590),
.Y(n_818)
);

OAI21xp5_ASAP7_75t_L g819 ( 
.A1(n_742),
.A2(n_591),
.B(n_499),
.Y(n_819)
);

BUFx8_ASAP7_75t_SL g820 ( 
.A(n_738),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_694),
.B(n_535),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_702),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_753),
.B(n_535),
.Y(n_823)
);

BUFx6f_ASAP7_75t_L g824 ( 
.A(n_718),
.Y(n_824)
);

BUFx6f_ASAP7_75t_L g825 ( 
.A(n_719),
.Y(n_825)
);

INVx3_ASAP7_75t_L g826 ( 
.A(n_725),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_728),
.B(n_535),
.Y(n_827)
);

AND2x2_ASAP7_75t_L g828 ( 
.A(n_741),
.B(n_536),
.Y(n_828)
);

BUFx6f_ASAP7_75t_L g829 ( 
.A(n_726),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_733),
.Y(n_830)
);

BUFx6f_ASAP7_75t_L g831 ( 
.A(n_734),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_753),
.B(n_536),
.Y(n_832)
);

AND2x4_ASAP7_75t_L g833 ( 
.A(n_740),
.B(n_743),
.Y(n_833)
);

INVxp33_ASAP7_75t_L g834 ( 
.A(n_747),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_756),
.Y(n_835)
);

AND2x6_ASAP7_75t_L g836 ( 
.A(n_746),
.B(n_749),
.Y(n_836)
);

BUFx3_ASAP7_75t_L g837 ( 
.A(n_705),
.Y(n_837)
);

OR2x2_ASAP7_75t_L g838 ( 
.A(n_748),
.B(n_515),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_757),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_750),
.B(n_536),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_752),
.B(n_538),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_722),
.Y(n_842)
);

NAND2x1_ASAP7_75t_SL g843 ( 
.A(n_788),
.B(n_759),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_826),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_780),
.B(n_745),
.Y(n_845)
);

BUFx6f_ASAP7_75t_L g846 ( 
.A(n_824),
.Y(n_846)
);

AND2x6_ASAP7_75t_L g847 ( 
.A(n_774),
.B(n_748),
.Y(n_847)
);

AND2x4_ASAP7_75t_L g848 ( 
.A(n_765),
.B(n_761),
.Y(n_848)
);

NOR2xp67_ASAP7_75t_L g849 ( 
.A(n_765),
.B(n_723),
.Y(n_849)
);

BUFx4f_ASAP7_75t_L g850 ( 
.A(n_793),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_807),
.B(n_689),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_803),
.Y(n_852)
);

OR2x2_ASAP7_75t_L g853 ( 
.A(n_817),
.B(n_760),
.Y(n_853)
);

OR2x6_ASAP7_75t_L g854 ( 
.A(n_837),
.B(n_738),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_780),
.B(n_739),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_L g856 ( 
.A(n_788),
.B(n_693),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_777),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_826),
.Y(n_858)
);

OR2x6_ASAP7_75t_L g859 ( 
.A(n_837),
.B(n_738),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_826),
.Y(n_860)
);

BUFx3_ASAP7_75t_L g861 ( 
.A(n_789),
.Y(n_861)
);

INVx2_ASAP7_75t_SL g862 ( 
.A(n_838),
.Y(n_862)
);

INVx3_ASAP7_75t_L g863 ( 
.A(n_824),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_777),
.Y(n_864)
);

INVx5_ASAP7_75t_L g865 ( 
.A(n_836),
.Y(n_865)
);

AND2x4_ASAP7_75t_L g866 ( 
.A(n_784),
.B(n_739),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_L g867 ( 
.A(n_767),
.B(n_680),
.Y(n_867)
);

BUFx6f_ASAP7_75t_L g868 ( 
.A(n_824),
.Y(n_868)
);

BUFx3_ASAP7_75t_L g869 ( 
.A(n_789),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_769),
.Y(n_870)
);

AND2x4_ASAP7_75t_L g871 ( 
.A(n_784),
.B(n_86),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_763),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_783),
.B(n_538),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_L g874 ( 
.A(n_786),
.B(n_754),
.Y(n_874)
);

OR2x6_ASAP7_75t_L g875 ( 
.A(n_842),
.B(n_706),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_830),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_830),
.Y(n_877)
);

INVx3_ASAP7_75t_L g878 ( 
.A(n_824),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_783),
.B(n_538),
.Y(n_879)
);

OR2x2_ASAP7_75t_L g880 ( 
.A(n_842),
.B(n_724),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_769),
.Y(n_881)
);

INVx4_ASAP7_75t_L g882 ( 
.A(n_787),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_775),
.Y(n_883)
);

AND2x2_ASAP7_75t_L g884 ( 
.A(n_827),
.B(n_706),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_L g885 ( 
.A(n_793),
.B(n_751),
.Y(n_885)
);

NOR2xp33_ASAP7_75t_SL g886 ( 
.A(n_820),
.B(n_546),
.Y(n_886)
);

CKINVDCx8_ASAP7_75t_R g887 ( 
.A(n_833),
.Y(n_887)
);

HB1xp67_ASAP7_75t_L g888 ( 
.A(n_812),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_802),
.B(n_545),
.Y(n_889)
);

BUFx2_ASAP7_75t_L g890 ( 
.A(n_787),
.Y(n_890)
);

NOR2xp33_ASAP7_75t_SL g891 ( 
.A(n_820),
.B(n_762),
.Y(n_891)
);

AND2x4_ASAP7_75t_L g892 ( 
.A(n_784),
.B(n_88),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_802),
.B(n_545),
.Y(n_893)
);

HB1xp67_ASAP7_75t_L g894 ( 
.A(n_833),
.Y(n_894)
);

AND2x4_ASAP7_75t_L g895 ( 
.A(n_866),
.B(n_833),
.Y(n_895)
);

INVx3_ASAP7_75t_L g896 ( 
.A(n_846),
.Y(n_896)
);

BUFx6f_ASAP7_75t_L g897 ( 
.A(n_846),
.Y(n_897)
);

BUFx3_ASAP7_75t_L g898 ( 
.A(n_861),
.Y(n_898)
);

NAND2x1p5_ASAP7_75t_L g899 ( 
.A(n_850),
.B(n_865),
.Y(n_899)
);

BUFx6f_ASAP7_75t_L g900 ( 
.A(n_846),
.Y(n_900)
);

BUFx3_ASAP7_75t_L g901 ( 
.A(n_869),
.Y(n_901)
);

INVx6_ASAP7_75t_SL g902 ( 
.A(n_854),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_844),
.Y(n_903)
);

INVx5_ASAP7_75t_L g904 ( 
.A(n_865),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_844),
.Y(n_905)
);

BUFx2_ASAP7_75t_SL g906 ( 
.A(n_887),
.Y(n_906)
);

INVx1_ASAP7_75t_SL g907 ( 
.A(n_888),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_845),
.B(n_793),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_854),
.Y(n_909)
);

BUFx10_ASAP7_75t_L g910 ( 
.A(n_856),
.Y(n_910)
);

BUFx10_ASAP7_75t_L g911 ( 
.A(n_867),
.Y(n_911)
);

BUFx3_ASAP7_75t_L g912 ( 
.A(n_859),
.Y(n_912)
);

BUFx6f_ASAP7_75t_L g913 ( 
.A(n_868),
.Y(n_913)
);

INVx1_ASAP7_75t_SL g914 ( 
.A(n_853),
.Y(n_914)
);

INVxp67_ASAP7_75t_SL g915 ( 
.A(n_868),
.Y(n_915)
);

BUFx3_ASAP7_75t_L g916 ( 
.A(n_859),
.Y(n_916)
);

INVx1_ASAP7_75t_SL g917 ( 
.A(n_866),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_858),
.Y(n_918)
);

INVx5_ASAP7_75t_L g919 ( 
.A(n_865),
.Y(n_919)
);

BUFx6f_ASAP7_75t_L g920 ( 
.A(n_868),
.Y(n_920)
);

INVx3_ASAP7_75t_SL g921 ( 
.A(n_875),
.Y(n_921)
);

INVx3_ASAP7_75t_L g922 ( 
.A(n_850),
.Y(n_922)
);

INVx1_ASAP7_75t_SL g923 ( 
.A(n_851),
.Y(n_923)
);

INVxp67_ASAP7_75t_SL g924 ( 
.A(n_863),
.Y(n_924)
);

INVx1_ASAP7_75t_SL g925 ( 
.A(n_880),
.Y(n_925)
);

INVx1_ASAP7_75t_SL g926 ( 
.A(n_843),
.Y(n_926)
);

BUFx12f_ASAP7_75t_L g927 ( 
.A(n_875),
.Y(n_927)
);

INVx4_ASAP7_75t_L g928 ( 
.A(n_882),
.Y(n_928)
);

INVx2_ASAP7_75t_SL g929 ( 
.A(n_898),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_903),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_905),
.Y(n_931)
);

INVx4_ASAP7_75t_SL g932 ( 
.A(n_897),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_918),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_908),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_914),
.B(n_855),
.Y(n_935)
);

INVx2_ASAP7_75t_SL g936 ( 
.A(n_898),
.Y(n_936)
);

BUFx12f_ASAP7_75t_L g937 ( 
.A(n_909),
.Y(n_937)
);

AOI22xp33_ASAP7_75t_L g938 ( 
.A1(n_926),
.A2(n_764),
.B1(n_816),
.B2(n_818),
.Y(n_938)
);

CKINVDCx11_ASAP7_75t_R g939 ( 
.A(n_921),
.Y(n_939)
);

NAND2x1p5_ASAP7_75t_L g940 ( 
.A(n_904),
.B(n_882),
.Y(n_940)
);

AOI22xp33_ASAP7_75t_L g941 ( 
.A1(n_910),
.A2(n_818),
.B1(n_816),
.B2(n_885),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_922),
.Y(n_942)
);

INVx3_ASAP7_75t_L g943 ( 
.A(n_904),
.Y(n_943)
);

AOI22xp33_ASAP7_75t_L g944 ( 
.A1(n_910),
.A2(n_879),
.B1(n_873),
.B2(n_815),
.Y(n_944)
);

AOI22xp33_ASAP7_75t_SL g945 ( 
.A1(n_927),
.A2(n_891),
.B1(n_874),
.B2(n_886),
.Y(n_945)
);

AOI22xp5_ASAP7_75t_L g946 ( 
.A1(n_923),
.A2(n_884),
.B1(n_787),
.B2(n_804),
.Y(n_946)
);

NAND2xp33_ASAP7_75t_SL g947 ( 
.A(n_922),
.B(n_890),
.Y(n_947)
);

AOI22xp5_ASAP7_75t_L g948 ( 
.A1(n_925),
.A2(n_834),
.B1(n_797),
.B2(n_849),
.Y(n_948)
);

AOI22xp33_ASAP7_75t_SL g949 ( 
.A1(n_927),
.A2(n_768),
.B1(n_770),
.B2(n_819),
.Y(n_949)
);

OAI22xp5_ASAP7_75t_L g950 ( 
.A1(n_904),
.A2(n_797),
.B1(n_863),
.B2(n_878),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_924),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_917),
.B(n_862),
.Y(n_952)
);

BUFx6f_ASAP7_75t_L g953 ( 
.A(n_897),
.Y(n_953)
);

BUFx3_ASAP7_75t_L g954 ( 
.A(n_901),
.Y(n_954)
);

OAI22xp5_ASAP7_75t_L g955 ( 
.A1(n_904),
.A2(n_878),
.B1(n_795),
.B2(n_793),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_896),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_896),
.Y(n_957)
);

AOI22xp33_ASAP7_75t_L g958 ( 
.A1(n_928),
.A2(n_815),
.B1(n_857),
.B2(n_864),
.Y(n_958)
);

OAI21xp5_ASAP7_75t_L g959 ( 
.A1(n_938),
.A2(n_773),
.B(n_823),
.Y(n_959)
);

OAI22xp5_ASAP7_75t_L g960 ( 
.A1(n_941),
.A2(n_794),
.B1(n_872),
.B2(n_876),
.Y(n_960)
);

OAI21xp5_ASAP7_75t_SL g961 ( 
.A1(n_945),
.A2(n_834),
.B(n_828),
.Y(n_961)
);

INVx2_ASAP7_75t_SL g962 ( 
.A(n_954),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_939),
.Y(n_963)
);

INVx4_ASAP7_75t_SL g964 ( 
.A(n_953),
.Y(n_964)
);

AOI22xp33_ASAP7_75t_L g965 ( 
.A1(n_941),
.A2(n_794),
.B1(n_911),
.B2(n_815),
.Y(n_965)
);

AND2x4_ASAP7_75t_SL g966 ( 
.A(n_952),
.B(n_928),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_935),
.B(n_895),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_930),
.Y(n_968)
);

NAND3xp33_ASAP7_75t_L g969 ( 
.A(n_949),
.B(n_776),
.C(n_827),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_934),
.B(n_895),
.Y(n_970)
);

OAI22xp5_ASAP7_75t_L g971 ( 
.A1(n_938),
.A2(n_794),
.B1(n_877),
.B2(n_871),
.Y(n_971)
);

BUFx12f_ASAP7_75t_L g972 ( 
.A(n_939),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_931),
.Y(n_973)
);

INVxp67_ASAP7_75t_L g974 ( 
.A(n_929),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_951),
.B(n_924),
.Y(n_975)
);

BUFx2_ASAP7_75t_L g976 ( 
.A(n_936),
.Y(n_976)
);

AOI211xp5_ASAP7_75t_L g977 ( 
.A1(n_946),
.A2(n_921),
.B(n_828),
.C(n_907),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_933),
.Y(n_978)
);

HB1xp67_ASAP7_75t_L g979 ( 
.A(n_942),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_956),
.Y(n_980)
);

NAND3xp33_ASAP7_75t_L g981 ( 
.A(n_949),
.B(n_821),
.C(n_808),
.Y(n_981)
);

BUFx6f_ASAP7_75t_L g982 ( 
.A(n_953),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_948),
.B(n_852),
.Y(n_983)
);

OAI21xp33_ASAP7_75t_L g984 ( 
.A1(n_945),
.A2(n_779),
.B(n_791),
.Y(n_984)
);

OAI21xp33_ASAP7_75t_L g985 ( 
.A1(n_944),
.A2(n_779),
.B(n_791),
.Y(n_985)
);

OAI22xp5_ASAP7_75t_L g986 ( 
.A1(n_958),
.A2(n_871),
.B1(n_892),
.B2(n_915),
.Y(n_986)
);

OAI222xp33_ASAP7_75t_L g987 ( 
.A1(n_944),
.A2(n_795),
.B1(n_770),
.B2(n_909),
.C1(n_893),
.C2(n_889),
.Y(n_987)
);

AOI22xp33_ASAP7_75t_SL g988 ( 
.A1(n_937),
.A2(n_911),
.B1(n_906),
.B2(n_916),
.Y(n_988)
);

OAI22xp5_ASAP7_75t_L g989 ( 
.A1(n_958),
.A2(n_892),
.B1(n_915),
.B2(n_899),
.Y(n_989)
);

AOI22xp33_ASAP7_75t_L g990 ( 
.A1(n_947),
.A2(n_815),
.B1(n_813),
.B2(n_847),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_957),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_953),
.Y(n_992)
);

OAI222xp33_ASAP7_75t_L g993 ( 
.A1(n_950),
.A2(n_798),
.B1(n_955),
.B2(n_940),
.C1(n_883),
.C2(n_781),
.Y(n_993)
);

OAI22xp5_ASAP7_75t_L g994 ( 
.A1(n_977),
.A2(n_912),
.B1(n_916),
.B2(n_902),
.Y(n_994)
);

AND2x2_ASAP7_75t_SL g995 ( 
.A(n_965),
.B(n_943),
.Y(n_995)
);

AOI22xp33_ASAP7_75t_L g996 ( 
.A1(n_984),
.A2(n_799),
.B1(n_814),
.B2(n_810),
.Y(n_996)
);

AOI22xp33_ASAP7_75t_SL g997 ( 
.A1(n_969),
.A2(n_912),
.B1(n_847),
.B2(n_805),
.Y(n_997)
);

AOI22xp5_ASAP7_75t_L g998 ( 
.A1(n_961),
.A2(n_847),
.B1(n_805),
.B2(n_799),
.Y(n_998)
);

AOI22xp33_ASAP7_75t_L g999 ( 
.A1(n_985),
.A2(n_813),
.B1(n_805),
.B2(n_847),
.Y(n_999)
);

OAI21xp5_ASAP7_75t_SL g1000 ( 
.A1(n_988),
.A2(n_940),
.B(n_841),
.Y(n_1000)
);

AOI22xp33_ASAP7_75t_L g1001 ( 
.A1(n_971),
.A2(n_813),
.B1(n_811),
.B2(n_801),
.Y(n_1001)
);

OAI22xp5_ASAP7_75t_SL g1002 ( 
.A1(n_972),
.A2(n_901),
.B1(n_835),
.B2(n_839),
.Y(n_1002)
);

OAI222xp33_ASAP7_75t_L g1003 ( 
.A1(n_971),
.A2(n_798),
.B1(n_883),
.B2(n_832),
.C1(n_806),
.C2(n_881),
.Y(n_1003)
);

OAI22xp5_ASAP7_75t_L g1004 ( 
.A1(n_983),
.A2(n_902),
.B1(n_899),
.B2(n_919),
.Y(n_1004)
);

AOI22xp33_ASAP7_75t_L g1005 ( 
.A1(n_967),
.A2(n_801),
.B1(n_809),
.B2(n_796),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_970),
.B(n_800),
.Y(n_1006)
);

AOI22xp33_ASAP7_75t_L g1007 ( 
.A1(n_981),
.A2(n_809),
.B1(n_785),
.B2(n_792),
.Y(n_1007)
);

AOI22xp33_ASAP7_75t_L g1008 ( 
.A1(n_960),
.A2(n_800),
.B1(n_782),
.B2(n_822),
.Y(n_1008)
);

HB1xp67_ASAP7_75t_L g1009 ( 
.A(n_968),
.Y(n_1009)
);

AOI22xp33_ASAP7_75t_L g1010 ( 
.A1(n_960),
.A2(n_782),
.B1(n_848),
.B2(n_841),
.Y(n_1010)
);

AOI22xp33_ASAP7_75t_L g1011 ( 
.A1(n_959),
.A2(n_848),
.B1(n_840),
.B2(n_545),
.Y(n_1011)
);

AOI22xp33_ASAP7_75t_L g1012 ( 
.A1(n_986),
.A2(n_782),
.B1(n_840),
.B2(n_775),
.Y(n_1012)
);

AOI22xp33_ASAP7_75t_SL g1013 ( 
.A1(n_986),
.A2(n_919),
.B1(n_943),
.B2(n_771),
.Y(n_1013)
);

AOI22xp33_ASAP7_75t_L g1014 ( 
.A1(n_989),
.A2(n_870),
.B1(n_831),
.B2(n_772),
.Y(n_1014)
);

AOI22xp33_ASAP7_75t_L g1015 ( 
.A1(n_989),
.A2(n_831),
.B1(n_766),
.B2(n_836),
.Y(n_1015)
);

AOI22xp33_ASAP7_75t_L g1016 ( 
.A1(n_959),
.A2(n_831),
.B1(n_836),
.B2(n_774),
.Y(n_1016)
);

OAI21xp33_ASAP7_75t_SL g1017 ( 
.A1(n_990),
.A2(n_860),
.B(n_858),
.Y(n_1017)
);

AOI22xp33_ASAP7_75t_SL g1018 ( 
.A1(n_966),
.A2(n_919),
.B1(n_774),
.B2(n_831),
.Y(n_1018)
);

AOI22xp33_ASAP7_75t_L g1019 ( 
.A1(n_976),
.A2(n_836),
.B1(n_790),
.B2(n_825),
.Y(n_1019)
);

BUFx3_ASAP7_75t_L g1020 ( 
.A(n_962),
.Y(n_1020)
);

AOI22xp5_ASAP7_75t_SL g1021 ( 
.A1(n_963),
.A2(n_790),
.B1(n_953),
.B2(n_836),
.Y(n_1021)
);

AOI22xp33_ASAP7_75t_L g1022 ( 
.A1(n_973),
.A2(n_548),
.B1(n_552),
.B2(n_570),
.Y(n_1022)
);

AOI22xp33_ASAP7_75t_L g1023 ( 
.A1(n_978),
.A2(n_548),
.B1(n_552),
.B2(n_570),
.Y(n_1023)
);

AND2x2_ASAP7_75t_L g1024 ( 
.A(n_979),
.B(n_894),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_975),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_980),
.Y(n_1026)
);

OAI22xp5_ASAP7_75t_L g1027 ( 
.A1(n_974),
.A2(n_919),
.B1(n_825),
.B2(n_829),
.Y(n_1027)
);

AOI22xp33_ASAP7_75t_L g1028 ( 
.A1(n_991),
.A2(n_836),
.B1(n_825),
.B2(n_829),
.Y(n_1028)
);

AOI22xp33_ASAP7_75t_L g1029 ( 
.A1(n_975),
.A2(n_548),
.B1(n_552),
.B2(n_570),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_992),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_982),
.B(n_778),
.Y(n_1031)
);

NAND3xp33_ASAP7_75t_L g1032 ( 
.A(n_1004),
.B(n_586),
.C(n_573),
.Y(n_1032)
);

OAI221xp5_ASAP7_75t_SL g1033 ( 
.A1(n_1000),
.A2(n_987),
.B1(n_778),
.B2(n_993),
.C(n_860),
.Y(n_1033)
);

NAND2xp33_ASAP7_75t_L g1034 ( 
.A(n_994),
.B(n_982),
.Y(n_1034)
);

NOR3xp33_ASAP7_75t_L g1035 ( 
.A(n_1006),
.B(n_964),
.C(n_932),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_1009),
.B(n_982),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_1025),
.B(n_964),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_1026),
.B(n_964),
.Y(n_1038)
);

AND2x2_ASAP7_75t_L g1039 ( 
.A(n_1030),
.B(n_932),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_1003),
.A2(n_920),
.B(n_913),
.Y(n_1040)
);

AND2x2_ASAP7_75t_L g1041 ( 
.A(n_1024),
.B(n_995),
.Y(n_1041)
);

NAND3xp33_ASAP7_75t_L g1042 ( 
.A(n_998),
.B(n_586),
.C(n_573),
.Y(n_1042)
);

OAI22xp5_ASAP7_75t_L g1043 ( 
.A1(n_996),
.A2(n_825),
.B1(n_829),
.B2(n_913),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_995),
.B(n_573),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_1020),
.B(n_997),
.Y(n_1045)
);

NAND3xp33_ASAP7_75t_L g1046 ( 
.A(n_1007),
.B(n_586),
.C(n_556),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_R g1047 ( 
.A(n_1031),
.B(n_897),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_1011),
.B(n_932),
.Y(n_1048)
);

AND2x2_ASAP7_75t_L g1049 ( 
.A(n_1013),
.B(n_897),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_1011),
.B(n_900),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_1017),
.Y(n_1051)
);

NAND3xp33_ASAP7_75t_L g1052 ( 
.A(n_996),
.B(n_593),
.C(n_556),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_1005),
.B(n_900),
.Y(n_1053)
);

AND2x2_ASAP7_75t_SL g1054 ( 
.A(n_1015),
.B(n_900),
.Y(n_1054)
);

AND2x2_ASAP7_75t_L g1055 ( 
.A(n_1021),
.B(n_900),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_1001),
.B(n_913),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_999),
.B(n_913),
.Y(n_1057)
);

NAND4xp25_ASAP7_75t_SL g1058 ( 
.A(n_1029),
.B(n_1016),
.C(n_1019),
.D(n_1018),
.Y(n_1058)
);

NOR3xp33_ASAP7_75t_L g1059 ( 
.A(n_1002),
.B(n_90),
.C(n_91),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_1008),
.B(n_920),
.Y(n_1060)
);

AND2x2_ASAP7_75t_L g1061 ( 
.A(n_1014),
.B(n_920),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_1012),
.B(n_920),
.Y(n_1062)
);

AOI221xp5_ASAP7_75t_L g1063 ( 
.A1(n_1033),
.A2(n_1059),
.B1(n_1058),
.B2(n_1042),
.C(n_1052),
.Y(n_1063)
);

AOI221xp5_ASAP7_75t_L g1064 ( 
.A1(n_1033),
.A2(n_1029),
.B1(n_1022),
.B2(n_1023),
.C(n_1010),
.Y(n_1064)
);

NAND3xp33_ASAP7_75t_L g1065 ( 
.A(n_1059),
.B(n_1023),
.C(n_1022),
.Y(n_1065)
);

HB1xp67_ASAP7_75t_L g1066 ( 
.A(n_1036),
.Y(n_1066)
);

OR2x2_ASAP7_75t_L g1067 ( 
.A(n_1041),
.B(n_1027),
.Y(n_1067)
);

NOR2xp33_ASAP7_75t_L g1068 ( 
.A(n_1045),
.B(n_93),
.Y(n_1068)
);

AND2x2_ASAP7_75t_L g1069 ( 
.A(n_1049),
.B(n_1039),
.Y(n_1069)
);

NAND4xp75_ASAP7_75t_L g1070 ( 
.A(n_1044),
.B(n_100),
.C(n_102),
.D(n_107),
.Y(n_1070)
);

NAND4xp75_ASAP7_75t_L g1071 ( 
.A(n_1055),
.B(n_108),
.C(n_109),
.D(n_110),
.Y(n_1071)
);

AND2x2_ASAP7_75t_L g1072 ( 
.A(n_1037),
.B(n_1028),
.Y(n_1072)
);

AND2x2_ASAP7_75t_L g1073 ( 
.A(n_1047),
.B(n_112),
.Y(n_1073)
);

OR2x2_ASAP7_75t_L g1074 ( 
.A(n_1051),
.B(n_507),
.Y(n_1074)
);

OA211x2_ASAP7_75t_L g1075 ( 
.A1(n_1032),
.A2(n_114),
.B(n_117),
.C(n_119),
.Y(n_1075)
);

NAND4xp75_ASAP7_75t_L g1076 ( 
.A(n_1038),
.B(n_1054),
.C(n_1048),
.D(n_1040),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_1061),
.Y(n_1077)
);

OR2x2_ASAP7_75t_L g1078 ( 
.A(n_1057),
.B(n_121),
.Y(n_1078)
);

OR2x2_ASAP7_75t_L g1079 ( 
.A(n_1050),
.B(n_122),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_1035),
.B(n_1054),
.Y(n_1080)
);

OR2x2_ASAP7_75t_L g1081 ( 
.A(n_1060),
.B(n_124),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_1035),
.Y(n_1082)
);

HB1xp67_ASAP7_75t_L g1083 ( 
.A(n_1062),
.Y(n_1083)
);

AND2x2_ASAP7_75t_L g1084 ( 
.A(n_1034),
.B(n_126),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_1066),
.Y(n_1085)
);

HB1xp67_ASAP7_75t_L g1086 ( 
.A(n_1083),
.Y(n_1086)
);

XNOR2xp5_ASAP7_75t_L g1087 ( 
.A(n_1069),
.B(n_1076),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_1077),
.B(n_1056),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_1074),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_1063),
.A2(n_1046),
.B(n_1043),
.Y(n_1090)
);

AND2x2_ASAP7_75t_L g1091 ( 
.A(n_1082),
.B(n_1053),
.Y(n_1091)
);

OR2x2_ASAP7_75t_L g1092 ( 
.A(n_1067),
.B(n_131),
.Y(n_1092)
);

XOR2x2_ASAP7_75t_L g1093 ( 
.A(n_1068),
.B(n_134),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_1080),
.Y(n_1094)
);

INVx3_ASAP7_75t_L g1095 ( 
.A(n_1072),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_1080),
.Y(n_1096)
);

INVxp67_ASAP7_75t_L g1097 ( 
.A(n_1081),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_1079),
.Y(n_1098)
);

NOR2xp33_ASAP7_75t_L g1099 ( 
.A(n_1078),
.B(n_137),
.Y(n_1099)
);

AND2x2_ASAP7_75t_L g1100 ( 
.A(n_1073),
.B(n_138),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_SL g1101 ( 
.A(n_1063),
.B(n_556),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_1084),
.B(n_593),
.Y(n_1102)
);

XOR2x2_ASAP7_75t_L g1103 ( 
.A(n_1071),
.B(n_141),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_1064),
.B(n_593),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_1086),
.Y(n_1105)
);

OA22x2_ASAP7_75t_L g1106 ( 
.A1(n_1087),
.A2(n_1101),
.B1(n_1096),
.B2(n_1094),
.Y(n_1106)
);

AND2x2_ASAP7_75t_L g1107 ( 
.A(n_1095),
.B(n_1070),
.Y(n_1107)
);

XOR2x2_ASAP7_75t_L g1108 ( 
.A(n_1093),
.B(n_1065),
.Y(n_1108)
);

XOR2x2_ASAP7_75t_L g1109 ( 
.A(n_1101),
.B(n_1065),
.Y(n_1109)
);

NOR2xp33_ASAP7_75t_L g1110 ( 
.A(n_1097),
.B(n_142),
.Y(n_1110)
);

XNOR2x1_ASAP7_75t_L g1111 ( 
.A(n_1103),
.B(n_1075),
.Y(n_1111)
);

AO22x2_ASAP7_75t_L g1112 ( 
.A1(n_1085),
.A2(n_1064),
.B1(n_147),
.B2(n_149),
.Y(n_1112)
);

AO22x1_ASAP7_75t_L g1113 ( 
.A1(n_1095),
.A2(n_829),
.B1(n_499),
.B2(n_156),
.Y(n_1113)
);

INVxp67_ASAP7_75t_L g1114 ( 
.A(n_1091),
.Y(n_1114)
);

OAI22x1_ASAP7_75t_L g1115 ( 
.A1(n_1097),
.A2(n_499),
.B1(n_152),
.B2(n_158),
.Y(n_1115)
);

HB1xp67_ASAP7_75t_L g1116 ( 
.A(n_1086),
.Y(n_1116)
);

OAI22x1_ASAP7_75t_L g1117 ( 
.A1(n_1098),
.A2(n_1089),
.B1(n_1088),
.B2(n_1092),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1089),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_1090),
.B(n_144),
.Y(n_1119)
);

NOR2x1_ASAP7_75t_R g1120 ( 
.A(n_1104),
.B(n_159),
.Y(n_1120)
);

INVx1_ASAP7_75t_SL g1121 ( 
.A(n_1100),
.Y(n_1121)
);

INVx2_ASAP7_75t_SL g1122 ( 
.A(n_1102),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_1099),
.B(n_161),
.Y(n_1123)
);

AOI22x1_ASAP7_75t_L g1124 ( 
.A1(n_1112),
.A2(n_1099),
.B1(n_164),
.B2(n_165),
.Y(n_1124)
);

AO22x2_ASAP7_75t_L g1125 ( 
.A1(n_1105),
.A2(n_162),
.B1(n_166),
.B2(n_169),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_1114),
.B(n_170),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1116),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_1118),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_1107),
.Y(n_1129)
);

AOI22x1_ASAP7_75t_L g1130 ( 
.A1(n_1112),
.A2(n_299),
.B1(n_172),
.B2(n_174),
.Y(n_1130)
);

INVx2_ASAP7_75t_SL g1131 ( 
.A(n_1122),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_1117),
.Y(n_1132)
);

XOR2x2_ASAP7_75t_L g1133 ( 
.A(n_1108),
.B(n_171),
.Y(n_1133)
);

XNOR2xp5_ASAP7_75t_L g1134 ( 
.A(n_1111),
.B(n_179),
.Y(n_1134)
);

INVx1_ASAP7_75t_SL g1135 ( 
.A(n_1121),
.Y(n_1135)
);

INVx1_ASAP7_75t_SL g1136 ( 
.A(n_1109),
.Y(n_1136)
);

AOI22xp5_ASAP7_75t_L g1137 ( 
.A1(n_1106),
.A2(n_180),
.B1(n_188),
.B2(n_190),
.Y(n_1137)
);

OA22x2_ASAP7_75t_L g1138 ( 
.A1(n_1119),
.A2(n_1115),
.B1(n_1123),
.B2(n_1120),
.Y(n_1138)
);

BUFx2_ASAP7_75t_L g1139 ( 
.A(n_1113),
.Y(n_1139)
);

OA22x2_ASAP7_75t_L g1140 ( 
.A1(n_1113),
.A2(n_193),
.B1(n_195),
.B2(n_200),
.Y(n_1140)
);

XOR2x2_ASAP7_75t_L g1141 ( 
.A(n_1110),
.B(n_207),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_1129),
.Y(n_1142)
);

INVx2_ASAP7_75t_SL g1143 ( 
.A(n_1131),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1127),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1128),
.Y(n_1145)
);

INVxp67_ASAP7_75t_L g1146 ( 
.A(n_1139),
.Y(n_1146)
);

OAI22xp5_ASAP7_75t_L g1147 ( 
.A1(n_1146),
.A2(n_1137),
.B1(n_1136),
.B2(n_1138),
.Y(n_1147)
);

NAND4xp25_ASAP7_75t_L g1148 ( 
.A(n_1146),
.B(n_1132),
.C(n_1135),
.D(n_1126),
.Y(n_1148)
);

AOI22xp5_ASAP7_75t_L g1149 ( 
.A1(n_1143),
.A2(n_1140),
.B1(n_1133),
.B2(n_1125),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1145),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1144),
.Y(n_1151)
);

OAI22xp5_ASAP7_75t_L g1152 ( 
.A1(n_1149),
.A2(n_1124),
.B1(n_1130),
.B2(n_1142),
.Y(n_1152)
);

OAI22xp5_ASAP7_75t_L g1153 ( 
.A1(n_1147),
.A2(n_1124),
.B1(n_1130),
.B2(n_1134),
.Y(n_1153)
);

AOI22x1_ASAP7_75t_SL g1154 ( 
.A1(n_1148),
.A2(n_1141),
.B1(n_1125),
.B2(n_213),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1150),
.Y(n_1155)
);

AOI22xp5_ASAP7_75t_L g1156 ( 
.A1(n_1153),
.A2(n_1151),
.B1(n_210),
.B2(n_217),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1155),
.Y(n_1157)
);

AND2x2_ASAP7_75t_L g1158 ( 
.A(n_1152),
.B(n_209),
.Y(n_1158)
);

AOI22xp5_ASAP7_75t_L g1159 ( 
.A1(n_1154),
.A2(n_219),
.B1(n_222),
.B2(n_224),
.Y(n_1159)
);

HB1xp67_ASAP7_75t_L g1160 ( 
.A(n_1158),
.Y(n_1160)
);

AOI22xp5_ASAP7_75t_L g1161 ( 
.A1(n_1159),
.A2(n_225),
.B1(n_226),
.B2(n_227),
.Y(n_1161)
);

AO211x2_ASAP7_75t_L g1162 ( 
.A1(n_1160),
.A2(n_1157),
.B(n_1156),
.C(n_232),
.Y(n_1162)
);

INVxp67_ASAP7_75t_L g1163 ( 
.A(n_1162),
.Y(n_1163)
);

AO22x2_ASAP7_75t_L g1164 ( 
.A1(n_1163),
.A2(n_1161),
.B1(n_229),
.B2(n_233),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1164),
.Y(n_1165)
);

AOI22xp5_ASAP7_75t_L g1166 ( 
.A1(n_1165),
.A2(n_228),
.B1(n_235),
.B2(n_236),
.Y(n_1166)
);

AO22x1_ASAP7_75t_SL g1167 ( 
.A1(n_1165),
.A2(n_237),
.B1(n_238),
.B2(n_243),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1167),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1166),
.Y(n_1169)
);

AOI22xp5_ASAP7_75t_L g1170 ( 
.A1(n_1168),
.A2(n_1169),
.B1(n_246),
.B2(n_247),
.Y(n_1170)
);

OAI22xp5_ASAP7_75t_L g1171 ( 
.A1(n_1168),
.A2(n_244),
.B1(n_248),
.B2(n_249),
.Y(n_1171)
);

HB1xp67_ASAP7_75t_L g1172 ( 
.A(n_1171),
.Y(n_1172)
);

AOI221xp5_ASAP7_75t_L g1173 ( 
.A1(n_1172),
.A2(n_1170),
.B1(n_253),
.B2(n_254),
.C(n_257),
.Y(n_1173)
);

AOI211xp5_ASAP7_75t_L g1174 ( 
.A1(n_1173),
.A2(n_250),
.B(n_283),
.C(n_286),
.Y(n_1174)
);


endmodule