module fake_jpeg_29923_n_72 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_72);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_72;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_44;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_62;
wire n_31;
wire n_25;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;
wire n_70;
wire n_66;

BUFx3_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

INVx3_ASAP7_75t_SL g28 ( 
.A(n_13),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_3),
.B(n_1),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_28),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_34),
.Y(n_44)
);

OR2x2_ASAP7_75t_SL g33 ( 
.A(n_29),
.B(n_0),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_33),
.A2(n_36),
.B(n_4),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_29),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_1),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_35),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g36 ( 
.A1(n_28),
.A2(n_14),
.B(n_23),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_28),
.A2(n_12),
.B1(n_22),
.B2(n_20),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_37),
.A2(n_31),
.B1(n_27),
.B2(n_25),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_27),
.B(n_2),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_38),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_41),
.A2(n_42),
.B(n_47),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_37),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_43),
.B(n_45),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_33),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_46),
.Y(n_48)
);

OA22x2_ASAP7_75t_L g47 ( 
.A1(n_37),
.A2(n_26),
.B1(n_31),
.B2(n_25),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_40),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g59 ( 
.A(n_51),
.B(n_52),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_4),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_5),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_53),
.B(n_6),
.C(n_7),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_47),
.A2(n_31),
.B1(n_26),
.B2(n_30),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_55),
.A2(n_24),
.B1(n_15),
.B2(n_8),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_26),
.C(n_30),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_16),
.C(n_18),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_54),
.B(n_6),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_57),
.B(n_58),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_61),
.A2(n_48),
.B1(n_49),
.B2(n_7),
.Y(n_67)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_63),
.B(n_17),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_65),
.B(n_63),
.C(n_60),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_67),
.B(n_59),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_68),
.B(n_69),
.Y(n_70)
);

OAI321xp33_ASAP7_75t_L g71 ( 
.A1(n_70),
.A2(n_67),
.A3(n_66),
.B1(n_64),
.B2(n_19),
.C(n_9),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_71),
.B(n_11),
.Y(n_72)
);


endmodule