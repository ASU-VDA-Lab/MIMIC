module real_aes_8001_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_717, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_717;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_635;
wire n_503;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_417;
wire n_182;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_502;
wire n_434;
wire n_527;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g170 ( .A1(n_0), .A2(n_171), .B(n_172), .C(n_176), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_1), .B(n_165), .Y(n_178) );
NAND3xp33_ASAP7_75t_SL g106 ( .A(n_2), .B(n_107), .C(n_108), .Y(n_106) );
INVx1_ASAP7_75t_L g423 ( .A(n_2), .Y(n_423) );
NAND2xp5_ASAP7_75t_SL g149 ( .A(n_3), .B(n_150), .Y(n_149) );
A2O1A1Ixp33_ASAP7_75t_L g465 ( .A1(n_4), .A2(n_139), .B(n_156), .C(n_466), .Y(n_465) );
AOI21xp5_ASAP7_75t_L g486 ( .A1(n_5), .A2(n_159), .B(n_487), .Y(n_486) );
AOI21xp5_ASAP7_75t_L g260 ( .A1(n_6), .A2(n_159), .B(n_261), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_7), .B(n_165), .Y(n_493) );
AO21x2_ASAP7_75t_L g217 ( .A1(n_8), .A2(n_131), .B(n_218), .Y(n_217) );
AND2x6_ASAP7_75t_L g156 ( .A(n_9), .B(n_157), .Y(n_156) );
A2O1A1Ixp33_ASAP7_75t_L g235 ( .A1(n_10), .A2(n_139), .B(n_156), .C(n_236), .Y(n_235) );
INVx1_ASAP7_75t_L g458 ( .A(n_11), .Y(n_458) );
NOR2xp33_ASAP7_75t_L g112 ( .A(n_12), .B(n_40), .Y(n_112) );
NAND2xp5_ASAP7_75t_SL g468 ( .A(n_13), .B(n_175), .Y(n_468) );
INVx1_ASAP7_75t_L g136 ( .A(n_14), .Y(n_136) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_15), .B(n_150), .Y(n_224) );
A2O1A1Ixp33_ASAP7_75t_L g476 ( .A1(n_16), .A2(n_151), .B(n_477), .C(n_479), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_17), .B(n_165), .Y(n_480) );
OAI22xp5_ASAP7_75t_SL g121 ( .A1(n_18), .A2(n_65), .B1(n_122), .B2(n_123), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_18), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_19), .B(n_208), .Y(n_527) );
A2O1A1Ixp33_ASAP7_75t_L g201 ( .A1(n_20), .A2(n_139), .B(n_202), .C(n_207), .Y(n_201) );
A2O1A1Ixp33_ASAP7_75t_L g447 ( .A1(n_21), .A2(n_174), .B(n_226), .C(n_448), .Y(n_447) );
NAND2xp5_ASAP7_75t_SL g500 ( .A(n_22), .B(n_175), .Y(n_500) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_23), .B(n_175), .Y(n_509) );
CKINVDCx16_ASAP7_75t_R g496 ( .A(n_24), .Y(n_496) );
INVx1_ASAP7_75t_L g508 ( .A(n_25), .Y(n_508) );
A2O1A1Ixp33_ASAP7_75t_L g220 ( .A1(n_26), .A2(n_139), .B(n_207), .C(n_221), .Y(n_220) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_27), .Y(n_143) );
CKINVDCx20_ASAP7_75t_R g464 ( .A(n_28), .Y(n_464) );
INVx1_ASAP7_75t_L g525 ( .A(n_29), .Y(n_525) );
AOI21xp5_ASAP7_75t_L g166 ( .A1(n_30), .A2(n_159), .B(n_167), .Y(n_166) );
INVx2_ASAP7_75t_L g141 ( .A(n_31), .Y(n_141) );
A2O1A1Ixp33_ASAP7_75t_L g185 ( .A1(n_32), .A2(n_154), .B(n_186), .C(n_187), .Y(n_185) );
CKINVDCx20_ASAP7_75t_R g471 ( .A(n_33), .Y(n_471) );
A2O1A1Ixp33_ASAP7_75t_L g489 ( .A1(n_34), .A2(n_174), .B(n_490), .C(n_492), .Y(n_489) );
AOI22xp33_ASAP7_75t_L g119 ( .A1(n_35), .A2(n_120), .B1(n_415), .B2(n_416), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g415 ( .A(n_35), .Y(n_415) );
INVxp67_ASAP7_75t_L g526 ( .A(n_36), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_37), .B(n_223), .Y(n_222) );
CKINVDCx14_ASAP7_75t_R g488 ( .A(n_38), .Y(n_488) );
A2O1A1Ixp33_ASAP7_75t_L g506 ( .A1(n_39), .A2(n_139), .B(n_207), .C(n_507), .Y(n_506) );
AOI222xp33_ASAP7_75t_L g429 ( .A1(n_41), .A2(n_430), .B1(n_698), .B2(n_699), .C1(n_705), .C2(n_709), .Y(n_429) );
A2O1A1Ixp33_ASAP7_75t_L g455 ( .A1(n_42), .A2(n_176), .B(n_456), .C(n_457), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_43), .B(n_200), .Y(n_199) );
CKINVDCx20_ASAP7_75t_R g240 ( .A(n_44), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_45), .B(n_150), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_46), .B(n_159), .Y(n_219) );
CKINVDCx20_ASAP7_75t_R g511 ( .A(n_47), .Y(n_511) );
CKINVDCx20_ASAP7_75t_R g522 ( .A(n_48), .Y(n_522) );
A2O1A1Ixp33_ASAP7_75t_L g246 ( .A1(n_49), .A2(n_154), .B(n_186), .C(n_247), .Y(n_246) );
INVx1_ASAP7_75t_L g173 ( .A(n_50), .Y(n_173) );
AOI22xp5_ASAP7_75t_L g699 ( .A1(n_51), .A2(n_700), .B1(n_701), .B2(n_702), .Y(n_699) );
CKINVDCx20_ASAP7_75t_R g700 ( .A(n_51), .Y(n_700) );
OAI22xp5_ASAP7_75t_L g702 ( .A1(n_52), .A2(n_84), .B1(n_703), .B2(n_704), .Y(n_702) );
CKINVDCx20_ASAP7_75t_R g704 ( .A(n_52), .Y(n_704) );
INVx1_ASAP7_75t_L g248 ( .A(n_53), .Y(n_248) );
INVx1_ASAP7_75t_L g446 ( .A(n_54), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_55), .B(n_159), .Y(n_245) );
CKINVDCx20_ASAP7_75t_R g211 ( .A(n_56), .Y(n_211) );
CKINVDCx14_ASAP7_75t_R g454 ( .A(n_57), .Y(n_454) );
INVx1_ASAP7_75t_L g157 ( .A(n_58), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_59), .B(n_159), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_60), .B(n_165), .Y(n_266) );
A2O1A1Ixp33_ASAP7_75t_L g263 ( .A1(n_61), .A2(n_146), .B(n_206), .C(n_264), .Y(n_263) );
INVx1_ASAP7_75t_L g135 ( .A(n_62), .Y(n_135) );
INVx1_ASAP7_75t_SL g491 ( .A(n_63), .Y(n_491) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_64), .Y(n_117) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_65), .Y(n_122) );
NAND2xp5_ASAP7_75t_SL g191 ( .A(n_66), .B(n_150), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_67), .B(n_165), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_68), .B(n_151), .Y(n_237) );
INVx1_ASAP7_75t_L g499 ( .A(n_69), .Y(n_499) );
CKINVDCx16_ASAP7_75t_R g168 ( .A(n_70), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_71), .B(n_190), .Y(n_203) );
A2O1A1Ixp33_ASAP7_75t_L g138 ( .A1(n_72), .A2(n_139), .B(n_144), .C(n_154), .Y(n_138) );
CKINVDCx16_ASAP7_75t_R g262 ( .A(n_73), .Y(n_262) );
INVx1_ASAP7_75t_L g110 ( .A(n_74), .Y(n_110) );
AOI22xp5_ASAP7_75t_L g103 ( .A1(n_75), .A2(n_104), .B1(n_113), .B2(n_714), .Y(n_103) );
AOI21xp5_ASAP7_75t_L g452 ( .A1(n_76), .A2(n_159), .B(n_453), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_77), .B(n_425), .Y(n_424) );
CKINVDCx20_ASAP7_75t_R g502 ( .A(n_78), .Y(n_502) );
AOI21xp5_ASAP7_75t_L g473 ( .A1(n_79), .A2(n_159), .B(n_474), .Y(n_473) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_80), .A2(n_200), .B(n_521), .Y(n_520) );
INVx1_ASAP7_75t_L g475 ( .A(n_81), .Y(n_475) );
CKINVDCx16_ASAP7_75t_R g505 ( .A(n_82), .Y(n_505) );
NAND2xp5_ASAP7_75t_SL g204 ( .A(n_83), .B(n_189), .Y(n_204) );
CKINVDCx20_ASAP7_75t_R g703 ( .A(n_84), .Y(n_703) );
CKINVDCx20_ASAP7_75t_R g195 ( .A(n_85), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g444 ( .A1(n_86), .A2(n_159), .B(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g478 ( .A(n_87), .Y(n_478) );
INVx2_ASAP7_75t_L g133 ( .A(n_88), .Y(n_133) );
INVx1_ASAP7_75t_L g467 ( .A(n_89), .Y(n_467) );
CKINVDCx20_ASAP7_75t_R g163 ( .A(n_90), .Y(n_163) );
NAND2xp5_ASAP7_75t_SL g238 ( .A(n_91), .B(n_175), .Y(n_238) );
INVx2_ASAP7_75t_L g107 ( .A(n_92), .Y(n_107) );
OR2x2_ASAP7_75t_L g420 ( .A(n_92), .B(n_421), .Y(n_420) );
OR2x2_ASAP7_75t_L g433 ( .A(n_92), .B(n_422), .Y(n_433) );
A2O1A1Ixp33_ASAP7_75t_L g497 ( .A1(n_93), .A2(n_139), .B(n_154), .C(n_498), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_94), .B(n_159), .Y(n_184) );
INVx1_ASAP7_75t_L g188 ( .A(n_95), .Y(n_188) );
INVxp67_ASAP7_75t_L g265 ( .A(n_96), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_97), .B(n_131), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_98), .B(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g145 ( .A(n_99), .Y(n_145) );
INVx1_ASAP7_75t_L g233 ( .A(n_100), .Y(n_233) );
INVx2_ASAP7_75t_L g449 ( .A(n_101), .Y(n_449) );
AND2x2_ASAP7_75t_L g250 ( .A(n_102), .B(n_193), .Y(n_250) );
INVx1_ASAP7_75t_SL g715 ( .A(n_104), .Y(n_715) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
OR2x2_ASAP7_75t_SL g105 ( .A(n_106), .B(n_111), .Y(n_105) );
OR2x2_ASAP7_75t_L g436 ( .A(n_107), .B(n_422), .Y(n_436) );
NOR2x2_ASAP7_75t_L g711 ( .A(n_107), .B(n_421), .Y(n_711) );
INVx1_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
INVxp67_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
AND2x2_ASAP7_75t_L g422 ( .A(n_112), .B(n_423), .Y(n_422) );
AO21x2_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_118), .B(n_428), .Y(n_113) );
HB1xp67_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx2_ASAP7_75t_SL g115 ( .A(n_116), .Y(n_115) );
BUFx2_ASAP7_75t_L g713 ( .A(n_116), .Y(n_713) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
OAI21xp5_ASAP7_75t_SL g118 ( .A1(n_119), .A2(n_417), .B(n_424), .Y(n_118) );
INVx1_ASAP7_75t_L g416 ( .A(n_120), .Y(n_416) );
XNOR2xp5_ASAP7_75t_L g120 ( .A(n_121), .B(n_124), .Y(n_120) );
INVx2_ASAP7_75t_L g434 ( .A(n_124), .Y(n_434) );
AOI22xp5_ASAP7_75t_L g706 ( .A1(n_124), .A2(n_432), .B1(n_707), .B2(n_708), .Y(n_706) );
NAND2x1p5_ASAP7_75t_L g124 ( .A(n_125), .B(n_358), .Y(n_124) );
AND4x1_ASAP7_75t_L g125 ( .A(n_126), .B(n_298), .C(n_313), .D(n_338), .Y(n_125) );
NOR2xp33_ASAP7_75t_SL g126 ( .A(n_127), .B(n_271), .Y(n_126) );
OAI21xp33_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_179), .B(n_251), .Y(n_127) );
AND2x2_ASAP7_75t_L g301 ( .A(n_128), .B(n_197), .Y(n_301) );
AND2x2_ASAP7_75t_L g314 ( .A(n_128), .B(n_196), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_128), .B(n_180), .Y(n_364) );
INVx1_ASAP7_75t_L g368 ( .A(n_128), .Y(n_368) );
AND2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_164), .Y(n_128) );
INVx2_ASAP7_75t_L g285 ( .A(n_129), .Y(n_285) );
BUFx2_ASAP7_75t_L g312 ( .A(n_129), .Y(n_312) );
AO21x2_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_137), .B(n_162), .Y(n_129) );
NOR2xp33_ASAP7_75t_L g162 ( .A(n_130), .B(n_163), .Y(n_162) );
INVx3_ASAP7_75t_L g165 ( .A(n_130), .Y(n_165) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_130), .B(n_195), .Y(n_194) );
AO21x2_ASAP7_75t_L g231 ( .A1(n_130), .A2(n_232), .B(n_239), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g470 ( .A(n_130), .B(n_471), .Y(n_470) );
AO21x2_ASAP7_75t_L g494 ( .A1(n_130), .A2(n_495), .B(n_501), .Y(n_494) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_130), .B(n_511), .Y(n_510) );
INVx4_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
AOI21xp5_ASAP7_75t_L g218 ( .A1(n_131), .A2(n_219), .B(n_220), .Y(n_218) );
HB1xp67_ASAP7_75t_L g259 ( .A(n_131), .Y(n_259) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx1_ASAP7_75t_L g241 ( .A(n_132), .Y(n_241) );
AND2x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_134), .Y(n_132) );
AND2x2_ASAP7_75t_SL g193 ( .A(n_133), .B(n_134), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_135), .B(n_136), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_138), .B(n_158), .Y(n_137) );
INVx5_ASAP7_75t_L g169 ( .A(n_139), .Y(n_169) );
AND2x6_ASAP7_75t_L g139 ( .A(n_140), .B(n_142), .Y(n_139) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_140), .Y(n_153) );
BUFx3_ASAP7_75t_L g177 ( .A(n_140), .Y(n_177) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx1_ASAP7_75t_L g161 ( .A(n_141), .Y(n_161) );
INVx1_ASAP7_75t_L g227 ( .A(n_141), .Y(n_227) );
INVx1_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_143), .Y(n_148) );
INVx3_ASAP7_75t_L g151 ( .A(n_143), .Y(n_151) );
AND2x2_ASAP7_75t_L g160 ( .A(n_143), .B(n_161), .Y(n_160) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_143), .Y(n_175) );
INVx1_ASAP7_75t_L g223 ( .A(n_143), .Y(n_223) );
O2A1O1Ixp33_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_146), .B(n_149), .C(n_152), .Y(n_144) );
INVx1_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
NOR2xp33_ASAP7_75t_L g448 ( .A(n_147), .B(n_449), .Y(n_448) );
NOR2xp33_ASAP7_75t_L g477 ( .A(n_147), .B(n_478), .Y(n_477) );
OAI22xp33_ASAP7_75t_L g524 ( .A1(n_147), .A2(n_150), .B1(n_525), .B2(n_526), .Y(n_524) );
INVx4_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g190 ( .A(n_148), .Y(n_190) );
INVx2_ASAP7_75t_L g171 ( .A(n_150), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g264 ( .A(n_150), .B(n_265), .Y(n_264) );
O2A1O1Ixp33_ASAP7_75t_L g507 ( .A1(n_150), .A2(n_205), .B(n_508), .C(n_509), .Y(n_507) );
INVx5_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
NOR2xp33_ASAP7_75t_L g457 ( .A(n_151), .B(n_458), .Y(n_457) );
HB1xp67_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx3_ASAP7_75t_L g492 ( .A(n_153), .Y(n_492) );
INVx1_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
O2A1O1Ixp33_ASAP7_75t_SL g167 ( .A1(n_155), .A2(n_168), .B(n_169), .C(n_170), .Y(n_167) );
O2A1O1Ixp33_ASAP7_75t_L g261 ( .A1(n_155), .A2(n_169), .B(n_262), .C(n_263), .Y(n_261) );
O2A1O1Ixp33_ASAP7_75t_SL g445 ( .A1(n_155), .A2(n_169), .B(n_446), .C(n_447), .Y(n_445) );
O2A1O1Ixp33_ASAP7_75t_SL g453 ( .A1(n_155), .A2(n_169), .B(n_454), .C(n_455), .Y(n_453) );
O2A1O1Ixp33_ASAP7_75t_SL g474 ( .A1(n_155), .A2(n_169), .B(n_475), .C(n_476), .Y(n_474) );
O2A1O1Ixp33_ASAP7_75t_L g487 ( .A1(n_155), .A2(n_169), .B(n_488), .C(n_489), .Y(n_487) );
O2A1O1Ixp33_ASAP7_75t_SL g521 ( .A1(n_155), .A2(n_169), .B(n_522), .C(n_523), .Y(n_521) );
INVx4_ASAP7_75t_SL g155 ( .A(n_156), .Y(n_155) );
AND2x4_ASAP7_75t_L g159 ( .A(n_156), .B(n_160), .Y(n_159) );
BUFx3_ASAP7_75t_L g207 ( .A(n_156), .Y(n_207) );
NAND2x1p5_ASAP7_75t_L g234 ( .A(n_156), .B(n_160), .Y(n_234) );
BUFx2_ASAP7_75t_L g200 ( .A(n_159), .Y(n_200) );
INVx1_ASAP7_75t_L g206 ( .A(n_161), .Y(n_206) );
AND2x2_ASAP7_75t_L g252 ( .A(n_164), .B(n_197), .Y(n_252) );
INVx2_ASAP7_75t_L g268 ( .A(n_164), .Y(n_268) );
AND2x2_ASAP7_75t_L g277 ( .A(n_164), .B(n_196), .Y(n_277) );
AND2x2_ASAP7_75t_L g356 ( .A(n_164), .B(n_285), .Y(n_356) );
OA21x2_ASAP7_75t_L g164 ( .A1(n_165), .A2(n_166), .B(n_178), .Y(n_164) );
INVx2_ASAP7_75t_L g186 ( .A(n_169), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g172 ( .A(n_173), .B(n_174), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g490 ( .A(n_174), .B(n_491), .Y(n_490) );
INVx4_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx2_ASAP7_75t_L g456 ( .A(n_175), .Y(n_456) );
INVx2_ASAP7_75t_L g469 ( .A(n_176), .Y(n_469) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
HB1xp67_ASAP7_75t_L g192 ( .A(n_177), .Y(n_192) );
INVx1_ASAP7_75t_L g479 ( .A(n_177), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_180), .B(n_213), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_180), .B(n_283), .Y(n_321) );
INVx1_ASAP7_75t_L g409 ( .A(n_180), .Y(n_409) );
AND2x2_ASAP7_75t_L g180 ( .A(n_181), .B(n_196), .Y(n_180) );
AND2x2_ASAP7_75t_L g267 ( .A(n_181), .B(n_268), .Y(n_267) );
OR2x2_ASAP7_75t_L g281 ( .A(n_181), .B(n_282), .Y(n_281) );
HB1xp67_ASAP7_75t_L g310 ( .A(n_181), .Y(n_310) );
OR2x2_ASAP7_75t_L g342 ( .A(n_181), .B(n_284), .Y(n_342) );
AND2x2_ASAP7_75t_L g350 ( .A(n_181), .B(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g383 ( .A(n_181), .B(n_352), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_181), .B(n_252), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_181), .B(n_312), .Y(n_408) );
AND2x2_ASAP7_75t_L g414 ( .A(n_181), .B(n_301), .Y(n_414) );
INVx5_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
BUFx2_ASAP7_75t_L g274 ( .A(n_182), .Y(n_274) );
AND2x2_ASAP7_75t_L g304 ( .A(n_182), .B(n_284), .Y(n_304) );
AND2x2_ASAP7_75t_L g337 ( .A(n_182), .B(n_297), .Y(n_337) );
AND2x2_ASAP7_75t_L g357 ( .A(n_182), .B(n_197), .Y(n_357) );
AND2x2_ASAP7_75t_L g391 ( .A(n_182), .B(n_257), .Y(n_391) );
OR2x6_ASAP7_75t_L g182 ( .A(n_183), .B(n_194), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g183 ( .A1(n_184), .A2(n_185), .B(n_193), .Y(n_183) );
O2A1O1Ixp33_ASAP7_75t_L g187 ( .A1(n_188), .A2(n_189), .B(n_191), .C(n_192), .Y(n_187) );
O2A1O1Ixp33_ASAP7_75t_L g247 ( .A1(n_189), .A2(n_192), .B(n_248), .C(n_249), .Y(n_247) );
O2A1O1Ixp5_ASAP7_75t_L g466 ( .A1(n_189), .A2(n_467), .B(n_468), .C(n_469), .Y(n_466) );
O2A1O1Ixp33_ASAP7_75t_L g498 ( .A1(n_189), .A2(n_469), .B(n_499), .C(n_500), .Y(n_498) );
INVx2_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
INVx2_ASAP7_75t_L g209 ( .A(n_193), .Y(n_209) );
INVx1_ASAP7_75t_L g212 ( .A(n_193), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g244 ( .A1(n_193), .A2(n_245), .B(n_246), .Y(n_244) );
OA21x2_ASAP7_75t_L g451 ( .A1(n_193), .A2(n_452), .B(n_459), .Y(n_451) );
O2A1O1Ixp33_ASAP7_75t_L g504 ( .A1(n_193), .A2(n_234), .B(n_505), .C(n_506), .Y(n_504) );
AND2x4_ASAP7_75t_L g297 ( .A(n_196), .B(n_268), .Y(n_297) );
AND2x2_ASAP7_75t_L g308 ( .A(n_196), .B(n_304), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_196), .B(n_284), .Y(n_347) );
INVx2_ASAP7_75t_L g362 ( .A(n_196), .Y(n_362) );
NOR2xp33_ASAP7_75t_L g385 ( .A(n_196), .B(n_296), .Y(n_385) );
AND2x2_ASAP7_75t_L g404 ( .A(n_196), .B(n_356), .Y(n_404) );
INVx5_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
HB1xp67_ASAP7_75t_L g303 ( .A(n_197), .Y(n_303) );
AND2x2_ASAP7_75t_L g311 ( .A(n_197), .B(n_312), .Y(n_311) );
AND2x4_ASAP7_75t_L g352 ( .A(n_197), .B(n_268), .Y(n_352) );
OR2x6_ASAP7_75t_L g197 ( .A(n_198), .B(n_210), .Y(n_197) );
AOI21xp5_ASAP7_75t_SL g198 ( .A1(n_199), .A2(n_201), .B(n_208), .Y(n_198) );
AOI21xp5_ASAP7_75t_L g202 ( .A1(n_203), .A2(n_204), .B(n_205), .Y(n_202) );
INVx2_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g523 ( .A(n_206), .B(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_209), .B(n_502), .Y(n_501) );
NOR2xp33_ASAP7_75t_L g210 ( .A(n_211), .B(n_212), .Y(n_210) );
AO21x2_ASAP7_75t_L g462 ( .A1(n_212), .A2(n_463), .B(n_470), .Y(n_462) );
INVx1_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_215), .B(n_228), .Y(n_214) );
AND2x2_ASAP7_75t_L g275 ( .A(n_215), .B(n_258), .Y(n_275) );
INVx1_ASAP7_75t_SL g215 ( .A(n_216), .Y(n_215) );
NAND2xp5_ASAP7_75t_SL g255 ( .A(n_216), .B(n_231), .Y(n_255) );
OR2x2_ASAP7_75t_L g288 ( .A(n_216), .B(n_258), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_216), .B(n_258), .Y(n_293) );
AND2x2_ASAP7_75t_L g320 ( .A(n_216), .B(n_257), .Y(n_320) );
AND2x2_ASAP7_75t_L g372 ( .A(n_216), .B(n_230), .Y(n_372) );
INVx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_217), .B(n_242), .Y(n_280) );
AND2x2_ASAP7_75t_L g316 ( .A(n_217), .B(n_231), .Y(n_316) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_222), .A2(n_224), .B(n_225), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g236 ( .A1(n_225), .A2(n_237), .B(n_238), .Y(n_236) );
INVx2_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
INVx3_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_228), .B(n_380), .Y(n_379) );
INVx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
OR2x2_ASAP7_75t_L g306 ( .A(n_229), .B(n_288), .Y(n_306) );
OR2x2_ASAP7_75t_L g229 ( .A(n_230), .B(n_242), .Y(n_229) );
OAI322xp33_ASAP7_75t_L g271 ( .A1(n_230), .A2(n_272), .A3(n_276), .B1(n_278), .B2(n_281), .C1(n_286), .C2(n_294), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_230), .B(n_257), .Y(n_279) );
OR2x2_ASAP7_75t_L g289 ( .A(n_230), .B(n_243), .Y(n_289) );
AND2x2_ASAP7_75t_L g291 ( .A(n_230), .B(n_243), .Y(n_291) );
NOR2xp33_ASAP7_75t_L g292 ( .A(n_230), .B(n_293), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_230), .B(n_258), .Y(n_353) );
NOR2xp33_ASAP7_75t_L g386 ( .A(n_230), .B(n_387), .Y(n_386) );
INVx5_ASAP7_75t_SL g230 ( .A(n_231), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_231), .B(n_275), .Y(n_401) );
OAI21xp5_ASAP7_75t_L g232 ( .A1(n_233), .A2(n_234), .B(n_235), .Y(n_232) );
OAI21xp5_ASAP7_75t_L g463 ( .A1(n_234), .A2(n_464), .B(n_465), .Y(n_463) );
OAI21xp5_ASAP7_75t_L g495 ( .A1(n_234), .A2(n_496), .B(n_497), .Y(n_495) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_240), .B(n_241), .Y(n_239) );
INVx2_ASAP7_75t_L g519 ( .A(n_241), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_242), .B(n_257), .Y(n_256) );
AND2x2_ASAP7_75t_L g269 ( .A(n_242), .B(n_270), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_242), .B(n_320), .Y(n_319) );
OR2x2_ASAP7_75t_L g331 ( .A(n_242), .B(n_258), .Y(n_331) );
AOI211xp5_ASAP7_75t_SL g359 ( .A1(n_242), .A2(n_360), .B(n_363), .C(n_375), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_242), .B(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g397 ( .A(n_242), .B(n_372), .Y(n_397) );
INVx5_ASAP7_75t_SL g242 ( .A(n_243), .Y(n_242) );
AND2x2_ASAP7_75t_L g325 ( .A(n_243), .B(n_258), .Y(n_325) );
HB1xp67_ASAP7_75t_L g334 ( .A(n_243), .Y(n_334) );
AND2x2_ASAP7_75t_L g374 ( .A(n_243), .B(n_372), .Y(n_374) );
AND2x2_ASAP7_75t_SL g405 ( .A(n_243), .B(n_275), .Y(n_405) );
AND2x2_ASAP7_75t_L g412 ( .A(n_243), .B(n_371), .Y(n_412) );
OR2x6_ASAP7_75t_L g243 ( .A(n_244), .B(n_250), .Y(n_243) );
AOI22xp33_ASAP7_75t_L g251 ( .A1(n_252), .A2(n_253), .B1(n_267), .B2(n_269), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_252), .B(n_274), .Y(n_322) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
OR2x2_ASAP7_75t_L g254 ( .A(n_255), .B(n_256), .Y(n_254) );
INVx1_ASAP7_75t_L g270 ( .A(n_255), .Y(n_270) );
OR2x2_ASAP7_75t_L g330 ( .A(n_255), .B(n_331), .Y(n_330) );
OAI221xp5_ASAP7_75t_SL g378 ( .A1(n_255), .A2(n_379), .B1(n_381), .B2(n_382), .C(n_384), .Y(n_378) );
INVx2_ASAP7_75t_L g317 ( .A(n_256), .Y(n_317) );
AND2x2_ASAP7_75t_L g290 ( .A(n_257), .B(n_291), .Y(n_290) );
INVx1_ASAP7_75t_L g380 ( .A(n_257), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_257), .B(n_372), .Y(n_393) );
INVx3_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
INVxp67_ASAP7_75t_L g335 ( .A(n_258), .Y(n_335) );
AND2x2_ASAP7_75t_L g371 ( .A(n_258), .B(n_372), .Y(n_371) );
OA21x2_ASAP7_75t_L g258 ( .A1(n_259), .A2(n_260), .B(n_266), .Y(n_258) );
OA21x2_ASAP7_75t_L g443 ( .A1(n_259), .A2(n_444), .B(n_450), .Y(n_443) );
OA21x2_ASAP7_75t_L g472 ( .A1(n_259), .A2(n_473), .B(n_480), .Y(n_472) );
OA21x2_ASAP7_75t_L g485 ( .A1(n_259), .A2(n_486), .B(n_493), .Y(n_485) );
AND2x2_ASAP7_75t_L g373 ( .A(n_267), .B(n_312), .Y(n_373) );
AND2x2_ASAP7_75t_L g283 ( .A(n_268), .B(n_284), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_268), .B(n_341), .Y(n_340) );
NOR2xp33_ASAP7_75t_SL g354 ( .A(n_270), .B(n_317), .Y(n_354) );
INVx1_ASAP7_75t_SL g272 ( .A(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g360 ( .A(n_273), .B(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
OR2x2_ASAP7_75t_L g346 ( .A(n_274), .B(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g411 ( .A(n_274), .B(n_356), .Y(n_411) );
INVx2_ASAP7_75t_L g344 ( .A(n_275), .Y(n_344) );
NAND4xp25_ASAP7_75t_SL g407 ( .A(n_276), .B(n_408), .C(n_409), .D(n_410), .Y(n_407) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_277), .B(n_341), .Y(n_376) );
OR2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
INVx1_ASAP7_75t_SL g413 ( .A(n_280), .Y(n_413) );
O2A1O1Ixp33_ASAP7_75t_SL g375 ( .A1(n_281), .A2(n_344), .B(n_348), .C(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g370 ( .A(n_283), .B(n_362), .Y(n_370) );
HB1xp67_ASAP7_75t_L g296 ( .A(n_284), .Y(n_296) );
INVx1_ASAP7_75t_L g351 ( .A(n_284), .Y(n_351) );
INVx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
HB1xp67_ASAP7_75t_L g328 ( .A(n_285), .Y(n_328) );
AOI211xp5_ASAP7_75t_L g286 ( .A1(n_287), .A2(n_289), .B(n_290), .C(n_292), .Y(n_286) );
AND2x2_ASAP7_75t_L g307 ( .A(n_287), .B(n_291), .Y(n_307) );
OAI322xp33_ASAP7_75t_SL g345 ( .A1(n_287), .A2(n_346), .A3(n_348), .B1(n_349), .B2(n_353), .C1(n_354), .C2(n_355), .Y(n_345) );
INVx1_ASAP7_75t_SL g287 ( .A(n_288), .Y(n_287) );
OR2x2_ASAP7_75t_L g367 ( .A(n_289), .B(n_293), .Y(n_367) );
INVx1_ASAP7_75t_L g348 ( .A(n_291), .Y(n_348) );
INVx1_ASAP7_75t_SL g366 ( .A(n_293), .Y(n_366) );
INVx2_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
AOI222xp33_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_305), .B1(n_307), .B2(n_308), .C1(n_309), .C2(n_717), .Y(n_298) );
NAND2xp5_ASAP7_75t_SL g299 ( .A(n_300), .B(n_302), .Y(n_299) );
OAI322xp33_ASAP7_75t_L g388 ( .A1(n_300), .A2(n_362), .A3(n_367), .B1(n_389), .B2(n_390), .C1(n_392), .C2(n_393), .Y(n_388) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
AOI221xp5_ASAP7_75t_L g338 ( .A1(n_301), .A2(n_315), .B1(n_339), .B2(n_343), .C(n_345), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
INVx1_ASAP7_75t_SL g305 ( .A(n_306), .Y(n_305) );
OAI222xp33_ASAP7_75t_L g318 ( .A1(n_306), .A2(n_319), .B1(n_321), .B2(n_322), .C1(n_323), .C2(n_326), .Y(n_318) );
AOI22xp5_ASAP7_75t_L g384 ( .A1(n_308), .A2(n_315), .B1(n_385), .B2(n_386), .Y(n_384) );
AND2x2_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
AOI211xp5_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_315), .B(n_318), .C(n_329), .Y(n_313) );
O2A1O1Ixp33_ASAP7_75t_L g394 ( .A1(n_315), .A2(n_352), .B(n_395), .C(n_398), .Y(n_394) );
AND2x4_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
AND2x2_ASAP7_75t_L g324 ( .A(n_316), .B(n_325), .Y(n_324) );
INVx1_ASAP7_75t_SL g387 ( .A(n_320), .Y(n_387) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_327), .B(n_352), .Y(n_381) );
BUFx2_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
AOI21xp33_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_332), .B(n_336), .Y(n_329) );
OAI221xp5_ASAP7_75t_SL g398 ( .A1(n_330), .A2(n_399), .B1(n_400), .B2(n_401), .C(n_402), .Y(n_398) );
INVxp33_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
NOR2xp33_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
NOR2xp33_ASAP7_75t_L g343 ( .A(n_334), .B(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_341), .B(n_352), .Y(n_392) );
INVx2_ASAP7_75t_SL g341 ( .A(n_342), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_350), .B(n_352), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_356), .B(n_357), .Y(n_355) );
AND2x2_ASAP7_75t_L g403 ( .A(n_356), .B(n_362), .Y(n_403) );
AND4x1_ASAP7_75t_L g358 ( .A(n_359), .B(n_377), .C(n_394), .D(n_406), .Y(n_358) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
OAI221xp5_ASAP7_75t_SL g363 ( .A1(n_364), .A2(n_365), .B1(n_367), .B2(n_368), .C(n_369), .Y(n_363) );
AOI22xp5_ASAP7_75t_L g369 ( .A1(n_370), .A2(n_371), .B1(n_373), .B2(n_374), .Y(n_369) );
INVx1_ASAP7_75t_L g399 ( .A(n_370), .Y(n_399) );
INVx1_ASAP7_75t_SL g389 ( .A(n_374), .Y(n_389) );
NOR2xp33_ASAP7_75t_SL g377 ( .A(n_378), .B(n_388), .Y(n_377) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
NOR2xp33_ASAP7_75t_L g395 ( .A(n_390), .B(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
AOI22xp33_ASAP7_75t_L g402 ( .A1(n_397), .A2(n_403), .B1(n_404), .B2(n_405), .Y(n_402) );
AOI22xp5_ASAP7_75t_L g406 ( .A1(n_407), .A2(n_412), .B1(n_413), .B2(n_414), .Y(n_406) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
BUFx2_ASAP7_75t_L g427 ( .A(n_420), .Y(n_427) );
INVx2_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
AOI21xp33_ASAP7_75t_L g428 ( .A1(n_424), .A2(n_429), .B(n_712), .Y(n_428) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
BUFx2_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
AOI22xp5_ASAP7_75t_L g431 ( .A1(n_432), .A2(n_434), .B1(n_435), .B2(n_437), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx6_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g707 ( .A(n_436), .Y(n_707) );
BUFx2_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g708 ( .A(n_438), .Y(n_708) );
AND2x2_ASAP7_75t_L g438 ( .A(n_439), .B(n_624), .Y(n_438) );
NOR4xp25_ASAP7_75t_L g439 ( .A(n_440), .B(n_566), .C(n_596), .D(n_606), .Y(n_439) );
OAI211xp5_ASAP7_75t_L g440 ( .A1(n_441), .A2(n_481), .B(n_529), .C(n_556), .Y(n_440) );
OAI222xp33_ASAP7_75t_L g651 ( .A1(n_441), .A2(n_571), .B1(n_652), .B2(n_653), .C1(n_654), .C2(n_655), .Y(n_651) );
OR2x2_ASAP7_75t_L g441 ( .A(n_442), .B(n_460), .Y(n_441) );
AOI33xp33_ASAP7_75t_L g577 ( .A1(n_442), .A2(n_564), .A3(n_565), .B1(n_578), .B2(n_583), .B3(n_585), .Y(n_577) );
OAI211xp5_ASAP7_75t_SL g634 ( .A1(n_442), .A2(n_635), .B(n_637), .C(n_639), .Y(n_634) );
OR2x2_ASAP7_75t_L g650 ( .A(n_442), .B(n_636), .Y(n_650) );
INVx1_ASAP7_75t_L g683 ( .A(n_442), .Y(n_683) );
OR2x2_ASAP7_75t_L g442 ( .A(n_443), .B(n_451), .Y(n_442) );
INVx2_ASAP7_75t_L g560 ( .A(n_443), .Y(n_560) );
AND2x2_ASAP7_75t_L g576 ( .A(n_443), .B(n_472), .Y(n_576) );
HB1xp67_ASAP7_75t_L g611 ( .A(n_443), .Y(n_611) );
AND2x2_ASAP7_75t_L g640 ( .A(n_443), .B(n_451), .Y(n_640) );
INVx2_ASAP7_75t_L g540 ( .A(n_451), .Y(n_540) );
BUFx3_ASAP7_75t_L g548 ( .A(n_451), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_451), .B(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g559 ( .A(n_451), .B(n_560), .Y(n_559) );
NOR2xp33_ASAP7_75t_L g588 ( .A(n_451), .B(n_461), .Y(n_588) );
AND2x2_ASAP7_75t_L g657 ( .A(n_451), .B(n_591), .Y(n_657) );
INVx2_ASAP7_75t_SL g551 ( .A(n_460), .Y(n_551) );
OR2x2_ASAP7_75t_L g460 ( .A(n_461), .B(n_472), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_461), .B(n_540), .Y(n_539) );
INVx1_ASAP7_75t_L g593 ( .A(n_461), .Y(n_593) );
AND2x2_ASAP7_75t_L g604 ( .A(n_461), .B(n_560), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_461), .B(n_589), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_461), .B(n_591), .Y(n_636) );
AND2x2_ASAP7_75t_L g695 ( .A(n_461), .B(n_640), .Y(n_695) );
INVx4_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
AND2x2_ASAP7_75t_L g565 ( .A(n_462), .B(n_472), .Y(n_565) );
AND2x2_ASAP7_75t_L g575 ( .A(n_462), .B(n_576), .Y(n_575) );
BUFx3_ASAP7_75t_L g597 ( .A(n_462), .Y(n_597) );
AND3x2_ASAP7_75t_L g656 ( .A(n_462), .B(n_657), .C(n_658), .Y(n_656) );
HB1xp67_ASAP7_75t_L g547 ( .A(n_472), .Y(n_547) );
INVx1_ASAP7_75t_SL g591 ( .A(n_472), .Y(n_591) );
NAND3xp33_ASAP7_75t_L g603 ( .A(n_472), .B(n_540), .C(n_604), .Y(n_603) );
NOR2xp33_ASAP7_75t_L g481 ( .A(n_482), .B(n_512), .Y(n_481) );
A2O1A1Ixp33_ASAP7_75t_L g626 ( .A1(n_482), .A2(n_575), .B(n_627), .C(n_629), .Y(n_626) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
NAND2xp5_ASAP7_75t_SL g483 ( .A(n_484), .B(n_503), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_484), .B(n_633), .Y(n_632) );
INVx2_ASAP7_75t_SL g643 ( .A(n_484), .Y(n_643) );
AND2x2_ASAP7_75t_L g664 ( .A(n_484), .B(n_514), .Y(n_664) );
NOR2xp33_ASAP7_75t_L g692 ( .A(n_484), .B(n_573), .Y(n_692) );
AND2x2_ASAP7_75t_L g484 ( .A(n_485), .B(n_494), .Y(n_484) );
AND2x2_ASAP7_75t_L g537 ( .A(n_485), .B(n_528), .Y(n_537) );
INVx2_ASAP7_75t_L g544 ( .A(n_485), .Y(n_544) );
AND2x2_ASAP7_75t_L g564 ( .A(n_485), .B(n_514), .Y(n_564) );
AND2x2_ASAP7_75t_L g614 ( .A(n_485), .B(n_503), .Y(n_614) );
INVx1_ASAP7_75t_L g618 ( .A(n_485), .Y(n_618) );
INVx2_ASAP7_75t_SL g528 ( .A(n_494), .Y(n_528) );
BUFx2_ASAP7_75t_L g554 ( .A(n_494), .Y(n_554) );
AND2x2_ASAP7_75t_L g681 ( .A(n_494), .B(n_503), .Y(n_681) );
INVx3_ASAP7_75t_SL g514 ( .A(n_503), .Y(n_514) );
AND2x2_ASAP7_75t_L g536 ( .A(n_503), .B(n_537), .Y(n_536) );
AND2x4_ASAP7_75t_L g543 ( .A(n_503), .B(n_544), .Y(n_543) );
OR2x2_ASAP7_75t_L g573 ( .A(n_503), .B(n_533), .Y(n_573) );
OR2x2_ASAP7_75t_L g582 ( .A(n_503), .B(n_528), .Y(n_582) );
HB1xp67_ASAP7_75t_L g600 ( .A(n_503), .Y(n_600) );
AND2x2_ASAP7_75t_L g605 ( .A(n_503), .B(n_558), .Y(n_605) );
AND2x2_ASAP7_75t_L g633 ( .A(n_503), .B(n_516), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_503), .B(n_669), .Y(n_668) );
OR2x2_ASAP7_75t_L g671 ( .A(n_503), .B(n_515), .Y(n_671) );
OR2x6_ASAP7_75t_L g503 ( .A(n_504), .B(n_510), .Y(n_503) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
OR2x2_ASAP7_75t_L g513 ( .A(n_514), .B(n_515), .Y(n_513) );
AND2x2_ASAP7_75t_L g595 ( .A(n_514), .B(n_544), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_514), .B(n_537), .Y(n_623) );
AND2x2_ASAP7_75t_L g641 ( .A(n_514), .B(n_558), .Y(n_641) );
OR2x2_ASAP7_75t_L g515 ( .A(n_516), .B(n_528), .Y(n_515) );
AND2x2_ASAP7_75t_L g542 ( .A(n_516), .B(n_528), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_516), .B(n_571), .Y(n_570) );
BUFx3_ASAP7_75t_L g580 ( .A(n_516), .Y(n_580) );
OR2x2_ASAP7_75t_L g628 ( .A(n_516), .B(n_548), .Y(n_628) );
OA21x2_ASAP7_75t_L g516 ( .A1(n_517), .A2(n_520), .B(n_527), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
AO21x2_ASAP7_75t_L g533 ( .A1(n_518), .A2(n_534), .B(n_535), .Y(n_533) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g534 ( .A(n_520), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_527), .Y(n_535) );
AND2x2_ASAP7_75t_L g563 ( .A(n_528), .B(n_533), .Y(n_563) );
INVx1_ASAP7_75t_L g571 ( .A(n_528), .Y(n_571) );
AND2x2_ASAP7_75t_L g666 ( .A(n_528), .B(n_544), .Y(n_666) );
AOI222xp33_ASAP7_75t_L g529 ( .A1(n_530), .A2(n_538), .B1(n_541), .B2(n_545), .C1(n_549), .C2(n_552), .Y(n_529) );
INVx1_ASAP7_75t_L g661 ( .A(n_530), .Y(n_661) );
AND2x2_ASAP7_75t_L g530 ( .A(n_531), .B(n_536), .Y(n_530) );
AND2x2_ASAP7_75t_L g557 ( .A(n_531), .B(n_558), .Y(n_557) );
AND2x2_ASAP7_75t_L g568 ( .A(n_531), .B(n_537), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_531), .B(n_559), .Y(n_584) );
OAI222xp33_ASAP7_75t_L g606 ( .A1(n_531), .A2(n_607), .B1(n_612), .B2(n_613), .C1(n_621), .C2(n_623), .Y(n_606) );
INVx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx1_ASAP7_75t_SL g532 ( .A(n_533), .Y(n_532) );
AND2x2_ASAP7_75t_L g594 ( .A(n_533), .B(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_533), .B(n_614), .Y(n_654) );
AND2x2_ASAP7_75t_L g665 ( .A(n_533), .B(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g673 ( .A(n_536), .Y(n_673) );
NAND2xp5_ASAP7_75t_SL g652 ( .A(n_538), .B(n_589), .Y(n_652) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
NOR2xp33_ASAP7_75t_L g592 ( .A(n_540), .B(n_593), .Y(n_592) );
AND2x2_ASAP7_75t_L g610 ( .A(n_540), .B(n_611), .Y(n_610) );
AND2x2_ASAP7_75t_L g541 ( .A(n_542), .B(n_543), .Y(n_541) );
INVx3_ASAP7_75t_L g555 ( .A(n_543), .Y(n_555) );
O2A1O1Ixp33_ASAP7_75t_L g645 ( .A1(n_543), .A2(n_646), .B(n_649), .C(n_651), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_543), .B(n_580), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_543), .B(n_563), .Y(n_685) );
AND2x2_ASAP7_75t_L g558 ( .A(n_544), .B(n_554), .Y(n_558) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_547), .B(n_548), .Y(n_546) );
INVx1_ASAP7_75t_L g585 ( .A(n_547), .Y(n_585) );
NAND2xp5_ASAP7_75t_SL g574 ( .A(n_548), .B(n_575), .Y(n_574) );
OR2x2_ASAP7_75t_L g637 ( .A(n_548), .B(n_638), .Y(n_637) );
AND2x2_ASAP7_75t_L g676 ( .A(n_548), .B(n_576), .Y(n_676) );
INVx1_ASAP7_75t_L g688 ( .A(n_548), .Y(n_688) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_551), .B(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
OR2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_555), .Y(n_553) );
INVx1_ASAP7_75t_L g669 ( .A(n_554), .Y(n_669) );
A2O1A1Ixp33_ASAP7_75t_SL g556 ( .A1(n_557), .A2(n_559), .B(n_561), .C(n_565), .Y(n_556) );
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_557), .A2(n_587), .B1(n_602), .B2(n_605), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_558), .B(n_572), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_558), .B(n_580), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_559), .B(n_617), .Y(n_616) );
INVx1_ASAP7_75t_SL g622 ( .A(n_559), .Y(n_622) );
AND2x2_ASAP7_75t_L g629 ( .A(n_559), .B(n_609), .Y(n_629) );
INVx2_ASAP7_75t_L g590 ( .A(n_560), .Y(n_590) );
INVxp67_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_563), .B(n_564), .Y(n_562) );
NOR4xp25_ASAP7_75t_L g567 ( .A(n_564), .B(n_568), .C(n_569), .D(n_572), .Y(n_567) );
INVx1_ASAP7_75t_SL g638 ( .A(n_565), .Y(n_638) );
AND2x2_ASAP7_75t_L g682 ( .A(n_565), .B(n_683), .Y(n_682) );
OAI211xp5_ASAP7_75t_SL g566 ( .A1(n_567), .A2(n_574), .B(n_577), .C(n_586), .Y(n_566) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx1_ASAP7_75t_SL g572 ( .A(n_573), .Y(n_572) );
NOR2xp33_ASAP7_75t_L g694 ( .A(n_573), .B(n_643), .Y(n_694) );
AOI22xp5_ASAP7_75t_L g693 ( .A1(n_575), .A2(n_694), .B1(n_695), .B2(n_696), .Y(n_693) );
INVx1_ASAP7_75t_SL g648 ( .A(n_576), .Y(n_648) );
AND2x2_ASAP7_75t_L g687 ( .A(n_576), .B(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_580), .B(n_581), .Y(n_579) );
NAND2xp5_ASAP7_75t_SL g680 ( .A(n_580), .B(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
NOR2xp33_ASAP7_75t_L g599 ( .A(n_584), .B(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_585), .B(n_610), .Y(n_670) );
OAI21xp5_ASAP7_75t_SL g586 ( .A1(n_587), .A2(n_592), .B(n_594), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_588), .B(n_589), .Y(n_587) );
INVx1_ASAP7_75t_L g662 ( .A(n_589), .Y(n_662) );
AND2x2_ASAP7_75t_L g589 ( .A(n_590), .B(n_591), .Y(n_589) );
INVx2_ASAP7_75t_L g690 ( .A(n_590), .Y(n_690) );
HB1xp67_ASAP7_75t_L g617 ( .A(n_591), .Y(n_617) );
OAI21xp33_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_598), .B(n_601), .Y(n_596) );
CKINVDCx16_ASAP7_75t_R g609 ( .A(n_597), .Y(n_609) );
OR2x2_ASAP7_75t_L g647 ( .A(n_597), .B(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
AOI21xp33_ASAP7_75t_SL g642 ( .A1(n_600), .A2(n_643), .B(n_644), .Y(n_642) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
AOI221xp5_ASAP7_75t_L g630 ( .A1(n_604), .A2(n_631), .B1(n_634), .B2(n_641), .C(n_642), .Y(n_630) );
INVx1_ASAP7_75t_SL g674 ( .A(n_605), .Y(n_674) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
AND2x2_ASAP7_75t_L g608 ( .A(n_609), .B(n_610), .Y(n_608) );
OR2x2_ASAP7_75t_L g621 ( .A(n_609), .B(n_622), .Y(n_621) );
INVxp67_ASAP7_75t_L g658 ( .A(n_611), .Y(n_658) );
AOI22xp5_ASAP7_75t_L g613 ( .A1(n_614), .A2(n_615), .B1(n_618), .B2(n_619), .Y(n_613) );
INVx1_ASAP7_75t_L g653 ( .A(n_614), .Y(n_653) );
INVxp67_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_617), .B(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
NOR4xp25_ASAP7_75t_L g624 ( .A(n_625), .B(n_659), .C(n_672), .D(n_684), .Y(n_624) );
NAND3xp33_ASAP7_75t_SL g625 ( .A(n_626), .B(n_630), .C(n_645), .Y(n_625) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
NOR2xp33_ASAP7_75t_L g646 ( .A(n_628), .B(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_635), .B(n_640), .Y(n_644) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
OAI221xp5_ASAP7_75t_SL g672 ( .A1(n_647), .A2(n_673), .B1(n_674), .B2(n_675), .C(n_677), .Y(n_672) );
O2A1O1Ixp33_ASAP7_75t_L g663 ( .A1(n_649), .A2(n_664), .B(n_665), .C(n_667), .Y(n_663) );
INVx2_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
OAI22xp5_ASAP7_75t_L g667 ( .A1(n_650), .A2(n_668), .B1(n_670), .B2(n_671), .Y(n_667) );
INVx2_ASAP7_75t_SL g655 ( .A(n_656), .Y(n_655) );
A2O1A1Ixp33_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_661), .B(n_662), .C(n_663), .Y(n_659) );
INVx1_ASAP7_75t_L g678 ( .A(n_671), .Y(n_678) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
OAI21xp5_ASAP7_75t_SL g677 ( .A1(n_678), .A2(n_679), .B(n_682), .Y(n_677) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
OAI221xp5_ASAP7_75t_SL g684 ( .A1(n_685), .A2(n_686), .B1(n_689), .B2(n_691), .C(n_693), .Y(n_684) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVxp67_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
CKINVDCx20_ASAP7_75t_R g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_SL g709 ( .A(n_710), .Y(n_709) );
INVx3_ASAP7_75t_SL g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_SL g712 ( .A(n_713), .Y(n_712) );
BUFx2_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
endmodule