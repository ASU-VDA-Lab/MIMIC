module fake_jpeg_17529_n_37 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_37);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_37;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_36;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_32;
wire n_15;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVx4_ASAP7_75t_SL g14 ( 
.A(n_6),
.Y(n_14)
);

INVx5_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_10),
.B(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_15),
.A2(n_12),
.B(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_16),
.B(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_15),
.A2(n_8),
.B1(n_7),
.B2(n_2),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_21),
.B(n_13),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_22),
.A2(n_21),
.B1(n_17),
.B2(n_2),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_18),
.B(n_13),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_3),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_27),
.A2(n_25),
.B1(n_5),
.B2(n_4),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_24),
.B(n_0),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_L g31 ( 
.A1(n_28),
.A2(n_29),
.B(n_30),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_26),
.B(n_1),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_27),
.A2(n_23),
.B1(n_14),
.B2(n_22),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_32),
.B(n_33),
.Y(n_35)
);

NOR2xp67_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_26),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_34),
.B(n_14),
.C(n_4),
.Y(n_36)
);

XOR2xp5_ASAP7_75t_L g37 ( 
.A(n_36),
.B(n_35),
.Y(n_37)
);


endmodule