module fake_jpeg_4805_n_332 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_332);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_332;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_20),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_38),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_16),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_37),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_27),
.B(n_15),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_42),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_45),
.Y(n_53)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_18),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_47),
.Y(n_94)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_27),
.Y(n_55)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

BUFx10_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_58),
.B(n_60),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_27),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_59),
.B(n_38),
.Y(n_77)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_44),
.A2(n_25),
.B1(n_19),
.B2(n_31),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_61),
.A2(n_25),
.B1(n_24),
.B2(n_33),
.Y(n_84)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_67),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_37),
.B(n_23),
.C(n_31),
.Y(n_68)
);

FAx1_ASAP7_75t_SL g74 ( 
.A(n_68),
.B(n_36),
.CI(n_37),
.CON(n_74),
.SN(n_74)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_70),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_56),
.A2(n_19),
.B1(n_43),
.B2(n_42),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_71),
.A2(n_87),
.B1(n_96),
.B2(n_98),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_74),
.B(n_90),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_77),
.B(n_93),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_52),
.A2(n_19),
.B1(n_25),
.B2(n_43),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_83),
.A2(n_86),
.B1(n_89),
.B2(n_92),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_84),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_52),
.A2(n_56),
.B1(n_60),
.B2(n_66),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_65),
.A2(n_42),
.B1(n_35),
.B2(n_28),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_53),
.A2(n_36),
.B1(n_39),
.B2(n_41),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_48),
.B(n_20),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_67),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_91),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_50),
.A2(n_21),
.B1(n_23),
.B2(n_22),
.Y(n_92)
);

A2O1A1Ixp33_ASAP7_75t_L g93 ( 
.A1(n_68),
.A2(n_22),
.B(n_32),
.C(n_28),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_58),
.A2(n_28),
.B1(n_35),
.B2(n_20),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_51),
.A2(n_21),
.B1(n_30),
.B2(n_33),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_97),
.A2(n_99),
.B1(n_24),
.B2(n_62),
.Y(n_115)
);

O2A1O1Ixp33_ASAP7_75t_SL g98 ( 
.A1(n_57),
.A2(n_41),
.B(n_35),
.C(n_26),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_51),
.A2(n_41),
.B1(n_32),
.B2(n_33),
.Y(n_99)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_101),
.B(n_103),
.Y(n_152)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_96),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_74),
.B(n_64),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_104),
.B(n_120),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_78),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_105),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_78),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_106),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_86),
.B(n_57),
.C(n_47),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_107),
.B(n_113),
.C(n_122),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_93),
.B(n_30),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_108),
.B(n_111),
.Y(n_135)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_94),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_109),
.B(n_110),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_71),
.B(n_57),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_30),
.Y(n_111)
);

INVx1_ASAP7_75t_SL g112 ( 
.A(n_94),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g137 ( 
.A(n_112),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_83),
.B(n_47),
.C(n_64),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_115),
.A2(n_84),
.B1(n_98),
.B2(n_99),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_85),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_116),
.B(n_119),
.Y(n_158)
);

OR2x2_ASAP7_75t_L g117 ( 
.A(n_85),
.B(n_63),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_117),
.A2(n_75),
.B(n_94),
.Y(n_150)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_87),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_74),
.B(n_64),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_89),
.B(n_47),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_121),
.B(n_125),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_73),
.B(n_49),
.C(n_69),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_81),
.B(n_29),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_81),
.B(n_29),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_126),
.B(n_127),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_77),
.B(n_29),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_124),
.A2(n_76),
.B1(n_72),
.B2(n_95),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_128),
.Y(n_163)
);

AO21x2_ASAP7_75t_L g129 ( 
.A1(n_110),
.A2(n_98),
.B(n_49),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_L g180 ( 
.A1(n_129),
.A2(n_110),
.B1(n_107),
.B2(n_117),
.Y(n_180)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_115),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_130),
.B(n_136),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_131),
.A2(n_132),
.B1(n_139),
.B2(n_147),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_124),
.A2(n_73),
.B1(n_62),
.B2(n_79),
.Y(n_132)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_115),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_118),
.A2(n_79),
.B1(n_95),
.B2(n_80),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_104),
.B(n_90),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_140),
.B(n_127),
.C(n_102),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_102),
.B(n_82),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_141),
.B(n_143),
.Y(n_164)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_123),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_142),
.B(n_144),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_105),
.Y(n_143)
);

BUFx2_ASAP7_75t_L g144 ( 
.A(n_101),
.Y(n_144)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_101),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_145),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_123),
.A2(n_88),
.B1(n_72),
.B2(n_76),
.Y(n_147)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_114),
.Y(n_148)
);

INVx1_ASAP7_75t_SL g176 ( 
.A(n_148),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_123),
.A2(n_80),
.B1(n_49),
.B2(n_82),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_149),
.A2(n_110),
.B1(n_113),
.B2(n_121),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_150),
.A2(n_111),
.B(n_125),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_106),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_151),
.B(n_108),
.Y(n_170)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_122),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_154),
.B(n_155),
.Y(n_177)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_122),
.Y(n_155)
);

XNOR2x1_ASAP7_75t_L g159 ( 
.A(n_134),
.B(n_120),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g214 ( 
.A(n_159),
.B(n_185),
.Y(n_214)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_152),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_160),
.B(n_162),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_157),
.B(n_100),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_161),
.B(n_175),
.Y(n_193)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_144),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_133),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_165),
.Y(n_192)
);

INVx2_ASAP7_75t_SL g167 ( 
.A(n_145),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_167),
.B(n_183),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_134),
.B(n_100),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_168),
.B(n_153),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_170),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_171),
.A2(n_180),
.B1(n_188),
.B2(n_131),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_172),
.B(n_150),
.C(n_130),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_174),
.A2(n_146),
.B(n_29),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_157),
.B(n_103),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_156),
.B(n_140),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_178),
.B(n_179),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_156),
.B(n_119),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_129),
.A2(n_107),
.B(n_113),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_181),
.A2(n_0),
.B(n_1),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_158),
.B(n_126),
.Y(n_182)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_182),
.Y(n_199)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_139),
.Y(n_183)
);

A2O1A1O1Ixp25_ASAP7_75t_L g185 ( 
.A1(n_129),
.A2(n_118),
.B(n_117),
.C(n_112),
.D(n_109),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_148),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_186),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_138),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_187),
.B(n_189),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_142),
.A2(n_129),
.B1(n_149),
.B2(n_136),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_132),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_135),
.B(n_155),
.Y(n_190)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_190),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_154),
.B(n_112),
.Y(n_191)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_191),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_159),
.A2(n_129),
.B(n_153),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_194),
.B(n_195),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_198),
.B(n_215),
.C(n_216),
.Y(n_229)
);

INVxp33_ASAP7_75t_L g200 ( 
.A(n_173),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_200),
.B(n_211),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_201),
.A2(n_205),
.B1(n_209),
.B2(n_212),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_188),
.A2(n_146),
.B1(n_137),
.B2(n_24),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_181),
.A2(n_146),
.B1(n_109),
.B2(n_70),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_206),
.A2(n_207),
.B1(n_171),
.B2(n_163),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_189),
.A2(n_183),
.B1(n_166),
.B2(n_177),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_208),
.B(n_160),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_169),
.A2(n_70),
.B1(n_26),
.B2(n_18),
.Y(n_209)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_164),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_174),
.A2(n_17),
.B(n_26),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_169),
.A2(n_26),
.B1(n_17),
.B2(n_2),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_213),
.A2(n_163),
.B1(n_187),
.B2(n_165),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_178),
.B(n_15),
.Y(n_215)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_191),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_217),
.B(n_220),
.Y(n_225)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_185),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_203),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_221),
.B(n_231),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_223),
.A2(n_192),
.B(n_202),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_219),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_224),
.B(n_230),
.Y(n_259)
);

OAI21xp33_ASAP7_75t_L g227 ( 
.A1(n_206),
.A2(n_179),
.B(n_175),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_227),
.B(n_195),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_210),
.B(n_168),
.Y(n_228)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_228),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_207),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_218),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_232),
.A2(n_241),
.B1(n_242),
.B2(n_243),
.Y(n_255)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_218),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_233),
.B(n_236),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_234),
.A2(n_235),
.B1(n_199),
.B2(n_193),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_220),
.A2(n_180),
.B1(n_161),
.B2(n_172),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_205),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_194),
.B(n_184),
.C(n_167),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_237),
.B(n_244),
.C(n_216),
.Y(n_250)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_213),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_238),
.B(n_240),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_210),
.B(n_186),
.Y(n_239)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_239),
.Y(n_249)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_209),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_201),
.A2(n_167),
.B1(n_162),
.B2(n_176),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_212),
.A2(n_176),
.B1(n_1),
.B2(n_2),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_198),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_204),
.B(n_3),
.C(n_4),
.Y(n_244)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_200),
.Y(n_246)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_246),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_223),
.A2(n_208),
.B(n_214),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_248),
.A2(n_256),
.B1(n_264),
.B2(n_265),
.Y(n_278)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_250),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_245),
.B(n_214),
.C(n_204),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_251),
.B(n_261),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_252),
.B(n_263),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_241),
.Y(n_253)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_253),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_226),
.B(n_211),
.Y(n_262)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_262),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_245),
.B(n_193),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_234),
.A2(n_196),
.B1(n_197),
.B2(n_215),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_230),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_237),
.B(n_5),
.C(n_6),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_266),
.B(n_267),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_235),
.B(n_228),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_253),
.A2(n_259),
.B1(n_255),
.B2(n_249),
.Y(n_270)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_270),
.Y(n_292)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_258),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_272),
.B(n_273),
.Y(n_294)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_259),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_264),
.B(n_244),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_274),
.B(n_279),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_260),
.A2(n_254),
.B1(n_225),
.B2(n_246),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_275),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_256),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_276),
.B(n_280),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_257),
.B(n_265),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_261),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_266),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_281),
.B(n_282),
.Y(n_287)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_250),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_269),
.B(n_263),
.C(n_251),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_285),
.B(n_289),
.C(n_298),
.Y(n_310)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_272),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_286),
.B(n_271),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_277),
.B(n_247),
.Y(n_288)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_288),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_284),
.B(n_252),
.C(n_267),
.Y(n_289)
);

AO221x1_ASAP7_75t_L g290 ( 
.A1(n_271),
.A2(n_224),
.B1(n_239),
.B2(n_232),
.C(n_222),
.Y(n_290)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_290),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_283),
.B(n_248),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_291),
.B(n_297),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_283),
.B(n_229),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_284),
.B(n_229),
.C(n_222),
.Y(n_298)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_299),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_293),
.B(n_278),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_300),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_287),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_301),
.B(n_304),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_293),
.A2(n_273),
.B(n_270),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_302),
.A2(n_305),
.B1(n_307),
.B2(n_242),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_298),
.B(n_275),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_285),
.B(n_243),
.Y(n_305)
);

OR2x2_ASAP7_75t_L g307 ( 
.A(n_292),
.B(n_295),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_294),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_308),
.A2(n_13),
.B(n_14),
.Y(n_318)
);

O2A1O1Ixp33_ASAP7_75t_SL g324 ( 
.A1(n_311),
.A2(n_309),
.B(n_310),
.C(n_6),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_309),
.B(n_297),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_312),
.B(n_310),
.Y(n_322)
);

AOI322xp5_ASAP7_75t_L g314 ( 
.A1(n_306),
.A2(n_296),
.A3(n_289),
.B1(n_268),
.B2(n_8),
.C1(n_11),
.C2(n_12),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_314),
.A2(n_317),
.B(n_301),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_303),
.A2(n_268),
.B1(n_12),
.B2(n_13),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_316),
.B(n_5),
.Y(n_321)
);

AOI322xp5_ASAP7_75t_L g317 ( 
.A1(n_307),
.A2(n_11),
.A3(n_14),
.B1(n_13),
.B2(n_8),
.C1(n_15),
.C2(n_7),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_318),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_320),
.B(n_321),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_322),
.A2(n_323),
.B(n_324),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_313),
.A2(n_6),
.B1(n_7),
.B2(n_319),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_325),
.A2(n_315),
.B(n_317),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_328),
.A2(n_314),
.B(n_323),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_326),
.Y(n_330)
);

XNOR2x2_ASAP7_75t_SL g331 ( 
.A(n_330),
.B(n_327),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_7),
.Y(n_332)
);


endmodule