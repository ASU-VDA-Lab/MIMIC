module real_jpeg_16762_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_578;
wire n_366;
wire n_149;
wire n_332;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_216;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_516;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_572;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_531;
wire n_285;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_568;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx5_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_0),
.B(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_1),
.B(n_203),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_1),
.B(n_206),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_1),
.B(n_306),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_1),
.B(n_328),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_1),
.B(n_366),
.Y(n_365)
);

AND2x2_ASAP7_75t_L g475 ( 
.A(n_1),
.B(n_476),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_1),
.B(n_479),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_1),
.B(n_496),
.Y(n_495)
);

BUFx5_ASAP7_75t_L g170 ( 
.A(n_2),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g252 ( 
.A(n_2),
.Y(n_252)
);

BUFx5_ASAP7_75t_L g299 ( 
.A(n_2),
.Y(n_299)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_2),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_3),
.Y(n_81)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_3),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g236 ( 
.A(n_3),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_4),
.B(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_4),
.B(n_39),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_4),
.B(n_92),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_4),
.B(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_4),
.B(n_238),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_4),
.B(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_4),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_4),
.B(n_170),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_5),
.B(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_5),
.B(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_5),
.B(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_5),
.B(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_5),
.B(n_156),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_5),
.B(n_254),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_5),
.B(n_259),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_5),
.A2(n_15),
.B1(n_297),
.B2(n_300),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g414 ( 
.A(n_5),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_6),
.B(n_66),
.Y(n_65)
);

INVxp33_ASAP7_75t_L g105 ( 
.A(n_6),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_6),
.B(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_6),
.B(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_6),
.B(n_201),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_6),
.B(n_308),
.Y(n_307)
);

AND2x4_ASAP7_75t_SL g325 ( 
.A(n_6),
.B(n_326),
.Y(n_325)
);

AND2x2_ASAP7_75t_SL g363 ( 
.A(n_6),
.B(n_170),
.Y(n_363)
);

BUFx5_ASAP7_75t_L g112 ( 
.A(n_7),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_7),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_7),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_7),
.Y(n_315)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_7),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_8),
.A2(n_20),
.B(n_22),
.Y(n_19)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_9),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g219 ( 
.A(n_9),
.Y(n_219)
);

BUFx4f_ASAP7_75t_L g256 ( 
.A(n_9),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_9),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_10),
.B(n_31),
.Y(n_30)
);

AND2x2_ASAP7_75t_SL g34 ( 
.A(n_10),
.B(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_10),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_10),
.B(n_71),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_10),
.B(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_10),
.B(n_574),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_11),
.B(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_11),
.B(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_11),
.B(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_11),
.B(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_11),
.B(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_11),
.B(n_161),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_11),
.B(n_217),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_11),
.B(n_250),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_12),
.Y(n_100)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_12),
.Y(n_151)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_12),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_13),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_13),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_13),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_13),
.Y(n_201)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_13),
.Y(n_323)
);

BUFx5_ASAP7_75t_L g510 ( 
.A(n_13),
.Y(n_510)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_14),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_14),
.B(n_63),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_14),
.B(n_242),
.Y(n_241)
);

AND2x2_ASAP7_75t_SL g264 ( 
.A(n_14),
.B(n_265),
.Y(n_264)
);

AND2x4_ASAP7_75t_SL g320 ( 
.A(n_14),
.B(n_321),
.Y(n_320)
);

AND2x4_ASAP7_75t_L g369 ( 
.A(n_14),
.B(n_370),
.Y(n_369)
);

AND2x4_ASAP7_75t_SL g422 ( 
.A(n_14),
.B(n_423),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_14),
.B(n_482),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_15),
.B(n_214),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_15),
.B(n_234),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g373 ( 
.A(n_15),
.B(n_374),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_15),
.B(n_407),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_15),
.B(n_450),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_15),
.B(n_259),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g471 ( 
.A(n_15),
.B(n_472),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_15),
.B(n_516),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_16),
.B(n_317),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_16),
.B(n_428),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_16),
.B(n_447),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_16),
.B(n_465),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_16),
.B(n_509),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_16),
.B(n_524),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_16),
.B(n_531),
.Y(n_530)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_17),
.Y(n_86)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_18),
.Y(n_63)
);

BUFx8_ASAP7_75t_L g68 ( 
.A(n_18),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g207 ( 
.A(n_18),
.Y(n_207)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_18),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

O2A1O1Ixp33_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_569),
.B(n_576),
.C(n_578),
.Y(n_23)
);

OAI21x1_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_120),
.B(n_568),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_74),
.Y(n_26)
);

OR2x2_ASAP7_75t_L g568 ( 
.A(n_27),
.B(n_74),
.Y(n_568)
);

XOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_55),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_42),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g577 ( 
.A(n_29),
.B(n_42),
.C(n_55),
.Y(n_577)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_34),
.C(n_38),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_30),
.A2(n_44),
.B1(n_49),
.B2(n_50),
.Y(n_43)
);

INVx1_ASAP7_75t_SL g49 ( 
.A(n_30),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_30),
.A2(n_34),
.B1(n_49),
.B2(n_59),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_SL g571 ( 
.A(n_30),
.B(n_44),
.C(n_51),
.Y(n_571)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_32),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_33),
.Y(n_94)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_33),
.Y(n_303)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_34),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_34),
.B(n_65),
.C(n_69),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_34),
.A2(n_59),
.B1(n_69),
.B2(n_70),
.Y(n_115)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_37),
.Y(n_159)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_37),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_41),
.Y(n_204)
);

INVx4_ASAP7_75t_L g429 ( 
.A(n_41),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_51),
.Y(n_42)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g572 ( 
.A1(n_44),
.A2(n_50),
.B1(n_573),
.B2(n_576),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_45),
.B(n_48),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

OR2x2_ASAP7_75t_SL g110 ( 
.A(n_48),
.B(n_111),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_48),
.B(n_132),
.Y(n_131)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_60),
.C(n_64),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_56),
.A2(n_57),
.B1(n_118),
.B2(n_119),
.Y(n_117)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_SL g119 ( 
.A(n_60),
.B(n_64),
.Y(n_119)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_65),
.B(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_68),
.Y(n_102)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_68),
.Y(n_575)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_69),
.A2(n_70),
.B1(n_110),
.B2(n_129),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_70),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_SL g103 ( 
.A(n_70),
.B(n_104),
.C(n_110),
.Y(n_103)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_116),
.C(n_117),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_75),
.B(n_186),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_103),
.C(n_113),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_76),
.B(n_184),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_87),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_82),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_78),
.B(n_82),
.C(n_87),
.Y(n_116)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_86),
.Y(n_266)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_86),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_95),
.C(n_101),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_88),
.A2(n_89),
.B1(n_95),
.B2(n_96),
.Y(n_165)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx4_ASAP7_75t_L g331 ( 
.A(n_94),
.Y(n_331)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx5_ASAP7_75t_L g306 ( 
.A(n_100),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_101),
.B(n_165),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_103),
.B(n_114),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g178 ( 
.A(n_104),
.B(n_179),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_109),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_110),
.A2(n_129),
.B1(n_130),
.B2(n_131),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g129 ( 
.A(n_110),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_110),
.B(n_130),
.C(n_135),
.Y(n_180)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_116),
.B(n_117),
.Y(n_186)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

AOI21x1_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_286),
.B(n_563),
.Y(n_120)
);

NOR3x1_ASAP7_75t_SL g121 ( 
.A(n_122),
.B(n_187),
.C(n_280),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g563 ( 
.A1(n_122),
.A2(n_564),
.B(n_567),
.Y(n_563)
);

NOR2xp67_ASAP7_75t_R g122 ( 
.A(n_123),
.B(n_185),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_123),
.B(n_185),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_177),
.C(n_182),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_124),
.B(n_283),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_163),
.C(n_166),
.Y(n_124)
);

INVxp33_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_126),
.B(n_277),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_138),
.C(n_152),
.Y(n_126)
);

XNOR2x2_ASAP7_75t_SL g225 ( 
.A(n_127),
.B(n_226),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_SL g127 ( 
.A(n_128),
.B(n_135),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_130),
.A2(n_131),
.B1(n_169),
.B2(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

MAJx2_ASAP7_75t_L g168 ( 
.A(n_131),
.B(n_169),
.C(n_171),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_134),
.Y(n_424)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_138),
.B(n_152),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_143),
.C(n_147),
.Y(n_138)
);

XNOR2x1_ASAP7_75t_L g211 ( 
.A(n_139),
.B(n_147),
.Y(n_211)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx4_ASAP7_75t_L g368 ( 
.A(n_141),
.Y(n_368)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_142),
.Y(n_451)
);

XNOR2x1_ASAP7_75t_L g210 ( 
.A(n_143),
.B(n_211),
.Y(n_210)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_145),
.Y(n_326)
);

INVx8_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_154),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_153),
.B(n_155),
.C(n_160),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_160),
.Y(n_154)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_164),
.B(n_166),
.Y(n_277)
);

MAJx2_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_175),
.C(n_176),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_167),
.A2(n_168),
.B1(n_192),
.B2(n_194),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_168),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_169),
.B(n_213),
.C(n_215),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_169),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_169),
.A2(n_216),
.B1(n_224),
.B2(n_231),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_171),
.A2(n_221),
.B1(n_222),
.B2(n_223),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_171),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_171),
.A2(n_221),
.B1(n_307),
.B2(n_358),
.Y(n_357)
);

OR2x2_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

INVx6_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_175),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_175),
.B(n_249),
.C(n_253),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_175),
.B(n_294),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_176),
.B(n_193),
.Y(n_192)
);

INVx2_ASAP7_75t_SL g208 ( 
.A(n_176),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_176),
.A2(n_205),
.B1(n_208),
.B2(n_269),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_177),
.B(n_183),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_180),
.C(n_181),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_178),
.B(n_275),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_180),
.B(n_181),
.Y(n_275)
);

INVxp67_ASAP7_75t_SL g182 ( 
.A(n_183),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_270),
.Y(n_187)
);

NOR2x1_ASAP7_75t_L g565 ( 
.A(n_188),
.B(n_270),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_225),
.C(n_227),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_189),
.B(n_225),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_209),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_195),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_191),
.B(n_195),
.C(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_192),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_205),
.C(n_208),
.Y(n_195)
);

XNOR2x1_ASAP7_75t_L g267 ( 
.A(n_196),
.B(n_268),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_200),
.C(n_202),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_197),
.B(n_202),
.Y(n_246)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_200),
.B(n_246),
.Y(n_245)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_201),
.Y(n_239)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_205),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

BUFx12f_ASAP7_75t_L g214 ( 
.A(n_207),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_209),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_212),
.C(n_220),
.Y(n_209)
);

XNOR2x1_ASAP7_75t_L g341 ( 
.A(n_210),
.B(n_212),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_213),
.B(n_230),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_216),
.Y(n_231)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx5_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_219),
.Y(n_308)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_219),
.Y(n_361)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_220),
.Y(n_340)
);

MAJx2_ASAP7_75t_L g304 ( 
.A(n_221),
.B(n_305),
.C(n_307),
.Y(n_304)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_227),
.B(n_385),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_247),
.C(n_267),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_228),
.B(n_338),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_232),
.C(n_245),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_229),
.B(n_232),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_237),
.C(n_240),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_233),
.A2(n_240),
.B1(n_241),
.B2(n_382),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_233),
.Y(n_382)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_237),
.B(n_381),
.Y(n_380)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_240),
.B(n_446),
.C(n_449),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_240),
.A2(n_241),
.B1(n_446),
.B2(n_490),
.Y(n_489)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx4_ASAP7_75t_L g467 ( 
.A(n_243),
.Y(n_467)
);

BUFx3_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_244),
.Y(n_375)
);

XNOR2x2_ASAP7_75t_L g350 ( 
.A(n_245),
.B(n_351),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_247),
.B(n_267),
.Y(n_338)
);

MAJx2_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_257),
.C(n_263),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_248),
.B(n_335),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_249),
.B(n_253),
.Y(n_294)
);

INVx6_ASAP7_75t_L g517 ( 
.A(n_250),
.Y(n_517)
);

INVx5_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_256),
.Y(n_480)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_258),
.B(n_264),
.Y(n_335)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g547 ( 
.A1(n_263),
.A2(n_264),
.B1(n_426),
.B2(n_427),
.Y(n_547)
);

INVx1_ASAP7_75t_SL g263 ( 
.A(n_264),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_264),
.B(n_421),
.C(n_426),
.Y(n_420)
);

INVx2_ASAP7_75t_SL g265 ( 
.A(n_266),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_273),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_271),
.B(n_274),
.C(n_285),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_276),
.B1(n_278),
.B2(n_279),
.Y(n_273)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_274),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_276),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g285 ( 
.A(n_279),
.Y(n_285)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g564 ( 
.A1(n_281),
.A2(n_565),
.B(n_566),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_284),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_282),
.B(n_284),
.Y(n_566)
);

AO21x2_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_390),
.B(n_560),
.Y(n_286)
);

NOR2xp67_ASAP7_75t_SL g287 ( 
.A(n_288),
.B(n_383),
.Y(n_287)
);

AND2x2_ASAP7_75t_SL g288 ( 
.A(n_289),
.B(n_344),
.Y(n_288)
);

OR2x2_ASAP7_75t_L g561 ( 
.A(n_289),
.B(n_344),
.Y(n_561)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_336),
.Y(n_289)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_290),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_309),
.C(n_332),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_292),
.B(n_348),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_295),
.C(n_304),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_293),
.B(n_431),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_295),
.A2(n_296),
.B1(n_304),
.B2(n_432),
.Y(n_431)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_296),
.A2(n_406),
.B(n_413),
.Y(n_405)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g476 ( 
.A(n_299),
.Y(n_476)
);

INVx3_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_303),
.Y(n_448)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_304),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_305),
.B(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_307),
.Y(n_358)
);

HB1xp67_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_310),
.A2(n_333),
.B1(n_334),
.B2(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_310),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_324),
.C(n_327),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_311),
.B(n_378),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_316),
.C(n_320),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_312),
.A2(n_320),
.B1(n_403),
.B2(n_404),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_312),
.Y(n_404)
);

INVx4_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx6_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_316),
.B(n_402),
.Y(n_401)
);

INVx6_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_320),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_320),
.B(n_463),
.Y(n_462)
);

INVx6_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_324),
.A2(n_325),
.B1(n_327),
.B2(n_379),
.Y(n_378)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_327),
.Y(n_379)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx4_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_337),
.A2(n_339),
.B1(n_342),
.B2(n_343),
.Y(n_336)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_337),
.Y(n_342)
);

INVx1_ASAP7_75t_SL g343 ( 
.A(n_339),
.Y(n_343)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_339),
.Y(n_389)
);

XOR2x2_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_341),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g387 ( 
.A(n_342),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_350),
.C(n_352),
.Y(n_344)
);

HB1xp67_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_346),
.A2(n_347),
.B1(n_350),
.B2(n_395),
.Y(n_394)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_350),
.Y(n_395)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_353),
.B(n_394),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_376),
.C(n_380),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_SL g398 ( 
.A(n_354),
.B(n_399),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_359),
.C(n_364),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

XNOR2x1_ASAP7_75t_L g454 ( 
.A(n_356),
.B(n_455),
.Y(n_454)
);

XNOR2x1_ASAP7_75t_L g455 ( 
.A(n_359),
.B(n_364),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_363),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_360),
.B(n_363),
.Y(n_453)
);

NOR2x1_ASAP7_75t_R g360 ( 
.A(n_361),
.B(n_362),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_369),
.C(n_373),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_365),
.B(n_441),
.Y(n_440)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_369),
.A2(n_373),
.B1(n_442),
.B2(n_443),
.Y(n_441)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_369),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_369),
.B(n_505),
.C(n_507),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_SL g520 ( 
.A1(n_369),
.A2(n_443),
.B1(n_507),
.B2(n_508),
.Y(n_520)
);

INVx8_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx3_ASAP7_75t_L g498 ( 
.A(n_371),
.Y(n_498)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_372),
.Y(n_526)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_373),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_377),
.B(n_380),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_L g560 ( 
.A1(n_383),
.A2(n_561),
.B(n_562),
.Y(n_560)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_386),
.Y(n_383)
);

OR2x2_ASAP7_75t_L g562 ( 
.A(n_384),
.B(n_386),
.Y(n_562)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_388),
.C(n_389),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_456),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_396),
.C(n_433),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_393),
.B(n_397),
.Y(n_559)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_400),
.C(n_430),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_398),
.B(n_435),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_400),
.B(n_430),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_405),
.C(n_420),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_401),
.B(n_405),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_403),
.B(n_464),
.C(n_468),
.Y(n_487)
);

INVx1_ASAP7_75t_SL g407 ( 
.A(n_408),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_415),
.Y(n_413)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_419),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_420),
.B(n_438),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_SL g546 ( 
.A(n_421),
.B(n_547),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_422),
.B(n_425),
.Y(n_421)
);

XNOR2x1_ASAP7_75t_L g494 ( 
.A(n_422),
.B(n_425),
.Y(n_494)
);

CKINVDCx14_ASAP7_75t_R g514 ( 
.A(n_422),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g527 ( 
.A1(n_422),
.A2(n_514),
.B1(n_515),
.B2(n_528),
.Y(n_527)
);

INVx4_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

NOR2xp67_ASAP7_75t_L g433 ( 
.A(n_434),
.B(n_436),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_434),
.B(n_436),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_437),
.B(n_439),
.C(n_454),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g555 ( 
.A(n_437),
.B(n_556),
.Y(n_555)
);

XNOR2xp5_ASAP7_75t_L g556 ( 
.A(n_439),
.B(n_454),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_440),
.B(n_444),
.C(n_452),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g541 ( 
.A(n_440),
.B(n_542),
.Y(n_541)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g542 ( 
.A(n_445),
.B(n_453),
.Y(n_542)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_446),
.Y(n_490)
);

INVx4_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_449),
.B(n_489),
.Y(n_488)
);

INVx5_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

NAND3xp33_ASAP7_75t_L g456 ( 
.A(n_457),
.B(n_558),
.C(n_559),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_SL g457 ( 
.A1(n_458),
.A2(n_553),
.B(n_557),
.Y(n_457)
);

AOI21xp5_ASAP7_75t_L g458 ( 
.A1(n_459),
.A2(n_538),
.B(n_552),
.Y(n_458)
);

OAI21x1_ASAP7_75t_L g459 ( 
.A1(n_460),
.A2(n_499),
.B(n_537),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_485),
.Y(n_460)
);

OR2x2_ASAP7_75t_L g537 ( 
.A(n_461),
.B(n_485),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_462),
.B(n_469),
.C(n_477),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_462),
.B(n_502),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_464),
.B(n_468),
.Y(n_463)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_469),
.A2(n_470),
.B1(n_477),
.B2(n_503),
.Y(n_502)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_471),
.B(n_475),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_SL g506 ( 
.A(n_471),
.B(n_475),
.Y(n_506)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

INVx3_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

BUFx3_ASAP7_75t_L g533 ( 
.A(n_474),
.Y(n_533)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_477),
.Y(n_503)
);

AO22x1_ASAP7_75t_SL g477 ( 
.A1(n_478),
.A2(n_481),
.B1(n_483),
.B2(n_484),
.Y(n_477)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_478),
.Y(n_483)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

INVx1_ASAP7_75t_SL g484 ( 
.A(n_481),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_481),
.B(n_483),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_484),
.B(n_530),
.Y(n_529)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_486),
.B(n_491),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_487),
.B(n_488),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_487),
.B(n_491),
.C(n_551),
.Y(n_550)
);

HB1xp67_ASAP7_75t_L g551 ( 
.A(n_488),
.Y(n_551)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_492),
.B(n_493),
.Y(n_491)
);

MAJx2_ASAP7_75t_L g549 ( 
.A(n_492),
.B(n_494),
.C(n_495),
.Y(n_549)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_494),
.B(n_495),
.Y(n_493)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_498),
.Y(n_497)
);

AOI21x1_ASAP7_75t_L g499 ( 
.A1(n_500),
.A2(n_511),
.B(n_536),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_501),
.B(n_504),
.Y(n_500)
);

NOR2xp67_ASAP7_75t_SL g536 ( 
.A(n_501),
.B(n_504),
.Y(n_536)
);

OAI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_505),
.A2(n_506),
.B1(n_519),
.B2(n_520),
.Y(n_518)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

OAI21xp5_ASAP7_75t_SL g511 ( 
.A1(n_512),
.A2(n_521),
.B(n_535),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_513),
.B(n_518),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_513),
.B(n_518),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_SL g513 ( 
.A(n_514),
.B(n_515),
.Y(n_513)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_515),
.Y(n_528)
);

INVx5_ASAP7_75t_L g516 ( 
.A(n_517),
.Y(n_516)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_520),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_SL g521 ( 
.A1(n_522),
.A2(n_529),
.B(n_534),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_523),
.B(n_527),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_523),
.B(n_527),
.Y(n_534)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_525),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_526),
.Y(n_525)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_532),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_533),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_539),
.B(n_550),
.Y(n_538)
);

NOR2xp67_ASAP7_75t_SL g552 ( 
.A(n_539),
.B(n_550),
.Y(n_552)
);

AOI22xp5_ASAP7_75t_L g539 ( 
.A1(n_540),
.A2(n_541),
.B1(n_543),
.B2(n_544),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_540),
.B(n_545),
.C(n_549),
.Y(n_554)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_541),
.Y(n_540)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_544),
.Y(n_543)
);

AOI22xp5_ASAP7_75t_L g544 ( 
.A1(n_545),
.A2(n_546),
.B1(n_548),
.B2(n_549),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_546),
.Y(n_545)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_549),
.Y(n_548)
);

NOR2xp67_ASAP7_75t_L g553 ( 
.A(n_554),
.B(n_555),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_554),
.B(n_555),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_570),
.B(n_577),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_570),
.B(n_577),
.Y(n_579)
);

XNOR2xp5_ASAP7_75t_L g570 ( 
.A(n_571),
.B(n_572),
.Y(n_570)
);

CKINVDCx20_ASAP7_75t_R g576 ( 
.A(n_573),
.Y(n_576)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_575),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g578 ( 
.A(n_579),
.Y(n_578)
);


endmodule