module fake_jpeg_4417_n_125 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_125);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_125;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_7),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_20),
.B(n_21),
.Y(n_28)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_28),
.A2(n_30),
.B(n_37),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_20),
.B(n_1),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_33),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_34),
.B(n_36),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_35),
.Y(n_57)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_17),
.B(n_3),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_23),
.Y(n_62)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_42),
.Y(n_64)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_37),
.A2(n_16),
.B1(n_24),
.B2(n_26),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_43),
.A2(n_47),
.B1(n_46),
.B2(n_55),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_32),
.A2(n_15),
.B1(n_14),
.B2(n_22),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_27),
.B(n_23),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_49),
.B(n_21),
.Y(n_63)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_53),
.B(n_54),
.Y(n_65)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_58),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_61),
.Y(n_72)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_63),
.B(n_71),
.Y(n_84)
);

A2O1A1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_52),
.A2(n_17),
.B(n_5),
.C(n_6),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_67),
.A2(n_77),
.B(n_66),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_51),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_68),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_44),
.B(n_18),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_70),
.B(n_75),
.Y(n_83)
);

FAx1_ASAP7_75t_SL g71 ( 
.A(n_47),
.B(n_3),
.CI(n_5),
.CON(n_71),
.SN(n_71)
);

AND2x4_ASAP7_75t_SL g73 ( 
.A(n_46),
.B(n_50),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_73),
.B(n_74),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_50),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_74),
.B(n_79),
.Y(n_80)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_45),
.B(n_11),
.Y(n_77)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_78),
.A2(n_75),
.B1(n_76),
.B2(n_73),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_73),
.B(n_57),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_81),
.B(n_86),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_64),
.B(n_59),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_87),
.B(n_88),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_56),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_63),
.B(n_58),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_89),
.B(n_90),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_65),
.Y(n_90)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_91),
.Y(n_94)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_92),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_71),
.B(n_68),
.Y(n_93)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_93),
.Y(n_101)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_86),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_96),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_102),
.B(n_71),
.Y(n_105)
);

BUFx12_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_103),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_105),
.B(n_100),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_94),
.A2(n_84),
.B(n_93),
.Y(n_107)
);

AO21x1_ASAP7_75t_L g112 ( 
.A1(n_107),
.A2(n_67),
.B(n_83),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_101),
.B(n_83),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_108),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_98),
.B(n_69),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_109),
.B(n_110),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_97),
.B(n_80),
.C(n_69),
.Y(n_110)
);

A2O1A1O1Ixp25_ASAP7_75t_L g111 ( 
.A1(n_106),
.A2(n_95),
.B(n_99),
.C(n_91),
.D(n_100),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_111),
.B(n_102),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_112),
.B(n_113),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_115),
.B(n_103),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_116),
.B(n_117),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_118),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_114),
.Y(n_121)
);

AO21x1_ASAP7_75t_L g123 ( 
.A1(n_121),
.A2(n_122),
.B(n_77),
.Y(n_123)
);

A2O1A1Ixp33_ASAP7_75t_L g122 ( 
.A1(n_119),
.A2(n_118),
.B(n_115),
.C(n_103),
.Y(n_122)
);

BUFx24_ASAP7_75t_SL g124 ( 
.A(n_123),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_124),
.B(n_104),
.Y(n_125)
);


endmodule