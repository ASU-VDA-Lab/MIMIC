module real_aes_6934_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_503;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_659;
wire n_547;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_754;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_505;
wire n_502;
wire n_434;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_385;
wire n_358;
wire n_214;
wire n_275;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g176 ( .A1(n_0), .A2(n_177), .B(n_178), .C(n_182), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_1), .B(n_172), .Y(n_183) );
INVx1_ASAP7_75t_L g435 ( .A(n_2), .Y(n_435) );
NAND2xp5_ASAP7_75t_SL g254 ( .A(n_3), .B(n_137), .Y(n_254) );
AOI21xp5_ASAP7_75t_L g478 ( .A1(n_4), .A2(n_118), .B(n_479), .Y(n_478) );
A2O1A1Ixp33_ASAP7_75t_L g514 ( .A1(n_5), .A2(n_123), .B(n_128), .C(n_515), .Y(n_514) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_6), .A2(n_118), .B(n_223), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_7), .B(n_172), .Y(n_485) );
AO21x2_ASAP7_75t_L g200 ( .A1(n_8), .A2(n_151), .B(n_201), .Y(n_200) );
AND2x6_ASAP7_75t_L g123 ( .A(n_9), .B(n_124), .Y(n_123) );
A2O1A1Ixp33_ASAP7_75t_L g190 ( .A1(n_10), .A2(n_123), .B(n_128), .C(n_191), .Y(n_190) );
INVx1_ASAP7_75t_L g540 ( .A(n_11), .Y(n_540) );
NOR2xp33_ASAP7_75t_L g436 ( .A(n_12), .B(n_41), .Y(n_436) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_13), .B(n_181), .Y(n_517) );
INVx1_ASAP7_75t_L g147 ( .A(n_14), .Y(n_147) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_15), .B(n_137), .Y(n_207) );
A2O1A1Ixp33_ASAP7_75t_L g524 ( .A1(n_16), .A2(n_138), .B(n_525), .C(n_527), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_17), .B(n_172), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_18), .B(n_165), .Y(n_569) );
A2O1A1Ixp33_ASAP7_75t_L g158 ( .A1(n_19), .A2(n_128), .B(n_159), .C(n_164), .Y(n_158) );
A2O1A1Ixp33_ASAP7_75t_L g504 ( .A1(n_20), .A2(n_180), .B(n_195), .C(n_505), .Y(n_504) );
NAND2xp5_ASAP7_75t_SL g470 ( .A(n_21), .B(n_181), .Y(n_470) );
OAI22xp5_ASAP7_75t_L g736 ( .A1(n_22), .A2(n_77), .B1(n_737), .B2(n_738), .Y(n_736) );
CKINVDCx20_ASAP7_75t_R g738 ( .A(n_22), .Y(n_738) );
NAND2xp5_ASAP7_75t_SL g492 ( .A(n_23), .B(n_181), .Y(n_492) );
CKINVDCx16_ASAP7_75t_R g466 ( .A(n_24), .Y(n_466) );
INVx1_ASAP7_75t_L g491 ( .A(n_25), .Y(n_491) );
A2O1A1Ixp33_ASAP7_75t_L g203 ( .A1(n_26), .A2(n_128), .B(n_164), .C(n_204), .Y(n_203) );
BUFx6f_ASAP7_75t_L g122 ( .A(n_27), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g513 ( .A(n_28), .Y(n_513) );
AOI22xp5_ASAP7_75t_L g733 ( .A1(n_29), .A2(n_734), .B1(n_735), .B2(n_736), .Y(n_733) );
CKINVDCx20_ASAP7_75t_R g734 ( .A(n_29), .Y(n_734) );
CKINVDCx20_ASAP7_75t_R g748 ( .A(n_30), .Y(n_748) );
INVx1_ASAP7_75t_L g567 ( .A(n_31), .Y(n_567) );
AOI21xp5_ASAP7_75t_L g173 ( .A1(n_32), .A2(n_118), .B(n_174), .Y(n_173) );
INVx2_ASAP7_75t_L g121 ( .A(n_33), .Y(n_121) );
A2O1A1Ixp33_ASAP7_75t_L g125 ( .A1(n_34), .A2(n_126), .B(n_131), .C(n_141), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g519 ( .A(n_35), .Y(n_519) );
A2O1A1Ixp33_ASAP7_75t_L g481 ( .A1(n_36), .A2(n_180), .B(n_482), .C(n_484), .Y(n_481) );
INVxp67_ASAP7_75t_L g568 ( .A(n_37), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_38), .B(n_206), .Y(n_205) );
CKINVDCx14_ASAP7_75t_R g480 ( .A(n_39), .Y(n_480) );
A2O1A1Ixp33_ASAP7_75t_L g489 ( .A1(n_40), .A2(n_128), .B(n_164), .C(n_490), .Y(n_489) );
A2O1A1Ixp33_ASAP7_75t_L g537 ( .A1(n_42), .A2(n_182), .B(n_538), .C(n_539), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_43), .B(n_157), .Y(n_156) );
CKINVDCx20_ASAP7_75t_R g198 ( .A(n_44), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_45), .B(n_137), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_46), .B(n_118), .Y(n_202) );
CKINVDCx20_ASAP7_75t_R g494 ( .A(n_47), .Y(n_494) );
CKINVDCx20_ASAP7_75t_R g438 ( .A(n_48), .Y(n_438) );
CKINVDCx20_ASAP7_75t_R g564 ( .A(n_49), .Y(n_564) );
A2O1A1Ixp33_ASAP7_75t_L g214 ( .A1(n_50), .A2(n_126), .B(n_141), .C(n_215), .Y(n_214) );
OAI22xp5_ASAP7_75t_SL g107 ( .A1(n_51), .A2(n_87), .B1(n_108), .B2(n_109), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g109 ( .A(n_51), .Y(n_109) );
INVx1_ASAP7_75t_L g179 ( .A(n_52), .Y(n_179) );
INVx1_ASAP7_75t_L g216 ( .A(n_53), .Y(n_216) );
INVx1_ASAP7_75t_L g503 ( .A(n_54), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_55), .B(n_118), .Y(n_213) );
CKINVDCx20_ASAP7_75t_R g168 ( .A(n_56), .Y(n_168) );
CKINVDCx14_ASAP7_75t_R g536 ( .A(n_57), .Y(n_536) );
INVx1_ASAP7_75t_L g124 ( .A(n_58), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_59), .B(n_118), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_60), .B(n_172), .Y(n_230) );
A2O1A1Ixp33_ASAP7_75t_L g225 ( .A1(n_61), .A2(n_163), .B(n_226), .C(n_228), .Y(n_225) );
INVx1_ASAP7_75t_L g146 ( .A(n_62), .Y(n_146) );
INVx1_ASAP7_75t_SL g483 ( .A(n_63), .Y(n_483) );
CKINVDCx20_ASAP7_75t_R g445 ( .A(n_64), .Y(n_445) );
NAND2xp5_ASAP7_75t_SL g136 ( .A(n_65), .B(n_137), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_66), .B(n_172), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_67), .B(n_138), .Y(n_192) );
INVx1_ASAP7_75t_L g469 ( .A(n_68), .Y(n_469) );
CKINVDCx16_ASAP7_75t_R g175 ( .A(n_69), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_70), .B(n_134), .Y(n_160) );
A2O1A1Ixp33_ASAP7_75t_L g251 ( .A1(n_71), .A2(n_128), .B(n_141), .C(n_252), .Y(n_251) );
CKINVDCx16_ASAP7_75t_R g224 ( .A(n_72), .Y(n_224) );
INVx1_ASAP7_75t_L g448 ( .A(n_73), .Y(n_448) );
AOI21xp5_ASAP7_75t_L g534 ( .A1(n_74), .A2(n_118), .B(n_535), .Y(n_534) );
CKINVDCx20_ASAP7_75t_R g473 ( .A(n_75), .Y(n_473) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_76), .A2(n_118), .B(n_522), .Y(n_521) );
CKINVDCx20_ASAP7_75t_R g737 ( .A(n_77), .Y(n_737) );
AOI21xp5_ASAP7_75t_L g562 ( .A1(n_78), .A2(n_157), .B(n_563), .Y(n_562) );
CKINVDCx16_ASAP7_75t_R g488 ( .A(n_79), .Y(n_488) );
INVx1_ASAP7_75t_L g523 ( .A(n_80), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g161 ( .A(n_81), .B(n_133), .Y(n_161) );
CKINVDCx20_ASAP7_75t_R g149 ( .A(n_82), .Y(n_149) );
AOI21xp5_ASAP7_75t_L g501 ( .A1(n_83), .A2(n_118), .B(n_502), .Y(n_501) );
INVx1_ASAP7_75t_L g526 ( .A(n_84), .Y(n_526) );
INVx2_ASAP7_75t_L g144 ( .A(n_85), .Y(n_144) );
INVx1_ASAP7_75t_L g516 ( .A(n_86), .Y(n_516) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_87), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g259 ( .A(n_88), .Y(n_259) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_89), .B(n_181), .Y(n_193) );
OR2x2_ASAP7_75t_L g432 ( .A(n_90), .B(n_433), .Y(n_432) );
OR2x2_ASAP7_75t_L g452 ( .A(n_90), .B(n_434), .Y(n_452) );
INVx2_ASAP7_75t_L g456 ( .A(n_90), .Y(n_456) );
A2O1A1Ixp33_ASAP7_75t_L g467 ( .A1(n_91), .A2(n_128), .B(n_141), .C(n_468), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g117 ( .A(n_92), .B(n_118), .Y(n_117) );
INVx1_ASAP7_75t_L g132 ( .A(n_93), .Y(n_132) );
INVxp67_ASAP7_75t_L g229 ( .A(n_94), .Y(n_229) );
AOI222xp33_ASAP7_75t_L g102 ( .A1(n_95), .A2(n_103), .B1(n_441), .B2(n_449), .C1(n_749), .C2(n_752), .Y(n_102) );
OAI22xp33_ASAP7_75t_SL g105 ( .A1(n_95), .A2(n_106), .B1(n_428), .B2(n_429), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g428 ( .A(n_95), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_96), .B(n_151), .Y(n_541) );
INVx2_ASAP7_75t_L g506 ( .A(n_97), .Y(n_506) );
INVx1_ASAP7_75t_L g188 ( .A(n_98), .Y(n_188) );
INVx1_ASAP7_75t_L g253 ( .A(n_99), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_100), .B(n_448), .Y(n_447) );
AND2x2_ASAP7_75t_L g218 ( .A(n_101), .B(n_143), .Y(n_218) );
INVxp67_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
AOI21xp5_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_430), .B(n_437), .Y(n_104) );
INVx1_ASAP7_75t_L g429 ( .A(n_106), .Y(n_429) );
XOR2xp5_ASAP7_75t_L g106 ( .A(n_107), .B(n_110), .Y(n_106) );
INVx2_ASAP7_75t_L g453 ( .A(n_110), .Y(n_453) );
AOI22xp5_ASAP7_75t_L g739 ( .A1(n_110), .A2(n_740), .B1(n_743), .B2(n_744), .Y(n_739) );
OR3x2_ASAP7_75t_L g110 ( .A(n_111), .B(n_342), .C(n_385), .Y(n_110) );
NAND5xp2_ASAP7_75t_L g111 ( .A(n_112), .B(n_269), .C(n_299), .D(n_316), .E(n_331), .Y(n_111) );
AOI221xp5_ASAP7_75t_SL g112 ( .A1(n_113), .A2(n_184), .B1(n_231), .B2(n_237), .C(n_241), .Y(n_112) );
AND2x2_ASAP7_75t_L g113 ( .A(n_114), .B(n_153), .Y(n_113) );
OR2x2_ASAP7_75t_L g246 ( .A(n_114), .B(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g286 ( .A(n_114), .B(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g304 ( .A(n_114), .B(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_114), .B(n_239), .Y(n_321) );
OR2x2_ASAP7_75t_L g333 ( .A(n_114), .B(n_334), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_114), .B(n_292), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_114), .B(n_366), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_114), .B(n_270), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_114), .B(n_278), .Y(n_384) );
AND2x2_ASAP7_75t_L g416 ( .A(n_114), .B(n_170), .Y(n_416) );
HB1xp67_ASAP7_75t_L g424 ( .A(n_114), .Y(n_424) );
INVx5_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_115), .B(n_239), .Y(n_238) );
AND2x2_ASAP7_75t_L g243 ( .A(n_115), .B(n_219), .Y(n_243) );
BUFx2_ASAP7_75t_L g266 ( .A(n_115), .Y(n_266) );
AND2x2_ASAP7_75t_L g295 ( .A(n_115), .B(n_154), .Y(n_295) );
AND2x2_ASAP7_75t_L g350 ( .A(n_115), .B(n_247), .Y(n_350) );
OR2x6_ASAP7_75t_L g115 ( .A(n_116), .B(n_148), .Y(n_115) );
AOI21xp5_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_125), .B(n_143), .Y(n_116) );
BUFx2_ASAP7_75t_L g157 ( .A(n_118), .Y(n_157) );
AND2x4_ASAP7_75t_L g118 ( .A(n_119), .B(n_123), .Y(n_118) );
NAND2x1p5_ASAP7_75t_L g189 ( .A(n_119), .B(n_123), .Y(n_189) );
AND2x2_ASAP7_75t_L g119 ( .A(n_120), .B(n_122), .Y(n_119) );
INVx1_ASAP7_75t_L g163 ( .A(n_120), .Y(n_163) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx2_ASAP7_75t_L g129 ( .A(n_121), .Y(n_129) );
INVx1_ASAP7_75t_L g196 ( .A(n_121), .Y(n_196) );
INVx1_ASAP7_75t_L g130 ( .A(n_122), .Y(n_130) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_122), .Y(n_135) );
INVx3_ASAP7_75t_L g138 ( .A(n_122), .Y(n_138) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_122), .Y(n_181) );
INVx1_ASAP7_75t_L g206 ( .A(n_122), .Y(n_206) );
INVx4_ASAP7_75t_SL g142 ( .A(n_123), .Y(n_142) );
BUFx3_ASAP7_75t_L g164 ( .A(n_123), .Y(n_164) );
INVx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
O2A1O1Ixp33_ASAP7_75t_SL g174 ( .A1(n_127), .A2(n_142), .B(n_175), .C(n_176), .Y(n_174) );
O2A1O1Ixp33_ASAP7_75t_L g223 ( .A1(n_127), .A2(n_142), .B(n_224), .C(n_225), .Y(n_223) );
O2A1O1Ixp33_ASAP7_75t_L g479 ( .A1(n_127), .A2(n_142), .B(n_480), .C(n_481), .Y(n_479) );
O2A1O1Ixp33_ASAP7_75t_SL g502 ( .A1(n_127), .A2(n_142), .B(n_503), .C(n_504), .Y(n_502) );
O2A1O1Ixp33_ASAP7_75t_SL g522 ( .A1(n_127), .A2(n_142), .B(n_523), .C(n_524), .Y(n_522) );
O2A1O1Ixp33_ASAP7_75t_SL g535 ( .A1(n_127), .A2(n_142), .B(n_536), .C(n_537), .Y(n_535) );
O2A1O1Ixp33_ASAP7_75t_SL g563 ( .A1(n_127), .A2(n_142), .B(n_564), .C(n_565), .Y(n_563) );
INVx5_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
AND2x6_ASAP7_75t_L g128 ( .A(n_129), .B(n_130), .Y(n_128) );
BUFx3_ASAP7_75t_L g140 ( .A(n_129), .Y(n_140) );
BUFx6f_ASAP7_75t_L g256 ( .A(n_129), .Y(n_256) );
O2A1O1Ixp33_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_133), .B(n_136), .C(n_139), .Y(n_131) );
O2A1O1Ixp33_ASAP7_75t_L g215 ( .A1(n_133), .A2(n_139), .B(n_216), .C(n_217), .Y(n_215) );
O2A1O1Ixp33_ASAP7_75t_L g468 ( .A1(n_133), .A2(n_469), .B(n_470), .C(n_471), .Y(n_468) );
O2A1O1Ixp5_ASAP7_75t_L g515 ( .A1(n_133), .A2(n_471), .B(n_516), .C(n_517), .Y(n_515) );
INVx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx4_ASAP7_75t_L g227 ( .A(n_135), .Y(n_227) );
INVx2_ASAP7_75t_L g177 ( .A(n_137), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_137), .B(n_229), .Y(n_228) );
O2A1O1Ixp33_ASAP7_75t_L g490 ( .A1(n_137), .A2(n_162), .B(n_491), .C(n_492), .Y(n_490) );
OAI22xp33_ASAP7_75t_L g566 ( .A1(n_137), .A2(n_227), .B1(n_567), .B2(n_568), .Y(n_566) );
INVx5_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
NOR2xp33_ASAP7_75t_L g539 ( .A(n_138), .B(n_540), .Y(n_539) );
HB1xp67_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx2_ASAP7_75t_L g182 ( .A(n_140), .Y(n_182) );
INVx1_ASAP7_75t_L g527 ( .A(n_140), .Y(n_527) );
INVx1_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx2_ASAP7_75t_L g166 ( .A(n_143), .Y(n_166) );
INVx1_ASAP7_75t_L g169 ( .A(n_143), .Y(n_169) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_143), .A2(n_213), .B(n_214), .Y(n_212) );
O2A1O1Ixp33_ASAP7_75t_L g487 ( .A1(n_143), .A2(n_189), .B(n_488), .C(n_489), .Y(n_487) );
OA21x2_ASAP7_75t_L g533 ( .A1(n_143), .A2(n_534), .B(n_541), .Y(n_533) );
AND2x2_ASAP7_75t_SL g143 ( .A(n_144), .B(n_145), .Y(n_143) );
AND2x2_ASAP7_75t_L g152 ( .A(n_144), .B(n_145), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_146), .B(n_147), .Y(n_145) );
NOR2xp33_ASAP7_75t_L g148 ( .A(n_149), .B(n_150), .Y(n_148) );
INVx3_ASAP7_75t_L g172 ( .A(n_150), .Y(n_172) );
AO21x2_ASAP7_75t_L g186 ( .A1(n_150), .A2(n_187), .B(n_197), .Y(n_186) );
AO21x2_ASAP7_75t_L g249 ( .A1(n_150), .A2(n_250), .B(n_258), .Y(n_249) );
NOR2xp33_ASAP7_75t_L g258 ( .A(n_150), .B(n_259), .Y(n_258) );
AO21x2_ASAP7_75t_L g464 ( .A1(n_150), .A2(n_465), .B(n_472), .Y(n_464) );
NOR2xp33_ASAP7_75t_L g493 ( .A(n_150), .B(n_494), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g518 ( .A(n_150), .B(n_519), .Y(n_518) );
INVx4_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
AOI21xp5_ASAP7_75t_L g201 ( .A1(n_151), .A2(n_202), .B(n_203), .Y(n_201) );
HB1xp67_ASAP7_75t_L g221 ( .A(n_151), .Y(n_221) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g199 ( .A(n_152), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_153), .B(n_304), .Y(n_313) );
OAI32xp33_ASAP7_75t_L g327 ( .A1(n_153), .A2(n_263), .A3(n_328), .B1(n_329), .B2(n_330), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_153), .B(n_329), .Y(n_359) );
NOR2xp33_ASAP7_75t_L g370 ( .A(n_153), .B(n_246), .Y(n_370) );
INVx1_ASAP7_75t_SL g399 ( .A(n_153), .Y(n_399) );
NAND4xp25_ASAP7_75t_L g408 ( .A(n_153), .B(n_186), .C(n_350), .D(n_409), .Y(n_408) );
AND2x4_ASAP7_75t_L g153 ( .A(n_154), .B(n_170), .Y(n_153) );
INVx5_ASAP7_75t_L g240 ( .A(n_154), .Y(n_240) );
AND2x2_ASAP7_75t_L g270 ( .A(n_154), .B(n_171), .Y(n_270) );
HB1xp67_ASAP7_75t_L g349 ( .A(n_154), .Y(n_349) );
AND2x2_ASAP7_75t_L g419 ( .A(n_154), .B(n_366), .Y(n_419) );
OR2x6_ASAP7_75t_L g154 ( .A(n_155), .B(n_167), .Y(n_154) );
AOI21xp5_ASAP7_75t_SL g155 ( .A1(n_156), .A2(n_158), .B(n_165), .Y(n_155) );
AOI21xp5_ASAP7_75t_L g159 ( .A1(n_160), .A2(n_161), .B(n_162), .Y(n_159) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
NAND2xp5_ASAP7_75t_SL g565 ( .A(n_163), .B(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
NOR2xp33_ASAP7_75t_L g472 ( .A(n_166), .B(n_473), .Y(n_472) );
NOR2xp33_ASAP7_75t_L g167 ( .A(n_168), .B(n_169), .Y(n_167) );
AO21x2_ASAP7_75t_L g511 ( .A1(n_169), .A2(n_512), .B(n_518), .Y(n_511) );
AND2x4_ASAP7_75t_L g292 ( .A(n_170), .B(n_240), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_170), .B(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g326 ( .A(n_170), .B(n_247), .Y(n_326) );
INVx2_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
AND2x2_ASAP7_75t_L g239 ( .A(n_171), .B(n_240), .Y(n_239) );
AND2x2_ASAP7_75t_L g278 ( .A(n_171), .B(n_249), .Y(n_278) );
AND2x2_ASAP7_75t_L g287 ( .A(n_171), .B(n_248), .Y(n_287) );
OA21x2_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_173), .B(n_183), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g178 ( .A(n_179), .B(n_180), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g482 ( .A(n_180), .B(n_483), .Y(n_482) );
INVx4_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx2_ASAP7_75t_L g538 ( .A(n_181), .Y(n_538) );
INVx2_ASAP7_75t_L g471 ( .A(n_182), .Y(n_471) );
AOI222xp33_ASAP7_75t_L g355 ( .A1(n_184), .A2(n_356), .B1(n_358), .B2(n_360), .C1(n_363), .C2(n_364), .Y(n_355) );
AND2x4_ASAP7_75t_L g184 ( .A(n_185), .B(n_208), .Y(n_184) );
AND2x2_ASAP7_75t_L g288 ( .A(n_185), .B(n_289), .Y(n_288) );
NAND3xp33_ASAP7_75t_L g405 ( .A(n_185), .B(n_266), .C(n_406), .Y(n_405) );
AND2x2_ASAP7_75t_L g185 ( .A(n_186), .B(n_200), .Y(n_185) );
INVx5_ASAP7_75t_SL g236 ( .A(n_186), .Y(n_236) );
OAI322xp33_ASAP7_75t_L g241 ( .A1(n_186), .A2(n_242), .A3(n_244), .B1(n_245), .B2(n_260), .C1(n_263), .C2(n_265), .Y(n_241) );
NAND2xp5_ASAP7_75t_SL g308 ( .A(n_186), .B(n_234), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_186), .B(n_220), .Y(n_414) );
OAI21xp5_ASAP7_75t_L g187 ( .A1(n_188), .A2(n_189), .B(n_190), .Y(n_187) );
OAI21xp5_ASAP7_75t_L g465 ( .A1(n_189), .A2(n_466), .B(n_467), .Y(n_465) );
OAI21xp5_ASAP7_75t_L g512 ( .A1(n_189), .A2(n_513), .B(n_514), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g191 ( .A1(n_192), .A2(n_193), .B(n_194), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_194), .A2(n_205), .B(n_207), .Y(n_204) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
INVx3_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_198), .B(n_199), .Y(n_197) );
INVx2_ASAP7_75t_L g561 ( .A(n_199), .Y(n_561) );
INVx2_ASAP7_75t_L g234 ( .A(n_200), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_200), .B(n_210), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_208), .B(n_273), .Y(n_328) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
OR2x2_ASAP7_75t_L g307 ( .A(n_209), .B(n_308), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_210), .B(n_219), .Y(n_209) );
OR2x2_ASAP7_75t_L g235 ( .A(n_210), .B(n_236), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_210), .B(n_243), .Y(n_242) );
OR2x2_ASAP7_75t_L g275 ( .A(n_210), .B(n_220), .Y(n_275) );
AND2x2_ASAP7_75t_L g298 ( .A(n_210), .B(n_234), .Y(n_298) );
NOR2xp33_ASAP7_75t_L g309 ( .A(n_210), .B(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g314 ( .A(n_210), .B(n_273), .Y(n_314) );
AND2x2_ASAP7_75t_L g322 ( .A(n_210), .B(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_210), .B(n_282), .Y(n_372) );
INVx5_ASAP7_75t_SL g210 ( .A(n_211), .Y(n_210) );
AND2x2_ASAP7_75t_L g262 ( .A(n_211), .B(n_236), .Y(n_262) );
OR2x2_ASAP7_75t_L g263 ( .A(n_211), .B(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g289 ( .A(n_211), .B(n_220), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_211), .B(n_336), .Y(n_377) );
OR2x2_ASAP7_75t_L g393 ( .A(n_211), .B(n_337), .Y(n_393) );
AND2x2_ASAP7_75t_SL g400 ( .A(n_211), .B(n_354), .Y(n_400) );
HB1xp67_ASAP7_75t_L g407 ( .A(n_211), .Y(n_407) );
OR2x6_ASAP7_75t_L g211 ( .A(n_212), .B(n_218), .Y(n_211) );
AND2x2_ASAP7_75t_L g261 ( .A(n_219), .B(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g311 ( .A(n_219), .B(n_234), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_219), .B(n_236), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_219), .B(n_273), .Y(n_395) );
INVx3_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_220), .B(n_236), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_220), .B(n_234), .Y(n_283) );
OR2x2_ASAP7_75t_L g337 ( .A(n_220), .B(n_234), .Y(n_337) );
AND2x2_ASAP7_75t_L g354 ( .A(n_220), .B(n_233), .Y(n_354) );
INVxp67_ASAP7_75t_L g376 ( .A(n_220), .Y(n_376) );
AND2x2_ASAP7_75t_L g403 ( .A(n_220), .B(n_273), .Y(n_403) );
HB1xp67_ASAP7_75t_L g410 ( .A(n_220), .Y(n_410) );
OA21x2_ASAP7_75t_L g220 ( .A1(n_221), .A2(n_222), .B(n_230), .Y(n_220) );
OA21x2_ASAP7_75t_L g477 ( .A1(n_221), .A2(n_478), .B(n_485), .Y(n_477) );
OA21x2_ASAP7_75t_L g500 ( .A1(n_221), .A2(n_501), .B(n_507), .Y(n_500) );
OA21x2_ASAP7_75t_L g520 ( .A1(n_221), .A2(n_521), .B(n_528), .Y(n_520) );
O2A1O1Ixp33_ASAP7_75t_L g252 ( .A1(n_226), .A2(n_253), .B(n_254), .C(n_255), .Y(n_252) );
INVx1_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g505 ( .A(n_227), .B(n_506), .Y(n_505) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_227), .B(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
OR2x2_ASAP7_75t_L g232 ( .A(n_233), .B(n_235), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_233), .B(n_284), .Y(n_357) );
INVx1_ASAP7_75t_SL g233 ( .A(n_234), .Y(n_233) );
AND2x2_ASAP7_75t_L g273 ( .A(n_234), .B(n_236), .Y(n_273) );
OR2x2_ASAP7_75t_L g340 ( .A(n_234), .B(n_341), .Y(n_340) );
INVx2_ASAP7_75t_L g284 ( .A(n_235), .Y(n_284) );
OR2x2_ASAP7_75t_L g345 ( .A(n_235), .B(n_337), .Y(n_345) );
INVx1_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
INVx1_ASAP7_75t_L g244 ( .A(n_239), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_239), .B(n_304), .Y(n_303) );
OR2x2_ASAP7_75t_L g245 ( .A(n_240), .B(n_246), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_240), .B(n_268), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_240), .B(n_247), .Y(n_280) );
INVx2_ASAP7_75t_L g325 ( .A(n_240), .Y(n_325) );
AND2x2_ASAP7_75t_L g338 ( .A(n_240), .B(n_278), .Y(n_338) );
AND2x2_ASAP7_75t_L g363 ( .A(n_240), .B(n_287), .Y(n_363) );
INVx1_ASAP7_75t_L g315 ( .A(n_245), .Y(n_315) );
INVx2_ASAP7_75t_SL g302 ( .A(n_246), .Y(n_302) );
INVx1_ASAP7_75t_L g305 ( .A(n_247), .Y(n_305) );
INVx2_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
HB1xp67_ASAP7_75t_L g268 ( .A(n_248), .Y(n_268) );
INVx2_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
BUFx2_ASAP7_75t_L g366 ( .A(n_249), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_251), .B(n_257), .Y(n_250) );
HB1xp67_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
INVx3_ASAP7_75t_L g484 ( .A(n_256), .Y(n_484) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g335 ( .A(n_262), .B(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g341 ( .A(n_262), .Y(n_341) );
AOI22xp5_ASAP7_75t_L g343 ( .A1(n_262), .A2(n_344), .B1(n_346), .B2(n_351), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_262), .B(n_354), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_263), .B(n_357), .Y(n_356) );
INVx1_ASAP7_75t_SL g297 ( .A(n_264), .Y(n_297) );
OR2x2_ASAP7_75t_L g265 ( .A(n_266), .B(n_267), .Y(n_265) );
OR2x2_ASAP7_75t_L g279 ( .A(n_266), .B(n_280), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_266), .B(n_270), .Y(n_330) );
AND2x2_ASAP7_75t_L g353 ( .A(n_266), .B(n_354), .Y(n_353) );
BUFx2_ASAP7_75t_L g329 ( .A(n_268), .Y(n_329) );
AOI211xp5_ASAP7_75t_L g269 ( .A1(n_270), .A2(n_271), .B(n_276), .C(n_290), .Y(n_269) );
INVx1_ASAP7_75t_L g293 ( .A(n_270), .Y(n_293) );
OAI221xp5_ASAP7_75t_SL g401 ( .A1(n_270), .A2(n_402), .B1(n_404), .B2(n_405), .C(n_408), .Y(n_401) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_273), .B(n_274), .Y(n_272) );
INVx1_ASAP7_75t_L g420 ( .A(n_273), .Y(n_420) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
OR2x2_ASAP7_75t_L g369 ( .A(n_275), .B(n_308), .Y(n_369) );
A2O1A1Ixp33_ASAP7_75t_L g276 ( .A1(n_277), .A2(n_279), .B(n_281), .C(n_285), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_282), .B(n_284), .Y(n_281) );
INVx1_ASAP7_75t_SL g282 ( .A(n_283), .Y(n_282) );
OAI32xp33_ASAP7_75t_L g394 ( .A1(n_283), .A2(n_284), .A3(n_347), .B1(n_384), .B2(n_395), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_286), .B(n_288), .Y(n_285) );
AND2x2_ASAP7_75t_L g426 ( .A(n_286), .B(n_325), .Y(n_426) );
AND2x2_ASAP7_75t_L g373 ( .A(n_287), .B(n_325), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_287), .B(n_295), .Y(n_391) );
AOI31xp33_ASAP7_75t_SL g290 ( .A1(n_291), .A2(n_293), .A3(n_294), .B(n_296), .Y(n_290) );
INVxp67_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_292), .B(n_304), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_292), .B(n_302), .Y(n_389) );
AOI221xp5_ASAP7_75t_L g411 ( .A1(n_292), .A2(n_322), .B1(n_412), .B2(n_415), .C(n_417), .Y(n_411) );
CKINVDCx16_ASAP7_75t_R g294 ( .A(n_295), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
AND2x2_ASAP7_75t_L g317 ( .A(n_297), .B(n_318), .Y(n_317) );
AOI222xp33_ASAP7_75t_L g299 ( .A1(n_300), .A2(n_306), .B1(n_309), .B2(n_312), .C1(n_314), .C2(n_315), .Y(n_299) );
NAND2xp5_ASAP7_75t_SL g300 ( .A(n_301), .B(n_303), .Y(n_300) );
INVx1_ASAP7_75t_L g382 ( .A(n_301), .Y(n_382) );
INVx1_ASAP7_75t_L g404 ( .A(n_304), .Y(n_404) );
INVx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
OAI22xp5_ASAP7_75t_L g417 ( .A1(n_307), .A2(n_418), .B1(n_420), .B2(n_421), .Y(n_417) );
INVx1_ASAP7_75t_L g323 ( .A(n_308), .Y(n_323) );
INVx1_ASAP7_75t_SL g310 ( .A(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
AOI221xp5_ASAP7_75t_L g316 ( .A1(n_317), .A2(n_320), .B1(n_322), .B2(n_324), .C(n_327), .Y(n_316) );
INVx1_ASAP7_75t_SL g318 ( .A(n_319), .Y(n_318) );
OR2x2_ASAP7_75t_L g361 ( .A(n_319), .B(n_362), .Y(n_361) );
OR2x2_ASAP7_75t_L g413 ( .A(n_319), .B(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g388 ( .A(n_324), .Y(n_388) );
AND2x2_ASAP7_75t_L g324 ( .A(n_325), .B(n_326), .Y(n_324) );
INVx1_ASAP7_75t_L g352 ( .A(n_325), .Y(n_352) );
INVx1_ASAP7_75t_L g334 ( .A(n_326), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_329), .B(n_416), .Y(n_421) );
AOI22xp33_ASAP7_75t_L g331 ( .A1(n_332), .A2(n_335), .B1(n_338), .B2(n_339), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx1_ASAP7_75t_SL g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_SL g425 ( .A(n_338), .Y(n_425) );
INVxp33_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
NOR2xp33_ASAP7_75t_L g383 ( .A(n_340), .B(n_384), .Y(n_383) );
OAI32xp33_ASAP7_75t_L g374 ( .A1(n_341), .A2(n_375), .A3(n_376), .B1(n_377), .B2(n_378), .Y(n_374) );
NAND4xp25_ASAP7_75t_L g342 ( .A(n_343), .B(n_355), .C(n_367), .D(n_379), .Y(n_342) );
INVx1_ASAP7_75t_SL g344 ( .A(n_345), .Y(n_344) );
NAND2xp33_ASAP7_75t_SL g346 ( .A(n_347), .B(n_348), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_349), .B(n_350), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_350), .B(n_399), .Y(n_398) );
AND2x2_ASAP7_75t_L g351 ( .A(n_352), .B(n_353), .Y(n_351) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
CKINVDCx16_ASAP7_75t_R g360 ( .A(n_361), .Y(n_360) );
AOI221xp5_ASAP7_75t_L g396 ( .A1(n_364), .A2(n_380), .B1(n_397), .B2(n_400), .C(n_401), .Y(n_396) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
AND2x2_ASAP7_75t_L g415 ( .A(n_366), .B(n_416), .Y(n_415) );
AOI221xp5_ASAP7_75t_L g367 ( .A1(n_368), .A2(n_370), .B1(n_371), .B2(n_373), .C(n_374), .Y(n_367) );
INVx1_ASAP7_75t_SL g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
NOR2xp33_ASAP7_75t_L g406 ( .A(n_376), .B(n_407), .Y(n_406) );
AOI21xp5_ASAP7_75t_L g379 ( .A1(n_380), .A2(n_382), .B(n_383), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
NAND4xp25_ASAP7_75t_L g385 ( .A(n_386), .B(n_396), .C(n_411), .D(n_422), .Y(n_385) );
O2A1O1Ixp33_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_390), .B(n_392), .C(n_394), .Y(n_386) );
NAND2xp5_ASAP7_75t_SL g387 ( .A(n_388), .B(n_389), .Y(n_387) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVxp67_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_SL g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g427 ( .A(n_414), .Y(n_427) );
INVx2_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
OAI21xp5_ASAP7_75t_L g422 ( .A1(n_423), .A2(n_426), .B(n_427), .Y(n_422) );
NOR2xp33_ASAP7_75t_L g423 ( .A(n_424), .B(n_425), .Y(n_423) );
NAND2xp33_ASAP7_75t_L g750 ( .A(n_430), .B(n_751), .Y(n_750) );
INVx1_ASAP7_75t_SL g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_SL g431 ( .A(n_432), .Y(n_431) );
INVx2_ASAP7_75t_L g440 ( .A(n_432), .Y(n_440) );
BUFx2_ASAP7_75t_L g754 ( .A(n_432), .Y(n_754) );
NOR2x2_ASAP7_75t_L g747 ( .A(n_433), .B(n_456), .Y(n_747) );
INVx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
OR2x2_ASAP7_75t_L g455 ( .A(n_434), .B(n_456), .Y(n_455) );
AND2x2_ASAP7_75t_L g434 ( .A(n_435), .B(n_436), .Y(n_434) );
NOR2xp33_ASAP7_75t_L g437 ( .A(n_438), .B(n_439), .Y(n_437) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
HB1xp67_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_443), .B(n_446), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
NOR2xp33_ASAP7_75t_SL g751 ( .A(n_445), .B(n_447), .Y(n_751) );
OA21x2_ASAP7_75t_L g753 ( .A1(n_445), .A2(n_446), .B(n_754), .Y(n_753) );
INVx1_ASAP7_75t_SL g446 ( .A(n_447), .Y(n_446) );
OAI222xp33_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_733), .B1(n_739), .B2(n_745), .C1(n_746), .C2(n_748), .Y(n_449) );
AOI22xp5_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_453), .B1(n_454), .B2(n_457), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g742 ( .A(n_452), .Y(n_742) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx6_ASAP7_75t_L g743 ( .A(n_455), .Y(n_743) );
INVx3_ASAP7_75t_L g744 ( .A(n_457), .Y(n_744) );
AND2x2_ASAP7_75t_SL g457 ( .A(n_458), .B(n_688), .Y(n_457) );
NOR4xp25_ASAP7_75t_L g458 ( .A(n_459), .B(n_625), .C(n_659), .D(n_675), .Y(n_458) );
NAND4xp25_ASAP7_75t_SL g459 ( .A(n_460), .B(n_554), .C(n_589), .D(n_605), .Y(n_459) );
AOI222xp33_ASAP7_75t_L g460 ( .A1(n_461), .A2(n_495), .B1(n_529), .B2(n_542), .C1(n_547), .C2(n_553), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
AOI31xp33_ASAP7_75t_L g721 ( .A1(n_462), .A2(n_722), .A3(n_723), .B(n_725), .Y(n_721) );
OR2x2_ASAP7_75t_L g462 ( .A(n_463), .B(n_474), .Y(n_462) );
AND2x2_ASAP7_75t_L g696 ( .A(n_463), .B(n_476), .Y(n_696) );
BUFx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx2_ASAP7_75t_SL g546 ( .A(n_464), .Y(n_546) );
AND2x2_ASAP7_75t_L g553 ( .A(n_464), .B(n_486), .Y(n_553) );
AND2x2_ASAP7_75t_L g610 ( .A(n_464), .B(n_477), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_474), .B(n_640), .Y(n_639) );
INVx3_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
NOR2xp33_ASAP7_75t_L g573 ( .A(n_475), .B(n_574), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_475), .B(n_557), .Y(n_600) );
AND2x2_ASAP7_75t_L g693 ( .A(n_475), .B(n_633), .Y(n_693) );
OAI321xp33_ASAP7_75t_L g727 ( .A1(n_475), .A2(n_546), .A3(n_700), .B1(n_728), .B2(n_730), .C(n_731), .Y(n_727) );
NAND4xp25_ASAP7_75t_L g731 ( .A(n_475), .B(n_532), .C(n_640), .D(n_732), .Y(n_731) );
AND2x4_ASAP7_75t_L g475 ( .A(n_476), .B(n_486), .Y(n_475) );
AND2x2_ASAP7_75t_L g595 ( .A(n_476), .B(n_544), .Y(n_595) );
AND2x2_ASAP7_75t_L g614 ( .A(n_476), .B(n_546), .Y(n_614) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
AND2x2_ASAP7_75t_L g545 ( .A(n_477), .B(n_546), .Y(n_545) );
AND2x2_ASAP7_75t_L g570 ( .A(n_477), .B(n_486), .Y(n_570) );
AND2x2_ASAP7_75t_L g656 ( .A(n_477), .B(n_544), .Y(n_656) );
INVx3_ASAP7_75t_SL g544 ( .A(n_486), .Y(n_544) );
AND2x2_ASAP7_75t_L g588 ( .A(n_486), .B(n_575), .Y(n_588) );
OR2x2_ASAP7_75t_L g621 ( .A(n_486), .B(n_546), .Y(n_621) );
HB1xp67_ASAP7_75t_L g628 ( .A(n_486), .Y(n_628) );
AND2x2_ASAP7_75t_L g657 ( .A(n_486), .B(n_545), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_486), .B(n_630), .Y(n_672) );
AND2x2_ASAP7_75t_L g704 ( .A(n_486), .B(n_696), .Y(n_704) );
AND2x2_ASAP7_75t_L g713 ( .A(n_486), .B(n_558), .Y(n_713) );
OR2x6_ASAP7_75t_L g486 ( .A(n_487), .B(n_493), .Y(n_486) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_497), .B(n_508), .Y(n_496) );
INVx1_ASAP7_75t_SL g681 ( .A(n_497), .Y(n_681) );
INVx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
AND2x2_ASAP7_75t_L g549 ( .A(n_498), .B(n_550), .Y(n_549) );
INVx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
AND2x2_ASAP7_75t_L g531 ( .A(n_499), .B(n_510), .Y(n_531) );
AND2x2_ASAP7_75t_L g617 ( .A(n_499), .B(n_533), .Y(n_617) );
INVx2_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
AND2x2_ASAP7_75t_L g587 ( .A(n_500), .B(n_520), .Y(n_587) );
OR2x2_ASAP7_75t_L g598 ( .A(n_500), .B(n_533), .Y(n_598) );
AND2x2_ASAP7_75t_L g624 ( .A(n_500), .B(n_533), .Y(n_624) );
HB1xp67_ASAP7_75t_L g669 ( .A(n_500), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_508), .B(n_624), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_508), .B(n_681), .Y(n_680) );
INVx2_ASAP7_75t_SL g508 ( .A(n_509), .Y(n_508) );
OR2x2_ASAP7_75t_L g597 ( .A(n_509), .B(n_598), .Y(n_597) );
AOI322xp5_ASAP7_75t_L g683 ( .A1(n_509), .A2(n_587), .A3(n_593), .B1(n_624), .B2(n_674), .C1(n_684), .C2(n_686), .Y(n_683) );
OR2x2_ASAP7_75t_L g509 ( .A(n_510), .B(n_520), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_510), .B(n_532), .Y(n_552) );
NOR2xp33_ASAP7_75t_L g580 ( .A(n_510), .B(n_533), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_510), .B(n_550), .Y(n_604) );
AND2x2_ASAP7_75t_L g658 ( .A(n_510), .B(n_624), .Y(n_658) );
INVx1_ASAP7_75t_L g662 ( .A(n_510), .Y(n_662) );
AND2x2_ASAP7_75t_L g674 ( .A(n_510), .B(n_520), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_510), .B(n_549), .Y(n_706) );
INVx4_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
AND2x2_ASAP7_75t_L g571 ( .A(n_511), .B(n_520), .Y(n_571) );
BUFx3_ASAP7_75t_L g585 ( .A(n_511), .Y(n_585) );
AND3x2_ASAP7_75t_L g667 ( .A(n_511), .B(n_647), .C(n_668), .Y(n_667) );
NAND3xp33_ASAP7_75t_L g530 ( .A(n_520), .B(n_531), .C(n_532), .Y(n_530) );
INVx1_ASAP7_75t_SL g550 ( .A(n_520), .Y(n_550) );
HB1xp67_ASAP7_75t_L g652 ( .A(n_520), .Y(n_652) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
AND2x2_ASAP7_75t_L g646 ( .A(n_531), .B(n_647), .Y(n_646) );
INVxp67_ASAP7_75t_L g653 ( .A(n_531), .Y(n_653) );
AND2x2_ASAP7_75t_L g691 ( .A(n_532), .B(n_669), .Y(n_691) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
BUFx3_ASAP7_75t_L g572 ( .A(n_533), .Y(n_572) );
AND2x2_ASAP7_75t_L g647 ( .A(n_533), .B(n_550), .Y(n_647) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_544), .B(n_545), .Y(n_543) );
OR2x2_ASAP7_75t_L g591 ( .A(n_544), .B(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g710 ( .A(n_544), .B(n_610), .Y(n_710) );
AND2x2_ASAP7_75t_L g724 ( .A(n_544), .B(n_546), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_545), .B(n_558), .Y(n_665) );
AND2x2_ASAP7_75t_L g712 ( .A(n_545), .B(n_713), .Y(n_712) );
AND2x2_ASAP7_75t_L g575 ( .A(n_546), .B(n_576), .Y(n_575) );
OR2x2_ASAP7_75t_L g592 ( .A(n_546), .B(n_558), .Y(n_592) );
INVx1_ASAP7_75t_L g602 ( .A(n_546), .Y(n_602) );
AND2x2_ASAP7_75t_L g633 ( .A(n_546), .B(n_558), .Y(n_633) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
OAI221xp5_ASAP7_75t_L g675 ( .A1(n_548), .A2(n_676), .B1(n_680), .B2(n_682), .C(n_683), .Y(n_675) );
NAND2xp5_ASAP7_75t_SL g548 ( .A(n_549), .B(n_551), .Y(n_548) );
AND2x2_ASAP7_75t_L g579 ( .A(n_549), .B(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
NOR2xp33_ASAP7_75t_L g729 ( .A(n_552), .B(n_586), .Y(n_729) );
AOI322xp5_ASAP7_75t_L g554 ( .A1(n_555), .A2(n_571), .A3(n_572), .B1(n_573), .B2(n_579), .C1(n_581), .C2(n_588), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_557), .B(n_570), .Y(n_556) );
NAND2x1p5_ASAP7_75t_L g609 ( .A(n_557), .B(n_610), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_557), .B(n_620), .Y(n_619) );
O2A1O1Ixp33_ASAP7_75t_L g643 ( .A1(n_557), .A2(n_570), .B(n_644), .C(n_645), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_557), .B(n_656), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_557), .B(n_614), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_557), .B(n_696), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_557), .B(n_724), .Y(n_723) );
BUFx3_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_558), .B(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_558), .B(n_602), .Y(n_601) );
OR2x2_ASAP7_75t_L g685 ( .A(n_558), .B(n_572), .Y(n_685) );
OA21x2_ASAP7_75t_L g558 ( .A1(n_559), .A2(n_562), .B(n_569), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
AO21x2_ASAP7_75t_L g576 ( .A1(n_560), .A2(n_577), .B(n_578), .Y(n_576) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx1_ASAP7_75t_L g577 ( .A(n_562), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_569), .Y(n_578) );
INVx1_ASAP7_75t_L g660 ( .A(n_570), .Y(n_660) );
OAI31xp33_ASAP7_75t_L g670 ( .A1(n_570), .A2(n_595), .A3(n_671), .B(n_673), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_570), .B(n_576), .Y(n_722) );
INVx1_ASAP7_75t_SL g583 ( .A(n_571), .Y(n_583) );
AND2x2_ASAP7_75t_L g616 ( .A(n_571), .B(n_617), .Y(n_616) );
AND2x2_ASAP7_75t_L g697 ( .A(n_571), .B(n_698), .Y(n_697) );
OR2x2_ASAP7_75t_L g582 ( .A(n_572), .B(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g607 ( .A(n_572), .Y(n_607) );
AND2x2_ASAP7_75t_L g634 ( .A(n_572), .B(n_587), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_572), .B(n_652), .Y(n_651) );
AND2x2_ASAP7_75t_L g726 ( .A(n_572), .B(n_674), .Y(n_726) );
NOR2xp33_ASAP7_75t_L g717 ( .A(n_574), .B(n_644), .Y(n_717) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g613 ( .A(n_576), .B(n_614), .Y(n_613) );
INVx1_ASAP7_75t_SL g631 ( .A(n_576), .Y(n_631) );
NAND2xp33_ASAP7_75t_SL g581 ( .A(n_582), .B(n_584), .Y(n_581) );
OAI211xp5_ASAP7_75t_SL g625 ( .A1(n_583), .A2(n_626), .B(n_632), .C(n_648), .Y(n_625) );
OR2x2_ASAP7_75t_L g700 ( .A(n_583), .B(n_681), .Y(n_700) );
OR2x2_ASAP7_75t_L g584 ( .A(n_585), .B(n_586), .Y(n_584) );
CKINVDCx16_ASAP7_75t_R g637 ( .A(n_585), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_585), .B(n_691), .Y(n_690) );
INVx1_ASAP7_75t_SL g586 ( .A(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g606 ( .A(n_587), .B(n_607), .Y(n_606) );
O2A1O1Ixp33_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_593), .B(n_596), .C(n_599), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
INVx1_ASAP7_75t_SL g640 ( .A(n_592), .Y(n_640) );
INVx1_ASAP7_75t_SL g593 ( .A(n_594), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_595), .B(n_633), .Y(n_638) );
INVx1_ASAP7_75t_L g644 ( .A(n_595), .Y(n_644) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
OR2x2_ASAP7_75t_L g603 ( .A(n_598), .B(n_604), .Y(n_603) );
OR2x2_ASAP7_75t_L g636 ( .A(n_598), .B(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g698 ( .A(n_598), .Y(n_698) );
AOI21xp33_ASAP7_75t_SL g599 ( .A1(n_600), .A2(n_601), .B(n_603), .Y(n_599) );
AOI21xp5_ASAP7_75t_L g611 ( .A1(n_601), .A2(n_612), .B(n_615), .Y(n_611) );
AOI211xp5_ASAP7_75t_L g605 ( .A1(n_606), .A2(n_608), .B(n_611), .C(n_618), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_606), .B(n_662), .Y(n_661) );
INVx1_ASAP7_75t_SL g608 ( .A(n_609), .Y(n_608) );
NOR2xp33_ASAP7_75t_L g699 ( .A(n_609), .B(n_700), .Y(n_699) );
INVx2_ASAP7_75t_SL g622 ( .A(n_610), .Y(n_622) );
OAI21xp5_ASAP7_75t_L g677 ( .A1(n_612), .A2(n_678), .B(n_679), .Y(n_677) );
INVx1_ASAP7_75t_SL g612 ( .A(n_613), .Y(n_612) );
INVx1_ASAP7_75t_SL g615 ( .A(n_616), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_617), .B(n_630), .Y(n_629) );
INVx1_ASAP7_75t_SL g642 ( .A(n_617), .Y(n_642) );
AOI21xp33_ASAP7_75t_SL g618 ( .A1(n_619), .A2(n_622), .B(n_623), .Y(n_618) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g673 ( .A(n_624), .B(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
NOR2xp33_ASAP7_75t_L g627 ( .A(n_628), .B(n_629), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_630), .B(n_656), .Y(n_682) );
AND2x2_ASAP7_75t_L g695 ( .A(n_630), .B(n_696), .Y(n_695) );
AND2x2_ASAP7_75t_L g709 ( .A(n_630), .B(n_710), .Y(n_709) );
AND2x2_ASAP7_75t_L g719 ( .A(n_630), .B(n_657), .Y(n_719) );
INVx2_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
AOI211xp5_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_634), .B(n_635), .C(n_643), .Y(n_632) );
INVx1_ASAP7_75t_L g679 ( .A(n_633), .Y(n_679) );
OAI22xp33_ASAP7_75t_L g635 ( .A1(n_636), .A2(n_638), .B1(n_639), .B2(n_641), .Y(n_635) );
OR2x2_ASAP7_75t_L g641 ( .A(n_637), .B(n_642), .Y(n_641) );
NAND2xp5_ASAP7_75t_SL g720 ( .A(n_637), .B(n_698), .Y(n_720) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g714 ( .A(n_647), .Y(n_714) );
AOI22xp33_ASAP7_75t_L g648 ( .A1(n_649), .A2(n_654), .B1(n_657), .B2(n_658), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
OR2x2_ASAP7_75t_L g650 ( .A(n_651), .B(n_653), .Y(n_650) );
INVx1_ASAP7_75t_L g732 ( .A(n_652), .Y(n_732) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g678 ( .A(n_656), .Y(n_678) );
OAI211xp5_ASAP7_75t_SL g659 ( .A1(n_660), .A2(n_661), .B(n_663), .C(n_670), .Y(n_659) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
NOR2xp33_ASAP7_75t_L g664 ( .A(n_665), .B(n_666), .Y(n_664) );
INVx2_ASAP7_75t_SL g666 ( .A(n_667), .Y(n_666) );
INVxp67_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVxp67_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
NOR2xp33_ASAP7_75t_L g684 ( .A(n_678), .B(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
NOR5xp2_ASAP7_75t_L g688 ( .A(n_689), .B(n_707), .C(n_715), .D(n_721), .E(n_727), .Y(n_688) );
OAI211xp5_ASAP7_75t_SL g689 ( .A1(n_690), .A2(n_692), .B(n_694), .C(n_701), .Y(n_689) );
INVxp67_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
AOI21xp5_ASAP7_75t_L g694 ( .A1(n_695), .A2(n_697), .B(n_699), .Y(n_694) );
OAI21xp33_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_704), .B(n_705), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
NOR2xp33_ASAP7_75t_L g716 ( .A(n_704), .B(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
AOI21xp33_ASAP7_75t_L g707 ( .A1(n_708), .A2(n_711), .B(n_714), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_SL g730 ( .A(n_710), .Y(n_730) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
AOI21xp5_ASAP7_75t_L g715 ( .A1(n_716), .A2(n_718), .B(n_720), .Y(n_715) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g745 ( .A(n_733), .Y(n_745) );
CKINVDCx16_ASAP7_75t_R g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_SL g740 ( .A(n_741), .Y(n_740) );
INVx2_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx3_ASAP7_75t_SL g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_SL g749 ( .A(n_750), .Y(n_749) );
CKINVDCx20_ASAP7_75t_R g752 ( .A(n_753), .Y(n_752) );
endmodule