module fake_jpeg_9305_n_295 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_295);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_295;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_288;
wire n_272;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_145;
wire n_20;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_213;
wire n_153;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_282;
wire n_96;

INVx4_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx8_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx8_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_42),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx3_ASAP7_75t_SL g50 ( 
.A(n_39),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_24),
.B(n_8),
.Y(n_42)
);

BUFx24_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_44),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_43),
.B(n_0),
.Y(n_45)
);

AOI32xp33_ASAP7_75t_L g83 ( 
.A1(n_45),
.A2(n_21),
.A3(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_83)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_47),
.B(n_51),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_36),
.A2(n_33),
.B1(n_31),
.B2(n_16),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_48),
.A2(n_68),
.B1(n_30),
.B2(n_29),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_43),
.A2(n_33),
.B1(n_31),
.B2(n_16),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_49),
.A2(n_28),
.B1(n_23),
.B2(n_21),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_26),
.Y(n_51)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_53),
.B(n_54),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_26),
.Y(n_54)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_56),
.B(n_64),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_26),
.Y(n_58)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_29),
.Y(n_59)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_29),
.Y(n_60)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_30),
.Y(n_63)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_22),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_34),
.B(n_27),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_65),
.B(n_67),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_34),
.B(n_27),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_36),
.A2(n_33),
.B1(n_16),
.B2(n_31),
.Y(n_68)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_70),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_68),
.A2(n_30),
.B1(n_27),
.B2(n_19),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_73),
.A2(n_63),
.B1(n_59),
.B2(n_58),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_45),
.A2(n_28),
.B1(n_19),
.B2(n_25),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_74),
.A2(n_46),
.B(n_60),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_75),
.Y(n_100)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_77),
.B(n_79),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_65),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_82),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_83),
.A2(n_46),
.B(n_51),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_67),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_84),
.B(n_47),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_85),
.A2(n_92),
.B1(n_50),
.B2(n_69),
.Y(n_111)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_87),
.Y(n_95)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_52),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_91),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_66),
.A2(n_23),
.B1(n_21),
.B2(n_32),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_80),
.A2(n_64),
.B1(n_53),
.B2(n_56),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_93),
.A2(n_90),
.B1(n_83),
.B2(n_87),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_94),
.A2(n_84),
.B(n_81),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_96),
.B(n_101),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_70),
.A2(n_66),
.B1(n_48),
.B2(n_69),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_98),
.A2(n_113),
.B1(n_99),
.B2(n_111),
.Y(n_122)
);

CKINVDCx14_ASAP7_75t_R g101 ( 
.A(n_86),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_102),
.B(n_103),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_80),
.B(n_45),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_104),
.B(n_109),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_89),
.A2(n_54),
.B(n_45),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_105),
.A2(n_111),
.B(n_17),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_74),
.B(n_50),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_107),
.B(n_90),
.C(n_78),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_86),
.B(n_57),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_89),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_110),
.B(n_114),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_79),
.A2(n_69),
.B1(n_44),
.B2(n_50),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_71),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_75),
.Y(n_115)
);

INVx4_ASAP7_75t_SL g125 ( 
.A(n_115),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_76),
.B(n_57),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_116),
.B(n_117),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_76),
.B(n_57),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_118),
.A2(n_94),
.B(n_105),
.Y(n_149)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_116),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_119),
.B(n_120),
.Y(n_158)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_117),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_109),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_121),
.B(n_123),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_122),
.A2(n_98),
.B1(n_107),
.B2(n_103),
.Y(n_146)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_97),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_114),
.B(n_78),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_126),
.B(n_128),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_101),
.B(n_81),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_127),
.B(n_142),
.Y(n_160)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_97),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_95),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_129),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_131),
.B(n_138),
.C(n_72),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_140),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_100),
.B(n_93),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_133),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_134),
.A2(n_23),
.B(n_82),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_99),
.A2(n_88),
.B1(n_77),
.B2(n_72),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_136),
.A2(n_44),
.B1(n_108),
.B2(n_106),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_104),
.B(n_23),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_113),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_96),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_141),
.B(n_102),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_110),
.B(n_17),
.Y(n_142)
);

BUFx2_ASAP7_75t_L g143 ( 
.A(n_100),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_143),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_125),
.A2(n_100),
.B1(n_112),
.B2(n_95),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_145),
.A2(n_146),
.B1(n_165),
.B2(n_132),
.Y(n_172)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_124),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_147),
.B(n_148),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_149),
.A2(n_167),
.B(n_170),
.Y(n_186)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_136),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_150),
.A2(n_152),
.B(n_155),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_151),
.B(n_91),
.C(n_82),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_121),
.B(n_0),
.Y(n_152)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_130),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_156),
.A2(n_120),
.B1(n_118),
.B2(n_125),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_112),
.Y(n_161)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_161),
.Y(n_171)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_137),
.Y(n_162)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_162),
.Y(n_177)
);

INVx13_ASAP7_75t_L g163 ( 
.A(n_129),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_163),
.Y(n_175)
);

AND2x6_ASAP7_75t_L g164 ( 
.A(n_139),
.B(n_14),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_164),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_140),
.A2(n_134),
.B1(n_122),
.B2(n_141),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_135),
.Y(n_166)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_166),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_119),
.B(n_0),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_128),
.B(n_15),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_169),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_172),
.A2(n_195),
.B(n_148),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_168),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_174),
.B(n_185),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_176),
.A2(n_178),
.B1(n_179),
.B2(n_182),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_150),
.A2(n_135),
.B1(n_131),
.B2(n_138),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_157),
.A2(n_143),
.B1(n_55),
.B2(n_62),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_144),
.A2(n_55),
.B1(n_62),
.B2(n_18),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_181),
.A2(n_187),
.B1(n_159),
.B2(n_163),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_157),
.A2(n_55),
.B1(n_62),
.B2(n_20),
.Y(n_182)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_158),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_184),
.B(n_191),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_154),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_144),
.A2(n_32),
.B1(n_20),
.B2(n_18),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_161),
.B(n_91),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_189),
.B(n_194),
.C(n_170),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_158),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_163),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_192),
.B(n_159),
.Y(n_200)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_156),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_193),
.B(n_167),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_149),
.A2(n_0),
.B(n_1),
.Y(n_195)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_196),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_190),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_197),
.B(n_202),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_198),
.B(n_201),
.C(n_204),
.Y(n_232)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_200),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_189),
.B(n_194),
.C(n_171),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_190),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_186),
.A2(n_176),
.B(n_195),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_203),
.B(n_186),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_178),
.B(n_146),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_179),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_205),
.B(n_208),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_172),
.B(n_151),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_206),
.B(n_216),
.C(n_198),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_184),
.B(n_166),
.Y(n_207)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_207),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_173),
.B(n_147),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_193),
.A2(n_164),
.B1(n_155),
.B2(n_162),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_209),
.A2(n_212),
.B1(n_215),
.B2(n_180),
.Y(n_222)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_192),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_210),
.B(n_214),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_175),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_182),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_181),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_217),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_221),
.B(n_227),
.C(n_229),
.Y(n_238)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_222),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g224 ( 
.A(n_210),
.Y(n_224)
);

BUFx2_ASAP7_75t_L g237 ( 
.A(n_224),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_225),
.B(n_11),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_204),
.B(n_188),
.Y(n_227)
);

BUFx24_ASAP7_75t_SL g228 ( 
.A(n_199),
.Y(n_228)
);

BUFx24_ASAP7_75t_SL g251 ( 
.A(n_228),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_206),
.B(n_188),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_201),
.B(n_183),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_230),
.A2(n_152),
.B(n_17),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_209),
.B(n_177),
.C(n_171),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_231),
.B(n_213),
.C(n_211),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_203),
.B(n_177),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_233),
.B(n_196),
.C(n_207),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_215),
.A2(n_183),
.B1(n_160),
.B2(n_175),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_234),
.A2(n_160),
.B1(n_169),
.B2(n_212),
.Y(n_239)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_239),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_240),
.B(n_244),
.C(n_249),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_236),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_241),
.B(n_247),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_242),
.B(n_243),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_232),
.B(n_187),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_232),
.B(n_207),
.C(n_153),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_218),
.A2(n_214),
.B1(n_153),
.B2(n_167),
.Y(n_245)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_245),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_246),
.A2(n_226),
.B(n_235),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_223),
.B(n_152),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_225),
.B(n_32),
.Y(n_249)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_250),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_253),
.A2(n_254),
.B(n_262),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_237),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_250),
.B(n_220),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_257),
.Y(n_264)
);

AO22x1_ASAP7_75t_L g259 ( 
.A1(n_248),
.A2(n_226),
.B1(n_219),
.B2(n_233),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_259),
.A2(n_9),
.B1(n_2),
.B2(n_3),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_244),
.A2(n_240),
.B(n_249),
.Y(n_262)
);

NOR2x1_ASAP7_75t_R g263 ( 
.A(n_238),
.B(n_230),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_263),
.B(n_10),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_260),
.A2(n_227),
.B1(n_237),
.B2(n_20),
.Y(n_265)
);

AOI322xp5_ASAP7_75t_L g280 ( 
.A1(n_265),
.A2(n_20),
.A3(n_18),
.B1(n_3),
.B2(n_5),
.C1(n_6),
.C2(n_7),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_263),
.A2(n_251),
.B(n_75),
.Y(n_266)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_266),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_258),
.B(n_17),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_268),
.B(n_270),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_10),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_258),
.B(n_17),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_252),
.B(n_32),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_271),
.B(n_252),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_257),
.B(n_9),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_272),
.A2(n_255),
.B(n_256),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_273),
.A2(n_253),
.B1(n_259),
.B2(n_3),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_275),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_267),
.B(n_262),
.C(n_261),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_276),
.A2(n_10),
.B(n_2),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_278),
.A2(n_273),
.B1(n_264),
.B2(n_269),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_279),
.A2(n_280),
.B1(n_281),
.B2(n_264),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_282),
.B(n_283),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_285),
.B(n_286),
.Y(n_289)
);

INVx11_ASAP7_75t_L g286 ( 
.A(n_281),
.Y(n_286)
);

OAI21xp33_ASAP7_75t_L g287 ( 
.A1(n_279),
.A2(n_5),
.B(n_7),
.Y(n_287)
);

NAND3xp33_ASAP7_75t_L g288 ( 
.A(n_287),
.B(n_15),
.C(n_7),
.Y(n_288)
);

AOI21x1_ASAP7_75t_L g291 ( 
.A1(n_288),
.A2(n_287),
.B(n_11),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_291),
.B(n_292),
.Y(n_293)
);

AOI21x1_ASAP7_75t_L g292 ( 
.A1(n_290),
.A2(n_276),
.B(n_289),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_293),
.A2(n_284),
.B(n_277),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_294),
.A2(n_274),
.B1(n_12),
.B2(n_15),
.Y(n_295)
);


endmodule