module fake_jpeg_9948_n_52 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_52);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_52;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx2_ASAP7_75t_L g7 ( 
.A(n_2),
.Y(n_7)
);

BUFx3_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

INVxp67_ASAP7_75t_SL g10 ( 
.A(n_3),
.Y(n_10)
);

BUFx16f_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

INVx5_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

INVx4_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_15),
.B(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_7),
.B(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

OR2x2_ASAP7_75t_L g18 ( 
.A(n_11),
.B(n_0),
.Y(n_18)
);

FAx1_ASAP7_75t_SL g25 ( 
.A(n_18),
.B(n_19),
.CI(n_22),
.CON(n_25),
.SN(n_25)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_7),
.B(n_2),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_SL g26 ( 
.A1(n_20),
.A2(n_24),
.B(n_8),
.Y(n_26)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_21),
.Y(n_30)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_L g23 ( 
.A1(n_13),
.A2(n_11),
.B1(n_10),
.B2(n_9),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_23),
.A2(n_14),
.B1(n_2),
.B2(n_5),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

AO21x1_ASAP7_75t_L g35 ( 
.A1(n_26),
.A2(n_29),
.B(n_18),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_19),
.A2(n_13),
.B1(n_14),
.B2(n_9),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_31),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_20),
.B(n_4),
.C(n_5),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_22),
.A2(n_6),
.B1(n_21),
.B2(n_24),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_24),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_35),
.B(n_38),
.Y(n_42)
);

HB1xp67_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_37),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_32),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_24),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_39),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_26),
.C(n_33),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_41),
.A2(n_33),
.B1(n_37),
.B2(n_31),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_SL g43 ( 
.A(n_34),
.B(n_35),
.Y(n_43)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_43),
.Y(n_48)
);

HB1xp67_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

OAI221xp5_ASAP7_75t_L g49 ( 
.A1(n_45),
.A2(n_47),
.B1(n_25),
.B2(n_44),
.C(n_27),
.Y(n_49)
);

MAJx2_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_25),
.C(n_42),
.Y(n_50)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

BUFx24_ASAP7_75t_SL g51 ( 
.A(n_49),
.Y(n_51)
);

OAI221xp5_ASAP7_75t_L g52 ( 
.A1(n_51),
.A2(n_50),
.B1(n_48),
.B2(n_25),
.C(n_45),
.Y(n_52)
);


endmodule