module fake_jpeg_2016_n_189 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_189);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_189;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx8_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_0),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_28),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_21),
.B(n_32),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_7),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_4),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_13),
.Y(n_59)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_10),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_62),
.Y(n_65)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

INVx6_ASAP7_75t_SL g66 ( 
.A(n_50),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_66),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_53),
.B(n_42),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_69),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_0),
.Y(n_68)
);

AOI21xp33_ASAP7_75t_L g77 ( 
.A1(n_68),
.A2(n_51),
.B(n_54),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_56),
.Y(n_69)
);

BUFx4f_ASAP7_75t_SL g70 ( 
.A(n_48),
.Y(n_70)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_71),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_72),
.Y(n_75)
);

NOR2x1_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_54),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_76),
.B(n_53),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_77),
.B(n_1),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_63),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_80),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_63),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_72),
.B(n_46),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_81),
.B(n_69),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_71),
.A2(n_55),
.B1(n_64),
.B2(n_48),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_83),
.A2(n_64),
.B1(n_55),
.B2(n_61),
.Y(n_96)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_85),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_88),
.B(n_89),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_82),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_82),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_91),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_73),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_93),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_57),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_94),
.Y(n_105)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_84),
.Y(n_95)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_95),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_96),
.B(n_97),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_78),
.B(n_59),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_98),
.B(n_100),
.Y(n_113)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_99),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_81),
.B(n_49),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_76),
.B(n_52),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_101),
.B(n_70),
.Y(n_117)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_74),
.Y(n_102)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_102),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_87),
.A2(n_80),
.B1(n_79),
.B2(n_75),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_107),
.A2(n_47),
.B1(n_44),
.B2(n_4),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_70),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_108),
.B(n_116),
.Y(n_132)
);

NAND3xp33_ASAP7_75t_SL g109 ( 
.A(n_93),
.B(n_66),
.C(n_52),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_109),
.B(n_112),
.Y(n_142)
);

AND2x2_ASAP7_75t_SL g110 ( 
.A(n_91),
.B(n_74),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_110),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_94),
.B(n_88),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_96),
.A2(n_73),
.B(n_58),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_115),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_102),
.B(n_75),
.Y(n_116)
);

NAND3xp33_ASAP7_75t_L g141 ( 
.A(n_117),
.B(n_3),
.C(n_5),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_95),
.B(n_60),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_119),
.B(n_41),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_99),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_120),
.B(n_2),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_114),
.B(n_86),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_122),
.B(n_125),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_105),
.A2(n_86),
.B1(n_61),
.B2(n_72),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_123),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_124),
.B(n_126),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_111),
.B(n_60),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_113),
.B(n_1),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_127),
.A2(n_135),
.B1(n_6),
.B2(n_7),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_104),
.B(n_47),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_128),
.B(n_133),
.Y(n_149)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_118),
.Y(n_129)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_129),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_107),
.A2(n_44),
.B1(n_40),
.B2(n_38),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_130),
.A2(n_128),
.B1(n_115),
.B2(n_131),
.Y(n_146)
);

BUFx24_ASAP7_75t_SL g133 ( 
.A(n_112),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_134),
.B(n_138),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_110),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_135)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_106),
.Y(n_137)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_137),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_110),
.B(n_121),
.Y(n_138)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_103),
.Y(n_139)
);

INVx13_ASAP7_75t_L g154 ( 
.A(n_139),
.Y(n_154)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_103),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_140),
.A2(n_141),
.B(n_6),
.Y(n_158)
);

HB1xp67_ASAP7_75t_SL g143 ( 
.A(n_142),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_143),
.A2(n_151),
.B(n_148),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_108),
.C(n_116),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_144),
.B(n_152),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_146),
.A2(n_159),
.B1(n_135),
.B2(n_139),
.Y(n_162)
);

NOR3xp33_ASAP7_75t_SL g147 ( 
.A(n_131),
.B(n_121),
.C(n_36),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_147),
.B(n_158),
.Y(n_164)
);

OAI22x1_ASAP7_75t_L g151 ( 
.A1(n_136),
.A2(n_31),
.B1(n_30),
.B2(n_27),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_151),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_132),
.B(n_26),
.C(n_25),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_130),
.B(n_20),
.C(n_19),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_155),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_127),
.B(n_9),
.C(n_10),
.Y(n_160)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_160),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_162),
.B(n_169),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_156),
.A2(n_9),
.B(n_11),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_163),
.A2(n_166),
.B(n_167),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_145),
.A2(n_149),
.B1(n_150),
.B2(n_156),
.Y(n_165)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_165),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_153),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_170),
.B(n_144),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_171),
.B(n_177),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_168),
.B(n_157),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_172),
.A2(n_161),
.B(n_155),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_164),
.B(n_152),
.Y(n_175)
);

AOI31xp67_ASAP7_75t_L g181 ( 
.A1(n_175),
.A2(n_12),
.A3(n_14),
.B(n_15),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_167),
.A2(n_147),
.B1(n_160),
.B2(n_154),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_178),
.B(n_181),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_171),
.B(n_161),
.C(n_163),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_179),
.B(n_176),
.C(n_173),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_183),
.B(n_180),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_184),
.B(n_182),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_185),
.B(n_177),
.C(n_174),
.Y(n_186)
);

AOI322xp5_ASAP7_75t_L g187 ( 
.A1(n_186),
.A2(n_15),
.A3(n_16),
.B1(n_17),
.B2(n_18),
.C1(n_154),
.C2(n_184),
.Y(n_187)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_187),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_188),
.B(n_16),
.Y(n_189)
);


endmodule