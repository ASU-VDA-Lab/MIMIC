module fake_jpeg_27794_n_168 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_168);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_168;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

OR2x2_ASAP7_75t_L g18 ( 
.A(n_12),
.B(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_18),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_38),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx3_ASAP7_75t_SL g36 ( 
.A(n_21),
.Y(n_36)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_39),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_41),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_18),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_46),
.Y(n_61)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_36),
.A2(n_28),
.B1(n_38),
.B2(n_22),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_47),
.A2(n_54),
.B1(n_58),
.B2(n_15),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_36),
.A2(n_28),
.B1(n_22),
.B2(n_20),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_51),
.A2(n_27),
.B1(n_19),
.B2(n_25),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_35),
.A2(n_28),
.B1(n_18),
.B2(n_26),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_33),
.B(n_30),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_41),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_23),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_57),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_23),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_33),
.A2(n_20),
.B1(n_29),
.B2(n_15),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_59),
.B(n_62),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_54),
.B(n_40),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_L g83 ( 
.A1(n_60),
.A2(n_65),
.B(n_25),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_56),
.Y(n_62)
);

CKINVDCx14_ASAP7_75t_R g81 ( 
.A(n_63),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_57),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_64),
.B(n_67),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g65 ( 
.A1(n_44),
.A2(n_29),
.B(n_30),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_66),
.A2(n_49),
.B1(n_48),
.B2(n_42),
.Y(n_89)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_68),
.B(n_70),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_43),
.B(n_19),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_43),
.B(n_27),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_73),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_58),
.A2(n_40),
.B1(n_39),
.B2(n_31),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_74),
.A2(n_49),
.B1(n_48),
.B2(n_42),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_46),
.B(n_39),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_75),
.B(n_50),
.Y(n_78)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_77),
.A2(n_74),
.B1(n_72),
.B2(n_73),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_78),
.B(n_79),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_69),
.B(n_31),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_83),
.A2(n_65),
.B(n_64),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_53),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_85),
.B(n_90),
.Y(n_99)
);

OAI21xp33_ASAP7_75t_L g87 ( 
.A1(n_61),
.A2(n_9),
.B(n_7),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_87),
.A2(n_60),
.B(n_75),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_89),
.A2(n_76),
.B1(n_59),
.B2(n_39),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_62),
.B(n_53),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_68),
.A2(n_17),
.B1(n_21),
.B2(n_24),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_91),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_61),
.B(n_24),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_92),
.B(n_79),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_63),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_95),
.B(n_109),
.Y(n_122)
);

HB1xp67_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_96),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_98),
.B(n_102),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_100),
.A2(n_105),
.B(n_84),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_101),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_84),
.B(n_60),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_107),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_106),
.A2(n_81),
.B1(n_77),
.B2(n_94),
.Y(n_113)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_108),
.A2(n_93),
.B1(n_37),
.B2(n_24),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_85),
.B(n_53),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_92),
.B(n_41),
.Y(n_110)
);

NAND3xp33_ASAP7_75t_L g115 ( 
.A(n_110),
.B(n_81),
.C(n_34),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_SL g126 ( 
.A(n_112),
.B(n_116),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_113),
.A2(n_124),
.B1(n_97),
.B2(n_16),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_115),
.B(n_117),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_86),
.C(n_94),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_100),
.A2(n_86),
.B(n_80),
.Y(n_117)
);

OR2x6_ASAP7_75t_L g118 ( 
.A(n_105),
.B(n_93),
.Y(n_118)
);

NAND2xp67_ASAP7_75t_SL g134 ( 
.A(n_118),
.B(n_97),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_99),
.B(n_37),
.C(n_34),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_121),
.B(n_104),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_104),
.A2(n_88),
.B(n_1),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_123),
.B(n_0),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_118),
.B(n_110),
.Y(n_125)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_125),
.Y(n_140)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_119),
.Y(n_127)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_127),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_128),
.B(n_16),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_118),
.A2(n_106),
.B1(n_99),
.B2(n_109),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_129),
.A2(n_131),
.B1(n_133),
.B2(n_134),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_114),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_130),
.Y(n_137)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_121),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_116),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_135),
.A2(n_136),
.B1(n_16),
.B2(n_6),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_126),
.B(n_122),
.C(n_118),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_138),
.B(n_141),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_126),
.B(n_122),
.C(n_120),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_128),
.B(n_111),
.C(n_115),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_142),
.B(n_145),
.Y(n_149)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_143),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_144),
.B(n_132),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_146),
.B(n_150),
.Y(n_157)
);

AOI31xp67_ASAP7_75t_L g150 ( 
.A1(n_140),
.A2(n_134),
.A3(n_125),
.B(n_129),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_138),
.B(n_0),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_151),
.B(n_145),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_139),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_152),
.B(n_2),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_149),
.B(n_142),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_153),
.B(n_148),
.C(n_10),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_150),
.A2(n_137),
.B(n_147),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_154),
.B(n_156),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_155),
.B(n_151),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_159),
.B(n_160),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_157),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_161),
.A2(n_3),
.B1(n_5),
.B2(n_153),
.Y(n_163)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_163),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_158),
.A2(n_161),
.B1(n_11),
.B2(n_13),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_164),
.B(n_3),
.Y(n_166)
);

A2O1A1Ixp33_ASAP7_75t_SL g167 ( 
.A1(n_166),
.A2(n_163),
.B(n_5),
.C(n_162),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_167),
.B(n_165),
.Y(n_168)
);


endmodule