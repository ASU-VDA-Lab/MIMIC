module real_jpeg_7257_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_288;
wire n_78;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_470;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_323;
wire n_176;
wire n_166;
wire n_215;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_438;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g56 ( 
.A(n_0),
.Y(n_56)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_1),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_1),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_2),
.B(n_191),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_2),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_2),
.B(n_234),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_2),
.B(n_392),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_2),
.B(n_409),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_2),
.B(n_251),
.Y(n_424)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_4),
.Y(n_141)
);

INVx8_ASAP7_75t_L g174 ( 
.A(n_4),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_4),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_5),
.B(n_176),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_5),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_5),
.B(n_238),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_5),
.B(n_286),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_5),
.B(n_438),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_6),
.B(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_6),
.B(n_223),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_6),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_6),
.B(n_288),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_6),
.B(n_304),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_6),
.B(n_339),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_6),
.B(n_374),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_6),
.B(n_405),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_7),
.B(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_7),
.B(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_7),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_7),
.B(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_7),
.B(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_7),
.B(n_172),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_7),
.Y(n_214)
);

AND2x2_ASAP7_75t_SL g270 ( 
.A(n_7),
.B(n_271),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_8),
.Y(n_89)
);

BUFx5_ASAP7_75t_L g145 ( 
.A(n_8),
.Y(n_145)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_8),
.Y(n_192)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_10),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_10),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_10),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_10),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_10),
.Y(n_286)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_10),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_11),
.B(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_11),
.B(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_11),
.B(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_11),
.B(n_62),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_11),
.B(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_11),
.B(n_188),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_11),
.B(n_251),
.Y(n_250)
);

AND2x2_ASAP7_75t_SL g266 ( 
.A(n_11),
.B(n_267),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_12),
.B(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_12),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_12),
.B(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_12),
.B(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_12),
.B(n_113),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_12),
.B(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_12),
.B(n_169),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_12),
.B(n_198),
.Y(n_197)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_13),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_13),
.Y(n_114)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_13),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_14),
.B(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_14),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_14),
.B(n_107),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_14),
.B(n_143),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_14),
.B(n_147),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_15),
.B(n_203),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_15),
.B(n_28),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_15),
.B(n_243),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_15),
.B(n_62),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_15),
.B(n_379),
.Y(n_378)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_15),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_15),
.B(n_426),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_15),
.B(n_384),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_158),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_157),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_97),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_20),
.B(n_97),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_79),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_45),
.B2(n_46),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_30),
.C(n_42),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_24),
.A2(n_25),
.B1(n_42),
.B2(n_83),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_29),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_SL g81 ( 
.A(n_30),
.B(n_82),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_36),
.C(n_39),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_31),
.A2(n_36),
.B1(n_135),
.B2(n_136),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_31),
.Y(n_136)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_35),
.Y(n_178)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_36),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_36),
.A2(n_135),
.B1(n_274),
.B2(n_275),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_36),
.B(n_140),
.C(n_183),
.Y(n_321)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_38),
.Y(n_126)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_38),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_39),
.A2(n_133),
.B1(n_134),
.B2(n_137),
.Y(n_132)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_39),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_40),
.B(n_41),
.Y(n_39)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_42),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_42),
.A2(n_83),
.B1(n_338),
.B2(n_342),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_42),
.B(n_342),
.C(n_359),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_42),
.A2(n_83),
.B1(n_146),
.B2(n_362),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_44),
.Y(n_104)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_44),
.Y(n_235)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_47),
.A2(n_48),
.B1(n_67),
.B2(n_68),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_51),
.B1(n_65),
.B2(n_66),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_49),
.Y(n_65)
);

CKINVDCx14_ASAP7_75t_R g66 ( 
.A(n_51),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_57),
.C(n_59),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_52),
.B(n_85),
.C(n_90),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_52),
.A2(n_59),
.B1(n_60),
.B2(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_52),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_52),
.A2(n_90),
.B1(n_91),
.B2(n_96),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_52),
.A2(n_96),
.B1(n_221),
.B2(n_226),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_52),
.B(n_112),
.C(n_222),
.Y(n_247)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_55),
.Y(n_381)
);

INVx5_ASAP7_75t_L g398 ( 
.A(n_55),
.Y(n_398)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_56),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_56),
.Y(n_182)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_56),
.Y(n_269)
);

BUFx5_ASAP7_75t_L g410 ( 
.A(n_56),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_57),
.B(n_95),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_59),
.A2(n_60),
.B1(n_71),
.B2(n_72),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_59),
.A2(n_60),
.B1(n_195),
.B2(n_196),
.Y(n_194)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_60),
.B(n_197),
.C(n_202),
.Y(n_283)
);

OR2x2_ASAP7_75t_SL g60 ( 
.A(n_61),
.B(n_64),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

OR2x2_ASAP7_75t_SL g72 ( 
.A(n_64),
.B(n_73),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_64),
.B(n_92),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g140 ( 
.A(n_64),
.B(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_69),
.A2(n_70),
.B1(n_75),
.B2(n_78),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_71),
.A2(n_72),
.B1(n_265),
.B2(n_272),
.Y(n_264)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_72),
.B(n_344),
.C(n_345),
.Y(n_343)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx5_ASAP7_75t_L g244 ( 
.A(n_74),
.Y(n_244)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_75),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_75),
.A2(n_78),
.B1(n_121),
.B2(n_122),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_75),
.B(n_123),
.C(n_131),
.Y(n_152)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_84),
.C(n_94),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_80),
.A2(n_81),
.B1(n_155),
.B2(n_156),
.Y(n_154)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_83),
.B(n_139),
.C(n_146),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g155 ( 
.A(n_84),
.B(n_94),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_85),
.B(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_90),
.A2(n_91),
.B1(n_106),
.B2(n_110),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_90),
.A2(n_91),
.B1(n_183),
.B2(n_276),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_91),
.B(n_102),
.C(n_106),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_91),
.B(n_180),
.C(n_183),
.Y(n_179)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_93),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_148),
.C(n_154),
.Y(n_97)
);

FAx1_ASAP7_75t_SL g482 ( 
.A(n_98),
.B(n_148),
.CI(n_154),
.CON(n_482),
.SN(n_482)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_132),
.C(n_138),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_99),
.A2(n_100),
.B1(n_485),
.B2(n_486),
.Y(n_484)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_111),
.C(n_120),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_101),
.B(n_353),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_105),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_104),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_106),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_106),
.B(n_140),
.C(n_142),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_106),
.B(n_302),
.C(n_306),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_106),
.A2(n_110),
.B1(n_140),
.B2(n_277),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_106),
.A2(n_110),
.B1(n_386),
.B2(n_387),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_107),
.Y(n_216)
);

INVx3_ASAP7_75t_L g440 ( 
.A(n_107),
.Y(n_440)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_108),
.Y(n_417)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_108),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_111),
.B(n_120),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_115),
.C(n_116),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_112),
.A2(n_222),
.B1(n_224),
.B2(n_225),
.Y(n_221)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_112),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_112),
.A2(n_224),
.B1(n_323),
.B2(n_324),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_SL g323 ( 
.A(n_115),
.B(n_116),
.Y(n_323)
);

INVx4_ASAP7_75t_SL g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_119),
.Y(n_129)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_127),
.B1(n_130),
.B2(n_131),
.Y(n_122)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_123),
.Y(n_130)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx8_ASAP7_75t_L g392 ( 
.A(n_125),
.Y(n_392)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_126),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g131 ( 
.A(n_127),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_127),
.B(n_250),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_127),
.B(n_250),
.C(n_254),
.Y(n_263)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_132),
.B(n_138),
.Y(n_485)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_139),
.B(n_361),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_140),
.A2(n_183),
.B1(n_276),
.B2(n_277),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_140),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_140),
.A2(n_277),
.B1(n_390),
.B2(n_391),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_142),
.A2(n_328),
.B1(n_329),
.B2(n_330),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_142),
.Y(n_328)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_144),
.B(n_218),
.Y(n_217)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx6_ASAP7_75t_L g289 ( 
.A(n_145),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_146),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_152),
.C(n_153),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_149),
.A2(n_150),
.B1(n_488),
.B2(n_489),
.Y(n_487)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_152),
.B(n_153),
.Y(n_489)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_155),
.Y(n_156)
);

AOI21x1_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_480),
.B(n_494),
.Y(n_158)
);

AO21x1_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_348),
.B(n_364),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_315),
.B(n_347),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_292),
.B(n_314),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_162),
.B(n_478),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_258),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_163),
.B(n_258),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_219),
.C(n_245),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_164),
.B(n_313),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_193),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_165),
.B(n_194),
.C(n_205),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_179),
.C(n_184),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_166),
.B(n_310),
.Y(n_309)
);

BUFx24_ASAP7_75t_SL g498 ( 
.A(n_166),
.Y(n_498)
);

FAx1_ASAP7_75t_SL g166 ( 
.A(n_167),
.B(n_171),
.CI(n_175),
.CON(n_166),
.SN(n_166)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_167),
.B(n_171),
.C(n_175),
.Y(n_257)
);

BUFx2_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

BUFx5_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

BUFx8_ASAP7_75t_L g376 ( 
.A(n_170),
.Y(n_376)
);

INVx8_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_174),
.Y(n_188)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_174),
.Y(n_200)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_174),
.Y(n_421)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_179),
.A2(n_184),
.B1(n_185),
.B2(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_179),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_180),
.B(n_300),
.Y(n_299)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_183),
.Y(n_276)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_189),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_186),
.A2(n_187),
.B1(n_189),
.B2(n_190),
.Y(n_308)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_205),
.Y(n_193)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_197),
.A2(n_201),
.B1(n_202),
.B2(n_204),
.Y(n_196)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_197),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_197),
.A2(n_204),
.B1(n_232),
.B2(n_233),
.Y(n_399)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_202),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_204),
.B(n_232),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_212),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_206),
.A2(n_207),
.B(n_208),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_206),
.B(n_213),
.C(n_217),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_209),
.B(n_211),
.Y(n_208)
);

INVx8_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_211),
.B(n_417),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_217),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_218),
.B(n_383),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_218),
.B(n_395),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_218),
.B(n_431),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_219),
.B(n_245),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_227),
.C(n_229),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_220),
.A2(n_227),
.B1(n_228),
.B2(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_220),
.Y(n_297)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_221),
.Y(n_226)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_222),
.Y(n_225)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_SL g295 ( 
.A(n_229),
.B(n_296),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_236),
.C(n_241),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_230),
.A2(n_231),
.B1(n_467),
.B2(n_468),
.Y(n_466)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_236),
.A2(n_237),
.B1(n_241),
.B2(n_242),
.Y(n_468)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx5_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx5_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx4_ASAP7_75t_SL g243 ( 
.A(n_244),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_257),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_247),
.B(n_248),
.C(n_257),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_249),
.B(n_254),
.Y(n_248)
);

INVx4_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx4_ASAP7_75t_L g271 ( 
.A(n_253),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_259),
.B(n_261),
.C(n_291),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_261),
.A2(n_278),
.B1(n_290),
.B2(n_291),
.Y(n_260)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_261),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_273),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_263),
.B(n_264),
.C(n_273),
.Y(n_332)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_265),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_270),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_266),
.Y(n_344)
);

INVx4_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx4_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_270),
.Y(n_345)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_277),
.B(n_390),
.Y(n_389)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_278),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_SL g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_279),
.B(n_281),
.C(n_282),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_283),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_287),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_285),
.B(n_287),
.C(n_335),
.Y(n_334)
);

INVx4_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_312),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_293),
.B(n_312),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_298),
.C(n_309),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_294),
.A2(n_295),
.B1(n_473),
.B2(n_474),
.Y(n_472)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_SL g473 ( 
.A(n_298),
.B(n_309),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_301),
.C(n_308),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_299),
.B(n_460),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_301),
.B(n_308),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_302),
.A2(n_303),
.B1(n_306),
.B2(n_307),
.Y(n_387)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx3_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx3_ASAP7_75t_L g384 ( 
.A(n_305),
.Y(n_384)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_316),
.B(n_348),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_318),
.Y(n_316)
);

OR2x2_ASAP7_75t_L g347 ( 
.A(n_317),
.B(n_318),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_318),
.B(n_349),
.Y(n_348)
);

OR2x2_ASAP7_75t_L g479 ( 
.A(n_318),
.B(n_349),
.Y(n_479)
);

FAx1_ASAP7_75t_SL g318 ( 
.A(n_319),
.B(n_331),
.CI(n_346),
.CON(n_318),
.SN(n_318)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_327),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_321),
.A2(n_322),
.B1(n_325),
.B2(n_326),
.Y(n_320)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_321),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_321),
.B(n_326),
.C(n_327),
.Y(n_356)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_322),
.Y(n_326)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_323),
.Y(n_324)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_329),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_SL g331 ( 
.A(n_332),
.B(n_333),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_332),
.B(n_334),
.C(n_336),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_336),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_343),
.Y(n_336)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_338),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_343),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_351),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_350),
.B(n_352),
.C(n_354),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_354),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_355),
.A2(n_356),
.B1(n_357),
.B2(n_363),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_355),
.B(n_358),
.C(n_360),
.Y(n_490)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_357),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_SL g357 ( 
.A(n_358),
.B(n_360),
.Y(n_357)
);

OAI31xp33_ASAP7_75t_L g364 ( 
.A1(n_365),
.A2(n_476),
.A3(n_477),
.B(n_479),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g365 ( 
.A1(n_366),
.A2(n_470),
.B(n_475),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_SL g366 ( 
.A1(n_367),
.A2(n_455),
.B(n_469),
.Y(n_366)
);

AOI21xp5_ASAP7_75t_L g367 ( 
.A1(n_368),
.A2(n_412),
.B(n_454),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_369),
.B(n_400),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_369),
.B(n_400),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_388),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_385),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_371),
.B(n_385),
.C(n_388),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_377),
.C(n_382),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_372),
.A2(n_373),
.B1(n_377),
.B2(n_378),
.Y(n_402)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx8_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx3_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_SL g401 ( 
.A(n_382),
.B(n_402),
.Y(n_401)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_SL g388 ( 
.A(n_389),
.B(n_393),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_389),
.B(n_464),
.C(n_465),
.Y(n_463)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_399),
.Y(n_393)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_394),
.Y(n_464)
);

INVx1_ASAP7_75t_SL g395 ( 
.A(n_396),
.Y(n_395)
);

BUFx3_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx5_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_399),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_403),
.C(n_411),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_401),
.B(n_451),
.Y(n_450)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_403),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_403),
.A2(n_411),
.B1(n_446),
.B2(n_452),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_SL g403 ( 
.A(n_404),
.B(n_408),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_404),
.Y(n_444)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx3_ASAP7_75t_L g431 ( 
.A(n_407),
.Y(n_431)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_408),
.Y(n_445)
);

INVx5_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_411),
.Y(n_452)
);

OAI21xp5_ASAP7_75t_L g412 ( 
.A1(n_413),
.A2(n_448),
.B(n_453),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_L g413 ( 
.A1(n_414),
.A2(n_433),
.B(n_447),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_L g414 ( 
.A1(n_415),
.A2(n_422),
.B(n_432),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_418),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_419),
.B(n_420),
.Y(n_418)
);

INVx4_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_SL g422 ( 
.A(n_423),
.B(n_430),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_423),
.B(n_430),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g423 ( 
.A1(n_424),
.A2(n_425),
.B(n_429),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_424),
.B(n_425),
.Y(n_429)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

INVx4_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_429),
.A2(n_435),
.B1(n_441),
.B2(n_442),
.Y(n_434)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_429),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_434),
.B(n_443),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_434),
.B(n_443),
.Y(n_447)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_435),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_SL g435 ( 
.A(n_436),
.B(n_437),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_SL g449 ( 
.A1(n_436),
.A2(n_437),
.B(n_441),
.Y(n_449)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

HB1xp67_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_SL g443 ( 
.A1(n_444),
.A2(n_445),
.B(n_446),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_449),
.B(n_450),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_449),
.B(n_450),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_456),
.B(n_457),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_456),
.B(n_457),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_L g457 ( 
.A1(n_458),
.A2(n_459),
.B1(n_461),
.B2(n_462),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_458),
.B(n_463),
.C(n_466),
.Y(n_471)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_463),
.B(n_466),
.Y(n_462)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_471),
.B(n_472),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_471),
.B(n_472),
.Y(n_475)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_473),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_481),
.B(n_491),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_SL g494 ( 
.A1(n_481),
.A2(n_495),
.B(n_496),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_482),
.B(n_483),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_482),
.B(n_483),
.Y(n_496)
);

BUFx24_ASAP7_75t_SL g497 ( 
.A(n_482),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_484),
.B(n_487),
.C(n_490),
.Y(n_483)
);

FAx1_ASAP7_75t_SL g493 ( 
.A(n_484),
.B(n_487),
.CI(n_490),
.CON(n_493),
.SN(n_493)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_485),
.Y(n_486)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_492),
.B(n_493),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_492),
.B(n_493),
.Y(n_495)
);

BUFx24_ASAP7_75t_SL g500 ( 
.A(n_493),
.Y(n_500)
);


endmodule