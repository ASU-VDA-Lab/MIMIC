module fake_jpeg_8947_n_79 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_79);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_79;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

INVx2_ASAP7_75t_SL g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_22),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

CKINVDCx14_ASAP7_75t_R g34 ( 
.A(n_25),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_27),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_37),
.A2(n_2),
.B(n_3),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_0),
.Y(n_38)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_1),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_40),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_33),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_44),
.Y(n_50)
);

INVx6_ASAP7_75t_SL g43 ( 
.A(n_27),
.Y(n_43)
);

CKINVDCx5p33_ASAP7_75t_R g63 ( 
.A(n_43),
.Y(n_63)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_8),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_36),
.B(n_34),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_64),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_37),
.A2(n_34),
.B1(n_29),
.B2(n_4),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_48),
.A2(n_52),
.B(n_61),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_45),
.A2(n_18),
.B1(n_26),
.B2(n_23),
.Y(n_49)
);

O2A1O1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_49),
.A2(n_53),
.B(n_55),
.C(n_62),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_41),
.A2(n_3),
.B1(n_4),
.B2(n_7),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_58),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_45),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_14),
.Y(n_57)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_15),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_38),
.B(n_17),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_19),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_38),
.B(n_21),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_66),
.B(n_59),
.Y(n_71)
);

NOR3xp33_ASAP7_75t_L g72 ( 
.A(n_71),
.B(n_67),
.C(n_47),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_72),
.B(n_50),
.C(n_68),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_73),
.A2(n_63),
.B1(n_65),
.B2(n_55),
.Y(n_74)
);

MAJx2_ASAP7_75t_L g75 ( 
.A(n_74),
.B(n_70),
.C(n_53),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_75),
.A2(n_60),
.B(n_51),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_65),
.C(n_69),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_56),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_78),
.B(n_60),
.Y(n_79)
);


endmodule