module real_jpeg_2269_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_167;
wire n_202;
wire n_128;
wire n_216;
wire n_179;
wire n_213;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

INVx2_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_1),
.A2(n_40),
.B1(n_42),
.B2(n_43),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_1),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_1),
.A2(n_43),
.B1(n_59),
.B2(n_60),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

OAI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_3),
.A2(n_25),
.B1(n_26),
.B2(n_66),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_3),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_3),
.A2(n_32),
.B1(n_66),
.B2(n_71),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_3),
.A2(n_59),
.B1(n_60),
.B2(n_66),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_3),
.A2(n_40),
.B1(n_42),
.B2(n_66),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_4),
.A2(n_59),
.B1(n_60),
.B2(n_86),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_4),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_4),
.A2(n_25),
.B1(n_26),
.B2(n_86),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_4),
.A2(n_40),
.B1(n_42),
.B2(n_86),
.Y(n_151)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_5),
.Y(n_58)
);

OAI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_6),
.A2(n_40),
.B1(n_42),
.B2(n_83),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_6),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_7),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_7),
.B(n_127),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_7),
.B(n_58),
.C(n_60),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_7),
.B(n_57),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_7),
.B(n_42),
.C(n_89),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_7),
.A2(n_36),
.B1(n_59),
.B2(n_60),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_7),
.B(n_46),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_7),
.B(n_93),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_7),
.A2(n_25),
.B1(n_26),
.B2(n_36),
.Y(n_221)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx16f_ASAP7_75t_L g89 ( 
.A(n_9),
.Y(n_89)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_11),
.A2(n_25),
.B1(n_26),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_11),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_11),
.A2(n_32),
.B1(n_54),
.B2(n_71),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_11),
.A2(n_54),
.B1(n_59),
.B2(n_60),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_11),
.A2(n_40),
.B1(n_42),
.B2(n_54),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_12),
.A2(n_40),
.B1(n_42),
.B2(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_12),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_13),
.A2(n_40),
.B1(n_42),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_13),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_13),
.A2(n_49),
.B1(n_59),
.B2(n_60),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_15),
.A2(n_32),
.B1(n_70),
.B2(n_71),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_15),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_15),
.A2(n_25),
.B1(n_26),
.B2(n_70),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_15),
.A2(n_59),
.B1(n_60),
.B2(n_70),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_15),
.A2(n_40),
.B1(n_42),
.B2(n_70),
.Y(n_206)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_16),
.Y(n_61)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_136),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_134),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_107),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_20),
.B(n_107),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_79),
.C(n_94),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_21),
.B(n_139),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_50),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_22),
.B(n_51),
.C(n_78),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_38),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_23),
.A2(n_24),
.B1(n_38),
.B2(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

AOI32xp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_29),
.A3(n_32),
.B1(n_34),
.B2(n_37),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_25),
.A2(n_26),
.B1(n_58),
.B2(n_62),
.Y(n_63)
);

OA22x2_ASAP7_75t_L g72 ( 
.A1(n_25),
.A2(n_26),
.B1(n_29),
.B2(n_30),
.Y(n_72)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp33_ASAP7_75t_SL g37 ( 
.A(n_26),
.B(n_30),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_26),
.B(n_167),
.Y(n_166)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_29),
.A2(n_30),
.B1(n_32),
.B2(n_71),
.Y(n_77)
);

INVx4_ASAP7_75t_SL g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_32),
.B(n_36),
.Y(n_35)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

O2A1O1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_32),
.A2(n_35),
.B(n_36),
.C(n_103),
.Y(n_102)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_36),
.A2(n_81),
.B(n_182),
.Y(n_203)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_38),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_44),
.B1(n_45),
.B2(n_47),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_39),
.A2(n_44),
.B1(n_45),
.B2(n_151),
.Y(n_150)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

OA22x2_ASAP7_75t_L g91 ( 
.A1(n_40),
.A2(n_42),
.B1(n_89),
.B2(n_90),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_42),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_42),
.B(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_44),
.A2(n_45),
.B1(n_114),
.B2(n_115),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_44),
.B(n_171),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_44),
.A2(n_180),
.B(n_181),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_44),
.A2(n_45),
.B1(n_180),
.B2(n_211),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_45),
.A2(n_151),
.B(n_169),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_45),
.B(n_171),
.Y(n_182)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_46),
.A2(n_48),
.B1(n_81),
.B2(n_82),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_46),
.A2(n_170),
.B(n_206),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_52),
.B1(n_67),
.B2(n_78),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_55),
.B(n_64),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_53),
.A2(n_55),
.B1(n_105),
.B2(n_106),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_55),
.A2(n_64),
.B(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_56),
.B(n_65),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_57),
.B(n_63),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_57),
.Y(n_106)
);

AO22x1_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_59),
.B1(n_60),
.B2(n_62),
.Y(n_57)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_58),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_L g88 ( 
.A1(n_59),
.A2(n_60),
.B1(n_89),
.B2(n_90),
.Y(n_88)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_60),
.B(n_194),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_72),
.B(n_73),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_69),
.A2(n_76),
.B1(n_126),
.B2(n_127),
.Y(n_125)
);

AND2x2_ASAP7_75t_SL g76 ( 
.A(n_72),
.B(n_77),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_72),
.B(n_75),
.Y(n_101)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_72),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_76),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_76),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_79),
.B(n_94),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_84),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_80),
.B(n_84),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_82),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_87),
.B1(n_92),
.B2(n_93),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_87),
.B(n_98),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_87),
.A2(n_92),
.B1(n_93),
.B2(n_118),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_87),
.A2(n_160),
.B(n_162),
.Y(n_159)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_87),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_91),
.Y(n_87)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_89),
.Y(n_90)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_91),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_91),
.A2(n_96),
.B(n_97),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_91),
.A2(n_97),
.B(n_188),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_91),
.A2(n_161),
.B1(n_188),
.B2(n_196),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_93),
.B(n_98),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_99),
.C(n_104),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_95),
.B(n_104),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_99),
.A2(n_100),
.B1(n_142),
.B2(n_143),
.Y(n_141)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_101),
.B(n_102),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_105),
.A2(n_106),
.B(n_131),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_106),
.A2(n_130),
.B(n_131),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_109),
.B1(n_110),
.B2(n_111),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_SL g111 ( 
.A(n_112),
.B(n_121),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_117),
.B1(n_119),
.B2(n_120),
.Y(n_112)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_113),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_117),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_123),
.B1(n_132),
.B2(n_133),
.Y(n_121)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_122),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_123),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_125),
.B1(n_128),
.B2(n_129),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_152),
.B(n_232),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_138),
.B(n_140),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_138),
.B(n_140),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_144),
.C(n_146),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_141),
.B(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_142),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_144),
.B(n_146),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_148),
.C(n_150),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_147),
.B(n_157),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_148),
.A2(n_149),
.B1(n_150),
.B2(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_150),
.Y(n_158)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_174),
.B(n_231),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_172),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_155),
.B(n_172),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_159),
.C(n_164),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_156),
.B(n_228),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_159),
.B(n_164),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_163),
.A2(n_196),
.B(n_197),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_168),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_165),
.A2(n_166),
.B1(n_168),
.B2(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_168),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_226),
.B(n_230),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_216),
.B(n_225),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_198),
.B(n_215),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_178),
.B(n_191),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_178),
.B(n_191),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_183),
.B1(n_189),
.B2(n_190),
.Y(n_178)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_179),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_183),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_185),
.B1(n_186),
.B2(n_187),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_185),
.B(n_186),
.C(n_189),
.Y(n_217)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_195),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_192),
.A2(n_193),
.B1(n_195),
.B2(n_213),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_195),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_209),
.B(n_214),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_204),
.B(n_208),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_203),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_205),
.B(n_207),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_205),
.B(n_207),
.Y(n_208)
);

CKINVDCx14_ASAP7_75t_R g211 ( 
.A(n_206),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_212),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_210),
.B(n_212),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_217),
.B(n_218),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_223),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_222),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_220),
.B(n_222),
.C(n_223),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_227),
.B(n_229),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_227),
.B(n_229),
.Y(n_230)
);


endmodule