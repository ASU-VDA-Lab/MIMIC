module fake_netlist_6_4625_n_1663 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1663);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1663;

wire n_992;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_1214;
wire n_928;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_683;
wire n_527;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1373;
wire n_1292;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g155 ( 
.A(n_90),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_80),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_50),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_137),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_39),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_79),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_76),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_106),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_38),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_133),
.Y(n_164)
);

BUFx10_ASAP7_75t_L g165 ( 
.A(n_130),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_121),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_140),
.Y(n_167)
);

BUFx10_ASAP7_75t_L g168 ( 
.A(n_103),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_5),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_123),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_66),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_33),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_126),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_64),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_55),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_112),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_138),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_41),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_129),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_113),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_44),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_111),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_149),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_41),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_45),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_25),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g187 ( 
.A(n_151),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_51),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_65),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_81),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_59),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_87),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_73),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_56),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_58),
.Y(n_195)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_43),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_93),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_31),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_75),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_34),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_28),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_125),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_23),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_46),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_97),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_143),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_52),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_5),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_108),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_102),
.Y(n_210)
);

BUFx2_ASAP7_75t_L g211 ( 
.A(n_148),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_94),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_47),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_48),
.Y(n_214)
);

BUFx10_ASAP7_75t_L g215 ( 
.A(n_14),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_31),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_35),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_96),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_82),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_4),
.Y(n_220)
);

BUFx10_ASAP7_75t_L g221 ( 
.A(n_109),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g222 ( 
.A(n_120),
.Y(n_222)
);

BUFx8_ASAP7_75t_SL g223 ( 
.A(n_86),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_45),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_124),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_26),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_43),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_15),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_127),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_11),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_85),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_144),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_35),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_49),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_117),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_100),
.Y(n_236)
);

BUFx10_ASAP7_75t_L g237 ( 
.A(n_71),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_21),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_132),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_78),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_107),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_42),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_34),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_135),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_15),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_77),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_12),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_26),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_25),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_146),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_17),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_20),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_119),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_21),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_61),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_70),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_29),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_22),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_57),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_83),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_48),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_24),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_152),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_3),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_116),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_84),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_36),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_29),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_33),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_40),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_30),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_50),
.Y(n_272)
);

BUFx10_ASAP7_75t_L g273 ( 
.A(n_23),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_6),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_131),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_4),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_104),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_27),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_0),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_0),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_40),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_101),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_39),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_63),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_92),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_6),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_46),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_42),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_62),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_14),
.Y(n_290)
);

BUFx5_ASAP7_75t_L g291 ( 
.A(n_99),
.Y(n_291)
);

BUFx2_ASAP7_75t_L g292 ( 
.A(n_122),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_67),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_128),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_8),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_134),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_20),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_53),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_91),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_7),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_98),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_22),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_95),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_19),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_89),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_154),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_139),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_283),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_188),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_227),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_227),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_196),
.Y(n_312)
);

INVxp67_ASAP7_75t_SL g313 ( 
.A(n_211),
.Y(n_313)
);

BUFx2_ASAP7_75t_L g314 ( 
.A(n_157),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_227),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_223),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_227),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_227),
.Y(n_318)
);

INVxp67_ASAP7_75t_SL g319 ( 
.A(n_292),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_215),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_158),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_238),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_238),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_238),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_238),
.Y(n_325)
);

BUFx2_ASAP7_75t_L g326 ( 
.A(n_157),
.Y(n_326)
);

BUFx3_ASAP7_75t_L g327 ( 
.A(n_175),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_188),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_193),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_238),
.Y(n_330)
);

INVxp33_ASAP7_75t_L g331 ( 
.A(n_163),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_193),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_196),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_161),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_196),
.Y(n_335)
);

INVx3_ASAP7_75t_L g336 ( 
.A(n_175),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_162),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_232),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_159),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_159),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_208),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_183),
.Y(n_342)
);

BUFx2_ASAP7_75t_L g343 ( 
.A(n_172),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_208),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_189),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_269),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_190),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_269),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_232),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_272),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_291),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_253),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_272),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_178),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_181),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_253),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_184),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_291),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_185),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_186),
.Y(n_360)
);

INVx1_ASAP7_75t_SL g361 ( 
.A(n_215),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_192),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_201),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_194),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_195),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_226),
.Y(n_366)
);

HB1xp67_ASAP7_75t_L g367 ( 
.A(n_172),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_228),
.Y(n_368)
);

BUFx2_ASAP7_75t_L g369 ( 
.A(n_290),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_242),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_197),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_243),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_248),
.Y(n_373)
);

BUFx3_ASAP7_75t_L g374 ( 
.A(n_222),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_251),
.Y(n_375)
);

CKINVDCx16_ASAP7_75t_R g376 ( 
.A(n_244),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_254),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_206),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_261),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_267),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_207),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_271),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_276),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_321),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_309),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_376),
.B(n_165),
.Y(n_386)
);

INVx3_ASAP7_75t_L g387 ( 
.A(n_342),
.Y(n_387)
);

CKINVDCx6p67_ASAP7_75t_R g388 ( 
.A(n_361),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_L g389 ( 
.A1(n_308),
.A2(n_169),
.B1(n_304),
.B2(n_270),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_310),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_367),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_342),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_310),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_342),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_342),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_351),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_311),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_311),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_315),
.Y(n_399)
);

BUFx3_ASAP7_75t_L g400 ( 
.A(n_327),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_333),
.B(n_222),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_351),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_315),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_317),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_317),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_358),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_318),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_318),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_336),
.B(n_156),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_322),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_322),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_358),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_323),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_323),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_324),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_336),
.B(n_156),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_324),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_336),
.B(n_164),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_334),
.Y(n_419)
);

HB1xp67_ASAP7_75t_L g420 ( 
.A(n_314),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_325),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_328),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_312),
.Y(n_423)
);

OAI21x1_ASAP7_75t_L g424 ( 
.A1(n_312),
.A2(n_209),
.B(n_170),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_329),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_325),
.Y(n_426)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_314),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_332),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_337),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_330),
.B(n_164),
.Y(n_430)
);

INVx3_ASAP7_75t_L g431 ( 
.A(n_330),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_354),
.Y(n_432)
);

HB1xp67_ASAP7_75t_L g433 ( 
.A(n_326),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g434 ( 
.A(n_333),
.B(n_170),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_335),
.B(n_166),
.Y(n_435)
);

HB1xp67_ASAP7_75t_L g436 ( 
.A(n_326),
.Y(n_436)
);

BUFx3_ASAP7_75t_L g437 ( 
.A(n_335),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_339),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_354),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_355),
.Y(n_440)
);

AND2x4_ASAP7_75t_L g441 ( 
.A(n_327),
.B(n_209),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_339),
.Y(n_442)
);

INVx3_ASAP7_75t_L g443 ( 
.A(n_340),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_355),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_357),
.Y(n_445)
);

INVx6_ASAP7_75t_L g446 ( 
.A(n_374),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_345),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_338),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_357),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_359),
.Y(n_450)
);

INVx3_ASAP7_75t_L g451 ( 
.A(n_340),
.Y(n_451)
);

OA21x2_ASAP7_75t_L g452 ( 
.A1(n_341),
.A2(n_288),
.B(n_278),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_374),
.B(n_236),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_384),
.B(n_347),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_437),
.Y(n_455)
);

AOI21x1_ASAP7_75t_L g456 ( 
.A1(n_424),
.A2(n_265),
.B(n_236),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_397),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_446),
.B(n_362),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_437),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_446),
.B(n_364),
.Y(n_460)
);

BUFx3_ASAP7_75t_L g461 ( 
.A(n_446),
.Y(n_461)
);

AND3x1_ASAP7_75t_L g462 ( 
.A(n_420),
.B(n_297),
.C(n_360),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_397),
.Y(n_463)
);

BUFx6f_ASAP7_75t_SL g464 ( 
.A(n_400),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_400),
.B(n_365),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_400),
.B(n_371),
.Y(n_466)
);

INVx8_ASAP7_75t_L g467 ( 
.A(n_419),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_453),
.B(n_313),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_429),
.B(n_378),
.Y(n_469)
);

INVx2_ASAP7_75t_SL g470 ( 
.A(n_446),
.Y(n_470)
);

INVx1_ASAP7_75t_SL g471 ( 
.A(n_388),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_446),
.B(n_381),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_447),
.B(n_316),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_446),
.B(n_319),
.Y(n_474)
);

INVx4_ASAP7_75t_L g475 ( 
.A(n_396),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_437),
.Y(n_476)
);

BUFx2_ASAP7_75t_L g477 ( 
.A(n_388),
.Y(n_477)
);

INVx2_ASAP7_75t_SL g478 ( 
.A(n_409),
.Y(n_478)
);

INVx3_ASAP7_75t_L g479 ( 
.A(n_394),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_390),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_388),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_453),
.B(n_341),
.Y(n_482)
);

INVx3_ASAP7_75t_L g483 ( 
.A(n_394),
.Y(n_483)
);

AND2x4_ASAP7_75t_L g484 ( 
.A(n_441),
.B(n_265),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_394),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_390),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_393),
.Y(n_487)
);

BUFx10_ASAP7_75t_L g488 ( 
.A(n_420),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_391),
.B(n_320),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_453),
.B(n_344),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_393),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_394),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_397),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_385),
.Y(n_494)
);

INVx2_ASAP7_75t_SL g495 ( 
.A(n_409),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_398),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_416),
.B(n_187),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_398),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_389),
.A2(n_169),
.B1(n_304),
.B2(n_295),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_391),
.B(n_343),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_394),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_399),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_416),
.B(n_343),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_407),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_399),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_403),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_403),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_427),
.B(n_369),
.Y(n_508)
);

OAI22xp33_ASAP7_75t_SL g509 ( 
.A1(n_435),
.A2(n_266),
.B1(n_289),
.B2(n_369),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_418),
.B(n_165),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_404),
.Y(n_511)
);

INVx3_ASAP7_75t_L g512 ( 
.A(n_394),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_418),
.B(n_386),
.Y(n_513)
);

INVx1_ASAP7_75t_SL g514 ( 
.A(n_385),
.Y(n_514)
);

INVxp33_ASAP7_75t_L g515 ( 
.A(n_433),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_407),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_404),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_405),
.Y(n_518)
);

OAI22xp33_ASAP7_75t_L g519 ( 
.A1(n_427),
.A2(n_252),
.B1(n_234),
.B2(n_233),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_408),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_408),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_394),
.Y(n_522)
);

INVxp33_ASAP7_75t_L g523 ( 
.A(n_433),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_422),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_408),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_386),
.B(n_331),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_411),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_405),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_411),
.Y(n_529)
);

INVx2_ASAP7_75t_SL g530 ( 
.A(n_436),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_410),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_410),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_411),
.Y(n_533)
);

CKINVDCx6p67_ASAP7_75t_R g534 ( 
.A(n_422),
.Y(n_534)
);

AOI22xp33_ASAP7_75t_L g535 ( 
.A1(n_452),
.A2(n_289),
.B1(n_266),
.B2(n_363),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_413),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_421),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_413),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_421),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_421),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_414),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_414),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_430),
.B(n_210),
.Y(n_543)
);

BUFx3_ASAP7_75t_L g544 ( 
.A(n_452),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_415),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_435),
.B(n_165),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_415),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_417),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_417),
.Y(n_549)
);

INVx3_ASAP7_75t_L g550 ( 
.A(n_394),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_441),
.B(n_168),
.Y(n_551)
);

AOI22xp5_ASAP7_75t_L g552 ( 
.A1(n_389),
.A2(n_290),
.B1(n_295),
.B2(n_300),
.Y(n_552)
);

NAND2xp33_ASAP7_75t_R g553 ( 
.A(n_452),
.B(n_441),
.Y(n_553)
);

BUFx6f_ASAP7_75t_L g554 ( 
.A(n_395),
.Y(n_554)
);

INVx4_ASAP7_75t_L g555 ( 
.A(n_396),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_426),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_441),
.B(n_168),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_426),
.Y(n_558)
);

BUFx3_ASAP7_75t_L g559 ( 
.A(n_452),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_430),
.B(n_231),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_425),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_441),
.B(n_168),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_452),
.Y(n_563)
);

AND2x4_ASAP7_75t_L g564 ( 
.A(n_434),
.B(n_155),
.Y(n_564)
);

BUFx3_ASAP7_75t_L g565 ( 
.A(n_401),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_424),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_424),
.Y(n_567)
);

BUFx3_ASAP7_75t_L g568 ( 
.A(n_401),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_431),
.Y(n_569)
);

NAND3xp33_ASAP7_75t_L g570 ( 
.A(n_434),
.B(n_284),
.C(n_359),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_431),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_431),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_436),
.B(n_221),
.Y(n_573)
);

NAND2xp33_ASAP7_75t_L g574 ( 
.A(n_401),
.B(n_183),
.Y(n_574)
);

NOR2x1p5_ASAP7_75t_L g575 ( 
.A(n_432),
.B(n_300),
.Y(n_575)
);

AO21x2_ASAP7_75t_L g576 ( 
.A1(n_434),
.A2(n_171),
.B(n_160),
.Y(n_576)
);

INVx2_ASAP7_75t_SL g577 ( 
.A(n_432),
.Y(n_577)
);

INVx1_ASAP7_75t_SL g578 ( 
.A(n_425),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_431),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_431),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_439),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_443),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_443),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_439),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_440),
.B(n_221),
.Y(n_585)
);

INVx3_ASAP7_75t_L g586 ( 
.A(n_395),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_443),
.Y(n_587)
);

AND2x6_ASAP7_75t_L g588 ( 
.A(n_396),
.B(n_183),
.Y(n_588)
);

BUFx3_ASAP7_75t_L g589 ( 
.A(n_387),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_443),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_444),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_444),
.Y(n_592)
);

INVx3_ASAP7_75t_L g593 ( 
.A(n_395),
.Y(n_593)
);

NAND2xp33_ASAP7_75t_R g594 ( 
.A(n_445),
.B(n_166),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_445),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_449),
.B(n_349),
.Y(n_596)
);

INVx2_ASAP7_75t_SL g597 ( 
.A(n_449),
.Y(n_597)
);

OAI22xp33_ASAP7_75t_L g598 ( 
.A1(n_450),
.A2(n_204),
.B1(n_203),
.B2(n_200),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_443),
.Y(n_599)
);

AND2x4_ASAP7_75t_L g600 ( 
.A(n_565),
.B(n_450),
.Y(n_600)
);

BUFx6f_ASAP7_75t_L g601 ( 
.A(n_461),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_581),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_478),
.B(n_183),
.Y(n_603)
);

AOI22x1_ASAP7_75t_L g604 ( 
.A1(n_563),
.A2(n_205),
.B1(n_255),
.B2(n_250),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_457),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_581),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_584),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_584),
.Y(n_608)
);

AOI22xp5_ASAP7_75t_L g609 ( 
.A1(n_478),
.A2(n_352),
.B1(n_356),
.B2(n_256),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_495),
.B(n_396),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_495),
.B(n_396),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_526),
.B(n_167),
.Y(n_612)
);

NOR2xp67_ASAP7_75t_L g613 ( 
.A(n_469),
.B(n_451),
.Y(n_613)
);

INVx2_ASAP7_75t_SL g614 ( 
.A(n_488),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_544),
.B(n_183),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_SL g616 ( 
.A(n_471),
.B(n_428),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_497),
.B(n_167),
.Y(n_617)
);

O2A1O1Ixp33_ASAP7_75t_L g618 ( 
.A1(n_509),
.A2(n_366),
.B(n_383),
.C(n_382),
.Y(n_618)
);

OR2x2_ASAP7_75t_L g619 ( 
.A(n_530),
.B(n_366),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_577),
.B(n_396),
.Y(n_620)
);

CKINVDCx11_ASAP7_75t_R g621 ( 
.A(n_524),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_457),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_544),
.B(n_241),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_577),
.B(n_396),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_503),
.B(n_174),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_597),
.B(n_396),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_559),
.B(n_509),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_513),
.B(n_174),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_597),
.B(n_402),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_559),
.B(n_241),
.Y(n_630)
);

OAI21xp33_ASAP7_75t_L g631 ( 
.A1(n_468),
.A2(n_370),
.B(n_368),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_565),
.B(n_402),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_463),
.Y(n_633)
);

INVxp67_ASAP7_75t_SL g634 ( 
.A(n_563),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_568),
.B(n_176),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_591),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_467),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_568),
.B(n_176),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_468),
.B(n_215),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_543),
.B(n_402),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_560),
.B(n_402),
.Y(n_641)
);

AOI21xp5_ASAP7_75t_L g642 ( 
.A1(n_474),
.A2(n_395),
.B(n_392),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_463),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_455),
.B(n_402),
.Y(n_644)
);

OR2x2_ASAP7_75t_L g645 ( 
.A(n_530),
.B(n_368),
.Y(n_645)
);

INVx2_ASAP7_75t_SL g646 ( 
.A(n_488),
.Y(n_646)
);

BUFx3_ASAP7_75t_L g647 ( 
.A(n_467),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_493),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_504),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_592),
.Y(n_650)
);

INVx2_ASAP7_75t_SL g651 ( 
.A(n_488),
.Y(n_651)
);

OAI22xp33_ASAP7_75t_L g652 ( 
.A1(n_499),
.A2(n_302),
.B1(n_230),
.B2(n_224),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_595),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_482),
.Y(n_654)
);

AO221x1_ASAP7_75t_L g655 ( 
.A1(n_519),
.A2(n_241),
.B1(n_294),
.B2(n_173),
.C(n_246),
.Y(n_655)
);

INVx3_ASAP7_75t_L g656 ( 
.A(n_589),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_459),
.B(n_241),
.Y(n_657)
);

NAND3xp33_ASAP7_75t_SL g658 ( 
.A(n_499),
.B(n_448),
.C(n_428),
.Y(n_658)
);

AOI22xp5_ASAP7_75t_L g659 ( 
.A1(n_575),
.A2(n_259),
.B1(n_307),
.B2(n_275),
.Y(n_659)
);

O2A1O1Ixp33_ASAP7_75t_L g660 ( 
.A1(n_510),
.A2(n_370),
.B(n_383),
.C(n_382),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_500),
.B(n_177),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_L g662 ( 
.A(n_508),
.B(n_177),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_476),
.B(n_564),
.Y(n_663)
);

INVx4_ASAP7_75t_L g664 ( 
.A(n_461),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_489),
.B(n_180),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_573),
.B(n_180),
.Y(n_666)
);

INVx4_ASAP7_75t_L g667 ( 
.A(n_589),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_476),
.B(n_564),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_546),
.B(n_239),
.Y(n_669)
);

AOI22xp5_ASAP7_75t_L g670 ( 
.A1(n_575),
.A2(n_260),
.B1(n_277),
.B2(n_263),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_465),
.B(n_239),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_516),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_466),
.B(n_240),
.Y(n_673)
);

BUFx3_ASAP7_75t_L g674 ( 
.A(n_467),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_454),
.B(n_240),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_490),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_490),
.Y(n_677)
);

NOR2xp67_ASAP7_75t_L g678 ( 
.A(n_481),
.B(n_451),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_564),
.B(n_406),
.Y(n_679)
);

AO22x2_ASAP7_75t_L g680 ( 
.A1(n_570),
.A2(n_218),
.B1(n_219),
.B2(n_225),
.Y(n_680)
);

OR2x6_ASAP7_75t_L g681 ( 
.A(n_467),
.B(n_372),
.Y(n_681)
);

INVx1_ASAP7_75t_SL g682 ( 
.A(n_514),
.Y(n_682)
);

OAI22xp5_ASAP7_75t_L g683 ( 
.A1(n_535),
.A2(n_282),
.B1(n_306),
.B2(n_179),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_484),
.B(n_241),
.Y(n_684)
);

INVx2_ASAP7_75t_SL g685 ( 
.A(n_488),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_598),
.B(n_293),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_564),
.B(n_406),
.Y(n_687)
);

NAND2xp33_ASAP7_75t_L g688 ( 
.A(n_458),
.B(n_291),
.Y(n_688)
);

AND2x6_ASAP7_75t_L g689 ( 
.A(n_566),
.B(n_294),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_480),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_520),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_596),
.B(n_293),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_486),
.B(n_406),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_487),
.B(n_406),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_487),
.B(n_491),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_491),
.B(n_406),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_496),
.B(n_406),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_462),
.B(n_298),
.Y(n_698)
);

INVx2_ASAP7_75t_SL g699 ( 
.A(n_585),
.Y(n_699)
);

INVx8_ASAP7_75t_L g700 ( 
.A(n_467),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_498),
.B(n_502),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_551),
.B(n_298),
.Y(n_702)
);

AOI22xp5_ASAP7_75t_L g703 ( 
.A1(n_553),
.A2(n_484),
.B1(n_464),
.B2(n_557),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_505),
.B(n_412),
.Y(n_704)
);

BUFx3_ASAP7_75t_L g705 ( 
.A(n_534),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_562),
.B(n_301),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_506),
.B(n_412),
.Y(n_707)
);

AOI221xp5_ASAP7_75t_L g708 ( 
.A1(n_552),
.A2(n_302),
.B1(n_279),
.B2(n_274),
.C(n_213),
.Y(n_708)
);

BUFx6f_ASAP7_75t_SL g709 ( 
.A(n_484),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_506),
.B(n_507),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_507),
.B(n_301),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_511),
.B(n_412),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_517),
.B(n_412),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_521),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_517),
.B(n_303),
.Y(n_715)
);

AND2x2_ASAP7_75t_L g716 ( 
.A(n_515),
.B(n_273),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_518),
.B(n_303),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_518),
.B(n_305),
.Y(n_718)
);

BUFx2_ASAP7_75t_L g719 ( 
.A(n_494),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_528),
.B(n_412),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_528),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_531),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_531),
.B(n_305),
.Y(n_723)
);

NAND2xp33_ASAP7_75t_L g724 ( 
.A(n_460),
.B(n_472),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_484),
.B(n_294),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_582),
.B(n_294),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_SL g727 ( 
.A(n_481),
.B(n_448),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_532),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_525),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_532),
.B(n_198),
.Y(n_730)
);

OR2x2_ASAP7_75t_L g731 ( 
.A(n_523),
.B(n_372),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_462),
.B(n_221),
.Y(n_732)
);

BUFx3_ASAP7_75t_L g733 ( 
.A(n_534),
.Y(n_733)
);

AOI22xp5_ASAP7_75t_L g734 ( 
.A1(n_464),
.A2(n_199),
.B1(n_299),
.B2(n_296),
.Y(n_734)
);

INVx3_ASAP7_75t_L g735 ( 
.A(n_582),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_536),
.B(n_412),
.Y(n_736)
);

BUFx6f_ASAP7_75t_L g737 ( 
.A(n_492),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_538),
.B(n_451),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_538),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_542),
.B(n_214),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_542),
.Y(n_741)
);

AND2x6_ASAP7_75t_L g742 ( 
.A(n_566),
.B(n_294),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_547),
.B(n_451),
.Y(n_743)
);

HB1xp67_ASAP7_75t_L g744 ( 
.A(n_594),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_525),
.Y(n_745)
);

BUFx6f_ASAP7_75t_L g746 ( 
.A(n_737),
.Y(n_746)
);

INVxp67_ASAP7_75t_L g747 ( 
.A(n_731),
.Y(n_747)
);

NOR2x1p5_ASAP7_75t_L g748 ( 
.A(n_658),
.B(n_494),
.Y(n_748)
);

AOI22xp5_ASAP7_75t_L g749 ( 
.A1(n_617),
.A2(n_576),
.B1(n_464),
.B2(n_547),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_735),
.Y(n_750)
);

INVx2_ASAP7_75t_SL g751 ( 
.A(n_619),
.Y(n_751)
);

NOR3xp33_ASAP7_75t_SL g752 ( 
.A(n_652),
.B(n_561),
.C(n_217),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_735),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_617),
.B(n_671),
.Y(n_754)
);

AOI22xp5_ASAP7_75t_L g755 ( 
.A1(n_671),
.A2(n_576),
.B1(n_556),
.B2(n_477),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_600),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_710),
.B(n_556),
.Y(n_757)
);

INVx1_ASAP7_75t_SL g758 ( 
.A(n_682),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_600),
.Y(n_759)
);

BUFx12f_ASAP7_75t_L g760 ( 
.A(n_621),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_602),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_605),
.Y(n_762)
);

AND2x4_ASAP7_75t_L g763 ( 
.A(n_654),
.B(n_477),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_606),
.Y(n_764)
);

INVx2_ASAP7_75t_SL g765 ( 
.A(n_645),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_607),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_710),
.B(n_576),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_703),
.B(n_583),
.Y(n_768)
);

INVx3_ASAP7_75t_L g769 ( 
.A(n_667),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_744),
.B(n_473),
.Y(n_770)
);

NOR3xp33_ASAP7_75t_SL g771 ( 
.A(n_652),
.B(n_561),
.C(n_220),
.Y(n_771)
);

BUFx6f_ASAP7_75t_L g772 ( 
.A(n_737),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_634),
.B(n_541),
.Y(n_773)
);

BUFx3_ASAP7_75t_L g774 ( 
.A(n_647),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_608),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_744),
.B(n_552),
.Y(n_776)
);

INVx3_ASAP7_75t_L g777 ( 
.A(n_667),
.Y(n_777)
);

NOR2x1p5_ASAP7_75t_L g778 ( 
.A(n_637),
.B(n_674),
.Y(n_778)
);

BUFx3_ASAP7_75t_L g779 ( 
.A(n_700),
.Y(n_779)
);

AND2x4_ASAP7_75t_L g780 ( 
.A(n_676),
.B(n_470),
.Y(n_780)
);

BUFx3_ASAP7_75t_L g781 ( 
.A(n_700),
.Y(n_781)
);

AOI22xp33_ASAP7_75t_L g782 ( 
.A1(n_627),
.A2(n_567),
.B1(n_541),
.B2(n_548),
.Y(n_782)
);

AOI22xp5_ASAP7_75t_L g783 ( 
.A1(n_661),
.A2(n_470),
.B1(n_549),
.B2(n_548),
.Y(n_783)
);

AO22x1_ASAP7_75t_L g784 ( 
.A1(n_686),
.A2(n_578),
.B1(n_216),
.B2(n_268),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_634),
.B(n_545),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_636),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_661),
.B(n_545),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_613),
.B(n_587),
.Y(n_788)
);

AOI22xp33_ASAP7_75t_L g789 ( 
.A1(n_627),
.A2(n_567),
.B1(n_549),
.B2(n_558),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_622),
.Y(n_790)
);

INVx2_ASAP7_75t_SL g791 ( 
.A(n_716),
.Y(n_791)
);

NOR2xp67_ASAP7_75t_L g792 ( 
.A(n_614),
.B(n_646),
.Y(n_792)
);

OAI22xp33_ASAP7_75t_L g793 ( 
.A1(n_677),
.A2(n_558),
.B1(n_262),
.B2(n_287),
.Y(n_793)
);

BUFx2_ASAP7_75t_L g794 ( 
.A(n_719),
.Y(n_794)
);

BUFx3_ASAP7_75t_L g795 ( 
.A(n_700),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_705),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_663),
.B(n_587),
.Y(n_797)
);

AOI21xp5_ASAP7_75t_L g798 ( 
.A1(n_640),
.A2(n_475),
.B(n_555),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_662),
.B(n_569),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_650),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_733),
.Y(n_801)
);

NAND2x1p5_ASAP7_75t_L g802 ( 
.A(n_656),
.B(n_590),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_653),
.B(n_569),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_612),
.B(n_590),
.Y(n_804)
);

AOI22xp5_ASAP7_75t_L g805 ( 
.A1(n_628),
.A2(n_574),
.B1(n_599),
.B2(n_475),
.Y(n_805)
);

OR2x2_ASAP7_75t_L g806 ( 
.A(n_609),
.B(n_373),
.Y(n_806)
);

OAI22xp5_ASAP7_75t_SL g807 ( 
.A1(n_686),
.A2(n_249),
.B1(n_245),
.B2(n_247),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_668),
.B(n_599),
.Y(n_808)
);

HB1xp67_ASAP7_75t_L g809 ( 
.A(n_639),
.Y(n_809)
);

INVx4_ASAP7_75t_L g810 ( 
.A(n_709),
.Y(n_810)
);

INVx3_ASAP7_75t_L g811 ( 
.A(n_656),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_690),
.B(n_479),
.Y(n_812)
);

CKINVDCx20_ASAP7_75t_R g813 ( 
.A(n_651),
.Y(n_813)
);

NOR3xp33_ASAP7_75t_SL g814 ( 
.A(n_698),
.B(n_257),
.C(n_281),
.Y(n_814)
);

AND2x6_ASAP7_75t_L g815 ( 
.A(n_721),
.B(n_571),
.Y(n_815)
);

AOI22xp33_ASAP7_75t_L g816 ( 
.A1(n_680),
.A2(n_291),
.B1(n_182),
.B2(n_191),
.Y(n_816)
);

CKINVDCx20_ASAP7_75t_R g817 ( 
.A(n_685),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_633),
.Y(n_818)
);

AOI22xp33_ASAP7_75t_L g819 ( 
.A1(n_680),
.A2(n_291),
.B1(n_202),
.B2(n_285),
.Y(n_819)
);

OAI22xp5_ASAP7_75t_SL g820 ( 
.A1(n_665),
.A2(n_258),
.B1(n_264),
.B2(n_280),
.Y(n_820)
);

OR2x6_ASAP7_75t_L g821 ( 
.A(n_681),
.B(n_373),
.Y(n_821)
);

OR2x2_ASAP7_75t_SL g822 ( 
.A(n_727),
.B(n_212),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_643),
.Y(n_823)
);

INVx2_ASAP7_75t_SL g824 ( 
.A(n_699),
.Y(n_824)
);

BUFx2_ASAP7_75t_L g825 ( 
.A(n_681),
.Y(n_825)
);

OAI22xp5_ASAP7_75t_SL g826 ( 
.A1(n_665),
.A2(n_286),
.B1(n_375),
.B2(n_377),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_722),
.B(n_479),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_728),
.B(n_479),
.Y(n_828)
);

AOI22xp33_ASAP7_75t_L g829 ( 
.A1(n_680),
.A2(n_604),
.B1(n_655),
.B2(n_615),
.Y(n_829)
);

BUFx3_ASAP7_75t_L g830 ( 
.A(n_681),
.Y(n_830)
);

BUFx2_ASAP7_75t_L g831 ( 
.A(n_739),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_741),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_695),
.B(n_483),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_628),
.B(n_571),
.Y(n_834)
);

AND2x4_ASAP7_75t_L g835 ( 
.A(n_678),
.B(n_375),
.Y(n_835)
);

INVx3_ASAP7_75t_SL g836 ( 
.A(n_732),
.Y(n_836)
);

BUFx12f_ASAP7_75t_L g837 ( 
.A(n_601),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_701),
.B(n_483),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_737),
.B(n_572),
.Y(n_839)
);

INVx5_ASAP7_75t_L g840 ( 
.A(n_737),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_648),
.Y(n_841)
);

OR2x2_ASAP7_75t_L g842 ( 
.A(n_692),
.B(n_377),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_SL g843 ( 
.A(n_679),
.B(n_572),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_711),
.B(n_485),
.Y(n_844)
);

OAI22xp5_ASAP7_75t_L g845 ( 
.A1(n_615),
.A2(n_623),
.B1(n_630),
.B2(n_611),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_687),
.B(n_579),
.Y(n_846)
);

BUFx6f_ASAP7_75t_L g847 ( 
.A(n_601),
.Y(n_847)
);

NOR2x2_ASAP7_75t_L g848 ( 
.A(n_708),
.B(n_579),
.Y(n_848)
);

INVx3_ASAP7_75t_L g849 ( 
.A(n_601),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_649),
.Y(n_850)
);

NOR3xp33_ASAP7_75t_L g851 ( 
.A(n_666),
.B(n_229),
.C(n_235),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_715),
.B(n_717),
.Y(n_852)
);

AND2x4_ASAP7_75t_L g853 ( 
.A(n_734),
.B(n_379),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_715),
.B(n_485),
.Y(n_854)
);

INVx2_ASAP7_75t_SL g855 ( 
.A(n_638),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_632),
.B(n_580),
.Y(n_856)
);

INVxp67_ASAP7_75t_L g857 ( 
.A(n_635),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_SL g858 ( 
.A(n_610),
.B(n_580),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_717),
.B(n_512),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_738),
.Y(n_860)
);

BUFx3_ASAP7_75t_L g861 ( 
.A(n_743),
.Y(n_861)
);

OR2x6_ASAP7_75t_L g862 ( 
.A(n_618),
.B(n_379),
.Y(n_862)
);

INVx2_ASAP7_75t_SL g863 ( 
.A(n_673),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_718),
.B(n_512),
.Y(n_864)
);

AND2x6_ASAP7_75t_SL g865 ( 
.A(n_675),
.B(n_380),
.Y(n_865)
);

BUFx5_ASAP7_75t_L g866 ( 
.A(n_689),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_675),
.Y(n_867)
);

AND2x2_ASAP7_75t_L g868 ( 
.A(n_625),
.B(n_273),
.Y(n_868)
);

OR2x2_ASAP7_75t_L g869 ( 
.A(n_625),
.B(n_380),
.Y(n_869)
);

INVx2_ASAP7_75t_SL g870 ( 
.A(n_666),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_718),
.B(n_512),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_693),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_672),
.Y(n_873)
);

HB1xp67_ASAP7_75t_L g874 ( 
.A(n_709),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_723),
.B(n_550),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_730),
.B(n_550),
.Y(n_876)
);

AOI22xp33_ASAP7_75t_L g877 ( 
.A1(n_623),
.A2(n_291),
.B1(n_273),
.B2(n_529),
.Y(n_877)
);

AND2x6_ASAP7_75t_L g878 ( 
.A(n_641),
.B(n_586),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_691),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_694),
.B(n_555),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_740),
.B(n_586),
.Y(n_881)
);

BUFx3_ASAP7_75t_L g882 ( 
.A(n_620),
.Y(n_882)
);

AND2x4_ASAP7_75t_L g883 ( 
.A(n_664),
.B(n_346),
.Y(n_883)
);

NAND3xp33_ASAP7_75t_SL g884 ( 
.A(n_669),
.B(n_346),
.C(n_348),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_696),
.Y(n_885)
);

AOI22xp5_ASAP7_75t_L g886 ( 
.A1(n_702),
.A2(n_475),
.B1(n_555),
.B2(n_586),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_697),
.Y(n_887)
);

INVx3_ASAP7_75t_L g888 ( 
.A(n_664),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_635),
.B(n_669),
.Y(n_889)
);

A2O1A1Ixp33_ASAP7_75t_L g890 ( 
.A1(n_631),
.A2(n_451),
.B(n_353),
.C(n_350),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_630),
.B(n_593),
.Y(n_891)
);

AOI22xp33_ASAP7_75t_L g892 ( 
.A1(n_683),
.A2(n_291),
.B1(n_540),
.B2(n_533),
.Y(n_892)
);

AND2x4_ASAP7_75t_L g893 ( 
.A(n_659),
.B(n_348),
.Y(n_893)
);

INVx2_ASAP7_75t_SL g894 ( 
.A(n_702),
.Y(n_894)
);

INVx2_ASAP7_75t_SL g895 ( 
.A(n_706),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_616),
.B(n_350),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_714),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_603),
.B(n_593),
.Y(n_898)
);

OR2x6_ASAP7_75t_L g899 ( 
.A(n_660),
.B(n_353),
.Y(n_899)
);

INVxp67_ASAP7_75t_L g900 ( 
.A(n_706),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_603),
.B(n_527),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_670),
.B(n_237),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_R g903 ( 
.A(n_724),
.B(n_456),
.Y(n_903)
);

INVx3_ASAP7_75t_L g904 ( 
.A(n_729),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_745),
.B(n_527),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_624),
.B(n_529),
.Y(n_906)
);

AOI22xp33_ASAP7_75t_L g907 ( 
.A1(n_742),
.A2(n_533),
.B1(n_540),
.B2(n_539),
.Y(n_907)
);

BUFx6f_ASAP7_75t_L g908 ( 
.A(n_626),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_644),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_629),
.A2(n_492),
.B(n_554),
.Y(n_910)
);

AOI22xp33_ASAP7_75t_L g911 ( 
.A1(n_689),
.A2(n_537),
.B1(n_539),
.B2(n_588),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_684),
.Y(n_912)
);

BUFx12f_ASAP7_75t_SL g913 ( 
.A(n_688),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_840),
.A2(n_845),
.B(n_798),
.Y(n_914)
);

O2A1O1Ixp33_ASAP7_75t_L g915 ( 
.A1(n_754),
.A2(n_657),
.B(n_684),
.C(n_725),
.Y(n_915)
);

A2O1A1Ixp33_ASAP7_75t_L g916 ( 
.A1(n_889),
.A2(n_725),
.B(n_642),
.C(n_736),
.Y(n_916)
);

INVx4_ASAP7_75t_L g917 ( 
.A(n_837),
.Y(n_917)
);

AND2x4_ASAP7_75t_L g918 ( 
.A(n_774),
.B(n_704),
.Y(n_918)
);

NAND2xp33_ASAP7_75t_L g919 ( 
.A(n_867),
.B(n_689),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_790),
.Y(n_920)
);

BUFx8_ASAP7_75t_SL g921 ( 
.A(n_760),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_796),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_L g923 ( 
.A(n_889),
.B(n_707),
.Y(n_923)
);

OAI22xp5_ASAP7_75t_L g924 ( 
.A1(n_852),
.A2(n_712),
.B1(n_713),
.B2(n_720),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_747),
.B(n_237),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_L g926 ( 
.A(n_857),
.B(n_657),
.Y(n_926)
);

OAI22xp5_ASAP7_75t_L g927 ( 
.A1(n_757),
.A2(n_726),
.B1(n_456),
.B2(n_537),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_747),
.B(n_237),
.Y(n_928)
);

NOR2xp33_ASAP7_75t_L g929 ( 
.A(n_857),
.B(n_554),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_900),
.B(n_742),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_761),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_R g932 ( 
.A(n_801),
.B(n_742),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_900),
.B(n_554),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_764),
.Y(n_934)
);

NOR3xp33_ASAP7_75t_SL g935 ( 
.A(n_776),
.B(n_1),
.C(n_2),
.Y(n_935)
);

A2O1A1Ixp33_ASAP7_75t_L g936 ( 
.A1(n_851),
.A2(n_442),
.B(n_438),
.C(n_392),
.Y(n_936)
);

OAI21xp5_ASAP7_75t_L g937 ( 
.A1(n_767),
.A2(n_789),
.B(n_782),
.Y(n_937)
);

AND2x2_ASAP7_75t_L g938 ( 
.A(n_809),
.B(n_438),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_790),
.Y(n_939)
);

NOR2xp67_ASAP7_75t_SL g940 ( 
.A(n_779),
.B(n_522),
.Y(n_940)
);

OAI22xp5_ASAP7_75t_L g941 ( 
.A1(n_816),
.A2(n_442),
.B1(n_438),
.B2(n_554),
.Y(n_941)
);

NAND2xp33_ASAP7_75t_R g942 ( 
.A(n_814),
.B(n_69),
.Y(n_942)
);

INVx5_ASAP7_75t_L g943 ( 
.A(n_746),
.Y(n_943)
);

INVx3_ASAP7_75t_L g944 ( 
.A(n_847),
.Y(n_944)
);

AOI22xp5_ASAP7_75t_L g945 ( 
.A1(n_870),
.A2(n_742),
.B1(n_689),
.B2(n_588),
.Y(n_945)
);

INVxp67_ASAP7_75t_L g946 ( 
.A(n_758),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_766),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_850),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_788),
.A2(n_881),
.B(n_876),
.Y(n_949)
);

AO32x2_ASAP7_75t_L g950 ( 
.A1(n_894),
.A2(n_895),
.A3(n_826),
.B1(n_807),
.B2(n_863),
.Y(n_950)
);

BUFx8_ASAP7_75t_L g951 ( 
.A(n_794),
.Y(n_951)
);

OAI22xp5_ASAP7_75t_SL g952 ( 
.A1(n_776),
.A2(n_822),
.B1(n_813),
.B2(n_817),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_873),
.Y(n_953)
);

INVx3_ASAP7_75t_L g954 ( 
.A(n_847),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_787),
.B(n_554),
.Y(n_955)
);

AOI22xp5_ASAP7_75t_L g956 ( 
.A1(n_770),
.A2(n_588),
.B1(n_522),
.B2(n_501),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_809),
.B(n_896),
.Y(n_957)
);

INVxp67_ASAP7_75t_L g958 ( 
.A(n_751),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_775),
.Y(n_959)
);

HB1xp67_ASAP7_75t_L g960 ( 
.A(n_765),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_SL g961 ( 
.A(n_763),
.B(n_522),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_860),
.B(n_501),
.Y(n_962)
);

AO32x2_ASAP7_75t_L g963 ( 
.A1(n_855),
.A2(n_1),
.A3(n_2),
.B1(n_3),
.B2(n_7),
.Y(n_963)
);

NAND3xp33_ASAP7_75t_SL g964 ( 
.A(n_851),
.B(n_8),
.C(n_9),
.Y(n_964)
);

NOR2xp67_ASAP7_75t_L g965 ( 
.A(n_791),
.B(n_60),
.Y(n_965)
);

INVx1_ASAP7_75t_SL g966 ( 
.A(n_848),
.Y(n_966)
);

A2O1A1Ixp33_ASAP7_75t_L g967 ( 
.A1(n_755),
.A2(n_387),
.B(n_423),
.C(n_492),
.Y(n_967)
);

O2A1O1Ixp33_ASAP7_75t_L g968 ( 
.A1(n_868),
.A2(n_869),
.B(n_793),
.C(n_806),
.Y(n_968)
);

BUFx6f_ASAP7_75t_L g969 ( 
.A(n_746),
.Y(n_969)
);

O2A1O1Ixp5_ASAP7_75t_L g970 ( 
.A1(n_768),
.A2(n_834),
.B(n_799),
.C(n_875),
.Y(n_970)
);

INVx4_ASAP7_75t_L g971 ( 
.A(n_779),
.Y(n_971)
);

A2O1A1Ixp33_ASAP7_75t_L g972 ( 
.A1(n_749),
.A2(n_423),
.B(n_395),
.C(n_11),
.Y(n_972)
);

INVx4_ASAP7_75t_L g973 ( 
.A(n_781),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_880),
.A2(n_423),
.B(n_588),
.Y(n_974)
);

INVxp67_ASAP7_75t_L g975 ( 
.A(n_763),
.Y(n_975)
);

NOR2xp67_ASAP7_75t_L g976 ( 
.A(n_824),
.B(n_54),
.Y(n_976)
);

OAI21xp33_ASAP7_75t_L g977 ( 
.A1(n_902),
.A2(n_423),
.B(n_10),
.Y(n_977)
);

O2A1O1Ixp5_ASAP7_75t_L g978 ( 
.A1(n_834),
.A2(n_588),
.B(n_118),
.C(n_153),
.Y(n_978)
);

NAND3xp33_ASAP7_75t_SL g979 ( 
.A(n_752),
.B(n_9),
.C(n_10),
.Y(n_979)
);

A2O1A1Ixp33_ASAP7_75t_L g980 ( 
.A1(n_804),
.A2(n_423),
.B(n_13),
.C(n_16),
.Y(n_980)
);

O2A1O1Ixp5_ASAP7_75t_L g981 ( 
.A1(n_844),
.A2(n_588),
.B(n_115),
.C(n_150),
.Y(n_981)
);

OR2x2_ASAP7_75t_L g982 ( 
.A(n_842),
.B(n_423),
.Y(n_982)
);

NOR2xp33_ASAP7_75t_L g983 ( 
.A(n_831),
.B(n_12),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_L g984 ( 
.A(n_836),
.B(n_13),
.Y(n_984)
);

NOR2xp67_ASAP7_75t_L g985 ( 
.A(n_810),
.B(n_147),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_786),
.Y(n_986)
);

AOI22xp33_ASAP7_75t_L g987 ( 
.A1(n_893),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_987)
);

OA21x2_ASAP7_75t_L g988 ( 
.A1(n_782),
.A2(n_145),
.B(n_142),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_R g989 ( 
.A(n_913),
.B(n_141),
.Y(n_989)
);

O2A1O1Ixp33_ASAP7_75t_L g990 ( 
.A1(n_793),
.A2(n_18),
.B(n_19),
.C(n_24),
.Y(n_990)
);

OAI22x1_ASAP7_75t_L g991 ( 
.A1(n_748),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_991)
);

A2O1A1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_804),
.A2(n_32),
.B(n_36),
.C(n_37),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_800),
.B(n_32),
.Y(n_993)
);

BUFx12f_ASAP7_75t_L g994 ( 
.A(n_810),
.Y(n_994)
);

O2A1O1Ixp33_ASAP7_75t_L g995 ( 
.A1(n_836),
.A2(n_37),
.B(n_38),
.C(n_44),
.Y(n_995)
);

AND2x4_ASAP7_75t_L g996 ( 
.A(n_774),
.B(n_88),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_756),
.B(n_47),
.Y(n_997)
);

AOI22xp33_ASAP7_75t_L g998 ( 
.A1(n_893),
.A2(n_49),
.B1(n_68),
.B2(n_72),
.Y(n_998)
);

A2O1A1Ixp33_ASAP7_75t_L g999 ( 
.A1(n_832),
.A2(n_74),
.B(n_105),
.C(n_110),
.Y(n_999)
);

OAI22xp5_ASAP7_75t_L g1000 ( 
.A1(n_816),
.A2(n_114),
.B1(n_136),
.B2(n_819),
.Y(n_1000)
);

INVx4_ASAP7_75t_L g1001 ( 
.A(n_795),
.Y(n_1001)
);

OAI22xp5_ASAP7_75t_L g1002 ( 
.A1(n_819),
.A2(n_912),
.B1(n_789),
.B2(n_829),
.Y(n_1002)
);

OAI21xp33_ASAP7_75t_L g1003 ( 
.A1(n_752),
.A2(n_771),
.B(n_853),
.Y(n_1003)
);

OAI22xp5_ASAP7_75t_L g1004 ( 
.A1(n_829),
.A2(n_785),
.B1(n_773),
.B2(n_907),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_L g1005 ( 
.A(n_759),
.B(n_865),
.Y(n_1005)
);

AND2x2_ASAP7_75t_L g1006 ( 
.A(n_853),
.B(n_835),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_872),
.B(n_885),
.Y(n_1007)
);

INVx3_ASAP7_75t_SL g1008 ( 
.A(n_848),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_833),
.A2(n_838),
.B(n_888),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_887),
.B(n_835),
.Y(n_1010)
);

AND2x2_ASAP7_75t_SL g1011 ( 
.A(n_825),
.B(n_874),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_904),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_R g1013 ( 
.A(n_795),
.B(n_849),
.Y(n_1013)
);

OR2x2_ASAP7_75t_L g1014 ( 
.A(n_784),
.B(n_874),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_904),
.Y(n_1015)
);

OAI22xp5_ASAP7_75t_L g1016 ( 
.A1(n_907),
.A2(n_911),
.B1(n_771),
.B2(n_877),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_SL g1017 ( 
.A(n_814),
.B(n_769),
.Y(n_1017)
);

HB1xp67_ASAP7_75t_L g1018 ( 
.A(n_883),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_762),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_888),
.A2(n_854),
.B(n_871),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_818),
.Y(n_1021)
);

NOR2xp33_ASAP7_75t_L g1022 ( 
.A(n_820),
.B(n_830),
.Y(n_1022)
);

INVx1_ASAP7_75t_SL g1023 ( 
.A(n_883),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_909),
.B(n_861),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_780),
.B(n_882),
.Y(n_1025)
);

BUFx6f_ASAP7_75t_L g1026 ( 
.A(n_746),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_859),
.A2(n_864),
.B(n_891),
.Y(n_1027)
);

BUFx12f_ASAP7_75t_L g1028 ( 
.A(n_778),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_SL g1029 ( 
.A(n_777),
.B(n_780),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_823),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_910),
.A2(n_906),
.B(n_856),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_882),
.B(n_908),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_797),
.A2(n_808),
.B(n_846),
.Y(n_1033)
);

O2A1O1Ixp33_ASAP7_75t_L g1034 ( 
.A1(n_884),
.A2(n_862),
.B(n_890),
.C(n_803),
.Y(n_1034)
);

CKINVDCx8_ASAP7_75t_R g1035 ( 
.A(n_821),
.Y(n_1035)
);

BUFx6f_ASAP7_75t_L g1036 ( 
.A(n_746),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_L g1037 ( 
.A(n_821),
.B(n_908),
.Y(n_1037)
);

INVx3_ASAP7_75t_L g1038 ( 
.A(n_847),
.Y(n_1038)
);

BUFx6f_ASAP7_75t_L g1039 ( 
.A(n_772),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_923),
.B(n_957),
.Y(n_1040)
);

AND2x6_ASAP7_75t_L g1041 ( 
.A(n_996),
.B(n_908),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_1007),
.B(n_908),
.Y(n_1042)
);

OAI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_970),
.A2(n_783),
.B(n_877),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_968),
.B(n_1010),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_931),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_1006),
.B(n_811),
.Y(n_1046)
);

OAI21x1_ASAP7_75t_L g1047 ( 
.A1(n_1031),
.A2(n_858),
.B(n_843),
.Y(n_1047)
);

NAND3xp33_ASAP7_75t_SL g1048 ( 
.A(n_1003),
.B(n_805),
.C(n_890),
.Y(n_1048)
);

OR2x2_ASAP7_75t_L g1049 ( 
.A(n_966),
.B(n_821),
.Y(n_1049)
);

INVxp67_ASAP7_75t_L g1050 ( 
.A(n_960),
.Y(n_1050)
);

OA21x2_ASAP7_75t_L g1051 ( 
.A1(n_967),
.A2(n_858),
.B(n_901),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_1024),
.B(n_811),
.Y(n_1052)
);

NAND2xp33_ASAP7_75t_R g1053 ( 
.A(n_932),
.B(n_903),
.Y(n_1053)
);

AND2x6_ASAP7_75t_L g1054 ( 
.A(n_996),
.B(n_969),
.Y(n_1054)
);

AO22x2_ASAP7_75t_L g1055 ( 
.A1(n_1002),
.A2(n_808),
.B1(n_797),
.B2(n_846),
.Y(n_1055)
);

NAND2x1_ASAP7_75t_L g1056 ( 
.A(n_940),
.B(n_772),
.Y(n_1056)
);

NOR2xp33_ASAP7_75t_L g1057 ( 
.A(n_1008),
.B(n_792),
.Y(n_1057)
);

AOI22xp5_ASAP7_75t_L g1058 ( 
.A1(n_966),
.A2(n_862),
.B1(n_899),
.B2(n_897),
.Y(n_1058)
);

OAI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_916),
.A2(n_843),
.B(n_886),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_949),
.A2(n_772),
.B(n_911),
.Y(n_1060)
);

OAI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_915),
.A2(n_898),
.B(n_828),
.Y(n_1061)
);

OAI21x1_ASAP7_75t_L g1062 ( 
.A1(n_914),
.A2(n_839),
.B(n_827),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_1020),
.A2(n_812),
.B(n_905),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_1027),
.A2(n_839),
.B(n_847),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_1009),
.A2(n_802),
.B(n_753),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_L g1066 ( 
.A(n_946),
.B(n_750),
.Y(n_1066)
);

AND2x2_ASAP7_75t_L g1067 ( 
.A(n_938),
.B(n_862),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_934),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_SL g1069 ( 
.A(n_1023),
.B(n_879),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_1024),
.B(n_841),
.Y(n_1070)
);

BUFx6f_ASAP7_75t_L g1071 ( 
.A(n_969),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_1023),
.B(n_815),
.Y(n_1072)
);

OAI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_1034),
.A2(n_892),
.B(n_878),
.Y(n_1073)
);

BUFx6f_ASAP7_75t_L g1074 ( 
.A(n_969),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_937),
.A2(n_866),
.B(n_878),
.Y(n_1075)
);

OA21x2_ASAP7_75t_L g1076 ( 
.A1(n_937),
.A2(n_878),
.B(n_815),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_1025),
.B(n_815),
.Y(n_1077)
);

NAND3xp33_ASAP7_75t_L g1078 ( 
.A(n_935),
.B(n_899),
.C(n_815),
.Y(n_1078)
);

AO31x2_ASAP7_75t_L g1079 ( 
.A1(n_1004),
.A2(n_878),
.A3(n_815),
.B(n_866),
.Y(n_1079)
);

BUFx10_ASAP7_75t_L g1080 ( 
.A(n_922),
.Y(n_1080)
);

OAI22xp5_ASAP7_75t_L g1081 ( 
.A1(n_1002),
.A2(n_899),
.B1(n_878),
.B2(n_866),
.Y(n_1081)
);

INVx3_ASAP7_75t_L g1082 ( 
.A(n_943),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_921),
.Y(n_1083)
);

OAI21xp5_ASAP7_75t_SL g1084 ( 
.A1(n_987),
.A2(n_866),
.B(n_984),
.Y(n_1084)
);

INVxp67_ASAP7_75t_L g1085 ( 
.A(n_1005),
.Y(n_1085)
);

OAI21xp5_ASAP7_75t_SL g1086 ( 
.A1(n_1022),
.A2(n_866),
.B(n_998),
.Y(n_1086)
);

NOR2xp67_ASAP7_75t_SL g1087 ( 
.A(n_1035),
.B(n_994),
.Y(n_1087)
);

CKINVDCx20_ASAP7_75t_R g1088 ( 
.A(n_951),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_920),
.Y(n_1089)
);

INVxp67_ASAP7_75t_L g1090 ( 
.A(n_951),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_1032),
.B(n_1037),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_947),
.B(n_959),
.Y(n_1092)
);

OAI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_930),
.A2(n_1004),
.B(n_926),
.Y(n_1093)
);

AND2x2_ASAP7_75t_L g1094 ( 
.A(n_925),
.B(n_928),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_986),
.Y(n_1095)
);

OR2x2_ASAP7_75t_L g1096 ( 
.A(n_975),
.B(n_1018),
.Y(n_1096)
);

AOI22xp5_ASAP7_75t_L g1097 ( 
.A1(n_964),
.A2(n_977),
.B1(n_979),
.B2(n_1000),
.Y(n_1097)
);

NAND3xp33_ASAP7_75t_L g1098 ( 
.A(n_990),
.B(n_992),
.C(n_995),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_SL g1099 ( 
.A1(n_1000),
.A2(n_972),
.B(n_988),
.Y(n_1099)
);

A2O1A1Ixp33_ASAP7_75t_L g1100 ( 
.A1(n_997),
.A2(n_1016),
.B(n_980),
.C(n_993),
.Y(n_1100)
);

AOI22xp5_ASAP7_75t_L g1101 ( 
.A1(n_952),
.A2(n_983),
.B1(n_942),
.B2(n_991),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_939),
.Y(n_1102)
);

A2O1A1Ixp33_ASAP7_75t_L g1103 ( 
.A1(n_1017),
.A2(n_978),
.B(n_933),
.C(n_929),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_955),
.A2(n_919),
.B(n_924),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_948),
.Y(n_1105)
);

A2O1A1Ixp33_ASAP7_75t_L g1106 ( 
.A1(n_965),
.A2(n_999),
.B(n_981),
.C(n_1019),
.Y(n_1106)
);

BUFx2_ASAP7_75t_L g1107 ( 
.A(n_958),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_918),
.B(n_1021),
.Y(n_1108)
);

OR2x2_ASAP7_75t_L g1109 ( 
.A(n_1014),
.B(n_1030),
.Y(n_1109)
);

AND2x2_ASAP7_75t_L g1110 ( 
.A(n_1011),
.B(n_950),
.Y(n_1110)
);

INVx1_ASAP7_75t_SL g1111 ( 
.A(n_989),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_924),
.A2(n_927),
.B(n_962),
.Y(n_1112)
);

AND2x4_ASAP7_75t_L g1113 ( 
.A(n_971),
.B(n_1001),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_SL g1114 ( 
.A(n_917),
.B(n_1015),
.Y(n_1114)
);

AOI22xp5_ASAP7_75t_L g1115 ( 
.A1(n_1029),
.A2(n_976),
.B1(n_985),
.B2(n_961),
.Y(n_1115)
);

AO31x2_ASAP7_75t_L g1116 ( 
.A1(n_941),
.A2(n_936),
.A3(n_974),
.B(n_953),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_943),
.A2(n_982),
.B(n_988),
.Y(n_1117)
);

INVx5_ASAP7_75t_L g1118 ( 
.A(n_1026),
.Y(n_1118)
);

AND2x4_ASAP7_75t_L g1119 ( 
.A(n_971),
.B(n_1001),
.Y(n_1119)
);

OAI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_956),
.A2(n_945),
.B(n_941),
.Y(n_1120)
);

AO21x1_ASAP7_75t_L g1121 ( 
.A1(n_963),
.A2(n_950),
.B(n_1012),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_1028),
.Y(n_1122)
);

A2O1A1Ixp33_ASAP7_75t_L g1123 ( 
.A1(n_950),
.A2(n_944),
.B(n_954),
.C(n_1038),
.Y(n_1123)
);

OAI21xp33_ASAP7_75t_L g1124 ( 
.A1(n_1013),
.A2(n_944),
.B(n_954),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_1038),
.A2(n_1026),
.B(n_1036),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_1036),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1039),
.Y(n_1127)
);

NOR2xp33_ASAP7_75t_L g1128 ( 
.A(n_917),
.B(n_973),
.Y(n_1128)
);

OAI22xp5_ASAP7_75t_L g1129 ( 
.A1(n_973),
.A2(n_889),
.B1(n_754),
.B2(n_867),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_1039),
.A2(n_949),
.B(n_1020),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_1039),
.B(n_963),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_963),
.B(n_889),
.Y(n_1132)
);

OR2x2_ASAP7_75t_L g1133 ( 
.A(n_966),
.B(n_514),
.Y(n_1133)
);

OAI21x1_ASAP7_75t_L g1134 ( 
.A1(n_1031),
.A2(n_914),
.B(n_1033),
.Y(n_1134)
);

OAI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_970),
.A2(n_754),
.B(n_889),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_923),
.B(n_889),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_931),
.Y(n_1137)
);

OR2x2_ASAP7_75t_L g1138 ( 
.A(n_966),
.B(n_514),
.Y(n_1138)
);

AND2x2_ASAP7_75t_L g1139 ( 
.A(n_957),
.B(n_966),
.Y(n_1139)
);

AOI211x1_ASAP7_75t_L g1140 ( 
.A1(n_937),
.A2(n_652),
.B(n_1002),
.C(n_1007),
.Y(n_1140)
);

INVx4_ASAP7_75t_L g1141 ( 
.A(n_943),
.Y(n_1141)
);

NAND3xp33_ASAP7_75t_L g1142 ( 
.A(n_968),
.B(n_889),
.C(n_754),
.Y(n_1142)
);

A2O1A1Ixp33_ASAP7_75t_L g1143 ( 
.A1(n_968),
.A2(n_889),
.B(n_754),
.C(n_852),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_931),
.Y(n_1144)
);

HB1xp67_ASAP7_75t_L g1145 ( 
.A(n_946),
.Y(n_1145)
);

BUFx6f_ASAP7_75t_L g1146 ( 
.A(n_969),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_923),
.B(n_889),
.Y(n_1147)
);

AOI221xp5_ASAP7_75t_SL g1148 ( 
.A1(n_968),
.A2(n_652),
.B1(n_807),
.B2(n_820),
.C(n_889),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_923),
.B(n_889),
.Y(n_1149)
);

NAND2x1_ASAP7_75t_L g1150 ( 
.A(n_940),
.B(n_746),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_923),
.B(n_889),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_931),
.Y(n_1152)
);

OAI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_970),
.A2(n_754),
.B(n_889),
.Y(n_1153)
);

BUFx2_ASAP7_75t_L g1154 ( 
.A(n_946),
.Y(n_1154)
);

BUFx2_ASAP7_75t_L g1155 ( 
.A(n_946),
.Y(n_1155)
);

A2O1A1Ixp33_ASAP7_75t_L g1156 ( 
.A1(n_968),
.A2(n_889),
.B(n_754),
.C(n_852),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_949),
.A2(n_1020),
.B(n_1027),
.Y(n_1157)
);

INVx3_ASAP7_75t_SL g1158 ( 
.A(n_922),
.Y(n_1158)
);

OA21x2_ASAP7_75t_L g1159 ( 
.A1(n_967),
.A2(n_949),
.B(n_937),
.Y(n_1159)
);

AND2x2_ASAP7_75t_L g1160 ( 
.A(n_957),
.B(n_966),
.Y(n_1160)
);

AO21x1_ASAP7_75t_L g1161 ( 
.A1(n_1002),
.A2(n_754),
.B(n_889),
.Y(n_1161)
);

INVx4_ASAP7_75t_L g1162 ( 
.A(n_943),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_923),
.B(n_889),
.Y(n_1163)
);

OAI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_970),
.A2(n_754),
.B(n_889),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_931),
.Y(n_1165)
);

INVx2_ASAP7_75t_SL g1166 ( 
.A(n_951),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_923),
.B(n_889),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1136),
.B(n_1147),
.Y(n_1168)
);

CKINVDCx20_ASAP7_75t_R g1169 ( 
.A(n_1083),
.Y(n_1169)
);

OAI21x1_ASAP7_75t_L g1170 ( 
.A1(n_1064),
.A2(n_1130),
.B(n_1047),
.Y(n_1170)
);

INVx6_ASAP7_75t_SL g1171 ( 
.A(n_1080),
.Y(n_1171)
);

CKINVDCx11_ASAP7_75t_R g1172 ( 
.A(n_1088),
.Y(n_1172)
);

AND2x4_ASAP7_75t_L g1173 ( 
.A(n_1113),
.B(n_1119),
.Y(n_1173)
);

OAI21x1_ASAP7_75t_L g1174 ( 
.A1(n_1065),
.A2(n_1062),
.B(n_1134),
.Y(n_1174)
);

AND2x4_ASAP7_75t_L g1175 ( 
.A(n_1113),
.B(n_1119),
.Y(n_1175)
);

INVx1_ASAP7_75t_SL g1176 ( 
.A(n_1139),
.Y(n_1176)
);

AO21x2_ASAP7_75t_L g1177 ( 
.A1(n_1075),
.A2(n_1073),
.B(n_1059),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1045),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1099),
.A2(n_1063),
.B(n_1060),
.Y(n_1179)
);

NOR2xp33_ASAP7_75t_SL g1180 ( 
.A(n_1149),
.B(n_1151),
.Y(n_1180)
);

AOI22xp33_ASAP7_75t_L g1181 ( 
.A1(n_1161),
.A2(n_1167),
.B1(n_1163),
.B2(n_1142),
.Y(n_1181)
);

AO31x2_ASAP7_75t_L g1182 ( 
.A1(n_1121),
.A2(n_1103),
.A3(n_1081),
.B(n_1100),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1068),
.Y(n_1183)
);

AO21x2_ASAP7_75t_L g1184 ( 
.A1(n_1093),
.A2(n_1153),
.B(n_1135),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1095),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_1143),
.B(n_1156),
.Y(n_1186)
);

AND2x2_ASAP7_75t_L g1187 ( 
.A(n_1160),
.B(n_1094),
.Y(n_1187)
);

OAI221xp5_ASAP7_75t_L g1188 ( 
.A1(n_1148),
.A2(n_1142),
.B1(n_1097),
.B2(n_1101),
.C(n_1098),
.Y(n_1188)
);

BUFx2_ASAP7_75t_L g1189 ( 
.A(n_1154),
.Y(n_1189)
);

NAND2x1p5_ASAP7_75t_L g1190 ( 
.A(n_1141),
.B(n_1162),
.Y(n_1190)
);

CKINVDCx20_ASAP7_75t_R g1191 ( 
.A(n_1158),
.Y(n_1191)
);

AOI22xp33_ASAP7_75t_L g1192 ( 
.A1(n_1098),
.A2(n_1097),
.B1(n_1164),
.B2(n_1101),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1140),
.B(n_1044),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_1080),
.Y(n_1194)
);

AO32x2_ASAP7_75t_L g1195 ( 
.A1(n_1129),
.A2(n_1140),
.A3(n_1132),
.B1(n_1055),
.B2(n_1131),
.Y(n_1195)
);

OAI22xp5_ASAP7_75t_L g1196 ( 
.A1(n_1040),
.A2(n_1086),
.B1(n_1058),
.B2(n_1084),
.Y(n_1196)
);

OAI22xp5_ASAP7_75t_L g1197 ( 
.A1(n_1058),
.A2(n_1144),
.B1(n_1137),
.B2(n_1152),
.Y(n_1197)
);

AO31x2_ASAP7_75t_L g1198 ( 
.A1(n_1123),
.A2(n_1117),
.A3(n_1106),
.B(n_1077),
.Y(n_1198)
);

NAND3xp33_ASAP7_75t_L g1199 ( 
.A(n_1085),
.B(n_1078),
.C(n_1133),
.Y(n_1199)
);

AOI22xp33_ASAP7_75t_L g1200 ( 
.A1(n_1048),
.A2(n_1055),
.B1(n_1067),
.B2(n_1110),
.Y(n_1200)
);

AOI21x1_ASAP7_75t_L g1201 ( 
.A1(n_1043),
.A2(n_1076),
.B(n_1061),
.Y(n_1201)
);

OR2x2_ASAP7_75t_L g1202 ( 
.A(n_1138),
.B(n_1109),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_1122),
.Y(n_1203)
);

AO22x2_ASAP7_75t_L g1204 ( 
.A1(n_1078),
.A2(n_1120),
.B1(n_1049),
.B2(n_1091),
.Y(n_1204)
);

AO31x2_ASAP7_75t_L g1205 ( 
.A1(n_1052),
.A2(n_1072),
.A3(n_1079),
.B(n_1076),
.Y(n_1205)
);

OR2x6_ASAP7_75t_L g1206 ( 
.A(n_1042),
.B(n_1141),
.Y(n_1206)
);

INVx2_ASAP7_75t_SL g1207 ( 
.A(n_1155),
.Y(n_1207)
);

O2A1O1Ixp33_ASAP7_75t_SL g1208 ( 
.A1(n_1056),
.A2(n_1150),
.B(n_1115),
.C(n_1108),
.Y(n_1208)
);

OAI21x1_ASAP7_75t_L g1209 ( 
.A1(n_1051),
.A2(n_1159),
.B(n_1125),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_1089),
.Y(n_1210)
);

OAI22xp5_ASAP7_75t_L g1211 ( 
.A1(n_1165),
.A2(n_1115),
.B1(n_1070),
.B2(n_1046),
.Y(n_1211)
);

AOI22xp33_ASAP7_75t_SL g1212 ( 
.A1(n_1041),
.A2(n_1054),
.B1(n_1145),
.B2(n_1057),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1041),
.B(n_1102),
.Y(n_1213)
);

OAI22xp33_ASAP7_75t_L g1214 ( 
.A1(n_1053),
.A2(n_1096),
.B1(n_1111),
.B2(n_1050),
.Y(n_1214)
);

INVxp67_ASAP7_75t_L g1215 ( 
.A(n_1107),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1105),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_1166),
.Y(n_1217)
);

OAI21x1_ASAP7_75t_L g1218 ( 
.A1(n_1082),
.A2(n_1069),
.B(n_1124),
.Y(n_1218)
);

INVx2_ASAP7_75t_L g1219 ( 
.A(n_1126),
.Y(n_1219)
);

BUFx2_ASAP7_75t_SL g1220 ( 
.A(n_1118),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1041),
.B(n_1054),
.Y(n_1221)
);

OAI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1124),
.A2(n_1041),
.B(n_1127),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1071),
.Y(n_1223)
);

OAI22xp33_ASAP7_75t_L g1224 ( 
.A1(n_1090),
.A2(n_1066),
.B1(n_1114),
.B2(n_1128),
.Y(n_1224)
);

OAI21x1_ASAP7_75t_L g1225 ( 
.A1(n_1116),
.A2(n_1079),
.B(n_1162),
.Y(n_1225)
);

NAND2x1p5_ASAP7_75t_L g1226 ( 
.A(n_1118),
.B(n_1087),
.Y(n_1226)
);

NOR2xp33_ASAP7_75t_L g1227 ( 
.A(n_1054),
.B(n_1071),
.Y(n_1227)
);

BUFx3_ASAP7_75t_L g1228 ( 
.A(n_1074),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1146),
.A2(n_1064),
.B(n_1130),
.Y(n_1229)
);

AOI22xp33_ASAP7_75t_SL g1230 ( 
.A1(n_1146),
.A2(n_328),
.B1(n_329),
.B2(n_309),
.Y(n_1230)
);

OAI21x1_ASAP7_75t_L g1231 ( 
.A1(n_1146),
.A2(n_1064),
.B(n_1130),
.Y(n_1231)
);

BUFx4f_ASAP7_75t_L g1232 ( 
.A(n_1158),
.Y(n_1232)
);

AO32x2_ASAP7_75t_L g1233 ( 
.A1(n_1081),
.A2(n_1002),
.A3(n_1129),
.B1(n_1004),
.B2(n_826),
.Y(n_1233)
);

AND2x2_ASAP7_75t_L g1234 ( 
.A(n_1139),
.B(n_966),
.Y(n_1234)
);

OA21x2_ASAP7_75t_L g1235 ( 
.A1(n_1112),
.A2(n_1104),
.B(n_1157),
.Y(n_1235)
);

INVx6_ASAP7_75t_L g1236 ( 
.A(n_1118),
.Y(n_1236)
);

AO21x1_ASAP7_75t_L g1237 ( 
.A1(n_1132),
.A2(n_889),
.B(n_754),
.Y(n_1237)
);

INVx2_ASAP7_75t_SL g1238 ( 
.A(n_1080),
.Y(n_1238)
);

BUFx6f_ASAP7_75t_L g1239 ( 
.A(n_1118),
.Y(n_1239)
);

AO21x2_ASAP7_75t_L g1240 ( 
.A1(n_1157),
.A2(n_1075),
.B(n_1112),
.Y(n_1240)
);

O2A1O1Ixp5_ASAP7_75t_L g1241 ( 
.A1(n_1161),
.A2(n_754),
.B(n_889),
.C(n_1143),
.Y(n_1241)
);

AOI22x1_ASAP7_75t_L g1242 ( 
.A1(n_1135),
.A2(n_867),
.B1(n_868),
.B2(n_1164),
.Y(n_1242)
);

HB1xp67_ASAP7_75t_L g1243 ( 
.A(n_1079),
.Y(n_1243)
);

AOI21xp33_ASAP7_75t_L g1244 ( 
.A1(n_1142),
.A2(n_754),
.B(n_889),
.Y(n_1244)
);

AND2x2_ASAP7_75t_SL g1245 ( 
.A(n_1132),
.B(n_889),
.Y(n_1245)
);

AND2x2_ASAP7_75t_L g1246 ( 
.A(n_1139),
.B(n_966),
.Y(n_1246)
);

OAI21x1_ASAP7_75t_SL g1247 ( 
.A1(n_1121),
.A2(n_1044),
.B(n_1161),
.Y(n_1247)
);

AOI22xp5_ASAP7_75t_L g1248 ( 
.A1(n_1101),
.A2(n_867),
.B1(n_889),
.B2(n_422),
.Y(n_1248)
);

INVx2_ASAP7_75t_L g1249 ( 
.A(n_1089),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_1089),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1092),
.Y(n_1251)
);

INVx2_ASAP7_75t_SL g1252 ( 
.A(n_1080),
.Y(n_1252)
);

HB1xp67_ASAP7_75t_L g1253 ( 
.A(n_1079),
.Y(n_1253)
);

INVx3_ASAP7_75t_L g1254 ( 
.A(n_1141),
.Y(n_1254)
);

HB1xp67_ASAP7_75t_L g1255 ( 
.A(n_1079),
.Y(n_1255)
);

OR2x6_ASAP7_75t_L g1256 ( 
.A(n_1099),
.B(n_700),
.Y(n_1256)
);

AOI22xp33_ASAP7_75t_L g1257 ( 
.A1(n_1161),
.A2(n_889),
.B1(n_754),
.B2(n_852),
.Y(n_1257)
);

AOI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1101),
.A2(n_867),
.B1(n_889),
.B2(n_422),
.Y(n_1258)
);

INVx2_ASAP7_75t_L g1259 ( 
.A(n_1089),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1092),
.Y(n_1260)
);

OAI22xp5_ASAP7_75t_L g1261 ( 
.A1(n_1136),
.A2(n_1149),
.B1(n_1151),
.B2(n_1147),
.Y(n_1261)
);

AO21x2_ASAP7_75t_L g1262 ( 
.A1(n_1157),
.A2(n_1075),
.B(n_1112),
.Y(n_1262)
);

BUFx3_ASAP7_75t_L g1263 ( 
.A(n_1107),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1092),
.Y(n_1264)
);

OAI21x1_ASAP7_75t_L g1265 ( 
.A1(n_1064),
.A2(n_1130),
.B(n_1047),
.Y(n_1265)
);

INVx3_ASAP7_75t_L g1266 ( 
.A(n_1141),
.Y(n_1266)
);

OAI21x1_ASAP7_75t_L g1267 ( 
.A1(n_1064),
.A2(n_1130),
.B(n_1047),
.Y(n_1267)
);

AO31x2_ASAP7_75t_L g1268 ( 
.A1(n_1161),
.A2(n_1112),
.A3(n_1157),
.B(n_1075),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1136),
.B(n_1147),
.Y(n_1269)
);

AOI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1157),
.A2(n_754),
.B(n_1099),
.Y(n_1270)
);

O2A1O1Ixp33_ASAP7_75t_SL g1271 ( 
.A1(n_1100),
.A2(n_1143),
.B(n_1156),
.C(n_992),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_1089),
.Y(n_1272)
);

OAI22xp5_ASAP7_75t_L g1273 ( 
.A1(n_1136),
.A2(n_1149),
.B1(n_1151),
.B2(n_1147),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1092),
.Y(n_1274)
);

O2A1O1Ixp33_ASAP7_75t_L g1275 ( 
.A1(n_1143),
.A2(n_1156),
.B(n_754),
.C(n_889),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1092),
.Y(n_1276)
);

O2A1O1Ixp33_ASAP7_75t_L g1277 ( 
.A1(n_1143),
.A2(n_1156),
.B(n_754),
.C(n_889),
.Y(n_1277)
);

AOI22xp33_ASAP7_75t_L g1278 ( 
.A1(n_1161),
.A2(n_889),
.B1(n_754),
.B2(n_852),
.Y(n_1278)
);

INVx2_ASAP7_75t_SL g1279 ( 
.A(n_1080),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1092),
.Y(n_1280)
);

OA21x2_ASAP7_75t_L g1281 ( 
.A1(n_1112),
.A2(n_1104),
.B(n_1157),
.Y(n_1281)
);

NOR2xp33_ASAP7_75t_L g1282 ( 
.A(n_1136),
.B(n_889),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1178),
.Y(n_1283)
);

CKINVDCx20_ASAP7_75t_R g1284 ( 
.A(n_1172),
.Y(n_1284)
);

HB1xp67_ASAP7_75t_L g1285 ( 
.A(n_1176),
.Y(n_1285)
);

O2A1O1Ixp33_ASAP7_75t_L g1286 ( 
.A1(n_1275),
.A2(n_1277),
.B(n_1244),
.C(n_1241),
.Y(n_1286)
);

OAI22xp5_ASAP7_75t_L g1287 ( 
.A1(n_1248),
.A2(n_1258),
.B1(n_1192),
.B2(n_1282),
.Y(n_1287)
);

AOI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_1270),
.A2(n_1179),
.B(n_1275),
.Y(n_1288)
);

HB1xp67_ASAP7_75t_L g1289 ( 
.A(n_1176),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1282),
.B(n_1261),
.Y(n_1290)
);

AND2x4_ASAP7_75t_L g1291 ( 
.A(n_1183),
.B(n_1185),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_1169),
.Y(n_1292)
);

O2A1O1Ixp33_ASAP7_75t_L g1293 ( 
.A1(n_1277),
.A2(n_1244),
.B(n_1241),
.C(n_1188),
.Y(n_1293)
);

AND2x2_ASAP7_75t_L g1294 ( 
.A(n_1187),
.B(n_1234),
.Y(n_1294)
);

NOR2xp33_ASAP7_75t_L g1295 ( 
.A(n_1180),
.B(n_1261),
.Y(n_1295)
);

INVxp33_ASAP7_75t_L g1296 ( 
.A(n_1202),
.Y(n_1296)
);

NOR2xp67_ASAP7_75t_L g1297 ( 
.A(n_1238),
.B(n_1252),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1273),
.B(n_1168),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_1246),
.B(n_1180),
.Y(n_1299)
);

O2A1O1Ixp33_ASAP7_75t_L g1300 ( 
.A1(n_1188),
.A2(n_1271),
.B(n_1224),
.C(n_1273),
.Y(n_1300)
);

A2O1A1Ixp33_ASAP7_75t_L g1301 ( 
.A1(n_1270),
.A2(n_1192),
.B(n_1179),
.C(n_1186),
.Y(n_1301)
);

CKINVDCx5p33_ASAP7_75t_R g1302 ( 
.A(n_1191),
.Y(n_1302)
);

INVxp33_ASAP7_75t_L g1303 ( 
.A(n_1189),
.Y(n_1303)
);

O2A1O1Ixp5_ASAP7_75t_L g1304 ( 
.A1(n_1186),
.A2(n_1237),
.B(n_1224),
.C(n_1196),
.Y(n_1304)
);

AOI21xp5_ASAP7_75t_SL g1305 ( 
.A1(n_1256),
.A2(n_1279),
.B(n_1226),
.Y(n_1305)
);

OR2x2_ASAP7_75t_L g1306 ( 
.A(n_1196),
.B(n_1200),
.Y(n_1306)
);

AND2x2_ASAP7_75t_L g1307 ( 
.A(n_1251),
.B(n_1260),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1264),
.B(n_1274),
.Y(n_1308)
);

CKINVDCx5p33_ASAP7_75t_R g1309 ( 
.A(n_1203),
.Y(n_1309)
);

HB1xp67_ASAP7_75t_L g1310 ( 
.A(n_1197),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1168),
.B(n_1269),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_1194),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1269),
.B(n_1276),
.Y(n_1313)
);

OAI31xp33_ASAP7_75t_L g1314 ( 
.A1(n_1214),
.A2(n_1199),
.A3(n_1257),
.B(n_1278),
.Y(n_1314)
);

A2O1A1Ixp33_ASAP7_75t_L g1315 ( 
.A1(n_1257),
.A2(n_1278),
.B(n_1181),
.C(n_1193),
.Y(n_1315)
);

O2A1O1Ixp33_ASAP7_75t_L g1316 ( 
.A1(n_1214),
.A2(n_1211),
.B(n_1208),
.C(n_1215),
.Y(n_1316)
);

OR2x2_ASAP7_75t_L g1317 ( 
.A(n_1200),
.B(n_1193),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1280),
.B(n_1173),
.Y(n_1318)
);

OR2x2_ASAP7_75t_L g1319 ( 
.A(n_1207),
.B(n_1215),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1175),
.B(n_1204),
.Y(n_1320)
);

OA21x2_ASAP7_75t_L g1321 ( 
.A1(n_1209),
.A2(n_1174),
.B(n_1225),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1181),
.B(n_1216),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1210),
.B(n_1249),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1204),
.B(n_1250),
.Y(n_1324)
);

AOI21x1_ASAP7_75t_SL g1325 ( 
.A1(n_1221),
.A2(n_1213),
.B(n_1253),
.Y(n_1325)
);

OR2x2_ASAP7_75t_L g1326 ( 
.A(n_1263),
.B(n_1182),
.Y(n_1326)
);

O2A1O1Ixp5_ASAP7_75t_L g1327 ( 
.A1(n_1201),
.A2(n_1222),
.B(n_1227),
.C(n_1254),
.Y(n_1327)
);

AND2x4_ASAP7_75t_L g1328 ( 
.A(n_1218),
.B(n_1222),
.Y(n_1328)
);

O2A1O1Ixp33_ASAP7_75t_L g1329 ( 
.A1(n_1247),
.A2(n_1184),
.B(n_1206),
.C(n_1177),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_1205),
.Y(n_1330)
);

O2A1O1Ixp33_ASAP7_75t_L g1331 ( 
.A1(n_1184),
.A2(n_1206),
.B(n_1177),
.C(n_1219),
.Y(n_1331)
);

OR2x2_ASAP7_75t_L g1332 ( 
.A(n_1182),
.B(n_1259),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1204),
.B(n_1272),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_1171),
.Y(n_1334)
);

OAI22xp5_ASAP7_75t_L g1335 ( 
.A1(n_1230),
.A2(n_1212),
.B1(n_1242),
.B2(n_1232),
.Y(n_1335)
);

O2A1O1Ixp33_ASAP7_75t_L g1336 ( 
.A1(n_1227),
.A2(n_1223),
.B(n_1253),
.C(n_1243),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1245),
.B(n_1212),
.Y(n_1337)
);

AND2x2_ASAP7_75t_L g1338 ( 
.A(n_1245),
.B(n_1228),
.Y(n_1338)
);

CKINVDCx16_ASAP7_75t_R g1339 ( 
.A(n_1220),
.Y(n_1339)
);

OAI22xp5_ASAP7_75t_L g1340 ( 
.A1(n_1230),
.A2(n_1232),
.B1(n_1217),
.B2(n_1171),
.Y(n_1340)
);

OAI22xp5_ASAP7_75t_L g1341 ( 
.A1(n_1236),
.A2(n_1190),
.B1(n_1254),
.B2(n_1266),
.Y(n_1341)
);

OAI22xp5_ASAP7_75t_L g1342 ( 
.A1(n_1236),
.A2(n_1266),
.B1(n_1243),
.B2(n_1255),
.Y(n_1342)
);

O2A1O1Ixp33_ASAP7_75t_L g1343 ( 
.A1(n_1240),
.A2(n_1262),
.B(n_1281),
.C(n_1235),
.Y(n_1343)
);

AND2x4_ASAP7_75t_L g1344 ( 
.A(n_1229),
.B(n_1231),
.Y(n_1344)
);

HB1xp67_ASAP7_75t_L g1345 ( 
.A(n_1205),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1195),
.B(n_1233),
.Y(n_1346)
);

A2O1A1Ixp33_ASAP7_75t_L g1347 ( 
.A1(n_1233),
.A2(n_1170),
.B(n_1267),
.C(n_1265),
.Y(n_1347)
);

OAI31xp33_ASAP7_75t_L g1348 ( 
.A1(n_1233),
.A2(n_1268),
.A3(n_1240),
.B(n_1195),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1195),
.B(n_1205),
.Y(n_1349)
);

AOI21x1_ASAP7_75t_SL g1350 ( 
.A1(n_1198),
.A2(n_754),
.B(n_1132),
.Y(n_1350)
);

AOI21xp5_ASAP7_75t_SL g1351 ( 
.A1(n_1275),
.A2(n_637),
.B(n_647),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1282),
.B(n_1261),
.Y(n_1352)
);

CKINVDCx5p33_ASAP7_75t_R g1353 ( 
.A(n_1172),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1282),
.B(n_1261),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1282),
.B(n_1261),
.Y(n_1355)
);

BUFx6f_ASAP7_75t_L g1356 ( 
.A(n_1239),
.Y(n_1356)
);

INVx3_ASAP7_75t_SL g1357 ( 
.A(n_1194),
.Y(n_1357)
);

CKINVDCx5p33_ASAP7_75t_R g1358 ( 
.A(n_1172),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1282),
.B(n_1261),
.Y(n_1359)
);

AOI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_1270),
.A2(n_1179),
.B(n_754),
.Y(n_1360)
);

NOR2xp67_ASAP7_75t_L g1361 ( 
.A(n_1238),
.B(n_1252),
.Y(n_1361)
);

AOI21xp5_ASAP7_75t_SL g1362 ( 
.A1(n_1275),
.A2(n_637),
.B(n_647),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1245),
.B(n_1195),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1282),
.B(n_1261),
.Y(n_1364)
);

OAI22xp5_ASAP7_75t_L g1365 ( 
.A1(n_1248),
.A2(n_867),
.B1(n_1101),
.B2(n_1258),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1245),
.B(n_1195),
.Y(n_1366)
);

AOI21xp5_ASAP7_75t_L g1367 ( 
.A1(n_1360),
.A2(n_1288),
.B(n_1301),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1298),
.B(n_1290),
.Y(n_1368)
);

HB1xp67_ASAP7_75t_L g1369 ( 
.A(n_1345),
.Y(n_1369)
);

BUFx3_ASAP7_75t_L g1370 ( 
.A(n_1328),
.Y(n_1370)
);

OR2x2_ASAP7_75t_L g1371 ( 
.A(n_1349),
.B(n_1330),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1363),
.B(n_1366),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1283),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1363),
.B(n_1366),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1352),
.B(n_1354),
.Y(n_1375)
);

AND2x2_ASAP7_75t_L g1376 ( 
.A(n_1346),
.B(n_1324),
.Y(n_1376)
);

INVx2_ASAP7_75t_SL g1377 ( 
.A(n_1344),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1333),
.B(n_1348),
.Y(n_1378)
);

NAND2x1_ASAP7_75t_L g1379 ( 
.A(n_1305),
.B(n_1351),
.Y(n_1379)
);

AO21x2_ASAP7_75t_L g1380 ( 
.A1(n_1347),
.A2(n_1301),
.B(n_1343),
.Y(n_1380)
);

INVx4_ASAP7_75t_L g1381 ( 
.A(n_1291),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1328),
.B(n_1320),
.Y(n_1382)
);

AO21x2_ASAP7_75t_L g1383 ( 
.A1(n_1331),
.A2(n_1329),
.B(n_1286),
.Y(n_1383)
);

HB1xp67_ASAP7_75t_L g1384 ( 
.A(n_1332),
.Y(n_1384)
);

HB1xp67_ASAP7_75t_L g1385 ( 
.A(n_1328),
.Y(n_1385)
);

HB1xp67_ASAP7_75t_L g1386 ( 
.A(n_1342),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1291),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_1321),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_1321),
.Y(n_1389)
);

OA21x2_ASAP7_75t_L g1390 ( 
.A1(n_1304),
.A2(n_1315),
.B(n_1327),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1291),
.Y(n_1391)
);

OR2x6_ASAP7_75t_L g1392 ( 
.A(n_1344),
.B(n_1362),
.Y(n_1392)
);

OA21x2_ASAP7_75t_L g1393 ( 
.A1(n_1322),
.A2(n_1295),
.B(n_1306),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1310),
.Y(n_1394)
);

AO21x2_ASAP7_75t_L g1395 ( 
.A1(n_1293),
.A2(n_1336),
.B(n_1364),
.Y(n_1395)
);

OAI21xp5_ASAP7_75t_L g1396 ( 
.A1(n_1300),
.A2(n_1287),
.B(n_1316),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_1321),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1355),
.B(n_1359),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1326),
.Y(n_1399)
);

AND2x4_ASAP7_75t_L g1400 ( 
.A(n_1337),
.B(n_1318),
.Y(n_1400)
);

CKINVDCx11_ASAP7_75t_R g1401 ( 
.A(n_1284),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1311),
.B(n_1317),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1323),
.Y(n_1403)
);

OR2x2_ASAP7_75t_L g1404 ( 
.A(n_1285),
.B(n_1289),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1372),
.B(n_1299),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1373),
.Y(n_1406)
);

OR2x2_ASAP7_75t_L g1407 ( 
.A(n_1371),
.B(n_1296),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1373),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_1388),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1388),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1372),
.B(n_1374),
.Y(n_1411)
);

NOR2xp67_ASAP7_75t_L g1412 ( 
.A(n_1377),
.B(n_1341),
.Y(n_1412)
);

AOI22xp33_ASAP7_75t_SL g1413 ( 
.A1(n_1396),
.A2(n_1365),
.B1(n_1335),
.B2(n_1340),
.Y(n_1413)
);

OR2x6_ASAP7_75t_L g1414 ( 
.A(n_1367),
.B(n_1392),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1372),
.B(n_1338),
.Y(n_1415)
);

BUFx6f_ASAP7_75t_L g1416 ( 
.A(n_1392),
.Y(n_1416)
);

INVx1_ASAP7_75t_SL g1417 ( 
.A(n_1404),
.Y(n_1417)
);

HB1xp67_ASAP7_75t_L g1418 ( 
.A(n_1369),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1368),
.B(n_1308),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1374),
.B(n_1294),
.Y(n_1420)
);

OAI22xp5_ASAP7_75t_L g1421 ( 
.A1(n_1396),
.A2(n_1313),
.B1(n_1319),
.B2(n_1303),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1374),
.B(n_1307),
.Y(n_1422)
);

HB1xp67_ASAP7_75t_L g1423 ( 
.A(n_1384),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1385),
.B(n_1303),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1370),
.B(n_1314),
.Y(n_1425)
);

AO21x2_ASAP7_75t_L g1426 ( 
.A1(n_1367),
.A2(n_1350),
.B(n_1325),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1370),
.B(n_1376),
.Y(n_1427)
);

OR2x2_ASAP7_75t_L g1428 ( 
.A(n_1371),
.B(n_1339),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1368),
.B(n_1361),
.Y(n_1429)
);

AOI22xp33_ASAP7_75t_L g1430 ( 
.A1(n_1413),
.A2(n_1393),
.B1(n_1395),
.B2(n_1390),
.Y(n_1430)
);

OAI211xp5_ASAP7_75t_SL g1431 ( 
.A1(n_1413),
.A2(n_1375),
.B(n_1398),
.C(n_1402),
.Y(n_1431)
);

OR2x2_ASAP7_75t_L g1432 ( 
.A(n_1417),
.B(n_1407),
.Y(n_1432)
);

OR2x2_ASAP7_75t_L g1433 ( 
.A(n_1417),
.B(n_1404),
.Y(n_1433)
);

OAI22xp5_ASAP7_75t_L g1434 ( 
.A1(n_1429),
.A2(n_1379),
.B1(n_1375),
.B2(n_1398),
.Y(n_1434)
);

OR2x2_ASAP7_75t_L g1435 ( 
.A(n_1407),
.B(n_1404),
.Y(n_1435)
);

BUFx2_ASAP7_75t_R g1436 ( 
.A(n_1429),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1423),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1406),
.Y(n_1438)
);

NAND4xp25_ASAP7_75t_L g1439 ( 
.A(n_1421),
.B(n_1402),
.C(n_1394),
.D(n_1378),
.Y(n_1439)
);

INVxp67_ASAP7_75t_L g1440 ( 
.A(n_1424),
.Y(n_1440)
);

AOI22xp5_ASAP7_75t_L g1441 ( 
.A1(n_1421),
.A2(n_1379),
.B1(n_1395),
.B2(n_1393),
.Y(n_1441)
);

AOI22xp33_ASAP7_75t_SL g1442 ( 
.A1(n_1425),
.A2(n_1390),
.B1(n_1393),
.B2(n_1395),
.Y(n_1442)
);

OAI221xp5_ASAP7_75t_SL g1443 ( 
.A1(n_1414),
.A2(n_1378),
.B1(n_1386),
.B2(n_1392),
.C(n_1399),
.Y(n_1443)
);

OA21x2_ASAP7_75t_L g1444 ( 
.A1(n_1409),
.A2(n_1389),
.B(n_1397),
.Y(n_1444)
);

OR2x6_ASAP7_75t_L g1445 ( 
.A(n_1414),
.B(n_1392),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1406),
.Y(n_1446)
);

OAI31xp33_ASAP7_75t_SL g1447 ( 
.A1(n_1425),
.A2(n_1378),
.A3(n_1382),
.B(n_1400),
.Y(n_1447)
);

AOI221xp5_ASAP7_75t_L g1448 ( 
.A1(n_1425),
.A2(n_1395),
.B1(n_1387),
.B2(n_1391),
.C(n_1399),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1419),
.B(n_1393),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1411),
.B(n_1382),
.Y(n_1450)
);

NAND4xp25_ASAP7_75t_L g1451 ( 
.A(n_1412),
.B(n_1394),
.C(n_1297),
.D(n_1403),
.Y(n_1451)
);

OAI211xp5_ASAP7_75t_L g1452 ( 
.A1(n_1412),
.A2(n_1390),
.B(n_1393),
.C(n_1386),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1423),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1411),
.B(n_1382),
.Y(n_1454)
);

BUFx3_ASAP7_75t_L g1455 ( 
.A(n_1424),
.Y(n_1455)
);

HB1xp67_ASAP7_75t_L g1456 ( 
.A(n_1418),
.Y(n_1456)
);

OAI22xp5_ASAP7_75t_L g1457 ( 
.A1(n_1428),
.A2(n_1390),
.B1(n_1419),
.B2(n_1414),
.Y(n_1457)
);

AOI22xp33_ASAP7_75t_L g1458 ( 
.A1(n_1414),
.A2(n_1395),
.B1(n_1390),
.B2(n_1381),
.Y(n_1458)
);

AO21x2_ASAP7_75t_L g1459 ( 
.A1(n_1410),
.A2(n_1397),
.B(n_1389),
.Y(n_1459)
);

NOR2x1_ASAP7_75t_L g1460 ( 
.A(n_1426),
.B(n_1383),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1408),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1418),
.Y(n_1462)
);

AOI22xp33_ASAP7_75t_L g1463 ( 
.A1(n_1414),
.A2(n_1381),
.B1(n_1400),
.B2(n_1383),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1407),
.Y(n_1464)
);

BUFx2_ASAP7_75t_L g1465 ( 
.A(n_1445),
.Y(n_1465)
);

INVx3_ASAP7_75t_L g1466 ( 
.A(n_1444),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1450),
.B(n_1411),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_SL g1468 ( 
.A(n_1430),
.B(n_1416),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1438),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1449),
.B(n_1422),
.Y(n_1470)
);

INVx3_ASAP7_75t_L g1471 ( 
.A(n_1459),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1438),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1446),
.Y(n_1473)
);

CKINVDCx5p33_ASAP7_75t_R g1474 ( 
.A(n_1436),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1462),
.B(n_1422),
.Y(n_1475)
);

NOR2x1_ASAP7_75t_L g1476 ( 
.A(n_1452),
.B(n_1426),
.Y(n_1476)
);

INVxp67_ASAP7_75t_SL g1477 ( 
.A(n_1456),
.Y(n_1477)
);

HB1xp67_ASAP7_75t_L g1478 ( 
.A(n_1461),
.Y(n_1478)
);

NOR2x1_ASAP7_75t_L g1479 ( 
.A(n_1460),
.B(n_1426),
.Y(n_1479)
);

INVx4_ASAP7_75t_L g1480 ( 
.A(n_1445),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1437),
.B(n_1422),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1461),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1464),
.Y(n_1483)
);

HB1xp67_ASAP7_75t_L g1484 ( 
.A(n_1432),
.Y(n_1484)
);

INVxp67_ASAP7_75t_L g1485 ( 
.A(n_1453),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1435),
.Y(n_1486)
);

INVx1_ASAP7_75t_SL g1487 ( 
.A(n_1433),
.Y(n_1487)
);

BUFx3_ASAP7_75t_L g1488 ( 
.A(n_1445),
.Y(n_1488)
);

INVx4_ASAP7_75t_SL g1489 ( 
.A(n_1445),
.Y(n_1489)
);

CKINVDCx20_ASAP7_75t_R g1490 ( 
.A(n_1434),
.Y(n_1490)
);

INVx3_ASAP7_75t_L g1491 ( 
.A(n_1480),
.Y(n_1491)
);

AND2x4_ASAP7_75t_L g1492 ( 
.A(n_1489),
.B(n_1450),
.Y(n_1492)
);

NAND3xp33_ASAP7_75t_L g1493 ( 
.A(n_1476),
.B(n_1441),
.C(n_1442),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1467),
.B(n_1454),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1487),
.B(n_1420),
.Y(n_1495)
);

OR2x2_ASAP7_75t_L g1496 ( 
.A(n_1487),
.B(n_1435),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_SL g1497 ( 
.A(n_1474),
.B(n_1447),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1466),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1478),
.Y(n_1499)
);

NOR3xp33_ASAP7_75t_L g1500 ( 
.A(n_1468),
.B(n_1431),
.C(n_1476),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1478),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1484),
.B(n_1420),
.Y(n_1502)
);

INVx1_ASAP7_75t_SL g1503 ( 
.A(n_1474),
.Y(n_1503)
);

OR2x2_ASAP7_75t_L g1504 ( 
.A(n_1470),
.B(n_1484),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1482),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1482),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1475),
.B(n_1448),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1482),
.Y(n_1508)
);

OAI321xp33_ASAP7_75t_L g1509 ( 
.A1(n_1468),
.A2(n_1439),
.A3(n_1443),
.B1(n_1457),
.B2(n_1458),
.C(n_1451),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1469),
.Y(n_1510)
);

OR2x2_ASAP7_75t_L g1511 ( 
.A(n_1486),
.B(n_1432),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1467),
.B(n_1454),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1469),
.Y(n_1513)
);

AND2x4_ASAP7_75t_L g1514 ( 
.A(n_1489),
.B(n_1416),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1467),
.B(n_1455),
.Y(n_1515)
);

INVx1_ASAP7_75t_SL g1516 ( 
.A(n_1490),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1465),
.B(n_1455),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1465),
.B(n_1440),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1465),
.B(n_1427),
.Y(n_1519)
);

BUFx3_ASAP7_75t_L g1520 ( 
.A(n_1490),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1481),
.B(n_1486),
.Y(n_1521)
);

OAI221xp5_ASAP7_75t_L g1522 ( 
.A1(n_1480),
.A2(n_1463),
.B1(n_1414),
.B2(n_1428),
.C(n_1416),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1472),
.Y(n_1523)
);

HB1xp67_ASAP7_75t_L g1524 ( 
.A(n_1485),
.Y(n_1524)
);

NOR2x1_ASAP7_75t_L g1525 ( 
.A(n_1479),
.B(n_1284),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1472),
.Y(n_1526)
);

NOR2xp33_ASAP7_75t_L g1527 ( 
.A(n_1480),
.B(n_1401),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1489),
.B(n_1427),
.Y(n_1528)
);

AOI22xp33_ASAP7_75t_L g1529 ( 
.A1(n_1488),
.A2(n_1416),
.B1(n_1383),
.B2(n_1380),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1492),
.B(n_1489),
.Y(n_1530)
);

OR2x2_ASAP7_75t_L g1531 ( 
.A(n_1504),
.B(n_1477),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1516),
.B(n_1485),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1505),
.Y(n_1533)
);

NOR2xp33_ASAP7_75t_SL g1534 ( 
.A(n_1503),
.B(n_1480),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1498),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1524),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1520),
.B(n_1483),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1505),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1492),
.B(n_1489),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1498),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1506),
.Y(n_1541)
);

INVxp67_ASAP7_75t_L g1542 ( 
.A(n_1520),
.Y(n_1542)
);

OR2x2_ASAP7_75t_L g1543 ( 
.A(n_1504),
.B(n_1477),
.Y(n_1543)
);

OR2x2_ASAP7_75t_L g1544 ( 
.A(n_1496),
.B(n_1473),
.Y(n_1544)
);

NOR2x1_ASAP7_75t_L g1545 ( 
.A(n_1497),
.B(n_1479),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1506),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1492),
.B(n_1489),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1515),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1510),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1510),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1500),
.B(n_1415),
.Y(n_1551)
);

OR2x2_ASAP7_75t_L g1552 ( 
.A(n_1496),
.B(n_1473),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1508),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1518),
.B(n_1415),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1515),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1528),
.B(n_1489),
.Y(n_1556)
);

OAI21xp33_ASAP7_75t_SL g1557 ( 
.A1(n_1525),
.A2(n_1480),
.B(n_1466),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1518),
.B(n_1405),
.Y(n_1558)
);

AO22x1_ASAP7_75t_L g1559 ( 
.A1(n_1527),
.A2(n_1358),
.B1(n_1353),
.B2(n_1357),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1528),
.B(n_1517),
.Y(n_1560)
);

NOR3xp33_ASAP7_75t_L g1561 ( 
.A(n_1509),
.B(n_1401),
.C(n_1488),
.Y(n_1561)
);

INVxp67_ASAP7_75t_L g1562 ( 
.A(n_1517),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1499),
.Y(n_1563)
);

AOI22xp33_ASAP7_75t_L g1564 ( 
.A1(n_1493),
.A2(n_1488),
.B1(n_1416),
.B2(n_1383),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1514),
.B(n_1488),
.Y(n_1565)
);

NAND3xp33_ASAP7_75t_SL g1566 ( 
.A(n_1561),
.B(n_1529),
.C(n_1522),
.Y(n_1566)
);

HB1xp67_ASAP7_75t_L g1567 ( 
.A(n_1542),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1560),
.B(n_1491),
.Y(n_1568)
);

OAI22xp5_ASAP7_75t_L g1569 ( 
.A1(n_1545),
.A2(n_1507),
.B1(n_1514),
.B2(n_1502),
.Y(n_1569)
);

CKINVDCx16_ASAP7_75t_R g1570 ( 
.A(n_1534),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1562),
.B(n_1519),
.Y(n_1571)
);

BUFx2_ASAP7_75t_L g1572 ( 
.A(n_1557),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1533),
.Y(n_1573)
);

AOI22xp33_ASAP7_75t_L g1574 ( 
.A1(n_1564),
.A2(n_1514),
.B1(n_1491),
.B2(n_1416),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1560),
.B(n_1491),
.Y(n_1575)
);

AND2x4_ASAP7_75t_L g1576 ( 
.A(n_1556),
.B(n_1499),
.Y(n_1576)
);

OR2x2_ASAP7_75t_L g1577 ( 
.A(n_1531),
.B(n_1511),
.Y(n_1577)
);

BUFx2_ASAP7_75t_L g1578 ( 
.A(n_1548),
.Y(n_1578)
);

NAND2x1p5_ASAP7_75t_L g1579 ( 
.A(n_1556),
.B(n_1519),
.Y(n_1579)
);

NAND2x1p5_ASAP7_75t_L g1580 ( 
.A(n_1530),
.B(n_1501),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1565),
.B(n_1494),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1536),
.B(n_1494),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1533),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1565),
.B(n_1512),
.Y(n_1584)
);

INVx2_ASAP7_75t_SL g1585 ( 
.A(n_1530),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1539),
.B(n_1547),
.Y(n_1586)
);

AO22x1_ASAP7_75t_L g1587 ( 
.A1(n_1563),
.A2(n_1358),
.B1(n_1353),
.B2(n_1357),
.Y(n_1587)
);

NOR2xp33_ASAP7_75t_L g1588 ( 
.A(n_1559),
.B(n_1302),
.Y(n_1588)
);

INVx3_ASAP7_75t_L g1589 ( 
.A(n_1539),
.Y(n_1589)
);

AOI22xp33_ASAP7_75t_L g1590 ( 
.A1(n_1551),
.A2(n_1416),
.B1(n_1383),
.B2(n_1380),
.Y(n_1590)
);

AOI222xp33_ASAP7_75t_L g1591 ( 
.A1(n_1566),
.A2(n_1532),
.B1(n_1537),
.B2(n_1559),
.C1(n_1555),
.C2(n_1548),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1578),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1578),
.Y(n_1593)
);

OAI22xp5_ASAP7_75t_L g1594 ( 
.A1(n_1570),
.A2(n_1572),
.B1(n_1579),
.B2(n_1569),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1586),
.B(n_1555),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_SL g1596 ( 
.A(n_1570),
.B(n_1547),
.Y(n_1596)
);

NAND3xp33_ASAP7_75t_L g1597 ( 
.A(n_1567),
.B(n_1563),
.C(n_1543),
.Y(n_1597)
);

NAND2xp33_ASAP7_75t_SL g1598 ( 
.A(n_1572),
.B(n_1334),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1573),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1586),
.B(n_1512),
.Y(n_1600)
);

AOI21xp33_ASAP7_75t_SL g1601 ( 
.A1(n_1587),
.A2(n_1543),
.B(n_1531),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1573),
.Y(n_1602)
);

AOI22xp5_ASAP7_75t_L g1603 ( 
.A1(n_1588),
.A2(n_1558),
.B1(n_1554),
.B2(n_1553),
.Y(n_1603)
);

INVx2_ASAP7_75t_SL g1604 ( 
.A(n_1579),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1581),
.B(n_1495),
.Y(n_1605)
);

NOR2xp33_ASAP7_75t_L g1606 ( 
.A(n_1587),
.B(n_1585),
.Y(n_1606)
);

OR2x2_ASAP7_75t_L g1607 ( 
.A(n_1571),
.B(n_1511),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1583),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1576),
.B(n_1549),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1576),
.B(n_1549),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1592),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1591),
.B(n_1576),
.Y(n_1612)
);

INVxp67_ASAP7_75t_L g1613 ( 
.A(n_1593),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1595),
.B(n_1576),
.Y(n_1614)
);

INVx1_ASAP7_75t_SL g1615 ( 
.A(n_1598),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1609),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1601),
.B(n_1585),
.Y(n_1617)
);

OR2x2_ASAP7_75t_L g1618 ( 
.A(n_1607),
.B(n_1582),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1610),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1600),
.B(n_1581),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1606),
.B(n_1589),
.Y(n_1621)
);

NOR4xp25_ASAP7_75t_SL g1622 ( 
.A(n_1611),
.B(n_1598),
.C(n_1596),
.D(n_1599),
.Y(n_1622)
);

OAI22xp5_ASAP7_75t_L g1623 ( 
.A1(n_1612),
.A2(n_1597),
.B1(n_1579),
.B2(n_1594),
.Y(n_1623)
);

OAI21xp5_ASAP7_75t_L g1624 ( 
.A1(n_1617),
.A2(n_1596),
.B(n_1606),
.Y(n_1624)
);

AOI221x1_ASAP7_75t_L g1625 ( 
.A1(n_1621),
.A2(n_1608),
.B1(n_1602),
.B2(n_1589),
.C(n_1583),
.Y(n_1625)
);

AOI21xp5_ASAP7_75t_L g1626 ( 
.A1(n_1615),
.A2(n_1604),
.B(n_1589),
.Y(n_1626)
);

AOI32xp33_ASAP7_75t_L g1627 ( 
.A1(n_1620),
.A2(n_1604),
.A3(n_1589),
.B1(n_1568),
.B2(n_1575),
.Y(n_1627)
);

NOR4xp25_ASAP7_75t_L g1628 ( 
.A(n_1613),
.B(n_1574),
.C(n_1577),
.D(n_1590),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1613),
.Y(n_1629)
);

OAI21xp5_ASAP7_75t_SL g1630 ( 
.A1(n_1614),
.A2(n_1603),
.B(n_1580),
.Y(n_1630)
);

XNOR2x1_ASAP7_75t_L g1631 ( 
.A(n_1623),
.B(n_1624),
.Y(n_1631)
);

AOI21xp33_ASAP7_75t_SL g1632 ( 
.A1(n_1628),
.A2(n_1630),
.B(n_1621),
.Y(n_1632)
);

OA22x2_ASAP7_75t_L g1633 ( 
.A1(n_1625),
.A2(n_1619),
.B1(n_1616),
.B2(n_1575),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1629),
.Y(n_1634)
);

AOI221xp5_ASAP7_75t_L g1635 ( 
.A1(n_1627),
.A2(n_1626),
.B1(n_1618),
.B2(n_1622),
.C(n_1568),
.Y(n_1635)
);

INVx1_ASAP7_75t_SL g1636 ( 
.A(n_1631),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1633),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_SL g1638 ( 
.A(n_1635),
.B(n_1577),
.Y(n_1638)
);

AOI22xp5_ASAP7_75t_L g1639 ( 
.A1(n_1634),
.A2(n_1580),
.B1(n_1584),
.B2(n_1605),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1632),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1635),
.B(n_1584),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1639),
.Y(n_1642)
);

AOI221xp5_ASAP7_75t_L g1643 ( 
.A1(n_1640),
.A2(n_1580),
.B1(n_1550),
.B2(n_1535),
.C(n_1540),
.Y(n_1643)
);

NOR2x1_ASAP7_75t_L g1644 ( 
.A(n_1637),
.B(n_1550),
.Y(n_1644)
);

OAI21xp5_ASAP7_75t_L g1645 ( 
.A1(n_1638),
.A2(n_1538),
.B(n_1541),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1641),
.Y(n_1646)
);

NOR2x1_ASAP7_75t_L g1647 ( 
.A(n_1644),
.B(n_1636),
.Y(n_1647)
);

AND2x4_ASAP7_75t_L g1648 ( 
.A(n_1642),
.B(n_1302),
.Y(n_1648)
);

OAI211xp5_ASAP7_75t_L g1649 ( 
.A1(n_1646),
.A2(n_1334),
.B(n_1312),
.C(n_1309),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1647),
.Y(n_1650)
);

OAI221xp5_ASAP7_75t_L g1651 ( 
.A1(n_1650),
.A2(n_1645),
.B1(n_1649),
.B2(n_1643),
.C(n_1648),
.Y(n_1651)
);

AOI22x1_ASAP7_75t_L g1652 ( 
.A1(n_1651),
.A2(n_1312),
.B1(n_1309),
.B2(n_1292),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1651),
.B(n_1535),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1652),
.Y(n_1654)
);

NAND2x1p5_ASAP7_75t_L g1655 ( 
.A(n_1653),
.B(n_1292),
.Y(n_1655)
);

OAI22xp5_ASAP7_75t_SL g1656 ( 
.A1(n_1655),
.A2(n_1546),
.B1(n_1538),
.B2(n_1541),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1654),
.Y(n_1657)
);

OAI22xp5_ASAP7_75t_L g1658 ( 
.A1(n_1657),
.A2(n_1540),
.B1(n_1546),
.B2(n_1544),
.Y(n_1658)
);

NAND2x1p5_ASAP7_75t_L g1659 ( 
.A(n_1658),
.B(n_1656),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1659),
.B(n_1544),
.Y(n_1660)
);

AOI22xp33_ASAP7_75t_SL g1661 ( 
.A1(n_1660),
.A2(n_1552),
.B1(n_1526),
.B2(n_1513),
.Y(n_1661)
);

AOI22xp5_ASAP7_75t_L g1662 ( 
.A1(n_1661),
.A2(n_1552),
.B1(n_1523),
.B2(n_1521),
.Y(n_1662)
);

AOI22xp33_ASAP7_75t_SL g1663 ( 
.A1(n_1662),
.A2(n_1356),
.B1(n_1471),
.B2(n_1466),
.Y(n_1663)
);


endmodule