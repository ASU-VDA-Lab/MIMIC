module fake_jpeg_14603_n_79 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_79);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_79;

wire n_10;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_8;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

INVx1_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

INVx2_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

INVx8_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_2),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_20),
.Y(n_25)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_21),
.B(n_22),
.Y(n_23)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_23),
.B(n_8),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_33),
.Y(n_38)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_29),
.B(n_30),
.Y(n_34)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g31 ( 
.A1(n_25),
.A2(n_19),
.B(n_15),
.Y(n_31)
);

XNOR2xp5_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_17),
.Y(n_36)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_32),
.B(n_26),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_10),
.Y(n_33)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_SL g43 ( 
.A1(n_36),
.A2(n_24),
.B(n_20),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_27),
.Y(n_37)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_32),
.A2(n_21),
.B1(n_26),
.B2(n_25),
.Y(n_39)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_39),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_8),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_40),
.B(n_13),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_27),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_41),
.B(n_43),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_45),
.B(n_12),
.Y(n_52)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_47),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_46),
.A2(n_36),
.B1(n_24),
.B2(n_38),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_50),
.A2(n_42),
.B1(n_24),
.B2(n_17),
.Y(n_57)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_53),
.Y(n_55)
);

BUFx24_ASAP7_75t_SL g58 ( 
.A(n_52),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_41),
.B(n_12),
.Y(n_53)
);

INVxp67_ASAP7_75t_SL g54 ( 
.A(n_42),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g56 ( 
.A(n_50),
.B(n_43),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_56),
.B(n_22),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_57),
.B(n_59),
.Y(n_62)
);

XOR2xp5_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_51),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_60),
.B(n_48),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_64),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_65),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_58),
.B(n_4),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_62),
.A2(n_0),
.B(n_1),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_66),
.A2(n_5),
.B(n_6),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g67 ( 
.A(n_61),
.B(n_15),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_67),
.B(n_18),
.Y(n_70)
);

AOI322xp5_ASAP7_75t_L g74 ( 
.A1(n_70),
.A2(n_72),
.A3(n_73),
.B1(n_22),
.B2(n_3),
.C1(n_0),
.C2(n_14),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_69),
.B(n_9),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_71),
.A2(n_16),
.B(n_11),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g73 ( 
.A1(n_68),
.A2(n_5),
.B(n_3),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_74),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_75),
.Y(n_77)
);

O2A1O1Ixp33_ASAP7_75t_SL g78 ( 
.A1(n_76),
.A2(n_0),
.B(n_3),
.C(n_11),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_78),
.B(n_77),
.Y(n_79)
);


endmodule