module fake_jpeg_32014_n_64 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_64);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_64;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_22;
wire n_51;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_43;
wire n_37;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

INVx1_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_4),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

INVxp67_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_5),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_11),
.B(n_0),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_18),
.B(n_19),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_11),
.B(n_0),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_20),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_8),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_21),
.B(n_1),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_25),
.A2(n_9),
.B1(n_12),
.B2(n_15),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_18),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_26),
.B(n_18),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_27),
.B(n_30),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_24),
.A2(n_17),
.B1(n_20),
.B2(n_13),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_29),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g29 ( 
.A1(n_24),
.A2(n_21),
.B(n_20),
.Y(n_29)
);

OR2x2_ASAP7_75t_L g30 ( 
.A(n_22),
.B(n_21),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_22),
.B(n_15),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_33),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_8),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_34),
.B(n_35),
.C(n_20),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_SL g35 ( 
.A(n_25),
.B(n_14),
.C(n_4),
.Y(n_35)
);

A2O1A1Ixp33_ASAP7_75t_L g36 ( 
.A1(n_24),
.A2(n_10),
.B(n_7),
.C(n_6),
.Y(n_36)
);

NOR3xp33_ASAP7_75t_L g38 ( 
.A(n_36),
.B(n_10),
.C(n_14),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_39),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_14),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_42),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_43),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_29),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_49),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_34),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_46),
.B(n_37),
.C(n_41),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_30),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_51),
.B(n_47),
.C(n_48),
.Y(n_57)
);

OAI21xp33_ASAP7_75t_L g53 ( 
.A1(n_49),
.A2(n_35),
.B(n_36),
.Y(n_53)
);

NAND2xp33_ASAP7_75t_SL g55 ( 
.A(n_53),
.B(n_50),
.Y(n_55)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_54),
.B(n_46),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_55),
.B(n_56),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_57),
.A2(n_52),
.B1(n_53),
.B2(n_44),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_L g60 ( 
.A1(n_58),
.A2(n_57),
.B(n_14),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_60),
.A2(n_61),
.B1(n_59),
.B2(n_5),
.Y(n_62)
);

AOI31xp67_ASAP7_75t_L g61 ( 
.A1(n_58),
.A2(n_43),
.A3(n_4),
.B(n_5),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_62),
.A2(n_2),
.B(n_17),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_63),
.Y(n_64)
);


endmodule