module real_jpeg_705_n_8 (n_5, n_4, n_0, n_1, n_2, n_6, n_7, n_3, n_8);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_8;

wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_49;
wire n_10;
wire n_68;
wire n_78;
wire n_83;
wire n_64;
wire n_47;
wire n_11;
wire n_22;
wire n_40;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_44;
wire n_28;
wire n_62;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_9;
wire n_72;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_61;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_24;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_85;
wire n_16;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_2),
.A2(n_16),
.B1(n_31),
.B2(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_2),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_2),
.A2(n_19),
.B1(n_26),
.B2(n_47),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_3),
.Y(n_80)
);

BUFx16f_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

MAJIxp5_ASAP7_75t_L g13 ( 
.A(n_5),
.B(n_14),
.C(n_16),
.Y(n_13)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_5),
.A2(n_19),
.B1(n_26),
.B2(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_5),
.B(n_44),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_5),
.A2(n_16),
.B1(n_31),
.B2(n_34),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_5),
.B(n_27),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_5),
.B(n_78),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_6),
.A2(n_19),
.B1(n_25),
.B2(n_26),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_6),
.A2(n_16),
.B1(n_25),
.B2(n_31),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g8 ( 
.A(n_9),
.B(n_63),
.Y(n_8)
);

OAI21xp5_ASAP7_75t_SL g9 ( 
.A1(n_10),
.A2(n_49),
.B(n_62),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_SL g10 ( 
.A(n_11),
.B(n_39),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_11),
.B(n_39),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g11 ( 
.A1(n_12),
.A2(n_22),
.B1(n_37),
.B2(n_38),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_12),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g12 ( 
.A(n_13),
.B(n_19),
.Y(n_12)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_14),
.A2(n_16),
.B1(n_30),
.B2(n_31),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_14),
.A2(n_19),
.B1(n_26),
.B2(n_30),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_16),
.B(n_43),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_16),
.B(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_19),
.A2(n_26),
.B1(n_80),
.B2(n_81),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_22),
.B(n_37),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_32),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_27),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_24),
.B(n_35),
.Y(n_76)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_29),
.B(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_35),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_45),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_41),
.B(n_54),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_42),
.B(n_43),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_48),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_43),
.B(n_46),
.Y(n_59)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_44),
.B(n_69),
.Y(n_68)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_48),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_55),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_56),
.B(n_61),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_53),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_57),
.B(n_60),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_57),
.B(n_60),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_58),
.B(n_59),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_86),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_85),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_66),
.B(n_85),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_71),
.B1(n_72),
.B2(n_84),
.Y(n_66)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_70),
.Y(n_67)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_73),
.A2(n_77),
.B1(n_82),
.B2(n_83),
.Y(n_72)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_76),
.Y(n_73)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_77),
.Y(n_83)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx3_ASAP7_75t_SL g81 ( 
.A(n_80),
.Y(n_81)
);


endmodule