module real_aes_6323_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_357;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_741;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g267 ( .A1(n_0), .A2(n_268), .B(n_269), .C(n_272), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_1), .B(n_209), .Y(n_273) );
NAND3xp33_ASAP7_75t_SL g110 ( .A(n_2), .B(n_92), .C(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g448 ( .A(n_2), .Y(n_448) );
NAND2xp5_ASAP7_75t_SL g245 ( .A(n_3), .B(n_179), .Y(n_245) );
A2O1A1Ixp33_ASAP7_75t_L g476 ( .A1(n_4), .A2(n_149), .B(n_152), .C(n_477), .Y(n_476) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_5), .A2(n_169), .B(n_517), .Y(n_516) );
AOI21xp5_ASAP7_75t_L g199 ( .A1(n_6), .A2(n_169), .B(n_200), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_7), .B(n_209), .Y(n_523) );
AO21x2_ASAP7_75t_L g188 ( .A1(n_8), .A2(n_136), .B(n_189), .Y(n_188) );
OAI22xp5_ASAP7_75t_SL g739 ( .A1(n_9), .A2(n_740), .B1(n_743), .B2(n_744), .Y(n_739) );
CKINVDCx20_ASAP7_75t_R g744 ( .A(n_9), .Y(n_744) );
AND2x6_ASAP7_75t_L g149 ( .A(n_10), .B(n_150), .Y(n_149) );
A2O1A1Ixp33_ASAP7_75t_L g151 ( .A1(n_11), .A2(n_149), .B(n_152), .C(n_155), .Y(n_151) );
INVx1_ASAP7_75t_L g493 ( .A(n_12), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g108 ( .A(n_13), .B(n_41), .Y(n_108) );
OAI22xp5_ASAP7_75t_L g740 ( .A1(n_14), .A2(n_45), .B1(n_741), .B2(n_742), .Y(n_740) );
CKINVDCx20_ASAP7_75t_R g741 ( .A(n_14), .Y(n_741) );
NAND2xp5_ASAP7_75t_SL g479 ( .A(n_15), .B(n_159), .Y(n_479) );
INVx1_ASAP7_75t_L g141 ( .A(n_16), .Y(n_141) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_17), .B(n_179), .Y(n_195) );
A2O1A1Ixp33_ASAP7_75t_L g500 ( .A1(n_18), .A2(n_157), .B(n_501), .C(n_503), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_19), .B(n_209), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_20), .B(n_233), .Y(n_536) );
A2O1A1Ixp33_ASAP7_75t_L g228 ( .A1(n_21), .A2(n_152), .B(n_196), .C(n_229), .Y(n_228) );
A2O1A1Ixp33_ASAP7_75t_L g509 ( .A1(n_22), .A2(n_161), .B(n_271), .C(n_510), .Y(n_509) );
NAND2xp5_ASAP7_75t_SL g555 ( .A(n_23), .B(n_159), .Y(n_555) );
NAND2xp5_ASAP7_75t_SL g544 ( .A(n_24), .B(n_159), .Y(n_544) );
CKINVDCx16_ASAP7_75t_R g551 ( .A(n_25), .Y(n_551) );
INVx1_ASAP7_75t_L g543 ( .A(n_26), .Y(n_543) );
A2O1A1Ixp33_ASAP7_75t_L g191 ( .A1(n_27), .A2(n_152), .B(n_192), .C(n_196), .Y(n_191) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_28), .Y(n_148) );
CKINVDCx20_ASAP7_75t_R g475 ( .A(n_29), .Y(n_475) );
INVx1_ASAP7_75t_L g534 ( .A(n_30), .Y(n_534) );
AOI21xp5_ASAP7_75t_L g264 ( .A1(n_31), .A2(n_169), .B(n_265), .Y(n_264) );
INVx2_ASAP7_75t_L g147 ( .A(n_32), .Y(n_147) );
A2O1A1Ixp33_ASAP7_75t_L g216 ( .A1(n_33), .A2(n_171), .B(n_182), .C(n_217), .Y(n_216) );
CKINVDCx20_ASAP7_75t_R g482 ( .A(n_34), .Y(n_482) );
A2O1A1Ixp33_ASAP7_75t_L g519 ( .A1(n_35), .A2(n_271), .B(n_520), .C(n_522), .Y(n_519) );
INVxp67_ASAP7_75t_L g535 ( .A(n_36), .Y(n_535) );
OAI22xp5_ASAP7_75t_SL g449 ( .A1(n_37), .A2(n_79), .B1(n_450), .B2(n_451), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_37), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_38), .B(n_194), .Y(n_193) );
CKINVDCx14_ASAP7_75t_R g518 ( .A(n_39), .Y(n_518) );
A2O1A1Ixp33_ASAP7_75t_L g541 ( .A1(n_40), .A2(n_152), .B(n_196), .C(n_542), .Y(n_541) );
A2O1A1Ixp33_ASAP7_75t_L g490 ( .A1(n_42), .A2(n_272), .B(n_491), .C(n_492), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_43), .B(n_227), .Y(n_226) );
CKINVDCx20_ASAP7_75t_R g164 ( .A(n_44), .Y(n_164) );
INVx1_ASAP7_75t_L g742 ( .A(n_45), .Y(n_742) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_46), .A2(n_105), .B1(n_114), .B2(n_753), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_47), .B(n_179), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_48), .B(n_169), .Y(n_190) );
CKINVDCx20_ASAP7_75t_R g546 ( .A(n_49), .Y(n_546) );
CKINVDCx20_ASAP7_75t_R g531 ( .A(n_50), .Y(n_531) );
A2O1A1Ixp33_ASAP7_75t_L g170 ( .A1(n_51), .A2(n_171), .B(n_173), .C(n_182), .Y(n_170) );
INVx1_ASAP7_75t_L g270 ( .A(n_52), .Y(n_270) );
INVx1_ASAP7_75t_L g174 ( .A(n_53), .Y(n_174) );
AOI222xp33_ASAP7_75t_L g460 ( .A1(n_54), .A2(n_461), .B1(n_735), .B2(n_736), .C1(n_745), .C2(n_748), .Y(n_460) );
INVx1_ASAP7_75t_L g508 ( .A(n_55), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_56), .B(n_169), .Y(n_168) );
OAI22xp5_ASAP7_75t_SL g123 ( .A1(n_57), .A2(n_60), .B1(n_124), .B2(n_125), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_57), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g236 ( .A(n_58), .Y(n_236) );
CKINVDCx14_ASAP7_75t_R g489 ( .A(n_59), .Y(n_489) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_60), .Y(n_124) );
INVx1_ASAP7_75t_L g150 ( .A(n_61), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_62), .B(n_169), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_63), .B(n_209), .Y(n_208) );
A2O1A1Ixp33_ASAP7_75t_L g202 ( .A1(n_64), .A2(n_203), .B(n_205), .C(n_207), .Y(n_202) );
INVx1_ASAP7_75t_L g140 ( .A(n_65), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_66), .B(n_457), .Y(n_456) );
INVx1_ASAP7_75t_SL g521 ( .A(n_67), .Y(n_521) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_68), .Y(n_119) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_69), .B(n_179), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_70), .B(n_209), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_71), .B(n_157), .Y(n_156) );
INVx1_ASAP7_75t_L g554 ( .A(n_72), .Y(n_554) );
CKINVDCx16_ASAP7_75t_R g266 ( .A(n_73), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_74), .B(n_176), .Y(n_230) );
A2O1A1Ixp33_ASAP7_75t_L g242 ( .A1(n_75), .A2(n_152), .B(n_182), .C(n_243), .Y(n_242) );
CKINVDCx16_ASAP7_75t_R g201 ( .A(n_76), .Y(n_201) );
INVx1_ASAP7_75t_L g113 ( .A(n_77), .Y(n_113) );
AOI21xp5_ASAP7_75t_L g487 ( .A1(n_78), .A2(n_169), .B(n_488), .Y(n_487) );
CKINVDCx20_ASAP7_75t_R g451 ( .A(n_79), .Y(n_451) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_80), .A2(n_169), .B(n_498), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_81), .A2(n_227), .B(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g499 ( .A(n_82), .Y(n_499) );
CKINVDCx16_ASAP7_75t_R g540 ( .A(n_83), .Y(n_540) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_84), .B(n_175), .Y(n_231) );
CKINVDCx20_ASAP7_75t_R g221 ( .A(n_85), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_86), .A2(n_169), .B(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g502 ( .A(n_87), .Y(n_502) );
INVx2_ASAP7_75t_L g138 ( .A(n_88), .Y(n_138) );
INVx1_ASAP7_75t_L g478 ( .A(n_89), .Y(n_478) );
CKINVDCx20_ASAP7_75t_R g250 ( .A(n_90), .Y(n_250) );
NAND2xp5_ASAP7_75t_SL g158 ( .A(n_91), .B(n_159), .Y(n_158) );
OR2x2_ASAP7_75t_L g445 ( .A(n_92), .B(n_446), .Y(n_445) );
OR2x2_ASAP7_75t_L g464 ( .A(n_92), .B(n_447), .Y(n_464) );
INVx2_ASAP7_75t_L g734 ( .A(n_92), .Y(n_734) );
A2O1A1Ixp33_ASAP7_75t_L g552 ( .A1(n_93), .A2(n_152), .B(n_182), .C(n_553), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_94), .B(n_169), .Y(n_215) );
AOI22xp5_ASAP7_75t_L g736 ( .A1(n_95), .A2(n_737), .B1(n_738), .B2(n_739), .Y(n_736) );
CKINVDCx20_ASAP7_75t_R g737 ( .A(n_95), .Y(n_737) );
INVx1_ASAP7_75t_L g218 ( .A(n_96), .Y(n_218) );
INVxp67_ASAP7_75t_L g206 ( .A(n_97), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_98), .B(n_136), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_99), .B(n_113), .Y(n_112) );
INVx1_ASAP7_75t_L g143 ( .A(n_100), .Y(n_143) );
INVx1_ASAP7_75t_L g244 ( .A(n_101), .Y(n_244) );
INVx2_ASAP7_75t_L g511 ( .A(n_102), .Y(n_511) );
AND2x2_ASAP7_75t_L g185 ( .A(n_103), .B(n_184), .Y(n_185) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
CKINVDCx12_ASAP7_75t_R g753 ( .A(n_107), .Y(n_753) );
AND2x2_ASAP7_75t_L g107 ( .A(n_108), .B(n_109), .Y(n_107) );
AND2x2_ASAP7_75t_L g447 ( .A(n_108), .B(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
INVx1_ASAP7_75t_SL g111 ( .A(n_112), .Y(n_111) );
OA21x2_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_120), .B(n_459), .Y(n_114) );
BUFx2_ASAP7_75t_SL g115 ( .A(n_116), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_117), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_SL g752 ( .A(n_118), .Y(n_752) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
OAI321xp33_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_443), .A3(n_449), .B1(n_452), .B2(n_453), .C(n_456), .Y(n_120) );
NAND2xp5_ASAP7_75t_SL g453 ( .A(n_121), .B(n_454), .Y(n_453) );
AOI22xp5_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_123), .B1(n_126), .B2(n_127), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
OAI22x1_ASAP7_75t_SL g461 ( .A1(n_126), .A2(n_462), .B1(n_465), .B2(n_731), .Y(n_461) );
INVx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
OAI22xp5_ASAP7_75t_SL g745 ( .A1(n_127), .A2(n_466), .B1(n_746), .B2(n_747), .Y(n_745) );
OR3x1_ASAP7_75t_L g127 ( .A(n_128), .B(n_341), .C(n_406), .Y(n_127) );
NAND4xp25_ASAP7_75t_SL g128 ( .A(n_129), .B(n_282), .C(n_308), .D(n_331), .Y(n_128) );
AOI221xp5_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_210), .B1(n_251), .B2(n_258), .C(n_274), .Y(n_129) );
CKINVDCx14_ASAP7_75t_R g130 ( .A(n_131), .Y(n_130) );
OAI22xp5_ASAP7_75t_L g429 ( .A1(n_131), .A2(n_275), .B1(n_299), .B2(n_430), .Y(n_429) );
OR2x2_ASAP7_75t_L g131 ( .A(n_132), .B(n_186), .Y(n_131) );
INVx1_ASAP7_75t_SL g335 ( .A(n_132), .Y(n_335) );
OR2x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_166), .Y(n_132) );
OR2x2_ASAP7_75t_L g256 ( .A(n_133), .B(n_257), .Y(n_256) );
AND2x2_ASAP7_75t_L g277 ( .A(n_133), .B(n_187), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_133), .B(n_197), .Y(n_290) );
AND2x2_ASAP7_75t_L g307 ( .A(n_133), .B(n_166), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_133), .B(n_254), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_133), .B(n_306), .Y(n_418) );
NOR2xp33_ASAP7_75t_L g428 ( .A(n_133), .B(n_186), .Y(n_428) );
AOI211xp5_ASAP7_75t_SL g439 ( .A1(n_133), .A2(n_345), .B(n_440), .C(n_441), .Y(n_439) );
INVx5_ASAP7_75t_SL g133 ( .A(n_134), .Y(n_133) );
NAND2xp5_ASAP7_75t_SL g311 ( .A(n_134), .B(n_187), .Y(n_311) );
AND2x2_ASAP7_75t_L g314 ( .A(n_134), .B(n_188), .Y(n_314) );
OR2x2_ASAP7_75t_L g359 ( .A(n_134), .B(n_187), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_134), .B(n_197), .Y(n_368) );
AO21x2_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_142), .B(n_163), .Y(n_134) );
INVx3_ASAP7_75t_L g209 ( .A(n_135), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g220 ( .A(n_135), .B(n_221), .Y(n_220) );
AO21x2_ASAP7_75t_L g240 ( .A1(n_135), .A2(n_241), .B(n_249), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g249 ( .A(n_135), .B(n_250), .Y(n_249) );
NOR2xp33_ASAP7_75t_L g481 ( .A(n_135), .B(n_482), .Y(n_481) );
NOR2xp33_ASAP7_75t_L g545 ( .A(n_135), .B(n_546), .Y(n_545) );
AO21x2_ASAP7_75t_L g549 ( .A1(n_135), .A2(n_550), .B(n_556), .Y(n_549) );
INVx4_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_136), .A2(n_190), .B(n_191), .Y(n_189) );
HB1xp67_ASAP7_75t_L g198 ( .A(n_136), .Y(n_198) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx1_ASAP7_75t_L g165 ( .A(n_137), .Y(n_165) );
AND2x2_ASAP7_75t_L g137 ( .A(n_138), .B(n_139), .Y(n_137) );
AND2x2_ASAP7_75t_SL g184 ( .A(n_138), .B(n_139), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_140), .B(n_141), .Y(n_139) );
OAI21xp5_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_144), .B(n_151), .Y(n_142) );
OAI21xp5_ASAP7_75t_L g474 ( .A1(n_144), .A2(n_475), .B(n_476), .Y(n_474) );
O2A1O1Ixp33_ASAP7_75t_L g539 ( .A1(n_144), .A2(n_184), .B(n_540), .C(n_541), .Y(n_539) );
OAI21xp5_ASAP7_75t_L g550 ( .A1(n_144), .A2(n_551), .B(n_552), .Y(n_550) );
NAND2x1p5_ASAP7_75t_L g144 ( .A(n_145), .B(n_149), .Y(n_144) );
AND2x4_ASAP7_75t_L g169 ( .A(n_145), .B(n_149), .Y(n_169) );
AND2x2_ASAP7_75t_L g145 ( .A(n_146), .B(n_148), .Y(n_145) );
INVx1_ASAP7_75t_L g207 ( .A(n_146), .Y(n_207) );
INVx1_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx2_ASAP7_75t_L g153 ( .A(n_147), .Y(n_153) );
INVx1_ASAP7_75t_L g162 ( .A(n_147), .Y(n_162) );
INVx1_ASAP7_75t_L g154 ( .A(n_148), .Y(n_154) );
INVx3_ASAP7_75t_L g157 ( .A(n_148), .Y(n_157) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_148), .Y(n_159) );
BUFx6f_ASAP7_75t_L g177 ( .A(n_148), .Y(n_177) );
INVx1_ASAP7_75t_L g194 ( .A(n_148), .Y(n_194) );
INVx4_ASAP7_75t_SL g183 ( .A(n_149), .Y(n_183) );
BUFx3_ASAP7_75t_L g196 ( .A(n_149), .Y(n_196) );
INVx5_ASAP7_75t_L g172 ( .A(n_152), .Y(n_172) );
AND2x6_ASAP7_75t_L g152 ( .A(n_153), .B(n_154), .Y(n_152) );
BUFx3_ASAP7_75t_L g181 ( .A(n_153), .Y(n_181) );
BUFx6f_ASAP7_75t_L g247 ( .A(n_153), .Y(n_247) );
AOI21xp5_ASAP7_75t_L g155 ( .A1(n_156), .A2(n_158), .B(n_160), .Y(n_155) );
INVx5_ASAP7_75t_L g179 ( .A(n_157), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_157), .B(n_493), .Y(n_492) );
INVx4_ASAP7_75t_L g271 ( .A(n_159), .Y(n_271) );
INVx2_ASAP7_75t_L g491 ( .A(n_159), .Y(n_491) );
AOI21xp5_ASAP7_75t_L g192 ( .A1(n_160), .A2(n_193), .B(n_195), .Y(n_192) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx3_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
NOR2xp33_ASAP7_75t_L g163 ( .A(n_164), .B(n_165), .Y(n_163) );
INVx2_ASAP7_75t_L g528 ( .A(n_165), .Y(n_528) );
INVx5_ASAP7_75t_SL g257 ( .A(n_166), .Y(n_257) );
AND2x2_ASAP7_75t_L g276 ( .A(n_166), .B(n_277), .Y(n_276) );
NOR2xp33_ASAP7_75t_L g358 ( .A(n_166), .B(n_359), .Y(n_358) );
AND2x2_ASAP7_75t_L g362 ( .A(n_166), .B(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_L g394 ( .A(n_166), .B(n_197), .Y(n_394) );
OR2x2_ASAP7_75t_L g400 ( .A(n_166), .B(n_290), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_166), .B(n_350), .Y(n_409) );
OR2x6_ASAP7_75t_L g166 ( .A(n_167), .B(n_185), .Y(n_166) );
AOI21xp5_ASAP7_75t_L g167 ( .A1(n_168), .A2(n_170), .B(n_184), .Y(n_167) );
BUFx2_ASAP7_75t_L g227 ( .A(n_169), .Y(n_227) );
INVx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
O2A1O1Ixp33_ASAP7_75t_L g200 ( .A1(n_172), .A2(n_183), .B(n_201), .C(n_202), .Y(n_200) );
O2A1O1Ixp33_ASAP7_75t_SL g265 ( .A1(n_172), .A2(n_183), .B(n_266), .C(n_267), .Y(n_265) );
O2A1O1Ixp33_ASAP7_75t_SL g488 ( .A1(n_172), .A2(n_183), .B(n_489), .C(n_490), .Y(n_488) );
O2A1O1Ixp33_ASAP7_75t_SL g498 ( .A1(n_172), .A2(n_183), .B(n_499), .C(n_500), .Y(n_498) );
O2A1O1Ixp33_ASAP7_75t_SL g507 ( .A1(n_172), .A2(n_183), .B(n_508), .C(n_509), .Y(n_507) );
O2A1O1Ixp33_ASAP7_75t_L g517 ( .A1(n_172), .A2(n_183), .B(n_518), .C(n_519), .Y(n_517) );
O2A1O1Ixp33_ASAP7_75t_SL g530 ( .A1(n_172), .A2(n_183), .B(n_531), .C(n_532), .Y(n_530) );
O2A1O1Ixp33_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_175), .B(n_178), .C(n_180), .Y(n_173) );
O2A1O1Ixp33_ASAP7_75t_L g217 ( .A1(n_175), .A2(n_180), .B(n_218), .C(n_219), .Y(n_217) );
O2A1O1Ixp5_ASAP7_75t_L g477 ( .A1(n_175), .A2(n_478), .B(n_479), .C(n_480), .Y(n_477) );
O2A1O1Ixp33_ASAP7_75t_L g553 ( .A1(n_175), .A2(n_480), .B(n_554), .C(n_555), .Y(n_553) );
INVx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx4_ASAP7_75t_L g204 ( .A(n_177), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g205 ( .A(n_179), .B(n_206), .Y(n_205) );
INVx2_ASAP7_75t_L g268 ( .A(n_179), .Y(n_268) );
OAI22xp33_ASAP7_75t_L g533 ( .A1(n_179), .A2(n_204), .B1(n_534), .B2(n_535), .Y(n_533) );
O2A1O1Ixp33_ASAP7_75t_L g542 ( .A1(n_179), .A2(n_232), .B(n_543), .C(n_544), .Y(n_542) );
HB1xp67_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx2_ASAP7_75t_L g272 ( .A(n_181), .Y(n_272) );
INVx1_ASAP7_75t_L g503 ( .A(n_181), .Y(n_503) );
INVx1_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_184), .A2(n_215), .B(n_216), .Y(n_214) );
INVx2_ASAP7_75t_L g234 ( .A(n_184), .Y(n_234) );
INVx1_ASAP7_75t_L g237 ( .A(n_184), .Y(n_237) );
OA21x2_ASAP7_75t_L g486 ( .A1(n_184), .A2(n_487), .B(n_494), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_187), .B(n_197), .Y(n_186) );
AND2x2_ASAP7_75t_L g291 ( .A(n_187), .B(n_257), .Y(n_291) );
INVx1_ASAP7_75t_SL g304 ( .A(n_187), .Y(n_304) );
OR2x2_ASAP7_75t_L g339 ( .A(n_187), .B(n_340), .Y(n_339) );
OR2x2_ASAP7_75t_L g345 ( .A(n_187), .B(n_197), .Y(n_345) );
AND2x2_ASAP7_75t_L g403 ( .A(n_187), .B(n_254), .Y(n_403) );
INVx2_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_188), .B(n_257), .Y(n_330) );
INVx3_ASAP7_75t_L g254 ( .A(n_197), .Y(n_254) );
OR2x2_ASAP7_75t_L g296 ( .A(n_197), .B(n_257), .Y(n_296) );
AND2x2_ASAP7_75t_L g306 ( .A(n_197), .B(n_304), .Y(n_306) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_197), .Y(n_354) );
AND2x2_ASAP7_75t_L g363 ( .A(n_197), .B(n_277), .Y(n_363) );
OA21x2_ASAP7_75t_L g197 ( .A1(n_198), .A2(n_199), .B(n_208), .Y(n_197) );
OA21x2_ASAP7_75t_L g496 ( .A1(n_198), .A2(n_497), .B(n_504), .Y(n_496) );
OA21x2_ASAP7_75t_L g505 ( .A1(n_198), .A2(n_506), .B(n_512), .Y(n_505) );
OA21x2_ASAP7_75t_L g515 ( .A1(n_198), .A2(n_516), .B(n_523), .Y(n_515) );
O2A1O1Ixp33_ASAP7_75t_L g243 ( .A1(n_203), .A2(n_244), .B(n_245), .C(n_246), .Y(n_243) );
INVx1_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_204), .B(n_502), .Y(n_501) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_204), .B(n_511), .Y(n_510) );
INVx2_ASAP7_75t_L g232 ( .A(n_207), .Y(n_232) );
NAND2xp5_ASAP7_75t_SL g532 ( .A(n_207), .B(n_533), .Y(n_532) );
OA21x2_ASAP7_75t_L g263 ( .A1(n_209), .A2(n_264), .B(n_273), .Y(n_263) );
AOI221xp5_ASAP7_75t_L g379 ( .A1(n_210), .A2(n_380), .B1(n_382), .B2(n_384), .C(n_387), .Y(n_379) );
INVx2_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
OR2x2_ASAP7_75t_L g211 ( .A(n_212), .B(n_222), .Y(n_211) );
AND2x2_ASAP7_75t_L g353 ( .A(n_212), .B(n_334), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_212), .B(n_412), .Y(n_416) );
OR2x2_ASAP7_75t_L g437 ( .A(n_212), .B(n_438), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_212), .B(n_442), .Y(n_441) );
BUFx2_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
INVx5_ASAP7_75t_L g284 ( .A(n_213), .Y(n_284) );
AND2x2_ASAP7_75t_L g361 ( .A(n_213), .B(n_224), .Y(n_361) );
AND2x2_ASAP7_75t_L g422 ( .A(n_213), .B(n_301), .Y(n_422) );
AND2x2_ASAP7_75t_L g435 ( .A(n_213), .B(n_254), .Y(n_435) );
OR2x6_ASAP7_75t_L g213 ( .A(n_214), .B(n_220), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_223), .B(n_238), .Y(n_222) );
AND2x4_ASAP7_75t_L g261 ( .A(n_223), .B(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g280 ( .A(n_223), .B(n_281), .Y(n_280) );
INVx2_ASAP7_75t_L g287 ( .A(n_223), .Y(n_287) );
AND2x2_ASAP7_75t_L g356 ( .A(n_223), .B(n_334), .Y(n_356) );
AND2x2_ASAP7_75t_L g366 ( .A(n_223), .B(n_284), .Y(n_366) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_223), .Y(n_374) );
AND2x2_ASAP7_75t_L g386 ( .A(n_223), .B(n_263), .Y(n_386) );
NOR2xp33_ASAP7_75t_L g390 ( .A(n_223), .B(n_318), .Y(n_390) );
AND2x2_ASAP7_75t_L g427 ( .A(n_223), .B(n_422), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_223), .B(n_301), .Y(n_438) );
OR2x2_ASAP7_75t_L g440 ( .A(n_223), .B(n_376), .Y(n_440) );
INVx5_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
AND2x2_ASAP7_75t_L g326 ( .A(n_224), .B(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g336 ( .A(n_224), .B(n_281), .Y(n_336) );
AND2x2_ASAP7_75t_L g348 ( .A(n_224), .B(n_263), .Y(n_348) );
HB1xp67_ASAP7_75t_L g378 ( .A(n_224), .Y(n_378) );
AND2x4_ASAP7_75t_L g412 ( .A(n_224), .B(n_262), .Y(n_412) );
OR2x6_ASAP7_75t_L g224 ( .A(n_225), .B(n_235), .Y(n_224) );
AOI21xp5_ASAP7_75t_SL g225 ( .A1(n_226), .A2(n_228), .B(n_233), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_230), .A2(n_231), .B(n_232), .Y(n_229) );
INVx1_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
NOR2xp33_ASAP7_75t_L g556 ( .A(n_234), .B(n_451), .Y(n_556) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_236), .B(n_237), .Y(n_235) );
AO21x2_ASAP7_75t_L g473 ( .A1(n_237), .A2(n_474), .B(n_481), .Y(n_473) );
BUFx2_ASAP7_75t_L g260 ( .A(n_238), .Y(n_260) );
HB1xp67_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
INVx2_ASAP7_75t_L g301 ( .A(n_239), .Y(n_301) );
AND2x2_ASAP7_75t_L g334 ( .A(n_239), .B(n_263), .Y(n_334) );
INVx2_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
AND2x2_ASAP7_75t_L g281 ( .A(n_240), .B(n_263), .Y(n_281) );
BUFx2_ASAP7_75t_L g327 ( .A(n_240), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_242), .B(n_248), .Y(n_241) );
HB1xp67_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
INVx3_ASAP7_75t_L g522 ( .A(n_247), .Y(n_522) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_253), .B(n_255), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_253), .B(n_335), .Y(n_414) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_254), .B(n_277), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_254), .B(n_257), .Y(n_316) );
AND2x2_ASAP7_75t_L g371 ( .A(n_254), .B(n_307), .Y(n_371) );
AOI221xp5_ASAP7_75t_SL g308 ( .A1(n_255), .A2(n_309), .B1(n_317), .B2(n_319), .C(n_323), .Y(n_308) );
INVx2_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
OR2x2_ASAP7_75t_L g303 ( .A(n_256), .B(n_304), .Y(n_303) );
OR2x2_ASAP7_75t_L g344 ( .A(n_256), .B(n_345), .Y(n_344) );
OAI321xp33_ASAP7_75t_L g351 ( .A1(n_256), .A2(n_310), .A3(n_352), .B1(n_354), .B2(n_355), .C(n_357), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_257), .B(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_260), .B(n_261), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_260), .B(n_412), .Y(n_430) );
AND2x2_ASAP7_75t_L g317 ( .A(n_261), .B(n_318), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_261), .B(n_321), .Y(n_320) );
HB1xp67_ASAP7_75t_L g293 ( .A(n_262), .Y(n_293) );
AND2x2_ASAP7_75t_L g300 ( .A(n_262), .B(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_262), .B(n_375), .Y(n_405) );
INVx1_ASAP7_75t_L g442 ( .A(n_262), .Y(n_442) );
INVx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
NOR2xp33_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_271), .B(n_521), .Y(n_520) );
INVx2_ASAP7_75t_L g480 ( .A(n_272), .Y(n_480) );
AOI21xp5_ASAP7_75t_L g274 ( .A1(n_275), .A2(n_278), .B(n_279), .Y(n_274) );
INVx1_ASAP7_75t_SL g275 ( .A(n_276), .Y(n_275) );
A2O1A1Ixp33_ASAP7_75t_L g434 ( .A1(n_276), .A2(n_386), .B(n_435), .C(n_436), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_277), .B(n_295), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_277), .B(n_315), .Y(n_381) );
INVx1_ASAP7_75t_SL g279 ( .A(n_280), .Y(n_279) );
INVx1_ASAP7_75t_L g324 ( .A(n_281), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_281), .B(n_284), .Y(n_338) );
NOR2xp33_ASAP7_75t_L g347 ( .A(n_281), .B(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_281), .B(n_366), .Y(n_365) );
AOI22xp33_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_285), .B1(n_297), .B2(n_302), .Y(n_282) );
HB1xp67_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
OR2x2_ASAP7_75t_L g298 ( .A(n_284), .B(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g321 ( .A(n_284), .B(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g333 ( .A(n_284), .B(n_334), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_284), .B(n_327), .Y(n_369) );
OR2x2_ASAP7_75t_L g376 ( .A(n_284), .B(n_301), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_284), .B(n_386), .Y(n_385) );
AND2x2_ASAP7_75t_L g426 ( .A(n_284), .B(n_412), .Y(n_426) );
OAI22xp33_ASAP7_75t_L g285 ( .A1(n_286), .A2(n_288), .B1(n_292), .B2(n_294), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g332 ( .A(n_287), .B(n_333), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_289), .B(n_291), .Y(n_288) );
INVx1_ASAP7_75t_SL g289 ( .A(n_290), .Y(n_289) );
OAI22xp33_ASAP7_75t_L g372 ( .A1(n_290), .A2(n_305), .B1(n_373), .B2(n_377), .Y(n_372) );
INVx1_ASAP7_75t_L g420 ( .A(n_291), .Y(n_420) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AOI221xp5_ASAP7_75t_L g331 ( .A1(n_295), .A2(n_332), .B1(n_335), .B2(n_336), .C(n_337), .Y(n_331) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
OR2x2_ASAP7_75t_L g310 ( .A(n_296), .B(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_300), .B(n_366), .Y(n_398) );
HB1xp67_ASAP7_75t_L g318 ( .A(n_301), .Y(n_318) );
INVx1_ASAP7_75t_L g322 ( .A(n_301), .Y(n_322) );
NAND2xp33_ASAP7_75t_L g302 ( .A(n_303), .B(n_305), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_306), .B(n_307), .Y(n_305) );
INVx1_ASAP7_75t_L g340 ( .A(n_307), .Y(n_340) );
AND2x2_ASAP7_75t_L g349 ( .A(n_307), .B(n_350), .Y(n_349) );
NAND2xp33_ASAP7_75t_L g309 ( .A(n_310), .B(n_312), .Y(n_309) );
INVx2_ASAP7_75t_SL g312 ( .A(n_313), .Y(n_312) );
AND2x4_ASAP7_75t_L g313 ( .A(n_314), .B(n_315), .Y(n_313) );
AND2x2_ASAP7_75t_L g393 ( .A(n_314), .B(n_394), .Y(n_393) );
INVx2_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
AOI221xp5_ASAP7_75t_L g342 ( .A1(n_317), .A2(n_343), .B1(n_346), .B2(n_349), .C(n_351), .Y(n_342) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_321), .B(n_378), .Y(n_377) );
AOI21xp33_ASAP7_75t_SL g323 ( .A1(n_324), .A2(n_325), .B(n_328), .Y(n_323) );
INVx2_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
CKINVDCx16_ASAP7_75t_R g425 ( .A(n_328), .Y(n_425) );
OR2x2_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
OR2x2_ASAP7_75t_L g367 ( .A(n_330), .B(n_368), .Y(n_367) );
INVx1_ASAP7_75t_SL g388 ( .A(n_333), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_333), .B(n_393), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_336), .B(n_358), .Y(n_357) );
NOR2xp33_ASAP7_75t_L g337 ( .A(n_338), .B(n_339), .Y(n_337) );
NAND4xp25_ASAP7_75t_L g341 ( .A(n_342), .B(n_360), .C(n_379), .D(n_392), .Y(n_341) );
INVx1_ASAP7_75t_SL g343 ( .A(n_344), .Y(n_343) );
INVx1_ASAP7_75t_SL g350 ( .A(n_345), .Y(n_350) );
INVxp67_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
OR2x2_ASAP7_75t_L g383 ( .A(n_354), .B(n_359), .Y(n_383) );
INVxp67_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
AOI211xp5_ASAP7_75t_L g360 ( .A1(n_361), .A2(n_362), .B(n_364), .C(n_372), .Y(n_360) );
AOI211xp5_ASAP7_75t_L g431 ( .A1(n_362), .A2(n_404), .B(n_432), .C(n_439), .Y(n_431) );
INVx1_ASAP7_75t_SL g391 ( .A(n_363), .Y(n_391) );
OAI22xp5_ASAP7_75t_L g364 ( .A1(n_365), .A2(n_367), .B1(n_369), .B2(n_370), .Y(n_364) );
INVx1_ASAP7_75t_L g395 ( .A(n_369), .Y(n_395) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_374), .B(n_375), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_375), .B(n_412), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_375), .B(n_386), .Y(n_419) );
INVx2_ASAP7_75t_SL g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_SL g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g396 ( .A(n_386), .Y(n_396) );
AOI21xp33_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_389), .B(n_391), .Y(n_387) );
INVxp33_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
AOI322xp5_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_395), .A3(n_396), .B1(n_397), .B2(n_399), .C1(n_401), .C2(n_404), .Y(n_392) );
INVxp67_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
NAND3xp33_ASAP7_75t_SL g406 ( .A(n_407), .B(n_424), .C(n_431), .Y(n_406) );
AOI221xp5_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_410), .B1(n_413), .B2(n_415), .C(n_417), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_SL g423 ( .A(n_412), .Y(n_423) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVxp67_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
OAI22xp33_ASAP7_75t_L g417 ( .A1(n_418), .A2(n_419), .B1(n_420), .B2(n_421), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_422), .B(n_423), .Y(n_421) );
AOI221xp5_ASAP7_75t_L g424 ( .A1(n_425), .A2(n_426), .B1(n_427), .B2(n_428), .C(n_429), .Y(n_424) );
NAND2xp33_ASAP7_75t_L g432 ( .A(n_433), .B(n_434), .Y(n_432) );
INVxp67_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
HB1xp67_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_SL g455 ( .A(n_445), .Y(n_455) );
HB1xp67_ASAP7_75t_L g458 ( .A(n_445), .Y(n_458) );
NOR2x2_ASAP7_75t_L g750 ( .A(n_446), .B(n_734), .Y(n_750) );
INVx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
OR2x2_ASAP7_75t_L g733 ( .A(n_447), .B(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g452 ( .A(n_449), .Y(n_452) );
INVx1_ASAP7_75t_SL g454 ( .A(n_455), .Y(n_454) );
NAND3xp33_ASAP7_75t_L g459 ( .A(n_456), .B(n_460), .C(n_751), .Y(n_459) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx2_ASAP7_75t_L g746 ( .A(n_463), .Y(n_746) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
OR2x2_ASAP7_75t_SL g466 ( .A(n_467), .B(n_686), .Y(n_466) );
NAND5xp2_ASAP7_75t_L g467 ( .A(n_468), .B(n_598), .C(n_636), .D(n_657), .E(n_674), .Y(n_467) );
NOR3xp33_ASAP7_75t_L g468 ( .A(n_469), .B(n_570), .C(n_591), .Y(n_468) );
OAI221xp5_ASAP7_75t_SL g469 ( .A1(n_470), .A2(n_513), .B1(n_537), .B2(n_557), .C(n_561), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_471), .B(n_483), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_472), .B(n_559), .Y(n_578) );
OR2x2_ASAP7_75t_L g605 ( .A(n_472), .B(n_496), .Y(n_605) );
AND2x2_ASAP7_75t_L g619 ( .A(n_472), .B(n_496), .Y(n_619) );
NOR2xp33_ASAP7_75t_L g633 ( .A(n_472), .B(n_486), .Y(n_633) );
AND2x2_ASAP7_75t_L g671 ( .A(n_472), .B(n_635), .Y(n_671) );
AND2x2_ASAP7_75t_L g700 ( .A(n_472), .B(n_610), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_472), .B(n_582), .Y(n_717) );
INVx4_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
AND2x2_ASAP7_75t_L g597 ( .A(n_473), .B(n_495), .Y(n_597) );
BUFx3_ASAP7_75t_L g622 ( .A(n_473), .Y(n_622) );
AND2x2_ASAP7_75t_L g651 ( .A(n_473), .B(n_496), .Y(n_651) );
AND3x2_ASAP7_75t_L g664 ( .A(n_473), .B(n_665), .C(n_666), .Y(n_664) );
INVx1_ASAP7_75t_L g587 ( .A(n_483), .Y(n_587) );
AND2x2_ASAP7_75t_L g483 ( .A(n_484), .B(n_495), .Y(n_483) );
AOI32xp33_ASAP7_75t_L g642 ( .A1(n_484), .A2(n_594), .A3(n_643), .B1(n_646), .B2(n_647), .Y(n_642) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
AND2x2_ASAP7_75t_L g569 ( .A(n_485), .B(n_495), .Y(n_569) );
NAND2xp5_ASAP7_75t_SL g640 ( .A(n_485), .B(n_597), .Y(n_640) );
AND2x2_ASAP7_75t_L g647 ( .A(n_485), .B(n_619), .Y(n_647) );
OR2x2_ASAP7_75t_L g653 ( .A(n_485), .B(n_654), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_485), .B(n_608), .Y(n_678) );
OR2x2_ASAP7_75t_L g696 ( .A(n_485), .B(n_525), .Y(n_696) );
BUFx3_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
AND2x2_ASAP7_75t_L g560 ( .A(n_486), .B(n_505), .Y(n_560) );
INVx2_ASAP7_75t_L g582 ( .A(n_486), .Y(n_582) );
OR2x2_ASAP7_75t_L g604 ( .A(n_486), .B(n_505), .Y(n_604) );
AND2x2_ASAP7_75t_L g609 ( .A(n_486), .B(n_610), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_486), .B(n_661), .Y(n_660) );
AND2x2_ASAP7_75t_L g665 ( .A(n_486), .B(n_559), .Y(n_665) );
INVx1_ASAP7_75t_SL g716 ( .A(n_495), .Y(n_716) );
AND2x2_ASAP7_75t_L g495 ( .A(n_496), .B(n_505), .Y(n_495) );
INVx1_ASAP7_75t_SL g559 ( .A(n_496), .Y(n_559) );
HB1xp67_ASAP7_75t_L g608 ( .A(n_496), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_496), .B(n_645), .Y(n_644) );
NAND3xp33_ASAP7_75t_L g711 ( .A(n_496), .B(n_582), .C(n_700), .Y(n_711) );
INVx2_ASAP7_75t_L g610 ( .A(n_505), .Y(n_610) );
HB1xp67_ASAP7_75t_L g624 ( .A(n_505), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_514), .B(n_524), .Y(n_513) );
INVx1_ASAP7_75t_L g646 ( .A(n_514), .Y(n_646) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
AND2x2_ASAP7_75t_L g564 ( .A(n_515), .B(n_548), .Y(n_564) );
INVx2_ASAP7_75t_L g581 ( .A(n_515), .Y(n_581) );
AND2x2_ASAP7_75t_L g586 ( .A(n_515), .B(n_549), .Y(n_586) );
AND2x2_ASAP7_75t_L g601 ( .A(n_515), .B(n_538), .Y(n_601) );
AND2x2_ASAP7_75t_L g613 ( .A(n_515), .B(n_585), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_524), .B(n_629), .Y(n_628) );
NAND2x1p5_ASAP7_75t_L g685 ( .A(n_524), .B(n_586), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_524), .B(n_705), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_524), .B(n_580), .Y(n_708) );
BUFx3_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
OR2x2_ASAP7_75t_L g547 ( .A(n_525), .B(n_548), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_525), .B(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g590 ( .A(n_525), .B(n_538), .Y(n_590) );
AND2x2_ASAP7_75t_L g616 ( .A(n_525), .B(n_548), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_525), .B(n_656), .Y(n_655) );
OA21x2_ASAP7_75t_L g525 ( .A1(n_526), .A2(n_529), .B(n_536), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
AO21x2_ASAP7_75t_L g574 ( .A1(n_527), .A2(n_575), .B(n_576), .Y(n_574) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g575 ( .A(n_529), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_536), .Y(n_576) );
OR2x2_ASAP7_75t_L g537 ( .A(n_538), .B(n_547), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_538), .B(n_567), .Y(n_566) );
AND2x4_ASAP7_75t_L g580 ( .A(n_538), .B(n_581), .Y(n_580) );
INVx3_ASAP7_75t_SL g585 ( .A(n_538), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_538), .B(n_572), .Y(n_638) );
OR2x2_ASAP7_75t_L g648 ( .A(n_538), .B(n_574), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_538), .B(n_616), .Y(n_676) );
OR2x2_ASAP7_75t_L g706 ( .A(n_538), .B(n_548), .Y(n_706) );
AND2x2_ASAP7_75t_L g710 ( .A(n_538), .B(n_549), .Y(n_710) );
NAND2xp5_ASAP7_75t_SL g723 ( .A(n_538), .B(n_586), .Y(n_723) );
AND2x2_ASAP7_75t_L g730 ( .A(n_538), .B(n_612), .Y(n_730) );
OR2x6_ASAP7_75t_L g538 ( .A(n_539), .B(n_545), .Y(n_538) );
INVx1_ASAP7_75t_SL g673 ( .A(n_547), .Y(n_673) );
AND2x2_ASAP7_75t_L g612 ( .A(n_548), .B(n_574), .Y(n_612) );
AND2x2_ASAP7_75t_L g626 ( .A(n_548), .B(n_581), .Y(n_626) );
AND2x2_ASAP7_75t_L g629 ( .A(n_548), .B(n_585), .Y(n_629) );
INVx1_ASAP7_75t_L g656 ( .A(n_548), .Y(n_656) );
INVx2_ASAP7_75t_SL g548 ( .A(n_549), .Y(n_548) );
BUFx2_ASAP7_75t_L g568 ( .A(n_549), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_558), .B(n_560), .Y(n_557) );
A2O1A1Ixp33_ASAP7_75t_L g727 ( .A1(n_558), .A2(n_604), .B(n_728), .C(n_729), .Y(n_727) );
HB1xp67_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g634 ( .A(n_559), .B(n_635), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_560), .B(n_577), .Y(n_592) );
AND2x2_ASAP7_75t_L g618 ( .A(n_560), .B(n_619), .Y(n_618) );
OAI21xp5_ASAP7_75t_SL g561 ( .A1(n_562), .A2(n_565), .B(n_569), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
NOR2xp33_ASAP7_75t_L g662 ( .A(n_563), .B(n_663), .Y(n_662) );
AND2x2_ASAP7_75t_L g589 ( .A(n_564), .B(n_590), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_564), .B(n_585), .Y(n_630) );
AND2x2_ASAP7_75t_L g721 ( .A(n_564), .B(n_572), .Y(n_721) );
INVxp67_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g594 ( .A(n_568), .B(n_581), .Y(n_594) );
OR2x2_ASAP7_75t_L g595 ( .A(n_568), .B(n_579), .Y(n_595) );
OAI322xp33_ASAP7_75t_L g570 ( .A1(n_571), .A2(n_578), .A3(n_579), .B1(n_582), .B2(n_583), .C1(n_587), .C2(n_588), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_572), .B(n_577), .Y(n_571) );
AND2x2_ASAP7_75t_L g682 ( .A(n_572), .B(n_594), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_572), .B(n_646), .Y(n_728) );
INVx2_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx1_ASAP7_75t_SL g573 ( .A(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g625 ( .A(n_574), .B(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
OR2x2_ASAP7_75t_L g691 ( .A(n_578), .B(n_604), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_579), .B(n_673), .Y(n_672) );
INVx3_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_580), .B(n_612), .Y(n_669) );
AND2x2_ASAP7_75t_L g615 ( .A(n_581), .B(n_585), .Y(n_615) );
AND2x2_ASAP7_75t_L g623 ( .A(n_582), .B(n_624), .Y(n_623) );
A2O1A1Ixp33_ASAP7_75t_L g720 ( .A1(n_582), .A2(n_661), .B(n_721), .C(n_722), .Y(n_720) );
AOI21xp33_ASAP7_75t_L g693 ( .A1(n_583), .A2(n_596), .B(n_694), .Y(n_693) );
INVx1_ASAP7_75t_SL g583 ( .A(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_585), .B(n_586), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_585), .B(n_612), .Y(n_652) );
AND2x2_ASAP7_75t_L g658 ( .A(n_585), .B(n_626), .Y(n_658) );
AND2x2_ASAP7_75t_L g692 ( .A(n_585), .B(n_594), .Y(n_692) );
NOR2xp33_ASAP7_75t_L g600 ( .A(n_586), .B(n_601), .Y(n_600) );
INVx2_ASAP7_75t_SL g702 ( .A(n_586), .Y(n_702) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
AOI22xp5_ASAP7_75t_L g617 ( .A1(n_590), .A2(n_618), .B1(n_620), .B2(n_625), .Y(n_617) );
OAI22xp5_ASAP7_75t_SL g591 ( .A1(n_592), .A2(n_593), .B1(n_595), .B2(n_596), .Y(n_591) );
OAI22xp33_ASAP7_75t_L g627 ( .A1(n_592), .A2(n_628), .B1(n_630), .B2(n_631), .Y(n_627) );
INVxp67_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx1_ASAP7_75t_SL g596 ( .A(n_597), .Y(n_596) );
AOI221xp5_ASAP7_75t_L g698 ( .A1(n_597), .A2(n_699), .B1(n_701), .B2(n_703), .C(n_707), .Y(n_698) );
AOI211xp5_ASAP7_75t_L g598 ( .A1(n_599), .A2(n_602), .B(n_606), .C(n_627), .Y(n_598) );
INVxp67_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
OR2x2_ASAP7_75t_L g603 ( .A(n_604), .B(n_605), .Y(n_603) );
OR2x2_ASAP7_75t_L g668 ( .A(n_604), .B(n_621), .Y(n_668) );
INVx1_ASAP7_75t_L g719 ( .A(n_604), .Y(n_719) );
OAI221xp5_ASAP7_75t_L g606 ( .A1(n_605), .A2(n_607), .B1(n_611), .B2(n_614), .C(n_617), .Y(n_606) );
INVx2_ASAP7_75t_SL g661 ( .A(n_605), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_608), .B(n_609), .Y(n_607) );
INVx1_ASAP7_75t_L g726 ( .A(n_608), .Y(n_726) );
AND2x2_ASAP7_75t_L g650 ( .A(n_609), .B(n_651), .Y(n_650) );
INVx2_ASAP7_75t_L g635 ( .A(n_610), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_612), .B(n_613), .Y(n_611) );
INVx1_ASAP7_75t_L g697 ( .A(n_613), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
AND2x2_ASAP7_75t_L g620 ( .A(n_621), .B(n_623), .Y(n_620) );
NOR2xp33_ASAP7_75t_L g722 ( .A(n_621), .B(n_723), .Y(n_722) );
CKINVDCx16_ASAP7_75t_R g621 ( .A(n_622), .Y(n_621) );
INVxp67_ASAP7_75t_L g666 ( .A(n_624), .Y(n_666) );
O2A1O1Ixp33_ASAP7_75t_L g636 ( .A1(n_625), .A2(n_637), .B(n_639), .C(n_641), .Y(n_636) );
INVx1_ASAP7_75t_L g714 ( .A(n_628), .Y(n_714) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
NOR2xp33_ASAP7_75t_L g689 ( .A(n_632), .B(n_690), .Y(n_689) );
AND2x2_ASAP7_75t_L g632 ( .A(n_633), .B(n_634), .Y(n_632) );
INVx2_ASAP7_75t_L g645 ( .A(n_635), .Y(n_645) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
OAI222xp33_ASAP7_75t_L g641 ( .A1(n_642), .A2(n_648), .B1(n_649), .B2(n_652), .C1(n_653), .C2(n_655), .Y(n_641) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_SL g681 ( .A(n_645), .Y(n_681) );
NOR2xp33_ASAP7_75t_L g701 ( .A(n_648), .B(n_702), .Y(n_701) );
NAND2xp33_ASAP7_75t_SL g679 ( .A(n_649), .B(n_680), .Y(n_679) );
INVx1_ASAP7_75t_SL g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_SL g654 ( .A(n_651), .Y(n_654) );
AND2x2_ASAP7_75t_L g718 ( .A(n_651), .B(n_719), .Y(n_718) );
OR2x2_ASAP7_75t_L g684 ( .A(n_654), .B(n_681), .Y(n_684) );
INVx1_ASAP7_75t_L g713 ( .A(n_655), .Y(n_713) );
AOI211xp5_ASAP7_75t_L g657 ( .A1(n_658), .A2(n_659), .B(n_662), .C(n_667), .Y(n_657) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_661), .B(n_681), .Y(n_680) );
INVx2_ASAP7_75t_SL g663 ( .A(n_664), .Y(n_663) );
AOI322xp5_ASAP7_75t_L g712 ( .A1(n_664), .A2(n_692), .A3(n_697), .B1(n_713), .B2(n_714), .C1(n_715), .C2(n_718), .Y(n_712) );
AND2x2_ASAP7_75t_L g699 ( .A(n_665), .B(n_700), .Y(n_699) );
OAI22xp33_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_669), .B1(n_670), .B2(n_672), .Y(n_667) );
INVxp33_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
AOI221xp5_ASAP7_75t_L g674 ( .A1(n_675), .A2(n_677), .B1(n_679), .B2(n_682), .C(n_683), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
NOR2xp33_ASAP7_75t_L g683 ( .A(n_684), .B(n_685), .Y(n_683) );
NAND5xp2_ASAP7_75t_L g686 ( .A(n_687), .B(n_698), .C(n_712), .D(n_720), .E(n_724), .Y(n_686) );
AOI21xp5_ASAP7_75t_L g687 ( .A1(n_688), .A2(n_692), .B(n_693), .Y(n_687) );
INVxp67_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx2_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVxp33_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
NOR2xp33_ASAP7_75t_L g695 ( .A(n_696), .B(n_697), .Y(n_695) );
A2O1A1Ixp33_ASAP7_75t_L g724 ( .A1(n_700), .A2(n_725), .B(n_726), .C(n_727), .Y(n_724) );
AOI31xp33_ASAP7_75t_L g707 ( .A1(n_702), .A2(n_708), .A3(n_709), .B(n_711), .Y(n_707) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
NOR2xp33_ASAP7_75t_L g715 ( .A(n_716), .B(n_717), .Y(n_715) );
INVx1_ASAP7_75t_L g725 ( .A(n_723), .Y(n_725) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx2_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx2_ASAP7_75t_L g747 ( .A(n_732), .Y(n_747) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
CKINVDCx20_ASAP7_75t_R g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g743 ( .A(n_740), .Y(n_743) );
INVx1_ASAP7_75t_SL g748 ( .A(n_749), .Y(n_748) );
INVx3_ASAP7_75t_SL g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_SL g751 ( .A(n_752), .Y(n_751) );
endmodule