module real_jpeg_25497_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_113;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_44;
wire n_28;
wire n_62;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

INVx6_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_0),
.B(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_0),
.Y(n_96)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_4),
.A2(n_18),
.B1(n_19),
.B2(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_4),
.A2(n_23),
.B1(n_24),
.B2(n_32),
.Y(n_46)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_4),
.A2(n_32),
.B1(n_51),
.B2(n_62),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g17 ( 
.A1(n_5),
.A2(n_18),
.B1(n_19),
.B2(n_21),
.Y(n_17)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_5),
.A2(n_21),
.B1(n_23),
.B2(n_24),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_6),
.A2(n_23),
.B1(n_24),
.B2(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_6),
.A2(n_18),
.B1(n_19),
.B2(n_43),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_8),
.A2(n_23),
.B1(n_24),
.B2(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_8),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_10),
.B(n_35),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_10),
.B(n_19),
.C(n_37),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_10),
.A2(n_51),
.B1(n_62),
.B2(n_63),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_10),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_10),
.A2(n_18),
.B1(n_19),
.B2(n_63),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_10),
.B(n_23),
.C(n_27),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_10),
.A2(n_40),
.B(n_44),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_75),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_74),
.Y(n_12)
);

INVxp67_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_47),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_15),
.B(n_47),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_33),
.C(n_39),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_16),
.A2(n_33),
.B1(n_34),
.B2(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_16),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_22),
.B(n_28),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_17),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_L g30 ( 
.A1(n_18),
.A2(n_19),
.B1(n_26),
.B2(n_27),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_18),
.A2(n_19),
.B1(n_37),
.B2(n_38),
.Y(n_36)
);

INVx5_ASAP7_75t_SL g18 ( 
.A(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_19),
.B(n_87),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_22),
.B(n_30),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_22),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_22),
.B(n_63),
.Y(n_102)
);

OA22x2_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_26),
.B2(n_27),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_23),
.B(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_SL g23 ( 
.A(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_24),
.B(n_107),
.Y(n_106)
);

INVx6_ASAP7_75t_SL g24 ( 
.A(n_25),
.Y(n_24)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_31),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_29),
.A2(n_69),
.B1(n_70),
.B2(n_71),
.Y(n_68)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_29),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_31),
.B(n_71),
.Y(n_85)
);

CKINVDCx14_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_35),
.B(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_36),
.B(n_65),
.Y(n_64)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_37),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_37),
.A2(n_38),
.B1(n_51),
.B2(n_62),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_39),
.B(n_78),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_42),
.B(n_44),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_46),
.Y(n_58)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_40),
.Y(n_91)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_41),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_42),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_59),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_SL g48 ( 
.A(n_49),
.B(n_53),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_50),
.B(n_51),
.Y(n_49)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_57),
.B(n_58),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_58),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_68),
.B1(n_72),
.B2(n_73),
.Y(n_59)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

OAI21xp33_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_64),
.B(n_66),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_63),
.B(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_68),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_76),
.A2(n_88),
.B(n_113),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_77),
.B(n_80),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_77),
.B(n_80),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_81),
.B(n_86),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_81),
.A2(n_82),
.B1(n_86),
.B2(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_83),
.A2(n_84),
.B(n_85),
.Y(n_82)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_100),
.B(n_112),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_98),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_98),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_92),
.B1(n_94),
.B2(n_97),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_93),
.A2(n_95),
.B(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_101),
.A2(n_105),
.B(n_111),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_102),
.B(n_103),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_110),
.Y(n_105)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);


endmodule