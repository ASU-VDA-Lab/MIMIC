module fake_jpeg_10805_n_105 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_29, n_12, n_8, n_15, n_7, n_105);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_105;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_9),
.B(n_24),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_0),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_43),
.B(n_0),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_45),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_1),
.Y(n_45)
);

CKINVDCx6p67_ASAP7_75t_R g46 ( 
.A(n_38),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_50),
.Y(n_55)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_33),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_51),
.B(n_41),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_53),
.B(n_54),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_37),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_50),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_59),
.B(n_35),
.Y(n_68)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_61),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_47),
.A2(n_34),
.B1(n_32),
.B2(n_36),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_SL g69 ( 
.A(n_62),
.B(n_42),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_52),
.B(n_40),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_66),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_55),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_68),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_70),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_1),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_58),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_74),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_58),
.B(n_2),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_52),
.B(n_2),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_75),
.A2(n_3),
.B1(n_4),
.B2(n_8),
.Y(n_80)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_76),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_65),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_83),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_80),
.B(n_89),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_82),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_64),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_63),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_87)
);

INVxp33_ASAP7_75t_L g92 ( 
.A(n_87),
.Y(n_92)
);

OAI21xp33_ASAP7_75t_L g96 ( 
.A1(n_90),
.A2(n_82),
.B(n_78),
.Y(n_96)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_84),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_93),
.B(n_94),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_21),
.C(n_22),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_96),
.B(n_98),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_91),
.B(n_88),
.C(n_86),
.Y(n_98)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_97),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_100),
.A2(n_95),
.B(n_92),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_101),
.A2(n_92),
.B1(n_99),
.B2(n_85),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_102),
.B(n_79),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_103),
.A2(n_79),
.B1(n_26),
.B2(n_28),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_23),
.Y(n_105)
);


endmodule