module real_jpeg_13340_n_12 (n_5, n_4, n_8, n_0, n_274, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_274;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_173;
wire n_40;
wire n_105;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_211;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_258;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_259;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_213;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_89;
wire n_16;

BUFx12f_ASAP7_75t_L g106 ( 
.A(n_0),
.Y(n_106)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx4f_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_4),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_5),
.A2(n_20),
.B1(n_23),
.B2(n_33),
.Y(n_32)
);

CKINVDCx14_ASAP7_75t_R g33 ( 
.A(n_5),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_5),
.A2(n_29),
.B1(n_30),
.B2(n_33),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_5),
.A2(n_33),
.B1(n_42),
.B2(n_43),
.Y(n_98)
);

O2A1O1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_5),
.A2(n_7),
.B(n_29),
.C(n_102),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_5),
.A2(n_33),
.B1(n_53),
.B2(n_54),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_5),
.B(n_34),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_5),
.B(n_51),
.C(n_54),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_5),
.B(n_41),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_5),
.B(n_26),
.C(n_30),
.Y(n_173)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

AO22x1_ASAP7_75t_L g41 ( 
.A1(n_7),
.A2(n_39),
.B1(n_42),
.B2(n_43),
.Y(n_41)
);

BUFx8_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_9),
.A2(n_29),
.B1(n_30),
.B2(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_9),
.A2(n_42),
.B1(n_43),
.B2(n_45),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_9),
.A2(n_45),
.B1(n_53),
.B2(n_54),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_10),
.A2(n_20),
.B1(n_22),
.B2(n_23),
.Y(n_19)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_10),
.A2(n_22),
.B1(n_29),
.B2(n_30),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_10),
.A2(n_22),
.B1(n_42),
.B2(n_43),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_10),
.A2(n_22),
.B1(n_53),
.B2(n_54),
.Y(n_120)
);

OAI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_11),
.A2(n_29),
.B1(n_30),
.B2(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_11),
.A2(n_20),
.B1(n_23),
.B2(n_37),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_11),
.A2(n_37),
.B1(n_53),
.B2(n_54),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_11),
.A2(n_37),
.B1(n_42),
.B2(n_43),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_82),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_80),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_67),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_15),
.B(n_67),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_59),
.Y(n_15)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_35),
.C(n_46),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_17),
.A2(n_69),
.B1(n_70),
.B2(n_71),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_17),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_17),
.A2(n_69),
.B1(n_113),
.B2(n_123),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_17),
.B(n_123),
.C(n_185),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_17),
.A2(n_69),
.B1(n_91),
.B2(n_92),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_24),
.B1(n_32),
.B2(n_34),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

OA21x2_ASAP7_75t_L g74 ( 
.A1(n_19),
.A2(n_28),
.B(n_62),
.Y(n_74)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_20),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_20),
.A2(n_23),
.B1(n_26),
.B2(n_27),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_23),
.B(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_24),
.B(n_32),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_24),
.B(n_34),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_28),
.Y(n_24)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_26),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_26),
.A2(n_27),
.B1(n_29),
.B2(n_30),
.Y(n_28)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_L g60 ( 
.A1(n_28),
.A2(n_61),
.B(n_62),
.Y(n_60)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

O2A1O1Ixp33_ASAP7_75t_L g38 ( 
.A1(n_30),
.A2(n_39),
.B(n_40),
.C(n_41),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_39),
.Y(n_40)
);

BUFx4f_ASAP7_75t_SL g30 ( 
.A(n_31),
.Y(n_30)
);

INVxp33_ASAP7_75t_L g242 ( 
.A(n_32),
.Y(n_242)
);

OAI21xp33_ASAP7_75t_SL g102 ( 
.A1(n_33),
.A2(n_39),
.B(n_42),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_33),
.B(n_109),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_33),
.B(n_57),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_35),
.A2(n_46),
.B1(n_72),
.B2(n_73),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_35),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_38),
.B1(n_41),
.B2(n_44),
.Y(n_35)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_36),
.Y(n_77)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_38),
.B(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_42),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_42),
.A2(n_43),
.B1(n_50),
.B2(n_51),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_43),
.B(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_64),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_46),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_46),
.B(n_74),
.C(n_76),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_46),
.A2(n_73),
.B1(n_76),
.B2(n_260),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_57),
.B(n_58),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_47),
.A2(n_57),
.B(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_48),
.B(n_98),
.Y(n_97)
);

AO22x1_ASAP7_75t_SL g128 ( 
.A1(n_48),
.A2(n_52),
.B1(n_96),
.B2(n_98),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_48),
.A2(n_52),
.B1(n_247),
.B2(n_248),
.Y(n_246)
);

NOR2x1_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_52),
.Y(n_48)
);

AO22x1_ASAP7_75t_L g52 ( 
.A1(n_50),
.A2(n_51),
.B1(n_53),
.B2(n_54),
.Y(n_52)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_52),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_53),
.B(n_152),
.Y(n_151)
);

INVx3_ASAP7_75t_SL g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_54),
.B(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

OA21x2_ASAP7_75t_L g94 ( 
.A1(n_57),
.A2(n_95),
.B(n_97),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_57),
.A2(n_97),
.B(n_226),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_58),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_63),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_65),
.B(n_66),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_65),
.A2(n_66),
.B1(n_93),
.B2(n_114),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_65),
.A2(n_66),
.B(n_114),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_66),
.A2(n_77),
.B(n_78),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_66),
.A2(n_78),
.B(n_93),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_74),
.C(n_75),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_68),
.A2(n_74),
.B1(n_175),
.B2(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_68),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_69),
.B(n_92),
.C(n_218),
.Y(n_250)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_74),
.A2(n_175),
.B1(n_176),
.B2(n_177),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_74),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_74),
.A2(n_175),
.B1(n_200),
.B2(n_201),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_74),
.A2(n_175),
.B1(n_258),
.B2(n_259),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_75),
.B(n_266),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_76),
.Y(n_260)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_79),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

AOI21xp33_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_252),
.B(n_269),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_85),
.A2(n_230),
.B(n_251),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_213),
.B(n_229),
.Y(n_85)
);

OAI321xp33_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_182),
.A3(n_208),
.B1(n_211),
.B2(n_212),
.C(n_274),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_165),
.B(n_181),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_131),
.B(n_164),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_110),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_90),
.B(n_110),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_94),
.C(n_99),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_91),
.A2(n_92),
.B1(n_94),
.B2(n_148),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_91),
.A2(n_92),
.B1(n_178),
.B2(n_179),
.Y(n_177)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_92),
.B(n_175),
.C(n_179),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_94),
.B(n_135),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_94),
.A2(n_135),
.B1(n_147),
.B2(n_148),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_94),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_94),
.A2(n_148),
.B1(n_188),
.B2(n_190),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_98),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_99),
.A2(n_100),
.B1(n_161),
.B2(n_162),
.Y(n_160)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_103),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_101),
.B(n_103),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_105),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_104),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_104),
.A2(n_108),
.B1(n_109),
.B2(n_120),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_105),
.B(n_206),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_107),
.Y(n_105)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_106),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_107),
.B(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_108),
.A2(n_109),
.B1(n_189),
.B2(n_206),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_109),
.A2(n_120),
.B(n_121),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_109),
.A2(n_121),
.B(n_189),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_111),
.A2(n_112),
.B1(n_125),
.B2(n_126),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_111),
.B(n_128),
.C(n_129),
.Y(n_166)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_115),
.B1(n_123),
.B2(n_124),
.Y(n_112)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_113),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_113),
.B(n_116),
.C(n_119),
.Y(n_169)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_115),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_117),
.B1(n_118),
.B2(n_119),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_118),
.B(n_146),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_118),
.B(n_146),
.Y(n_156)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_119),
.B(n_151),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_123),
.A2(n_246),
.B(n_249),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_123),
.B(n_246),
.Y(n_249)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_127),
.A2(n_128),
.B1(n_129),
.B2(n_130),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_127),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_128),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_128),
.A2(n_130),
.B1(n_139),
.B2(n_140),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_128),
.B(n_140),
.C(n_142),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_128),
.A2(n_130),
.B1(n_204),
.B2(n_205),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_128),
.B(n_205),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_158),
.B(n_163),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_144),
.B(n_157),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_137),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_134),
.B(n_137),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_135),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_141),
.B1(n_142),
.B2(n_143),
.Y(n_137)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_138),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_139),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_141),
.A2(n_142),
.B1(n_171),
.B2(n_172),
.Y(n_170)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_142),
.B(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_142),
.B(n_154),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_142),
.B(n_171),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_149),
.B(n_156),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_148),
.B(n_188),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_153),
.B(n_155),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_159),
.B(n_160),
.Y(n_163)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_167),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_166),
.B(n_167),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_174),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_169),
.B(n_170),
.C(n_174),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_172),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_175),
.B(n_196),
.C(n_201),
.Y(n_215)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_192),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_183),
.B(n_192),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_187),
.C(n_191),
.Y(n_183)
);

FAx1_ASAP7_75t_SL g210 ( 
.A(n_184),
.B(n_187),
.CI(n_191),
.CON(n_210),
.SN(n_210)
);

XNOR2xp5_ASAP7_75t_SL g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_188),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_207),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_194),
.A2(n_195),
.B1(n_202),
.B2(n_203),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_194),
.B(n_203),
.C(n_207),
.Y(n_228)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_197),
.B1(n_198),
.B2(n_199),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_209),
.B(n_210),
.Y(n_211)
);

BUFx24_ASAP7_75t_SL g272 ( 
.A(n_210),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_214),
.B(n_228),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_214),
.B(n_228),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_215),
.B(n_217),
.C(n_222),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_222),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_219),
.B1(n_220),
.B2(n_221),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_224),
.B1(n_225),
.B2(n_227),
.Y(n_222)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_223),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_225),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_223),
.A2(n_227),
.B1(n_240),
.B2(n_241),
.Y(n_239)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_226),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_227),
.A2(n_236),
.B(n_241),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_231),
.B(n_232),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_250),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_234),
.A2(n_235),
.B1(n_244),
.B2(n_245),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_235),
.B(n_244),
.C(n_250),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_237),
.B1(n_238),
.B2(n_239),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_237),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_249),
.A2(n_256),
.B1(n_257),
.B2(n_261),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_249),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_264),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_254),
.B(n_263),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_254),
.B(n_263),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_262),
.Y(n_254)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_257),
.B(n_261),
.C(n_262),
.Y(n_268)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_264),
.A2(n_270),
.B(n_271),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_265),
.B(n_268),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_265),
.B(n_268),
.Y(n_271)
);


endmodule