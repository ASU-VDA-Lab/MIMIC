module real_aes_11905_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_800;
wire n_778;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_528;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_860;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_874;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_505;
wire n_434;
wire n_502;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_880;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
INVx1_ASAP7_75t_L g197 ( .A(n_0), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_1), .B(n_253), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_2), .B(n_178), .Y(n_608) );
CKINVDCx5p33_ASAP7_75t_R g208 ( .A(n_3), .Y(n_208) );
NAND2xp5_ASAP7_75t_SL g257 ( .A(n_4), .B(n_177), .Y(n_257) );
INVx1_ASAP7_75t_L g108 ( .A(n_5), .Y(n_108) );
NOR2xp67_ASAP7_75t_L g122 ( .A(n_5), .B(n_85), .Y(n_122) );
NAND2xp5_ASAP7_75t_SL g606 ( .A(n_6), .B(n_151), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_7), .B(n_144), .Y(n_599) );
CKINVDCx5p33_ASAP7_75t_R g319 ( .A(n_8), .Y(n_319) );
CKINVDCx5p33_ASAP7_75t_R g327 ( .A(n_9), .Y(n_327) );
NAND2x1p5_ASAP7_75t_L g553 ( .A(n_10), .B(n_144), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_11), .B(n_275), .Y(n_623) );
CKINVDCx5p33_ASAP7_75t_R g877 ( .A(n_12), .Y(n_877) );
AOI22xp5_ASAP7_75t_L g872 ( .A1(n_13), .A2(n_98), .B1(n_873), .B2(n_874), .Y(n_872) );
INVx1_ASAP7_75t_L g873 ( .A(n_13), .Y(n_873) );
NAND2xp5_ASAP7_75t_SL g238 ( .A(n_14), .B(n_239), .Y(n_238) );
AND2x2_ASAP7_75t_L g580 ( .A(n_15), .B(n_581), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_16), .B(n_160), .Y(n_159) );
CKINVDCx5p33_ASAP7_75t_R g278 ( .A(n_17), .Y(n_278) );
CKINVDCx5p33_ASAP7_75t_R g189 ( .A(n_18), .Y(n_189) );
NAND2xp5_ASAP7_75t_SL g243 ( .A(n_19), .B(n_151), .Y(n_243) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_20), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_21), .B(n_154), .Y(n_153) );
NAND2xp5_ASAP7_75t_SL g531 ( .A(n_22), .B(n_169), .Y(n_531) );
CKINVDCx5p33_ASAP7_75t_R g224 ( .A(n_23), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_24), .B(n_191), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_25), .B(n_160), .Y(n_256) );
NAND2xp33_ASAP7_75t_L g549 ( .A(n_26), .B(n_177), .Y(n_549) );
NAND2xp33_ASAP7_75t_L g598 ( .A(n_27), .B(n_177), .Y(n_598) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_28), .Y(n_152) );
OAI21xp33_ASAP7_75t_L g274 ( .A1(n_29), .A2(n_185), .B(n_275), .Y(n_274) );
CKINVDCx5p33_ASAP7_75t_R g562 ( .A(n_30), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_31), .A2(n_102), .B1(n_103), .B2(n_114), .Y(n_101) );
NAND2xp5_ASAP7_75t_SL g251 ( .A(n_32), .B(n_151), .Y(n_251) );
CKINVDCx5p33_ASAP7_75t_R g187 ( .A(n_33), .Y(n_187) );
NAND2xp5_ASAP7_75t_SL g552 ( .A(n_34), .B(n_188), .Y(n_552) );
NOR2xp33_ASAP7_75t_L g109 ( .A(n_35), .B(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g121 ( .A(n_35), .Y(n_121) );
OAI21x1_ASAP7_75t_L g146 ( .A1(n_36), .A2(n_67), .B(n_147), .Y(n_146) );
A2O1A1Ixp33_ASAP7_75t_L g583 ( .A1(n_37), .A2(n_156), .B(n_584), .C(n_586), .Y(n_583) );
CKINVDCx5p33_ASAP7_75t_R g221 ( .A(n_38), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_39), .B(n_151), .Y(n_150) );
CKINVDCx5p33_ASAP7_75t_R g322 ( .A(n_40), .Y(n_322) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_41), .B(n_161), .Y(n_527) );
CKINVDCx5p33_ASAP7_75t_R g529 ( .A(n_42), .Y(n_529) );
NAND2xp33_ASAP7_75t_L g626 ( .A(n_43), .B(n_239), .Y(n_626) );
AND2x6_ASAP7_75t_L g166 ( .A(n_44), .B(n_167), .Y(n_166) );
AOI22xp33_ASAP7_75t_L g276 ( .A1(n_45), .A2(n_81), .B1(n_177), .B2(n_241), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_46), .B(n_191), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_47), .B(n_160), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_48), .B(n_585), .Y(n_597) );
NAND2xp33_ASAP7_75t_L g609 ( .A(n_49), .B(n_239), .Y(n_609) );
CKINVDCx5p33_ASAP7_75t_R g179 ( .A(n_50), .Y(n_179) );
INVx1_ASAP7_75t_L g167 ( .A(n_51), .Y(n_167) );
CKINVDCx5p33_ASAP7_75t_R g570 ( .A(n_52), .Y(n_570) );
OAI22x1_ASAP7_75t_R g860 ( .A1(n_53), .A2(n_89), .B1(n_861), .B2(n_862), .Y(n_860) );
INVx1_ASAP7_75t_L g862 ( .A(n_53), .Y(n_862) );
CKINVDCx5p33_ASAP7_75t_R g222 ( .A(n_54), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_55), .B(n_241), .Y(n_244) );
NAND2xp5_ASAP7_75t_SL g622 ( .A(n_56), .B(n_239), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_57), .B(n_241), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_58), .B(n_169), .Y(n_168) );
CKINVDCx5p33_ASAP7_75t_R g181 ( .A(n_59), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_60), .B(n_191), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_61), .B(n_253), .Y(n_252) );
CKINVDCx5p33_ASAP7_75t_R g524 ( .A(n_62), .Y(n_524) );
AND2x2_ASAP7_75t_L g111 ( .A(n_63), .B(n_112), .Y(n_111) );
AND2x2_ASAP7_75t_L g588 ( .A(n_64), .B(n_191), .Y(n_588) );
INVx2_ASAP7_75t_L g209 ( .A(n_65), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_66), .B(n_241), .Y(n_539) );
CKINVDCx5p33_ASAP7_75t_R g551 ( .A(n_68), .Y(n_551) );
NAND2xp33_ASAP7_75t_L g538 ( .A(n_69), .B(n_207), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g162 ( .A(n_70), .B(n_161), .Y(n_162) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_71), .Y(n_116) );
INVx1_ASAP7_75t_L g201 ( .A(n_72), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_73), .B(n_253), .Y(n_625) );
CKINVDCx5p33_ASAP7_75t_R g330 ( .A(n_74), .Y(n_330) );
BUFx10_ASAP7_75t_L g128 ( .A(n_75), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_76), .B(n_526), .Y(n_595) );
NAND2xp33_ASAP7_75t_L g542 ( .A(n_77), .B(n_151), .Y(n_542) );
INVx1_ASAP7_75t_L g324 ( .A(n_78), .Y(n_324) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_79), .B(n_161), .Y(n_226) );
NAND2xp5_ASAP7_75t_SL g594 ( .A(n_80), .B(n_177), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_82), .B(n_191), .Y(n_246) );
INVx1_ASAP7_75t_L g212 ( .A(n_83), .Y(n_212) );
CKINVDCx5p33_ASAP7_75t_R g587 ( .A(n_84), .Y(n_587) );
INVx1_ASAP7_75t_L g107 ( .A(n_85), .Y(n_107) );
INVx2_ASAP7_75t_L g147 ( .A(n_86), .Y(n_147) );
INVx1_ASAP7_75t_L g113 ( .A(n_87), .Y(n_113) );
OR2x2_ASAP7_75t_L g118 ( .A(n_87), .B(n_119), .Y(n_118) );
BUFx2_ASAP7_75t_L g512 ( .A(n_87), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g880 ( .A(n_87), .B(n_120), .Y(n_880) );
CKINVDCx5p33_ASAP7_75t_R g567 ( .A(n_88), .Y(n_567) );
INVx1_ASAP7_75t_L g861 ( .A(n_89), .Y(n_861) );
NAND2xp5_ASAP7_75t_SL g530 ( .A(n_90), .B(n_188), .Y(n_530) );
CKINVDCx5p33_ASAP7_75t_R g604 ( .A(n_91), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_92), .B(n_169), .Y(n_628) );
INVx1_ASAP7_75t_L g112 ( .A(n_93), .Y(n_112) );
INVx1_ASAP7_75t_L g579 ( .A(n_94), .Y(n_579) );
CKINVDCx5p33_ASAP7_75t_R g564 ( .A(n_95), .Y(n_564) );
NOR2xp67_ASAP7_75t_L g271 ( .A(n_96), .B(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g571 ( .A(n_97), .B(n_144), .Y(n_571) );
INVx1_ASAP7_75t_L g874 ( .A(n_98), .Y(n_874) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_99), .B(n_191), .Y(n_543) );
NAND2xp33_ASAP7_75t_L g217 ( .A(n_100), .B(n_191), .Y(n_217) );
INVx1_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
BUFx6f_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
AND2x2_ASAP7_75t_L g105 ( .A(n_106), .B(n_109), .Y(n_105) );
NOR2xp33_ASAP7_75t_SL g106 ( .A(n_107), .B(n_108), .Y(n_106) );
NAND2xp5_ASAP7_75t_SL g110 ( .A(n_111), .B(n_113), .Y(n_110) );
OR2x6_ASAP7_75t_L g114 ( .A(n_115), .B(n_123), .Y(n_114) );
INVx1_ASAP7_75t_L g875 ( .A(n_115), .Y(n_875) );
NOR2xp67_ASAP7_75t_SL g115 ( .A(n_116), .B(n_117), .Y(n_115) );
INVx4_ASAP7_75t_L g870 ( .A(n_117), .Y(n_870) );
BUFx6f_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
OR2x6_ASAP7_75t_L g126 ( .A(n_120), .B(n_127), .Y(n_126) );
AND2x4_ASAP7_75t_L g120 ( .A(n_121), .B(n_122), .Y(n_120) );
OAI21xp5_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_129), .B(n_864), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
OR2x2_ASAP7_75t_L g879 ( .A(n_127), .B(n_880), .Y(n_879) );
INVx2_ASAP7_75t_SL g127 ( .A(n_128), .Y(n_127) );
BUFx12f_ASAP7_75t_L g868 ( .A(n_128), .Y(n_868) );
INVx2_ASAP7_75t_SL g129 ( .A(n_130), .Y(n_129) );
OAI22x1_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_859), .B1(n_860), .B2(n_863), .Y(n_130) );
INVx2_ASAP7_75t_L g863 ( .A(n_131), .Y(n_863) );
OAI22x1_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_511), .B1(n_513), .B2(n_858), .Y(n_131) );
XNOR2x1_ASAP7_75t_L g871 ( .A(n_132), .B(n_872), .Y(n_871) );
AND2x4_ASAP7_75t_L g132 ( .A(n_133), .B(n_448), .Y(n_132) );
NOR2x1_ASAP7_75t_L g133 ( .A(n_134), .B(n_375), .Y(n_133) );
NAND3xp33_ASAP7_75t_L g134 ( .A(n_135), .B(n_308), .C(n_355), .Y(n_134) );
NOR2xp33_ASAP7_75t_L g135 ( .A(n_136), .B(n_290), .Y(n_135) );
OAI21xp33_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_214), .B(n_260), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
AOI322xp5_ASAP7_75t_L g456 ( .A1(n_138), .A2(n_305), .A3(n_457), .B1(n_459), .B2(n_461), .C1(n_465), .C2(n_467), .Y(n_456) );
AND2x2_ASAP7_75t_L g138 ( .A(n_139), .B(n_171), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
AOI322xp5_ASAP7_75t_L g308 ( .A1(n_140), .A2(n_309), .A3(n_333), .B1(n_336), .B2(n_338), .C1(n_343), .C2(n_347), .Y(n_308) );
AND2x2_ASAP7_75t_L g425 ( .A(n_140), .B(n_171), .Y(n_425) );
AND2x2_ASAP7_75t_L g427 ( .A(n_140), .B(n_428), .Y(n_427) );
INVx2_ASAP7_75t_L g477 ( .A(n_140), .Y(n_477) );
OR2x2_ASAP7_75t_L g495 ( .A(n_140), .B(n_471), .Y(n_495) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
AND2x4_ASAP7_75t_L g299 ( .A(n_141), .B(n_300), .Y(n_299) );
AND2x4_ASAP7_75t_L g344 ( .A(n_141), .B(n_268), .Y(n_344) );
BUFx3_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx2_ASAP7_75t_L g263 ( .A(n_142), .Y(n_263) );
OAI21x1_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_148), .B(n_168), .Y(n_142) );
OAI21x1_ASAP7_75t_SL g248 ( .A1(n_143), .A2(n_249), .B(n_259), .Y(n_248) );
OAI21x1_ASAP7_75t_L g521 ( .A1(n_143), .A2(n_522), .B(n_531), .Y(n_521) );
OA21x2_ASAP7_75t_L g545 ( .A1(n_143), .A2(n_546), .B(n_553), .Y(n_545) );
OA21x2_ASAP7_75t_L g601 ( .A1(n_143), .A2(n_602), .B(n_610), .Y(n_601) );
OAI21x1_ASAP7_75t_L g618 ( .A1(n_143), .A2(n_522), .B(n_531), .Y(n_618) );
OAI21x1_ASAP7_75t_L g647 ( .A1(n_143), .A2(n_546), .B(n_553), .Y(n_647) );
BUFx4f_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
NOR2xp33_ASAP7_75t_L g182 ( .A(n_144), .B(n_183), .Y(n_182) );
INVx3_ASAP7_75t_L g235 ( .A(n_144), .Y(n_235) );
OA21x2_ASAP7_75t_L g535 ( .A1(n_144), .A2(n_536), .B(n_543), .Y(n_535) );
INVx4_ASAP7_75t_L g558 ( .A(n_144), .Y(n_558) );
OA21x2_ASAP7_75t_L g641 ( .A1(n_144), .A2(n_536), .B(n_543), .Y(n_641) );
OA21x2_ASAP7_75t_L g673 ( .A1(n_144), .A2(n_536), .B(n_543), .Y(n_673) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx2_ASAP7_75t_L g170 ( .A(n_145), .Y(n_170) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx1_ASAP7_75t_L g192 ( .A(n_146), .Y(n_192) );
OAI21x1_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_158), .B(n_164), .Y(n_148) );
AOI21xp5_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_153), .B(n_156), .Y(n_149) );
INVx2_ASAP7_75t_L g199 ( .A(n_151), .Y(n_199) );
INVx2_ASAP7_75t_L g253 ( .A(n_151), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g561 ( .A(n_151), .B(n_562), .Y(n_561) );
INVx2_ASAP7_75t_SL g585 ( .A(n_151), .Y(n_585) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_152), .Y(n_155) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_152), .Y(n_161) );
INVx2_ASAP7_75t_L g178 ( .A(n_152), .Y(n_178) );
BUFx6f_ASAP7_75t_L g207 ( .A(n_152), .Y(n_207) );
INVx1_ASAP7_75t_L g321 ( .A(n_152), .Y(n_321) );
NOR2xp33_ASAP7_75t_L g200 ( .A(n_154), .B(n_201), .Y(n_200) );
INVxp67_ASAP7_75t_L g225 ( .A(n_154), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g329 ( .A(n_154), .B(n_330), .Y(n_329) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx2_ASAP7_75t_L g180 ( .A(n_155), .Y(n_180) );
INVx2_ASAP7_75t_L g569 ( .A(n_155), .Y(n_569) );
INVx2_ASAP7_75t_SL g163 ( .A(n_156), .Y(n_163) );
CKINVDCx6p67_ASAP7_75t_R g219 ( .A(n_156), .Y(n_219) );
INVx2_ASAP7_75t_SL g227 ( .A(n_156), .Y(n_227) );
INVx5_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx5_ASAP7_75t_L g175 ( .A(n_157), .Y(n_175) );
BUFx12f_ASAP7_75t_L g185 ( .A(n_157), .Y(n_185) );
O2A1O1Ixp33_ASAP7_75t_L g523 ( .A1(n_157), .A2(n_524), .B(n_525), .C(n_527), .Y(n_523) );
AOI21xp5_ASAP7_75t_L g158 ( .A1(n_159), .A2(n_162), .B(n_163), .Y(n_158) );
OAI22xp5_ASAP7_75t_L g204 ( .A1(n_160), .A2(n_205), .B1(n_208), .B2(n_209), .Y(n_204) );
OAI22xp5_ASAP7_75t_L g220 ( .A1(n_160), .A2(n_177), .B1(n_221), .B2(n_222), .Y(n_220) );
NOR2xp67_ASAP7_75t_L g563 ( .A(n_160), .B(n_564), .Y(n_563) );
INVx5_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
OR2x2_ASAP7_75t_L g326 ( .A(n_161), .B(n_327), .Y(n_326) );
OAI21xp5_ASAP7_75t_L g560 ( .A1(n_163), .A2(n_561), .B(n_563), .Y(n_560) );
INVx2_ASAP7_75t_SL g164 ( .A(n_165), .Y(n_164) );
INVx8_ASAP7_75t_L g245 ( .A(n_165), .Y(n_245) );
OAI21xp5_ASAP7_75t_L g331 ( .A1(n_165), .A2(n_169), .B(n_332), .Y(n_331) );
AOI21xp5_ASAP7_75t_L g559 ( .A1(n_165), .A2(n_560), .B(n_565), .Y(n_559) );
NOR2xp67_ASAP7_75t_L g574 ( .A(n_165), .B(n_575), .Y(n_574) );
INVx8_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx1_ASAP7_75t_L g183 ( .A(n_166), .Y(n_183) );
AOI21xp33_ASAP7_75t_L g213 ( .A1(n_166), .A2(n_170), .B(n_211), .Y(n_213) );
INVx1_ASAP7_75t_L g229 ( .A(n_166), .Y(n_229) );
BUFx2_ASAP7_75t_L g627 ( .A(n_166), .Y(n_627) );
INVx3_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g211 ( .A(n_170), .B(n_212), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g323 ( .A(n_170), .B(n_324), .Y(n_323) );
AND2x4_ASAP7_75t_SL g298 ( .A(n_171), .B(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g171 ( .A(n_172), .B(n_193), .Y(n_171) );
AND2x2_ASAP7_75t_L g262 ( .A(n_172), .B(n_263), .Y(n_262) );
INVx2_ASAP7_75t_SL g172 ( .A(n_173), .Y(n_172) );
AND2x4_ASAP7_75t_L g284 ( .A(n_173), .B(n_267), .Y(n_284) );
AND2x2_ASAP7_75t_L g335 ( .A(n_173), .B(n_282), .Y(n_335) );
OR2x2_ASAP7_75t_L g346 ( .A(n_173), .B(n_283), .Y(n_346) );
INVx1_ASAP7_75t_L g366 ( .A(n_173), .Y(n_366) );
AND2x2_ASAP7_75t_L g374 ( .A(n_173), .B(n_283), .Y(n_374) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_173), .Y(n_384) );
AND2x2_ASAP7_75t_L g437 ( .A(n_173), .B(n_263), .Y(n_437) );
OA21x2_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_184), .B(n_190), .Y(n_173) );
OAI21xp33_ASAP7_75t_L g174 ( .A1(n_175), .A2(n_176), .B(n_182), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_175), .A2(n_243), .B(n_244), .Y(n_242) );
INVx1_ASAP7_75t_L g258 ( .A(n_175), .Y(n_258) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_175), .A2(n_541), .B(n_542), .Y(n_540) );
AOI21x1_ASAP7_75t_L g621 ( .A1(n_175), .A2(n_622), .B(n_623), .Y(n_621) );
OAI22xp33_ASAP7_75t_L g176 ( .A1(n_177), .A2(n_179), .B1(n_180), .B2(n_181), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g586 ( .A(n_177), .B(n_587), .Y(n_586) );
INVx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVx1_ASAP7_75t_L g188 ( .A(n_178), .Y(n_188) );
INVx2_ASAP7_75t_L g239 ( .A(n_178), .Y(n_239) );
AOI22xp5_ASAP7_75t_L g186 ( .A1(n_180), .A2(n_187), .B1(n_188), .B2(n_189), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g184 ( .A(n_185), .B(n_186), .Y(n_184) );
BUFx2_ASAP7_75t_L g202 ( .A(n_185), .Y(n_202) );
CKINVDCx5p33_ASAP7_75t_R g210 ( .A(n_185), .Y(n_210) );
INVx3_ASAP7_75t_L g254 ( .A(n_185), .Y(n_254) );
OAI22xp5_ASAP7_75t_L g270 ( .A1(n_185), .A2(n_271), .B1(n_274), .B2(n_276), .Y(n_270) );
AOI21xp5_ASAP7_75t_L g624 ( .A1(n_185), .A2(n_625), .B(n_626), .Y(n_624) );
NOR2x1p5_ASAP7_75t_SL g228 ( .A(n_191), .B(n_229), .Y(n_228) );
INVx2_ASAP7_75t_L g269 ( .A(n_191), .Y(n_269) );
BUFx5_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
INVx1_ASAP7_75t_L g279 ( .A(n_192), .Y(n_279) );
INVx2_ASAP7_75t_L g265 ( .A(n_193), .Y(n_265) );
AND2x2_ASAP7_75t_L g364 ( .A(n_193), .B(n_263), .Y(n_364) );
AND2x2_ASAP7_75t_L g441 ( .A(n_193), .B(n_405), .Y(n_441) );
INVx2_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
INVx2_ASAP7_75t_L g283 ( .A(n_194), .Y(n_283) );
AO21x2_ASAP7_75t_L g194 ( .A1(n_195), .A2(n_203), .B(n_213), .Y(n_194) );
OAI21xp5_ASAP7_75t_L g195 ( .A1(n_196), .A2(n_200), .B(n_202), .Y(n_195) );
NOR2x1_ASAP7_75t_L g196 ( .A(n_197), .B(n_198), .Y(n_196) );
O2A1O1Ixp33_ASAP7_75t_L g528 ( .A1(n_198), .A2(n_254), .B(n_529), .C(n_530), .Y(n_528) );
O2A1O1Ixp5_ASAP7_75t_L g550 ( .A1(n_198), .A2(n_254), .B(n_551), .C(n_552), .Y(n_550) );
INVx2_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
OAI22xp5_ASAP7_75t_L g318 ( .A1(n_199), .A2(n_319), .B1(n_320), .B2(n_322), .Y(n_318) );
OAI21x1_ASAP7_75t_L g577 ( .A1(n_202), .A2(n_578), .B(n_580), .Y(n_577) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_204), .A2(n_210), .B(n_211), .Y(n_203) );
INVx2_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
INVx2_ASAP7_75t_L g241 ( .A(n_207), .Y(n_241) );
INVx2_ASAP7_75t_L g273 ( .A(n_207), .Y(n_273) );
INVx2_ASAP7_75t_L g275 ( .A(n_207), .Y(n_275) );
INVx1_ASAP7_75t_L g526 ( .A(n_207), .Y(n_526) );
AO21x1_ASAP7_75t_L g317 ( .A1(n_210), .A2(n_318), .B(n_323), .Y(n_317) );
AOI21x1_ASAP7_75t_L g325 ( .A1(n_210), .A2(n_326), .B(n_328), .Y(n_325) );
OAI21xp33_ASAP7_75t_L g565 ( .A1(n_210), .A2(n_566), .B(n_568), .Y(n_565) );
AOI21xp5_ASAP7_75t_L g593 ( .A1(n_210), .A2(n_594), .B(n_595), .Y(n_593) );
OAI21xp5_ASAP7_75t_L g469 ( .A1(n_214), .A2(n_470), .B(n_472), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_215), .B(n_230), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_215), .B(n_307), .Y(n_361) );
HB1xp67_ASAP7_75t_SL g215 ( .A(n_216), .Y(n_215) );
INVx1_ASAP7_75t_L g287 ( .A(n_216), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_216), .B(n_296), .Y(n_295) );
INVx2_ASAP7_75t_L g342 ( .A(n_216), .Y(n_342) );
AND2x2_ASAP7_75t_L g354 ( .A(n_216), .B(n_288), .Y(n_354) );
INVx1_ASAP7_75t_L g370 ( .A(n_216), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_216), .B(n_340), .Y(n_447) );
INVx1_ASAP7_75t_L g463 ( .A(n_216), .Y(n_463) );
AND2x2_ASAP7_75t_L g480 ( .A(n_216), .B(n_314), .Y(n_480) );
AND2x4_ASAP7_75t_L g216 ( .A(n_217), .B(n_218), .Y(n_216) );
A2O1A1Ixp33_ASAP7_75t_L g218 ( .A1(n_219), .A2(n_220), .B(n_223), .C(n_228), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_219), .A2(n_238), .B(n_240), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g537 ( .A1(n_219), .A2(n_538), .B(n_539), .Y(n_537) );
AOI21xp5_ASAP7_75t_L g547 ( .A1(n_219), .A2(n_548), .B(n_549), .Y(n_547) );
AOI21xp5_ASAP7_75t_L g607 ( .A1(n_219), .A2(n_608), .B(n_609), .Y(n_607) );
O2A1O1Ixp33_ASAP7_75t_L g223 ( .A1(n_224), .A2(n_225), .B(n_226), .C(n_227), .Y(n_223) );
AND2x2_ASAP7_75t_L g479 ( .A(n_230), .B(n_480), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_230), .B(n_499), .Y(n_498) );
AND2x4_ASAP7_75t_L g230 ( .A(n_231), .B(n_247), .Y(n_230) );
BUFx2_ASAP7_75t_L g289 ( .A(n_231), .Y(n_289) );
INVx1_ASAP7_75t_L g350 ( .A(n_231), .Y(n_350) );
AND2x4_ASAP7_75t_L g395 ( .A(n_231), .B(n_396), .Y(n_395) );
AND2x2_ASAP7_75t_L g415 ( .A(n_231), .B(n_342), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_231), .B(n_359), .Y(n_452) );
INVx3_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
AND2x4_ASAP7_75t_L g379 ( .A(n_232), .B(n_380), .Y(n_379) );
INVx2_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
INVx1_ASAP7_75t_L g296 ( .A(n_233), .Y(n_296) );
OAI21x1_ASAP7_75t_SL g233 ( .A1(n_234), .A2(n_236), .B(n_246), .Y(n_233) );
OAI21x1_ASAP7_75t_L g591 ( .A1(n_234), .A2(n_592), .B(n_599), .Y(n_591) );
OAI21xp5_ASAP7_75t_L g619 ( .A1(n_234), .A2(n_620), .B(n_628), .Y(n_619) );
OAI21x1_ASAP7_75t_L g653 ( .A1(n_234), .A2(n_620), .B(n_628), .Y(n_653) );
INVx2_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
OAI21xp5_ASAP7_75t_L g236 ( .A1(n_237), .A2(n_242), .B(n_245), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_239), .B(n_567), .Y(n_566) );
OAI21x1_ASAP7_75t_SL g249 ( .A1(n_245), .A2(n_250), .B(n_255), .Y(n_249) );
AO31x2_ASAP7_75t_L g268 ( .A1(n_245), .A2(n_269), .A3(n_270), .B(n_277), .Y(n_268) );
OAI21x1_ASAP7_75t_L g522 ( .A1(n_245), .A2(n_523), .B(n_528), .Y(n_522) );
OAI21x1_ASAP7_75t_L g536 ( .A1(n_245), .A2(n_537), .B(n_540), .Y(n_536) );
OAI21x1_ASAP7_75t_L g546 ( .A1(n_245), .A2(n_547), .B(n_550), .Y(n_546) );
OAI21x1_ASAP7_75t_L g592 ( .A1(n_245), .A2(n_593), .B(n_596), .Y(n_592) );
OAI21xp5_ASAP7_75t_L g602 ( .A1(n_245), .A2(n_603), .B(n_607), .Y(n_602) );
AND2x2_ASAP7_75t_L g312 ( .A(n_247), .B(n_296), .Y(n_312) );
AND2x2_ASAP7_75t_L g339 ( .A(n_247), .B(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g351 ( .A(n_247), .B(n_342), .Y(n_351) );
BUFx2_ASAP7_75t_L g378 ( .A(n_247), .Y(n_378) );
INVx2_ASAP7_75t_L g396 ( .A(n_247), .Y(n_396) );
BUFx3_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
INVx1_ASAP7_75t_L g288 ( .A(n_248), .Y(n_288) );
AOI21x1_ASAP7_75t_L g250 ( .A1(n_251), .A2(n_252), .B(n_254), .Y(n_250) );
O2A1O1Ixp5_ASAP7_75t_L g603 ( .A1(n_254), .A2(n_604), .B(n_605), .C(n_606), .Y(n_603) );
AOI21xp5_ASAP7_75t_L g255 ( .A1(n_256), .A2(n_257), .B(n_258), .Y(n_255) );
AOI21xp5_ASAP7_75t_L g596 ( .A1(n_258), .A2(n_597), .B(n_598), .Y(n_596) );
OAI21xp5_ASAP7_75t_L g260 ( .A1(n_261), .A2(n_280), .B(n_285), .Y(n_260) );
AND2x4_ASAP7_75t_L g261 ( .A(n_262), .B(n_264), .Y(n_261) );
AND2x2_ASAP7_75t_L g336 ( .A(n_262), .B(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_L g303 ( .A(n_263), .B(n_268), .Y(n_303) );
INVx1_ASAP7_75t_L g410 ( .A(n_263), .Y(n_410) );
HB1xp67_ASAP7_75t_L g440 ( .A(n_263), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_263), .B(n_265), .Y(n_510) );
AND2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
INVx2_ASAP7_75t_L g302 ( .A(n_265), .Y(n_302) );
HB1xp67_ASAP7_75t_L g372 ( .A(n_266), .Y(n_372) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
INVx2_ASAP7_75t_SL g267 ( .A(n_268), .Y(n_267) );
INVx2_ASAP7_75t_L g300 ( .A(n_268), .Y(n_300) );
AND2x2_ASAP7_75t_L g365 ( .A(n_268), .B(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g401 ( .A(n_268), .Y(n_401) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
INVx1_ASAP7_75t_L g605 ( .A(n_275), .Y(n_605) );
NOR2xp33_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
AND2x2_ASAP7_75t_L g280 ( .A(n_281), .B(n_284), .Y(n_280) );
INVx1_ASAP7_75t_L g429 ( .A(n_281), .Y(n_429) );
INVxp67_ASAP7_75t_SL g281 ( .A(n_282), .Y(n_281) );
AND2x4_ASAP7_75t_L g337 ( .A(n_282), .B(n_300), .Y(n_337) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g428 ( .A(n_284), .B(n_429), .Y(n_428) );
INVx2_ASAP7_75t_L g471 ( .A(n_284), .Y(n_471) );
AND2x4_ASAP7_75t_L g285 ( .A(n_286), .B(n_289), .Y(n_285) );
AND2x4_ASAP7_75t_L g305 ( .A(n_286), .B(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g434 ( .A(n_286), .B(n_404), .Y(n_434) );
AND2x4_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
INVx1_ASAP7_75t_L g294 ( .A(n_288), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_288), .B(n_296), .Y(n_391) );
OR2x2_ASAP7_75t_L g386 ( .A(n_289), .B(n_341), .Y(n_386) );
INVx1_ASAP7_75t_L g445 ( .A(n_289), .Y(n_445) );
OAI22xp5_ASAP7_75t_L g290 ( .A1(n_291), .A2(n_297), .B1(n_301), .B2(n_304), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_293), .B(n_295), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_294), .B(n_389), .Y(n_464) );
BUFx2_ASAP7_75t_L g491 ( .A(n_294), .Y(n_491) );
OR2x2_ASAP7_75t_L g506 ( .A(n_295), .B(n_313), .Y(n_506) );
INVx2_ASAP7_75t_L g307 ( .A(n_296), .Y(n_307) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
AOI221xp5_ASAP7_75t_L g496 ( .A1(n_298), .A2(n_381), .B1(n_446), .B2(n_497), .C(n_500), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_299), .B(n_383), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_302), .B(n_303), .Y(n_301) );
AOI322xp5_ASAP7_75t_L g503 ( .A1(n_302), .A2(n_365), .A3(n_476), .B1(n_504), .B2(n_505), .C1(n_507), .C2(n_508), .Y(n_503) );
INVx1_ASAP7_75t_L g421 ( .A(n_303), .Y(n_421) );
AOI22xp5_ASAP7_75t_L g439 ( .A1(n_303), .A2(n_388), .B1(n_440), .B2(n_441), .Y(n_439) );
NAND3xp33_ASAP7_75t_L g472 ( .A(n_303), .B(n_335), .C(n_473), .Y(n_472) );
AND2x2_ASAP7_75t_L g507 ( .A(n_303), .B(n_374), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_304), .B(n_413), .Y(n_412) );
INVx2_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g353 ( .A(n_307), .B(n_354), .Y(n_353) );
OR2x2_ASAP7_75t_L g367 ( .A(n_307), .B(n_368), .Y(n_367) );
AND2x4_ASAP7_75t_L g481 ( .A(n_307), .B(n_369), .Y(n_481) );
INVx2_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx2_ASAP7_75t_SL g310 ( .A(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g508 ( .A(n_311), .B(n_509), .Y(n_508) );
AND2x2_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_312), .B(n_341), .Y(n_406) );
INVx2_ASAP7_75t_L g394 ( .A(n_313), .Y(n_394) );
INVx2_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
HB1xp67_ASAP7_75t_L g359 ( .A(n_315), .Y(n_359) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g340 ( .A(n_316), .Y(n_340) );
BUFx3_ASAP7_75t_L g380 ( .A(n_316), .Y(n_380) );
OAI21x1_ASAP7_75t_L g316 ( .A1(n_317), .A2(n_325), .B(n_331), .Y(n_316) );
INVx2_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx2_ASAP7_75t_L g582 ( .A(n_321), .Y(n_582) );
INVxp67_ASAP7_75t_L g332 ( .A(n_323), .Y(n_332) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
AOI21xp33_ASAP7_75t_L g355 ( .A1(n_333), .A2(n_356), .B(n_360), .Y(n_355) );
AOI22xp5_ASAP7_75t_L g450 ( .A1(n_333), .A2(n_419), .B1(n_451), .B2(n_453), .Y(n_450) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
OR2x2_ASAP7_75t_L g420 ( .A(n_334), .B(n_421), .Y(n_420) );
INVx2_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx2_ASAP7_75t_SL g502 ( .A(n_336), .Y(n_502) );
AND2x4_ASAP7_75t_L g408 ( .A(n_337), .B(n_409), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_337), .B(n_437), .Y(n_436) );
NOR2x1_ASAP7_75t_L g486 ( .A(n_338), .B(n_487), .Y(n_486) );
AND2x4_ASAP7_75t_SL g338 ( .A(n_339), .B(n_341), .Y(n_338) );
INVx1_ASAP7_75t_L g423 ( .A(n_339), .Y(n_423) );
AND2x2_ASAP7_75t_L g369 ( .A(n_340), .B(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g389 ( .A(n_340), .Y(n_389) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
AND2x4_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
AND2x2_ASAP7_75t_L g397 ( .A(n_344), .B(n_373), .Y(n_397) );
INVx1_ASAP7_75t_L g418 ( .A(n_344), .Y(n_418) );
HB1xp67_ASAP7_75t_L g432 ( .A(n_344), .Y(n_432) );
INVx2_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
OR2x2_ASAP7_75t_L g458 ( .A(n_346), .B(n_404), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_348), .B(n_352), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
AND2x4_ASAP7_75t_L g349 ( .A(n_350), .B(n_351), .Y(n_349) );
AND2x2_ASAP7_75t_L g403 ( .A(n_351), .B(n_404), .Y(n_403) );
INVx2_ASAP7_75t_L g455 ( .A(n_351), .Y(n_455) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_353), .B(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g467 ( .A(n_358), .B(n_390), .Y(n_467) );
INVx1_ASAP7_75t_L g499 ( .A(n_358), .Y(n_499) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
OAI22xp5_ASAP7_75t_L g360 ( .A1(n_361), .A2(n_362), .B1(n_367), .B2(n_371), .Y(n_360) );
INVx2_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
AND2x4_ASAP7_75t_L g363 ( .A(n_364), .B(n_365), .Y(n_363) );
INVx1_ASAP7_75t_L g478 ( .A(n_365), .Y(n_478) );
AND2x2_ASAP7_75t_L g400 ( .A(n_366), .B(n_401), .Y(n_400) );
OAI21xp5_ASAP7_75t_L g430 ( .A1(n_367), .A2(n_431), .B(n_433), .Y(n_430) );
INVx1_ASAP7_75t_L g504 ( .A(n_367), .Y(n_504) );
INVx2_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_372), .B(n_373), .Y(n_371) );
BUFx3_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_374), .B(n_409), .Y(n_466) );
NAND3xp33_ASAP7_75t_L g375 ( .A(n_376), .B(n_411), .C(n_426), .Y(n_375) );
AOI221xp5_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_381), .B1(n_385), .B2(n_397), .C(n_398), .Y(n_376) );
AOI221xp5_ASAP7_75t_L g411 ( .A1(n_377), .A2(n_412), .B1(n_416), .B2(n_419), .C(n_422), .Y(n_411) );
AND2x4_ASAP7_75t_L g377 ( .A(n_378), .B(n_379), .Y(n_377) );
AND2x4_ASAP7_75t_L g414 ( .A(n_378), .B(n_415), .Y(n_414) );
AOI211xp5_ASAP7_75t_L g426 ( .A1(n_379), .A2(n_427), .B(n_430), .C(n_438), .Y(n_426) );
INVx2_ASAP7_75t_L g405 ( .A(n_380), .Y(n_405) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
OR2x2_ASAP7_75t_L g417 ( .A(n_383), .B(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
NAND3xp33_ASAP7_75t_L g385 ( .A(n_386), .B(n_387), .C(n_392), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_388), .B(n_390), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_389), .B(n_415), .Y(n_501) );
INVx1_ASAP7_75t_L g488 ( .A(n_390), .Y(n_488) );
INVx2_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_394), .B(n_395), .Y(n_393) );
OR2x6_ASAP7_75t_L g454 ( .A(n_394), .B(n_455), .Y(n_454) );
INVx2_ASAP7_75t_L g442 ( .A(n_395), .Y(n_442) );
OAI22xp33_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_402), .B1(n_406), .B2(n_407), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx2_ASAP7_75t_L g460 ( .A(n_401), .Y(n_460) );
INVx2_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx2_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
AOI21xp33_ASAP7_75t_L g422 ( .A1(n_406), .A2(n_423), .B(n_424), .Y(n_422) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
OR2x2_ASAP7_75t_L g470 ( .A(n_409), .B(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx2_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx2_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
OAI22xp5_ASAP7_75t_L g474 ( .A1(n_427), .A2(n_475), .B1(n_479), .B2(n_481), .Y(n_474) );
INVx2_ASAP7_75t_SL g443 ( .A(n_428), .Y(n_443) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
NAND2xp5_ASAP7_75t_SL g433 ( .A(n_434), .B(n_435), .Y(n_433) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
OAI22xp5_ASAP7_75t_L g438 ( .A1(n_439), .A2(n_442), .B1(n_443), .B2(n_444), .Y(n_438) );
BUFx2_ASAP7_75t_L g493 ( .A(n_441), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_445), .B(n_446), .Y(n_444) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
NOR2xp67_ASAP7_75t_L g448 ( .A(n_449), .B(n_482), .Y(n_448) );
NAND4xp25_ASAP7_75t_SL g449 ( .A(n_450), .B(n_456), .C(n_468), .D(n_474), .Y(n_449) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g473 ( .A(n_455), .Y(n_473) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
OR2x2_ASAP7_75t_L g462 ( .A(n_463), .B(n_464), .Y(n_462) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx3_ASAP7_75t_L g484 ( .A(n_470), .Y(n_484) );
NOR2xp33_ASAP7_75t_L g475 ( .A(n_476), .B(n_478), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx2_ASAP7_75t_L g489 ( .A(n_480), .Y(n_489) );
NAND3xp33_ASAP7_75t_L g482 ( .A(n_483), .B(n_496), .C(n_503), .Y(n_482) );
AOI22xp5_ASAP7_75t_L g483 ( .A1(n_484), .A2(n_485), .B1(n_490), .B2(n_492), .Y(n_483) );
INVxp67_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
NOR2xp67_ASAP7_75t_L g487 ( .A(n_488), .B(n_489), .Y(n_487) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
AND2x2_ASAP7_75t_L g492 ( .A(n_493), .B(n_494), .Y(n_492) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
NOR2xp67_ASAP7_75t_L g500 ( .A(n_501), .B(n_502), .Y(n_500) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g858 ( .A(n_511), .Y(n_858) );
BUFx8_ASAP7_75t_SL g511 ( .A(n_512), .Y(n_511) );
AND2x4_ASAP7_75t_L g513 ( .A(n_514), .B(n_766), .Y(n_513) );
NOR4xp25_ASAP7_75t_L g514 ( .A(n_515), .B(n_663), .C(n_707), .D(n_726), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_516), .B(n_648), .Y(n_515) );
AOI222xp33_ASAP7_75t_L g516 ( .A1(n_517), .A2(n_554), .B1(n_589), .B2(n_614), .C1(n_629), .C2(n_638), .Y(n_516) );
AOI221xp5_ASAP7_75t_L g845 ( .A1(n_517), .A2(n_671), .B1(n_791), .B2(n_846), .C(n_848), .Y(n_845) );
AND2x2_ASAP7_75t_L g517 ( .A(n_518), .B(n_532), .Y(n_517) );
BUFx2_ASAP7_75t_L g782 ( .A(n_518), .Y(n_782) );
INVx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
AND2x4_ASAP7_75t_L g682 ( .A(n_519), .B(n_667), .Y(n_682) );
AND2x4_ASAP7_75t_L g760 ( .A(n_519), .B(n_761), .Y(n_760) );
AND2x2_ASAP7_75t_L g817 ( .A(n_519), .B(n_757), .Y(n_817) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx2_ASAP7_75t_L g643 ( .A(n_521), .Y(n_643) );
HB1xp67_ASAP7_75t_L g763 ( .A(n_521), .Y(n_763) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
AND2x2_ASAP7_75t_L g722 ( .A(n_532), .B(n_723), .Y(n_722) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVxp67_ASAP7_75t_SL g785 ( .A(n_533), .Y(n_785) );
NAND2x1p5_ASAP7_75t_L g533 ( .A(n_534), .B(n_544), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
OR2x2_ASAP7_75t_L g733 ( .A(n_535), .B(n_645), .Y(n_733) );
AND2x2_ASAP7_75t_L g790 ( .A(n_535), .B(n_645), .Y(n_790) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_535), .B(n_698), .Y(n_799) );
INVx1_ASAP7_75t_L g615 ( .A(n_544), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_544), .B(n_643), .Y(n_686) );
INVx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
AND2x2_ASAP7_75t_L g674 ( .A(n_545), .B(n_651), .Y(n_674) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g764 ( .A(n_556), .B(n_765), .Y(n_764) );
AND2x2_ASAP7_75t_L g809 ( .A(n_556), .B(n_810), .Y(n_809) );
AND2x2_ASAP7_75t_L g556 ( .A(n_557), .B(n_572), .Y(n_556) );
AND2x2_ASAP7_75t_L g655 ( .A(n_557), .B(n_613), .Y(n_655) );
OR2x2_ASAP7_75t_L g662 ( .A(n_557), .B(n_591), .Y(n_662) );
AND2x2_ASAP7_75t_L g815 ( .A(n_557), .B(n_601), .Y(n_815) );
AO21x2_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_559), .B(n_571), .Y(n_557) );
INVx3_ASAP7_75t_L g575 ( .A(n_558), .Y(n_575) );
AO21x2_ASAP7_75t_L g636 ( .A1(n_558), .A2(n_559), .B(n_571), .Y(n_636) );
NOR2xp33_ASAP7_75t_SL g568 ( .A(n_569), .B(n_570), .Y(n_568) );
NOR2xp33_ASAP7_75t_L g578 ( .A(n_569), .B(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g613 ( .A(n_572), .Y(n_613) );
AND2x2_ASAP7_75t_L g715 ( .A(n_572), .B(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g794 ( .A(n_572), .Y(n_794) );
INVx2_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g633 ( .A(n_573), .Y(n_633) );
AOI21x1_ASAP7_75t_L g573 ( .A1(n_574), .A2(n_576), .B(n_588), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_577), .B(n_583), .Y(n_576) );
INVx2_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx2_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
AOI221xp5_ASAP7_75t_L g727 ( .A1(n_589), .A2(n_728), .B1(n_730), .B2(n_734), .C(n_739), .Y(n_727) );
AND2x2_ASAP7_75t_L g589 ( .A(n_590), .B(n_611), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_590), .B(n_745), .Y(n_744) );
NAND2xp67_ASAP7_75t_L g781 ( .A(n_590), .B(n_655), .Y(n_781) );
AND2x4_ASAP7_75t_L g836 ( .A(n_590), .B(n_715), .Y(n_836) );
AND2x2_ASAP7_75t_L g590 ( .A(n_591), .B(n_600), .Y(n_590) );
INVx1_ASAP7_75t_L g637 ( .A(n_591), .Y(n_637) );
HB1xp67_ASAP7_75t_L g658 ( .A(n_591), .Y(n_658) );
INVx1_ASAP7_75t_L g703 ( .A(n_591), .Y(n_703) );
INVx1_ASAP7_75t_L g752 ( .A(n_591), .Y(n_752) );
AND2x2_ASAP7_75t_L g793 ( .A(n_591), .B(n_794), .Y(n_793) );
NOR2xp33_ASAP7_75t_L g693 ( .A(n_600), .B(n_636), .Y(n_693) );
OR2x2_ASAP7_75t_L g751 ( .A(n_600), .B(n_752), .Y(n_751) );
BUFx3_ASAP7_75t_L g840 ( .A(n_600), .Y(n_840) );
INVx2_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx2_ASAP7_75t_L g634 ( .A(n_601), .Y(n_634) );
AOI22xp33_ASAP7_75t_SL g841 ( .A1(n_611), .A2(n_682), .B1(n_842), .B2(n_843), .Y(n_841) );
INVx2_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g800 ( .A(n_612), .B(n_736), .Y(n_800) );
OR2x2_ASAP7_75t_L g844 ( .A(n_612), .B(n_662), .Y(n_844) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
AOI22xp5_ASAP7_75t_L g648 ( .A1(n_614), .A2(n_649), .B1(n_654), .B2(n_659), .Y(n_648) );
AND2x2_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
OR2x2_ASAP7_75t_L g826 ( .A(n_615), .B(n_742), .Y(n_826) );
BUFx3_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx2_ASAP7_75t_L g720 ( .A(n_617), .Y(n_720) );
AND2x2_ASAP7_75t_L g617 ( .A(n_618), .B(n_619), .Y(n_617) );
INVx1_ASAP7_75t_L g698 ( .A(n_618), .Y(n_698) );
OR2x2_ASAP7_75t_L g711 ( .A(n_618), .B(n_652), .Y(n_711) );
AND2x2_ASAP7_75t_L g808 ( .A(n_618), .B(n_645), .Y(n_808) );
BUFx2_ASAP7_75t_L g743 ( .A(n_619), .Y(n_743) );
OAI21x1_ASAP7_75t_L g620 ( .A1(n_621), .A2(n_624), .B(n_627), .Y(n_620) );
INVx2_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
OR2x2_ASAP7_75t_L g630 ( .A(n_631), .B(n_635), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_632), .B(n_634), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_632), .B(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g661 ( .A(n_633), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_633), .B(n_634), .Y(n_689) );
INVxp67_ASAP7_75t_SL g746 ( .A(n_633), .Y(n_746) );
OR2x2_ASAP7_75t_L g657 ( .A(n_634), .B(n_658), .Y(n_657) );
INVx2_ASAP7_75t_L g737 ( .A(n_634), .Y(n_737) );
AND2x2_ASAP7_75t_L g787 ( .A(n_634), .B(n_703), .Y(n_787) );
NAND2xp5_ASAP7_75t_L g812 ( .A(n_634), .B(n_738), .Y(n_812) );
OR2x2_ASAP7_75t_L g688 ( .A(n_635), .B(n_689), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_636), .B(n_637), .Y(n_635) );
INVx1_ASAP7_75t_L g705 ( .A(n_636), .Y(n_705) );
INVx2_ASAP7_75t_SL g716 ( .A(n_636), .Y(n_716) );
INVx1_ASAP7_75t_L g772 ( .A(n_637), .Y(n_772) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
OR2x2_ASAP7_75t_L g639 ( .A(n_640), .B(n_642), .Y(n_639) );
OR2x2_ASAP7_75t_L g824 ( .A(n_640), .B(n_699), .Y(n_824) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx2_ASAP7_75t_SL g670 ( .A(n_641), .Y(n_670) );
INVx1_ASAP7_75t_SL g681 ( .A(n_641), .Y(n_681) );
BUFx2_ASAP7_75t_L g830 ( .A(n_641), .Y(n_830) );
NAND2xp5_ASAP7_75t_L g834 ( .A(n_642), .B(n_835), .Y(n_834) );
NAND2x1_ASAP7_75t_L g642 ( .A(n_643), .B(n_644), .Y(n_642) );
AND2x4_ASAP7_75t_SL g666 ( .A(n_643), .B(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g723 ( .A(n_643), .Y(n_723) );
BUFx2_ASAP7_75t_L g731 ( .A(n_643), .Y(n_731) );
INVx1_ASAP7_75t_L g779 ( .A(n_644), .Y(n_779) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_645), .B(n_651), .Y(n_650) );
OR2x2_ASAP7_75t_L g669 ( .A(n_645), .B(n_670), .Y(n_669) );
INVx2_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
AND2x2_ASAP7_75t_L g761 ( .A(n_646), .B(n_652), .Y(n_761) );
INVx2_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
AND2x2_ASAP7_75t_L g757 ( .A(n_647), .B(n_652), .Y(n_757) );
AND2x2_ASAP7_75t_L g706 ( .A(n_649), .B(n_673), .Y(n_706) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
OR2x2_ASAP7_75t_L g762 ( .A(n_650), .B(n_763), .Y(n_762) );
INVx2_ASAP7_75t_L g667 ( .A(n_651), .Y(n_667) );
INVx2_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx2_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
AOI22xp5_ASAP7_75t_L g768 ( .A1(n_654), .A2(n_672), .B1(n_769), .B2(n_774), .Y(n_768) );
AND2x4_ASAP7_75t_L g654 ( .A(n_655), .B(n_656), .Y(n_654) );
INVx1_ASAP7_75t_L g724 ( .A(n_655), .Y(n_724) );
INVx1_ASAP7_75t_L g857 ( .A(n_655), .Y(n_857) );
INVx1_ASAP7_75t_L g803 ( .A(n_656), .Y(n_803) );
INVx2_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx2_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
OAI211xp5_ASAP7_75t_L g663 ( .A1(n_660), .A2(n_664), .B(n_675), .C(n_690), .Y(n_663) );
OR2x2_ASAP7_75t_L g660 ( .A(n_661), .B(n_662), .Y(n_660) );
INVx1_ASAP7_75t_L g821 ( .A(n_661), .Y(n_821) );
INVx2_ASAP7_75t_L g738 ( .A(n_662), .Y(n_738) );
INVxp67_ASAP7_75t_SL g664 ( .A(n_665), .Y(n_664) );
AO21x1_ASAP7_75t_L g665 ( .A1(n_666), .A2(n_668), .B(n_671), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_666), .B(n_678), .Y(n_677) );
INVx2_ASAP7_75t_L g729 ( .A(n_666), .Y(n_729) );
INVx1_ASAP7_75t_L g807 ( .A(n_667), .Y(n_807) );
BUFx2_ASAP7_75t_L g842 ( .A(n_667), .Y(n_842) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
NOR2x1_ASAP7_75t_SL g719 ( .A(n_669), .B(n_720), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_670), .B(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g750 ( .A(n_670), .Y(n_750) );
AND2x2_ASAP7_75t_L g671 ( .A(n_672), .B(n_674), .Y(n_671) );
OR2x6_ASAP7_75t_SL g710 ( .A(n_672), .B(n_711), .Y(n_710) );
NOR2xp33_ASAP7_75t_L g728 ( .A(n_672), .B(n_729), .Y(n_728) );
INVx2_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx2_ASAP7_75t_L g678 ( .A(n_673), .Y(n_678) );
INVx2_ASAP7_75t_L g699 ( .A(n_674), .Y(n_699) );
OAI31xp33_ASAP7_75t_L g675 ( .A1(n_676), .A2(n_679), .A3(n_683), .B(n_687), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
AND2x2_ASAP7_75t_L g839 ( .A(n_678), .B(n_840), .Y(n_839) );
AND2x2_ASAP7_75t_L g679 ( .A(n_680), .B(n_682), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
NOR2x1p5_ASAP7_75t_L g804 ( .A(n_681), .B(n_759), .Y(n_804) );
INVx2_ASAP7_75t_L g773 ( .A(n_682), .Y(n_773) );
INVxp67_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx2_ASAP7_75t_SL g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g847 ( .A(n_689), .Y(n_847) );
AOI22xp33_ASAP7_75t_SL g690 ( .A1(n_691), .A2(n_694), .B1(n_700), .B2(n_706), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
OR2x2_ASAP7_75t_L g831 ( .A(n_692), .B(n_702), .Y(n_831) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
AOI21xp5_ASAP7_75t_L g739 ( .A1(n_695), .A2(n_740), .B(n_744), .Y(n_739) );
OR2x2_ASAP7_75t_L g695 ( .A(n_696), .B(n_699), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_696), .B(n_776), .Y(n_775) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
AND2x2_ASAP7_75t_SL g756 ( .A(n_697), .B(n_757), .Y(n_756) );
BUFx2_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_702), .B(n_704), .Y(n_701) );
INVx1_ASAP7_75t_L g725 ( .A(n_702), .Y(n_725) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
BUFx2_ASAP7_75t_SL g704 ( .A(n_705), .Y(n_704) );
AND2x2_ASAP7_75t_L g792 ( .A(n_705), .B(n_793), .Y(n_792) );
O2A1O1Ixp5_ASAP7_75t_L g707 ( .A1(n_708), .A2(n_712), .B(n_717), .C(n_725), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVxp67_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_710), .B(n_775), .Y(n_774) );
OR2x2_ASAP7_75t_L g849 ( .A(n_711), .B(n_750), .Y(n_849) );
OAI21xp5_ASAP7_75t_L g851 ( .A1(n_711), .A2(n_852), .B(n_854), .Y(n_851) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
AND2x2_ASAP7_75t_L g771 ( .A(n_715), .B(n_772), .Y(n_771) );
HB1xp67_ASAP7_75t_L g755 ( .A(n_716), .Y(n_755) );
AO21x1_ASAP7_75t_L g717 ( .A1(n_718), .A2(n_721), .B(n_724), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
OAI22xp5_ASAP7_75t_L g769 ( .A1(n_720), .A2(n_724), .B1(n_770), .B2(n_773), .Y(n_769) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
OAI21xp5_ASAP7_75t_L g796 ( .A1(n_722), .A2(n_797), .B(n_800), .Y(n_796) );
AND2x2_ASAP7_75t_L g789 ( .A(n_723), .B(n_790), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_727), .B(n_747), .Y(n_726) );
AND2x2_ASAP7_75t_L g730 ( .A(n_731), .B(n_732), .Y(n_730) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g833 ( .A(n_733), .Y(n_833) );
INVx2_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx3_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
AND2x4_ASAP7_75t_L g736 ( .A(n_737), .B(n_738), .Y(n_736) );
AND2x4_ASAP7_75t_L g791 ( .A(n_737), .B(n_792), .Y(n_791) );
OR2x2_ASAP7_75t_L g856 ( .A(n_737), .B(n_857), .Y(n_856) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g835 ( .A(n_743), .Y(n_835) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
AOI32xp33_ASAP7_75t_L g747 ( .A1(n_748), .A2(n_753), .A3(n_756), .B1(n_758), .B2(n_764), .Y(n_747) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
OR2x2_ASAP7_75t_L g749 ( .A(n_750), .B(n_751), .Y(n_749) );
INVx1_ASAP7_75t_L g776 ( .A(n_750), .Y(n_776) );
INVx1_ASAP7_75t_L g765 ( .A(n_751), .Y(n_765) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_754), .B(n_787), .Y(n_786) );
INVx2_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
OAI21xp33_ASAP7_75t_L g854 ( .A1(n_756), .A2(n_809), .B(n_855), .Y(n_854) );
AND2x2_ASAP7_75t_L g829 ( .A(n_757), .B(n_830), .Y(n_829) );
NAND2xp33_ASAP7_75t_SL g758 ( .A(n_759), .B(n_762), .Y(n_758) );
INVx3_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
NOR4xp75_ASAP7_75t_L g766 ( .A(n_767), .B(n_795), .C(n_837), .D(n_851), .Y(n_766) );
NAND3xp33_ASAP7_75t_L g767 ( .A(n_768), .B(n_777), .C(n_788), .Y(n_767) );
INVx1_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
INVx1_ASAP7_75t_L g810 ( .A(n_772), .Y(n_810) );
A2O1A1Ixp33_ASAP7_75t_L g777 ( .A1(n_778), .A2(n_780), .B(n_782), .C(n_783), .Y(n_777) );
INVx1_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
INVx1_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
OAI21xp5_ASAP7_75t_L g783 ( .A1(n_782), .A2(n_784), .B(n_786), .Y(n_783) );
INVx1_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
INVx1_ASAP7_75t_L g822 ( .A(n_787), .Y(n_822) );
NAND2x1_ASAP7_75t_L g788 ( .A(n_789), .B(n_791), .Y(n_788) );
AND2x4_ASAP7_75t_L g814 ( .A(n_793), .B(n_815), .Y(n_814) );
NAND4xp75_ASAP7_75t_L g795 ( .A(n_796), .B(n_801), .C(n_818), .D(n_827), .Y(n_795) );
INVx1_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
HB1xp67_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
AOI211x1_ASAP7_75t_L g801 ( .A1(n_802), .A2(n_804), .B(n_805), .C(n_811), .Y(n_801) );
AOI22xp5_ASAP7_75t_L g818 ( .A1(n_802), .A2(n_819), .B1(n_823), .B2(n_825), .Y(n_818) );
INVx1_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
NOR3xp33_ASAP7_75t_L g848 ( .A(n_803), .B(n_849), .C(n_850), .Y(n_848) );
AND2x2_ASAP7_75t_L g805 ( .A(n_806), .B(n_809), .Y(n_805) );
AND2x4_ASAP7_75t_L g806 ( .A(n_807), .B(n_808), .Y(n_806) );
AOI21xp5_ASAP7_75t_L g811 ( .A1(n_812), .A2(n_813), .B(n_816), .Y(n_811) );
NOR2xp67_ASAP7_75t_L g853 ( .A(n_813), .B(n_830), .Y(n_853) );
INVx2_ASAP7_75t_SL g813 ( .A(n_814), .Y(n_813) );
INVx2_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
INVx2_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
OR2x2_ASAP7_75t_L g820 ( .A(n_821), .B(n_822), .Y(n_820) );
INVx1_ASAP7_75t_L g850 ( .A(n_821), .Y(n_850) );
INVx1_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
INVx1_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
OA21x2_ASAP7_75t_L g827 ( .A1(n_828), .A2(n_831), .B(n_832), .Y(n_827) );
INVx1_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
OAI21xp5_ASAP7_75t_L g832 ( .A1(n_833), .A2(n_834), .B(n_836), .Y(n_832) );
OAI21xp5_ASAP7_75t_L g837 ( .A1(n_838), .A2(n_841), .B(n_845), .Y(n_837) );
INVx1_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
INVx2_ASAP7_75t_L g843 ( .A(n_844), .Y(n_843) );
HB1xp67_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
INVxp67_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
INVx1_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
INVx2_ASAP7_75t_SL g859 ( .A(n_860), .Y(n_859) );
AOI21xp5_ASAP7_75t_L g864 ( .A1(n_865), .A2(n_869), .B(n_876), .Y(n_864) );
CKINVDCx5p33_ASAP7_75t_R g865 ( .A(n_866), .Y(n_865) );
CKINVDCx5p33_ASAP7_75t_R g866 ( .A(n_867), .Y(n_866) );
CKINVDCx5p33_ASAP7_75t_R g867 ( .A(n_868), .Y(n_867) );
OAI21xp5_ASAP7_75t_L g869 ( .A1(n_870), .A2(n_871), .B(n_875), .Y(n_869) );
NOR2xp33_ASAP7_75t_L g876 ( .A(n_877), .B(n_878), .Y(n_876) );
BUFx12f_ASAP7_75t_L g878 ( .A(n_879), .Y(n_878) );
endmodule