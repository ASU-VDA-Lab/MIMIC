module real_jpeg_6497_n_17 (n_108, n_8, n_0, n_111, n_2, n_10, n_9, n_12, n_107, n_6, n_104, n_106, n_11, n_14, n_110, n_7, n_3, n_5, n_4, n_102, n_105, n_109, n_1, n_16, n_15, n_13, n_103, n_17);

input n_108;
input n_8;
input n_0;
input n_111;
input n_2;
input n_10;
input n_9;
input n_12;
input n_107;
input n_6;
input n_104;
input n_106;
input n_11;
input n_14;
input n_110;
input n_7;
input n_3;
input n_5;
input n_4;
input n_102;
input n_105;
input n_109;
input n_1;
input n_16;
input n_15;
input n_13;
input n_103;

output n_17;

wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_78;
wire n_83;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_85;
wire n_96;
wire n_89;

INVx5_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_0),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_0),
.B(n_73),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_2),
.B(n_55),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_2),
.B(n_55),
.Y(n_82)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_3),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_4),
.B(n_30),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_4),
.B(n_30),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_5),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_5),
.B(n_45),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_6),
.B(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_6),
.B(n_77),
.Y(n_79)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_7),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

OR2x2_ASAP7_75t_L g19 ( 
.A(n_9),
.B(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_9),
.B(n_20),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_10),
.B(n_36),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_10),
.B(n_36),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_11),
.B(n_58),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_11),
.B(n_58),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_12),
.B(n_69),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_13),
.B(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_13),
.B(n_90),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_14),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_15),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_16),
.B(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_16),
.B(n_42),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_26),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_25),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_22),
.Y(n_20)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_22),
.B(n_86),
.Y(n_85)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_49),
.B(n_93),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NOR4xp25_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_35),
.C(n_41),
.D(n_44),
.Y(n_28)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_29),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_32),
.Y(n_30)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_34),
.B(n_59),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_34),
.B(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_35),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_38),
.Y(n_36)
);

BUFx8_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_39),
.B(n_43),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_56),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_40),
.B(n_70),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_41),
.A2(n_96),
.B(n_97),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_47),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_47),
.B(n_91),
.Y(n_90)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_89),
.B(n_92),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_84),
.B(n_88),
.Y(n_51)
);

AO221x1_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_60),
.B1(n_81),
.B2(n_82),
.C(n_83),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_57),
.Y(n_53)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

AO21x1_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_66),
.B(n_80),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_62),
.B(n_65),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_65),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_64),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_SL g66 ( 
.A1(n_67),
.A2(n_76),
.B(n_79),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_71),
.B(n_75),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_72),
.B(n_74),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_72),
.B(n_74),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_85),
.B(n_87),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_85),
.B(n_87),
.Y(n_88)
);

A2O1A1O1Ixp25_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_95),
.B(n_98),
.C(n_99),
.D(n_100),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_102),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_103),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_104),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_105),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_106),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_107),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_108),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_109),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_110),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_111),
.Y(n_91)
);


endmodule