module fake_jpeg_25487_n_276 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_276);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_276;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_57;
wire n_21;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_240;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx2_ASAP7_75t_R g15 ( 
.A(n_14),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

INVx11_ASAP7_75t_SL g30 ( 
.A(n_4),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_35),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_15),
.B(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_23),
.B(n_0),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_40),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_15),
.B(n_7),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_39),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

BUFx12f_ASAP7_75t_SL g39 ( 
.A(n_30),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_23),
.B(n_0),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_36),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_42),
.Y(n_67)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_15),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_48),
.B(n_50),
.Y(n_66)
);

BUFx10_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_15),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_23),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_51),
.B(n_55),
.Y(n_58)
);

CKINVDCx14_ASAP7_75t_R g54 ( 
.A(n_39),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_54),
.A2(n_24),
.B1(n_18),
.B2(n_28),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_17),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_34),
.A2(n_20),
.B1(n_19),
.B2(n_30),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_56),
.A2(n_34),
.B1(n_20),
.B2(n_31),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_23),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_33),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_59),
.A2(n_60),
.B1(n_68),
.B2(n_71),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_42),
.A2(n_31),
.B1(n_34),
.B2(n_19),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_62),
.Y(n_89)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_63),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_64),
.B(n_70),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_42),
.A2(n_57),
.B1(n_51),
.B2(n_55),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_49),
.A2(n_20),
.B1(n_19),
.B2(n_29),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_23),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_41),
.A2(n_57),
.B1(n_51),
.B2(n_44),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_72),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_56),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_73),
.Y(n_84)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_74),
.B(n_77),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_44),
.A2(n_16),
.B1(n_22),
.B2(n_28),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_75),
.A2(n_26),
.B1(n_22),
.B2(n_16),
.Y(n_105)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_76),
.B(n_78),
.Y(n_91)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_80),
.A2(n_82),
.B(n_48),
.Y(n_103)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_81),
.B(n_18),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_44),
.A2(n_16),
.B(n_22),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_73),
.A2(n_54),
.B1(n_53),
.B2(n_52),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_86),
.A2(n_94),
.B1(n_100),
.B2(n_65),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_79),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_90),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_80),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_92),
.B(n_97),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_60),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_93),
.B(n_96),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_74),
.A2(n_53),
.B1(n_52),
.B2(n_50),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_66),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_67),
.Y(n_97)
);

BUFx8_ASAP7_75t_L g99 ( 
.A(n_62),
.Y(n_99)
);

BUFx24_ASAP7_75t_L g129 ( 
.A(n_99),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_67),
.A2(n_53),
.B1(n_52),
.B2(n_49),
.Y(n_100)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_61),
.Y(n_101)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_101),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_64),
.B(n_33),
.C(n_32),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_102),
.B(n_33),
.C(n_72),
.Y(n_110)
);

AO21x1_ASAP7_75t_L g122 ( 
.A1(n_103),
.A2(n_24),
.B(n_29),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_66),
.B(n_49),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_104),
.B(n_108),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_105),
.A2(n_107),
.B1(n_65),
.B2(n_81),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_58),
.A2(n_47),
.B1(n_46),
.B2(n_49),
.Y(n_107)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_101),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_109),
.B(n_113),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_110),
.B(n_130),
.C(n_102),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_111),
.A2(n_124),
.B1(n_89),
.B2(n_88),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_97),
.B(n_58),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_112),
.B(n_126),
.Y(n_138)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_91),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_114),
.B(n_120),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_70),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_SL g139 ( 
.A(n_115),
.B(n_128),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_87),
.A2(n_82),
.B(n_77),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_116),
.A2(n_117),
.B(n_118),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_87),
.A2(n_75),
.B(n_49),
.Y(n_117)
);

HAxp5_ASAP7_75t_SL g118 ( 
.A(n_106),
.B(n_27),
.CON(n_118),
.SN(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_106),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_122),
.B(n_17),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_93),
.A2(n_63),
.B1(n_78),
.B2(n_76),
.Y(n_124)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_99),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_125),
.B(n_129),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_98),
.B(n_33),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_96),
.B(n_23),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_127),
.B(n_38),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_SL g128 ( 
.A(n_103),
.B(n_25),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_85),
.B(n_21),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_84),
.A2(n_0),
.B(n_47),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_132),
.Y(n_134)
);

AND2x6_ASAP7_75t_L g135 ( 
.A(n_128),
.B(n_85),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_135),
.B(n_157),
.Y(n_162)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_124),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_136),
.B(n_148),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_141),
.B(n_38),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_110),
.B(n_107),
.C(n_104),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_142),
.B(n_144),
.C(n_130),
.Y(n_172)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_121),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_143),
.B(n_147),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_115),
.B(n_94),
.C(n_95),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_111),
.A2(n_84),
.B1(n_105),
.B2(n_95),
.Y(n_145)
);

OAI21xp33_ASAP7_75t_SL g174 ( 
.A1(n_145),
.A2(n_117),
.B(n_118),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_123),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_146),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_112),
.A2(n_86),
.B1(n_100),
.B2(n_90),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_126),
.Y(n_148)
);

O2A1O1Ixp33_ASAP7_75t_L g150 ( 
.A1(n_132),
.A2(n_88),
.B(n_83),
.C(n_89),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_150),
.A2(n_131),
.B(n_99),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_151),
.B(n_152),
.Y(n_171)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_127),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_119),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_153),
.B(n_154),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g154 ( 
.A(n_133),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_155),
.B(n_114),
.Y(n_173)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_156),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_125),
.B(n_83),
.Y(n_157)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_158),
.Y(n_166)
);

CKINVDCx10_ASAP7_75t_R g159 ( 
.A(n_129),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_159),
.B(n_160),
.Y(n_169)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_119),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_137),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_161),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_158),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_165),
.B(n_181),
.Y(n_189)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_138),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_167),
.B(n_175),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_139),
.B(n_116),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_168),
.B(n_184),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_172),
.B(n_185),
.C(n_186),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_173),
.A2(n_174),
.B1(n_150),
.B2(n_140),
.Y(n_194)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_138),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_143),
.B(n_129),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_176),
.B(n_178),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_147),
.B(n_131),
.Y(n_178)
);

OA21x2_ASAP7_75t_L g206 ( 
.A1(n_179),
.A2(n_142),
.B(n_159),
.Y(n_206)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_155),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_180),
.B(n_145),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_153),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_134),
.A2(n_122),
.B(n_29),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_183),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_139),
.B(n_99),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_141),
.B(n_38),
.Y(n_185)
);

OA21x2_ASAP7_75t_SL g187 ( 
.A1(n_161),
.A2(n_171),
.B(n_168),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_187),
.B(n_201),
.Y(n_209)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_190),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_182),
.A2(n_180),
.B1(n_162),
.B2(n_134),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_192),
.A2(n_28),
.B1(n_26),
.B2(n_25),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_185),
.B(n_172),
.C(n_186),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_193),
.B(n_184),
.C(n_166),
.Y(n_211)
);

CKINVDCx14_ASAP7_75t_R g217 ( 
.A(n_194),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_173),
.A2(n_148),
.B1(n_149),
.B2(n_152),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_195),
.A2(n_179),
.B1(n_166),
.B2(n_173),
.Y(n_210)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_177),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_196),
.B(n_202),
.Y(n_213)
);

NAND3xp33_ASAP7_75t_L g201 ( 
.A(n_163),
.B(n_135),
.C(n_140),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_169),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_167),
.B(n_175),
.Y(n_203)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_203),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_170),
.B(n_144),
.Y(n_204)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_204),
.Y(n_222)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_182),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_205),
.B(n_207),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_206),
.A2(n_183),
.B(n_164),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_164),
.B(n_17),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_210),
.A2(n_219),
.B1(n_199),
.B2(n_200),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_211),
.B(n_221),
.C(n_197),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_215),
.A2(n_206),
.B(n_190),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_216),
.A2(n_220),
.B1(n_199),
.B2(n_202),
.Y(n_227)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_206),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_218),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_196),
.A2(n_26),
.B1(n_2),
.B2(n_3),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_205),
.A2(n_32),
.B1(n_21),
.B2(n_3),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_191),
.B(n_32),
.C(n_25),
.Y(n_221)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_189),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_223),
.A2(n_198),
.B1(n_192),
.B2(n_195),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_214),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_224),
.B(n_223),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_225),
.A2(n_231),
.B1(n_232),
.B2(n_216),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_226),
.B(n_229),
.Y(n_238)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_227),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_221),
.B(n_191),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_228),
.B(n_213),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_211),
.B(n_193),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_215),
.B(n_204),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_233),
.B(n_234),
.C(n_236),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_222),
.B(n_197),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_209),
.A2(n_198),
.B(n_203),
.Y(n_235)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_235),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_222),
.B(n_188),
.C(n_194),
.Y(n_236)
);

OR2x2_ASAP7_75t_L g254 ( 
.A(n_239),
.B(n_240),
.Y(n_254)
);

FAx1_ASAP7_75t_L g240 ( 
.A(n_230),
.B(n_218),
.CI(n_217),
.CON(n_240),
.SN(n_240)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_229),
.B(n_212),
.C(n_213),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_243),
.B(n_244),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_236),
.B(n_214),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_245),
.A2(n_188),
.B1(n_226),
.B2(n_25),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_246),
.B(n_247),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_233),
.B(n_208),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_242),
.A2(n_232),
.B1(n_230),
.B2(n_212),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_248),
.A2(n_252),
.B1(n_256),
.B2(n_1),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_237),
.B(n_234),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_250),
.B(n_255),
.Y(n_257)
);

NOR2x1_ASAP7_75t_L g252 ( 
.A(n_240),
.B(n_220),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_253),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_241),
.A2(n_240),
.B(n_243),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_237),
.A2(n_1),
.B1(n_2),
.B2(n_5),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_251),
.B(n_238),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_258),
.B(n_259),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_249),
.B(n_238),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_260),
.B(n_262),
.Y(n_264)
);

AOI322xp5_ASAP7_75t_L g262 ( 
.A1(n_252),
.A2(n_5),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.C1(n_9),
.C2(n_10),
.Y(n_262)
);

AOI322xp5_ASAP7_75t_L g263 ( 
.A1(n_254),
.A2(n_6),
.A3(n_8),
.B1(n_10),
.B2(n_11),
.C1(n_12),
.C2(n_13),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_263),
.B(n_254),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_265),
.B(n_268),
.Y(n_269)
);

NOR3xp33_ASAP7_75t_L g266 ( 
.A(n_261),
.B(n_250),
.C(n_10),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_266),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_257),
.A2(n_6),
.B(n_11),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_267),
.A2(n_261),
.B1(n_13),
.B2(n_12),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_271),
.B(n_264),
.Y(n_272)
);

OAI31xp33_ASAP7_75t_SL g274 ( 
.A1(n_272),
.A2(n_273),
.A3(n_25),
.B(n_21),
.Y(n_274)
);

MAJx2_ASAP7_75t_L g273 ( 
.A(n_269),
.B(n_270),
.C(n_13),
.Y(n_273)
);

OAI21x1_ASAP7_75t_L g275 ( 
.A1(n_274),
.A2(n_21),
.B(n_25),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_275),
.B(n_21),
.Y(n_276)
);


endmodule