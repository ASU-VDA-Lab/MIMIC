module fake_jpeg_25556_n_31 (n_3, n_2, n_1, n_0, n_4, n_5, n_31);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_31;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_29;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

INVx6_ASAP7_75t_L g6 ( 
.A(n_0),
.Y(n_6)
);

BUFx5_ASAP7_75t_L g7 ( 
.A(n_5),
.Y(n_7)
);

INVx13_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

BUFx12f_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

BUFx4f_ASAP7_75t_SL g10 ( 
.A(n_3),
.Y(n_10)
);

BUFx12f_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_10),
.Y(n_12)
);

AOI22xp5_ASAP7_75t_L g13 ( 
.A1(n_6),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_13)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_13),
.A2(n_8),
.B1(n_10),
.B2(n_4),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g14 ( 
.A(n_11),
.B(n_0),
.C(n_2),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_15),
.B(n_16),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_9),
.B(n_2),
.Y(n_16)
);

INVx5_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_17),
.A2(n_18),
.B1(n_10),
.B2(n_7),
.Y(n_21)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_L g22 ( 
.A1(n_19),
.A2(n_16),
.B(n_14),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_21),
.B(n_9),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g26 ( 
.A1(n_22),
.A2(n_23),
.B(n_24),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_20),
.B(n_12),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_19),
.B(n_17),
.Y(n_25)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_15),
.C(n_24),
.Y(n_27)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

AO21x1_ASAP7_75t_L g30 ( 
.A1(n_29),
.A2(n_28),
.B(n_27),
.Y(n_30)
);

BUFx24_ASAP7_75t_SL g31 ( 
.A(n_30),
.Y(n_31)
);


endmodule