module real_jpeg_4563_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_372;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_148;
wire n_373;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_14;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx8_ASAP7_75t_L g57 ( 
.A(n_0),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_1),
.A2(n_25),
.B1(n_28),
.B2(n_29),
.Y(n_24)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_1),
.A2(n_28),
.B1(n_147),
.B2(n_149),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_1),
.A2(n_28),
.B1(n_54),
.B2(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_1),
.B(n_89),
.Y(n_232)
);

O2A1O1Ixp33_ASAP7_75t_L g255 ( 
.A1(n_1),
.A2(n_92),
.B(n_256),
.C(n_258),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_1),
.B(n_52),
.C(n_283),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_1),
.B(n_123),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_1),
.B(n_155),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_1),
.B(n_45),
.Y(n_321)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_3),
.A2(n_103),
.B1(n_105),
.B2(n_106),
.Y(n_102)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_3),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_3),
.A2(n_105),
.B1(n_218),
.B2(n_221),
.Y(n_217)
);

OAI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_3),
.A2(n_105),
.B1(n_269),
.B2(n_271),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_L g291 ( 
.A1(n_3),
.A2(n_105),
.B1(n_292),
.B2(n_294),
.Y(n_291)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_4),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_5),
.Y(n_155)
);

INVx8_ASAP7_75t_L g174 ( 
.A(n_5),
.Y(n_174)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_6),
.Y(n_91)
);

BUFx5_ASAP7_75t_L g113 ( 
.A(n_6),
.Y(n_113)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_6),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_7),
.A2(n_54),
.B1(n_58),
.B2(n_59),
.Y(n_53)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_7),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_7),
.A2(n_58),
.B1(n_165),
.B2(n_167),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_7),
.A2(n_58),
.B1(n_380),
.B2(n_384),
.Y(n_379)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_8),
.Y(n_95)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_9),
.Y(n_86)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_9),
.Y(n_88)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_9),
.Y(n_104)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_9),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_9),
.Y(n_111)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_9),
.Y(n_118)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_10),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_11),
.A2(n_38),
.B1(n_41),
.B2(n_42),
.Y(n_37)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_11),
.A2(n_41),
.B1(n_66),
.B2(n_68),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_11),
.A2(n_41),
.B1(n_93),
.B2(n_122),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_11),
.A2(n_41),
.B1(n_104),
.B2(n_111),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_360),
.Y(n_12)
);

OAI21xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_223),
.B(n_358),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_185),
.Y(n_14)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_15),
.B(n_185),
.Y(n_359)
);

BUFx24_ASAP7_75t_SL g391 ( 
.A(n_15),
.Y(n_391)
);

FAx1_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_150),
.CI(n_161),
.CON(n_15),
.SN(n_15)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_16),
.B(n_150),
.C(n_161),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_80),
.B2(n_81),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_17),
.B(n_82),
.C(n_119),
.Y(n_389)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_43),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_19),
.B(n_43),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_30),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_20),
.B(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_23),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_24),
.A2(n_32),
.B(n_152),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_24),
.B(n_32),
.Y(n_234)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_26),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_27),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_28),
.A2(n_85),
.B(n_87),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_28),
.B(n_88),
.Y(n_87)
);

OAI21xp33_ASAP7_75t_L g258 ( 
.A1(n_28),
.A2(n_259),
.B(n_261),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_30),
.B(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_31),
.A2(n_153),
.B(n_164),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_37),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_32),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_32),
.B(n_291),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_36),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_35),
.Y(n_169)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_35),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_37),
.B(n_172),
.Y(n_171)
);

BUFx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_39),
.Y(n_316)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

AO22x1_ASAP7_75t_SL g45 ( 
.A1(n_42),
.A2(n_46),
.B1(n_49),
.B2(n_51),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_53),
.B(n_64),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_44),
.A2(n_158),
.B(n_248),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_44),
.B(n_248),
.Y(n_266)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NOR2x1_ASAP7_75t_L g70 ( 
.A(n_45),
.B(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_45),
.B(n_65),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_45),
.B(n_268),
.Y(n_286)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx3_ASAP7_75t_SL g49 ( 
.A(n_50),
.Y(n_49)
);

INVx4_ASAP7_75t_SL g51 ( 
.A(n_52),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_52),
.A2(n_72),
.B1(n_74),
.B2(n_77),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_53),
.A2(n_158),
.B(n_159),
.Y(n_157)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

INVx6_ASAP7_75t_L g273 ( 
.A(n_56),
.Y(n_273)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g129 ( 
.A(n_57),
.Y(n_129)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_57),
.Y(n_270)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_62),
.Y(n_178)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g262 ( 
.A(n_63),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_64),
.B(n_286),
.Y(n_330)
);

INVxp67_ASAP7_75t_SL g387 ( 
.A(n_64),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_70),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_70),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_70),
.B(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_70),
.B(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_78),
.A2(n_125),
.B1(n_129),
.B2(n_130),
.Y(n_124)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx4_ASAP7_75t_L g281 ( 
.A(n_79),
.Y(n_281)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_119),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_101),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_84),
.B(n_89),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_84),
.B(n_109),
.Y(n_239)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_84),
.Y(n_375)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVxp33_ASAP7_75t_L g204 ( 
.A(n_87),
.Y(n_204)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_88),
.Y(n_203)
);

NOR2x1_ASAP7_75t_L g109 ( 
.A(n_89),
.B(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_89),
.B(n_102),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_89),
.B(n_183),
.Y(n_191)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_89),
.Y(n_373)
);

AO22x2_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_92),
.B1(n_96),
.B2(n_99),
.Y(n_89)
);

INVx6_ASAP7_75t_L g211 ( 
.A(n_90),
.Y(n_211)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_91),
.Y(n_100)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx5_ASAP7_75t_L g145 ( 
.A(n_94),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_94),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_94),
.Y(n_220)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_95),
.Y(n_98)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_95),
.Y(n_141)
);

BUFx5_ASAP7_75t_L g148 ( 
.A(n_95),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_95),
.Y(n_383)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_96),
.Y(n_122)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_101),
.B(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_109),
.Y(n_101)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_109),
.B(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_109),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_112),
.B1(n_114),
.B2(n_116),
.Y(n_110)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_113),
.Y(n_115)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_132),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_120),
.B(n_216),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_121),
.B(n_123),
.Y(n_120)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_121),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_123),
.A2(n_133),
.B(n_146),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_123),
.B(n_217),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g378 ( 
.A1(n_123),
.A2(n_243),
.B(n_379),
.Y(n_378)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_124),
.B(n_135),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_124),
.B(n_215),
.Y(n_214)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_127),
.Y(n_257)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_128),
.Y(n_131)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_128),
.Y(n_139)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_128),
.Y(n_260)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_132),
.B(n_245),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_133),
.B(n_146),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_133),
.B(n_217),
.Y(n_216)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_134),
.B(n_244),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_140),
.B1(n_142),
.B2(n_145),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_139),
.Y(n_144)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVxp67_ASAP7_75t_SL g215 ( 
.A(n_146),
.Y(n_215)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_147),
.Y(n_149)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx6_ASAP7_75t_L g209 ( 
.A(n_148),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_156),
.B1(n_157),
.B2(n_160),
.Y(n_150)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_151),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_151),
.B(n_255),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_151),
.A2(n_160),
.B1(n_255),
.B2(n_333),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_151),
.B(n_157),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_151),
.A2(n_160),
.B1(n_371),
.B2(n_372),
.Y(n_370)
);

INVx1_ASAP7_75t_SL g152 ( 
.A(n_153),
.Y(n_152)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

AND2x2_ASAP7_75t_SL g175 ( 
.A(n_159),
.B(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_159),
.B(n_267),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_179),
.C(n_181),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_162),
.B(n_187),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_175),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_163),
.B(n_175),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_170),
.B(n_171),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_167),
.Y(n_294)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx6_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

OR2x2_ASAP7_75t_L g233 ( 
.A(n_171),
.B(n_234),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_171),
.B(n_290),
.Y(n_320)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_174),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_176),
.B(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_177),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_179),
.A2(n_180),
.B1(n_181),
.B2(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_181),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_182),
.B(n_184),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_184),
.B(n_239),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_189),
.C(n_222),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_186),
.B(n_222),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_189),
.B(n_353),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_192),
.C(n_212),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_190),
.B(n_212),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_SL g349 ( 
.A(n_192),
.B(n_350),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_193),
.B(n_194),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_193),
.B(n_194),
.Y(n_236)
);

AOI32xp33_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_199),
.A3(n_202),
.B1(n_204),
.B2(n_205),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx4_ASAP7_75t_SL g196 ( 
.A(n_197),
.Y(n_196)
);

INVx5_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

NAND2xp33_ASAP7_75t_SL g205 ( 
.A(n_206),
.B(n_210),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_216),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_218),
.Y(n_221)
);

INVx6_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx5_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_220),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_342),
.B(n_355),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_274),
.B(n_341),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_226),
.B(n_250),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_226),
.B(n_250),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_237),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_228),
.A2(n_229),
.B1(n_235),
.B2(n_236),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_229),
.B(n_235),
.C(n_237),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.C(n_233),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_230),
.B(n_252),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_231),
.A2(n_232),
.B1(n_233),
.B2(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_233),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_234),
.B(n_306),
.Y(n_318)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_238),
.B(n_240),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_238),
.B(n_241),
.C(n_247),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_246),
.B1(n_247),
.B2(n_249),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_241),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_242),
.B(n_245),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_254),
.C(n_263),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_251),
.B(n_337),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_254),
.A2(n_263),
.B1(n_264),
.B2(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_254),
.Y(n_338)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_255),
.Y(n_333)
);

INVx8_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx6_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_267),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_266),
.B(n_387),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx5_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_335),
.B(n_340),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_276),
.A2(n_325),
.B(n_334),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_300),
.B(n_324),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_287),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_278),
.B(n_287),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_285),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_279),
.A2(n_280),
.B1(n_285),
.B2(n_303),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_280),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_285),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_295),
.Y(n_287)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_288),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_291),
.B(n_307),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_296),
.A2(n_297),
.B1(n_298),
.B2(n_299),
.Y(n_295)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_296),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_297),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_297),
.B(n_298),
.C(n_327),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_301),
.A2(n_309),
.B(n_323),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_302),
.B(n_304),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_302),
.B(n_304),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx4_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_310),
.A2(n_319),
.B(n_322),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_318),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_317),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_SL g313 ( 
.A(n_314),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_320),
.B(n_321),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_320),
.B(n_321),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_328),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_326),
.B(n_328),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_332),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_331),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_330),
.B(n_331),
.C(n_332),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_336),
.B(n_339),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_336),
.B(n_339),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_351),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_345),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_344),
.B(n_345),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_349),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_348),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_347),
.B(n_348),
.C(n_349),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_L g355 ( 
.A1(n_351),
.A2(n_356),
.B(n_357),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_SL g351 ( 
.A(n_352),
.B(n_354),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_352),
.B(n_354),
.Y(n_357)
);

CKINVDCx16_ASAP7_75t_R g358 ( 
.A(n_359),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_390),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_363),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_362),
.B(n_363),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_389),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_365),
.A2(n_366),
.B1(n_376),
.B2(n_377),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_367),
.A2(n_368),
.B1(n_369),
.B2(n_370),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

AOI21xp5_ASAP7_75t_SL g372 ( 
.A1(n_373),
.A2(n_374),
.B(n_375),
.Y(n_372)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_L g377 ( 
.A1(n_378),
.A2(n_386),
.B(n_388),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_378),
.B(n_386),
.Y(n_388)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx3_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);


endmodule