module fake_jpeg_4662_n_60 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_60);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_60;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

BUFx12f_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_6),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_2),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_6),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_0),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_1),
.B(n_7),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx2_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_14),
.B(n_10),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_17),
.B(n_12),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

AND2x2_ASAP7_75t_SL g22 ( 
.A(n_18),
.B(n_20),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_14),
.B(n_12),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_19),
.B(n_11),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

OAI22xp33_ASAP7_75t_L g23 ( 
.A1(n_17),
.A2(n_11),
.B1(n_13),
.B2(n_10),
.Y(n_23)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_24),
.B(n_25),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_21),
.B(n_17),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_29),
.Y(n_32)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_22),
.B(n_19),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_31),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_22),
.B(n_15),
.Y(n_31)
);

AOI21xp5_ASAP7_75t_L g33 ( 
.A1(n_28),
.A2(n_20),
.B(n_8),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_33),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_28),
.A2(n_16),
.B1(n_18),
.B2(n_20),
.Y(n_34)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_20),
.C(n_16),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_37),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_16),
.C(n_18),
.Y(n_37)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g44 ( 
.A(n_40),
.Y(n_44)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_43),
.Y(n_48)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_SL g45 ( 
.A1(n_42),
.A2(n_37),
.B(n_29),
.Y(n_45)
);

A2O1A1O1Ixp25_ASAP7_75t_L g49 ( 
.A1(n_45),
.A2(n_46),
.B(n_47),
.C(n_38),
.D(n_0),
.Y(n_49)
);

NOR2xp67_ASAP7_75t_SL g46 ( 
.A(n_40),
.B(n_8),
.Y(n_46)
);

AO22x1_ASAP7_75t_L g47 ( 
.A1(n_39),
.A2(n_18),
.B1(n_1),
.B2(n_2),
.Y(n_47)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_45),
.Y(n_53)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_48),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_50),
.B(n_51),
.Y(n_52)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_53),
.B(n_54),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_50),
.B(n_42),
.C(n_39),
.Y(n_54)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_52),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_56),
.B(n_3),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_57),
.Y(n_58)
);

OAI321xp33_ASAP7_75t_L g59 ( 
.A1(n_58),
.A2(n_55),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C(n_7),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_L g60 ( 
.A(n_59),
.B(n_0),
.Y(n_60)
);


endmodule