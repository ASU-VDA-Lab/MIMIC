module fake_ariane_1577_n_2522 (n_83, n_8, n_233, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_240, n_167, n_90, n_195, n_38, n_213, n_47, n_110, n_153, n_18, n_197, n_221, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_237, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_236, n_71, n_24, n_7, n_109, n_208, n_96, n_156, n_209, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_225, n_235, n_200, n_51, n_166, n_76, n_218, n_103, n_79, n_26, n_226, n_3, n_46, n_220, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_217, n_44, n_224, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_229, n_70, n_222, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_214, n_227, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_212, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_232, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_228, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_241, n_29, n_238, n_41, n_219, n_140, n_55, n_191, n_151, n_136, n_231, n_192, n_28, n_80, n_146, n_234, n_230, n_211, n_194, n_97, n_154, n_215, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_216, n_16, n_5, n_155, n_127, n_239, n_223, n_35, n_54, n_25, n_2522);

input n_83;
input n_8;
input n_233;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_240;
input n_167;
input n_90;
input n_195;
input n_38;
input n_213;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_221;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_237;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_236;
input n_71;
input n_24;
input n_7;
input n_109;
input n_208;
input n_96;
input n_156;
input n_209;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_225;
input n_235;
input n_200;
input n_51;
input n_166;
input n_76;
input n_218;
input n_103;
input n_79;
input n_26;
input n_226;
input n_3;
input n_46;
input n_220;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_217;
input n_44;
input n_224;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_229;
input n_70;
input n_222;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_214;
input n_227;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_232;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_228;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_241;
input n_29;
input n_238;
input n_41;
input n_219;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_231;
input n_192;
input n_28;
input n_80;
input n_146;
input n_234;
input n_230;
input n_211;
input n_194;
input n_97;
input n_154;
input n_215;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_216;
input n_16;
input n_5;
input n_155;
input n_127;
input n_239;
input n_223;
input n_35;
input n_54;
input n_25;

output n_2522;

wire n_913;
wire n_1681;
wire n_2163;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_2484;
wire n_1174;
wire n_2346;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_2131;
wire n_2500;
wire n_2509;
wire n_423;
wire n_1383;
wire n_2182;
wire n_603;
wire n_373;
wire n_2135;
wire n_2334;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_2407;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_2446;
wire n_1096;
wire n_1379;
wire n_2436;
wire n_2376;
wire n_2367;
wire n_1706;
wire n_2461;
wire n_2207;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_2238;
wire n_2374;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_2380;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_2084;
wire n_568;
wire n_2278;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_2482;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_2248;
wire n_813;
wire n_419;
wire n_1985;
wire n_2288;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_2323;
wire n_1073;
wire n_402;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_2221;
wire n_672;
wire n_740;
wire n_1283;
wire n_2317;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_2342;
wire n_2200;
wire n_259;
wire n_2442;
wire n_953;
wire n_1364;
wire n_2390;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_625;
wire n_557;
wire n_2322;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_242;
wire n_1944;
wire n_331;
wire n_559;
wire n_2370;
wire n_2233;
wire n_495;
wire n_267;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_2359;
wire n_2201;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_2232;
wire n_1847;
wire n_2458;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_2227;
wire n_2301;
wire n_1539;
wire n_884;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_2433;
wire n_352;
wire n_899;
wire n_1703;
wire n_2332;
wire n_2391;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_365;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_2427;
wire n_661;
wire n_2098;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_2456;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_2341;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2094;
wire n_2512;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_2382;
wire n_2043;
wire n_780;
wire n_2349;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_2466;
wire n_676;
wire n_2038;
wire n_2263;
wire n_2116;
wire n_2271;
wire n_2145;
wire n_2326;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_249;
wire n_1108;
wire n_355;
wire n_851;
wire n_444;
wire n_1590;
wire n_1351;
wire n_2216;
wire n_1274;
wire n_257;
wire n_2426;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_2134;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_2499;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_2166;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_2185;
wire n_2398;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_306;
wire n_2415;
wire n_436;
wire n_324;
wire n_2087;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_2462;
wire n_1389;
wire n_2155;
wire n_615;
wire n_1139;
wire n_2439;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_2172;
wire n_892;
wire n_1880;
wire n_959;
wire n_2365;
wire n_2257;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_2219;
wire n_1855;
wire n_2100;
wire n_2333;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_2435;
wire n_1226;
wire n_2224;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_2167;
wire n_2293;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_2400;
wire n_632;
wire n_477;
wire n_650;
wire n_2388;
wire n_425;
wire n_2273;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_964;
wire n_1627;
wire n_2220;
wire n_382;
wire n_489;
wire n_2294;
wire n_2274;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_2378;
wire n_397;
wire n_2467;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_2253;
wire n_934;
wire n_2213;
wire n_1447;
wire n_2363;
wire n_1220;
wire n_356;
wire n_2019;
wire n_698;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_2507;
wire n_2142;
wire n_1633;
wire n_404;
wire n_1913;
wire n_2069;
wire n_2495;
wire n_1058;
wire n_2328;
wire n_347;
wire n_2434;
wire n_1042;
wire n_1234;
wire n_2311;
wire n_479;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_2287;
wire n_299;
wire n_836;
wire n_2223;
wire n_1279;
wire n_2473;
wire n_2144;
wire n_2511;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_2438;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_2262;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_2335;
wire n_370;
wire n_706;
wire n_2120;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_2404;
wire n_2168;
wire n_348;
wire n_552;
wire n_2312;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_2483;
wire n_441;
wire n_1951;
wire n_2490;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_2296;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_2241;
wire n_2373;
wire n_1173;
wire n_2350;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_2099;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2481;
wire n_2129;
wire n_855;
wire n_2327;
wire n_808;
wire n_1365;
wire n_2476;
wire n_553;
wire n_2059;
wire n_2437;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_2122;
wire n_2399;
wire n_320;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_1906;
wire n_529;
wire n_1899;
wire n_2195;
wire n_502;
wire n_2194;
wire n_1467;
wire n_247;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_2267;
wire n_1105;
wire n_547;
wire n_604;
wire n_439;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_326;
wire n_681;
wire n_874;
wire n_2286;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_2075;
wire n_1945;
wire n_545;
wire n_1015;
wire n_2418;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_2496;
wire n_2118;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_2338;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_887;
wire n_729;
wire n_2057;
wire n_2218;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_2125;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_2184;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_2254;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_1402;
wire n_957;
wire n_388;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_2217;
wire n_321;
wire n_2226;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_2256;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_1883;
wire n_2516;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_2379;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_2300;
wire n_1649;
wire n_2452;
wire n_1677;
wire n_2470;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_2284;
wire n_1844;
wire n_2283;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_2508;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_2266;
wire n_2449;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_769;
wire n_1797;
wire n_2366;
wire n_2493;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_2474;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_2460;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_2448;
wire n_2211;
wire n_2292;
wire n_2480;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_2306;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_2424;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2414;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_2389;
wire n_1309;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_2468;
wire n_1400;
wire n_342;
wire n_2035;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_2494;
wire n_1538;
wire n_2457;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_2486;
wire n_1897;
wire n_2520;
wire n_2137;
wire n_1161;
wire n_2489;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_2492;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_2337;
wire n_2265;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_2106;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_2272;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_2264;
wire n_805;
wire n_2032;
wire n_2090;
wire n_295;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_2348;
wire n_1281;
wire n_516;
wire n_2364;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_2307;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_2412;
wire n_374;
wire n_1352;
wire n_2405;
wire n_1824;
wire n_643;
wire n_1492;
wire n_2383;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_2416;
wire n_819;
wire n_2386;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_2353;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_2325;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_2022;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_1505;
wire n_2408;
wire n_2320;
wire n_979;
wire n_2329;
wire n_1642;
wire n_2417;
wire n_1815;
wire n_897;
wire n_949;
wire n_2454;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_2354;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_2368;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_2352;
wire n_2502;
wire n_1256;
wire n_714;
wire n_2170;
wire n_790;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_354;
wire n_725;
wire n_2377;
wire n_1577;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_2410;
wire n_2314;
wire n_2477;
wire n_2279;
wire n_594;
wire n_2222;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2203;
wire n_2133;
wire n_833;
wire n_1426;
wire n_2250;
wire n_2497;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_2506;
wire n_1472;
wire n_2413;
wire n_1593;
wire n_1050;
wire n_566;
wire n_2158;
wire n_2285;
wire n_1288;
wire n_1201;
wire n_858;
wire n_1185;
wire n_2475;
wire n_2173;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_2070;
wire n_2136;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_2403;
wire n_1367;
wire n_2044;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_2310;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_689;
wire n_400;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_2177;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_2343;
wire n_775;
wire n_667;
wire n_2419;
wire n_1049;
wire n_2330;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_2450;
wire n_2411;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_2309;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_2431;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_2401;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_2331;
wire n_935;
wire n_2478;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_2396;
wire n_543;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_2459;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_2196;
wire n_1038;
wire n_2371;
wire n_1978;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_2313;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_2303;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_2154;
wire n_2441;
wire n_2236;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_540;
wire n_692;
wire n_2054;
wire n_1857;
wire n_2315;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_2498;
wire n_800;
wire n_2046;
wire n_1910;
wire n_1816;
wire n_1756;
wire n_1606;
wire n_2189;
wire n_395;
wire n_621;
wire n_1587;
wire n_2093;
wire n_2340;
wire n_2018;
wire n_1772;
wire n_2444;
wire n_1014;
wire n_724;
wire n_2204;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_2199;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_2455;
wire n_827;
wire n_2231;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_2305;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_2289;
wire n_2299;
wire n_751;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_2180;
wire n_580;
wire n_1579;
wire n_494;
wire n_2181;
wire n_434;
wire n_2014;
wire n_975;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_2276;
wire n_1805;
wire n_2282;
wire n_981;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_2503;
wire n_2270;
wire n_243;
wire n_2443;
wire n_1407;
wire n_2465;
wire n_1204;
wire n_1554;
wire n_994;
wire n_2428;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_2251;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_2126;
wire n_1952;
wire n_2425;
wire n_2394;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_2356;
wire n_1601;
wire n_1057;
wire n_2487;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_2488;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_2197;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_2385;
wire n_2387;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_2291;
wire n_1980;
wire n_2518;
wire n_987;
wire n_936;
wire n_2510;
wire n_1620;
wire n_2501;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_2165;
wire n_541;
wire n_499;
wire n_1775;
wire n_908;
wire n_788;
wire n_1036;
wire n_2169;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_2402;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_663;
wire n_1720;
wire n_2409;
wire n_443;
wire n_2176;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_2453;
wire n_2344;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_2392;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_2321;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_385;
wire n_2395;
wire n_917;
wire n_1271;
wire n_372;
wire n_2096;
wire n_2440;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_631;
wire n_399;
wire n_1170;
wire n_2258;
wire n_1261;
wire n_2471;
wire n_702;
wire n_898;
wire n_857;
wire n_968;
wire n_1067;
wire n_363;
wire n_1235;
wire n_1323;
wire n_2375;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_761;
wire n_733;
wire n_2212;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_2268;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_2252;
wire n_2111;
wire n_2420;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_2445;
wire n_1770;
wire n_701;
wire n_1003;
wire n_2469;
wire n_1125;
wire n_2103;
wire n_2358;
wire n_1710;
wire n_1865;
wire n_2463;
wire n_309;
wire n_1344;
wire n_2355;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_2062;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_2153;
wire n_2324;
wire n_1510;
wire n_2505;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_2397;
wire n_2521;
wire n_369;
wire n_1727;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_2351;
wire n_2260;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_2206;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_2347;
wire n_248;
wire n_1152;
wire n_2447;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_2101;
wire n_921;
wire n_2362;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_2372;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_2422;
wire n_1334;
wire n_654;
wire n_2290;
wire n_2088;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2429;
wire n_2108;
wire n_1039;
wire n_2246;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_2339;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2191;
wire n_1497;
wire n_1866;
wire n_2472;
wire n_2056;
wire n_459;
wire n_1136;
wire n_2515;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_2519;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_2360;
wire n_723;
wire n_1393;
wire n_2240;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_2085;
wire n_2432;
wire n_1686;
wire n_1964;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_2188;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_2430;
wire n_2504;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_2297;
wire n_371;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_1223;
wire n_308;
wire n_1768;
wire n_2513;
wire n_2193;
wire n_2369;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2451;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_2148;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_415;
wire n_2381;
wire n_1967;
wire n_2384;
wire n_2179;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_2485;
wire n_537;
wire n_1063;
wire n_991;
wire n_2183;
wire n_2275;
wire n_2205;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1799;
wire n_1707;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2357;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_2209;
wire n_2421;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_2269;
wire n_472;
wire n_937;
wire n_1474;
wire n_2081;
wire n_265;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_2318;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_2361;
wire n_1115;
wire n_2229;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_2255;
wire n_1129;
wire n_1252;
wire n_2239;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_2316;
wire n_2464;
wire n_1010;
wire n_882;
wire n_2304;
wire n_1249;
wire n_803;
wire n_1871;
wire n_2514;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_289;
wire n_548;
wire n_2336;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_2491;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_2517;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_484;
wire n_411;
wire n_2259;
wire n_849;
wire n_2095;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_2208;
wire n_2423;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_2479;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_2345;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_SL g242 ( 
.A(n_208),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_191),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_210),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g245 ( 
.A(n_96),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_107),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_20),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_162),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_240),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_7),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_143),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_92),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_36),
.Y(n_253)
);

BUFx10_ASAP7_75t_L g254 ( 
.A(n_94),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_132),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_226),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_163),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_36),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_118),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_91),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_137),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_188),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_18),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_151),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_203),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_56),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_43),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_199),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_204),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_78),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_88),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_232),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_72),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_158),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_6),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_235),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_229),
.Y(n_277)
);

INVx1_ASAP7_75t_SL g278 ( 
.A(n_175),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_121),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_45),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_157),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_10),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_99),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_40),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_98),
.Y(n_285)
);

BUFx8_ASAP7_75t_SL g286 ( 
.A(n_57),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_8),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_202),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_3),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_170),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_178),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_110),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_144),
.Y(n_293)
);

INVx1_ASAP7_75t_SL g294 ( 
.A(n_105),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_221),
.Y(n_295)
);

INVx2_ASAP7_75t_SL g296 ( 
.A(n_166),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_207),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_91),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_23),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_239),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_98),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_27),
.Y(n_302)
);

INVx2_ASAP7_75t_SL g303 ( 
.A(n_32),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_176),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_123),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_65),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_48),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_171),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_5),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_120),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_79),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_47),
.Y(n_312)
);

INVx1_ASAP7_75t_SL g313 ( 
.A(n_172),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_112),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_194),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_100),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_146),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_56),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_94),
.Y(n_319)
);

BUFx3_ASAP7_75t_L g320 ( 
.A(n_82),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_187),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_19),
.Y(n_322)
);

INVx1_ASAP7_75t_SL g323 ( 
.A(n_150),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_218),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_238),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_113),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_136),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_46),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_73),
.Y(n_329)
);

INVx2_ASAP7_75t_SL g330 ( 
.A(n_160),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_55),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_111),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_139),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_42),
.Y(n_334)
);

BUFx3_ASAP7_75t_L g335 ( 
.A(n_149),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_100),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_119),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_109),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_193),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_124),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_105),
.Y(n_341)
);

CKINVDCx16_ASAP7_75t_R g342 ( 
.A(n_63),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_48),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_89),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_95),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_206),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_18),
.Y(n_347)
);

BUFx3_ASAP7_75t_L g348 ( 
.A(n_213),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_79),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_45),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_73),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_103),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_201),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_148),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_85),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_190),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_10),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_177),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_99),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_25),
.Y(n_360)
);

CKINVDCx16_ASAP7_75t_R g361 ( 
.A(n_80),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_211),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_184),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_169),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_47),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_11),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_165),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_101),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_186),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_159),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_237),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_127),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_227),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_64),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_233),
.Y(n_375)
);

BUFx3_ASAP7_75t_L g376 ( 
.A(n_97),
.Y(n_376)
);

INVx1_ASAP7_75t_SL g377 ( 
.A(n_197),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_54),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_156),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_19),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_0),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_58),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_114),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_35),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_22),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_78),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_53),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_102),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_101),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_25),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_134),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_224),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_155),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_2),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_62),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_225),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_168),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_2),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_21),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_67),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_234),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_116),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_198),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_81),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_128),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_28),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_102),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_161),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_34),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_40),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_154),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_181),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_44),
.Y(n_413)
);

BUFx10_ASAP7_75t_L g414 ( 
.A(n_220),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_58),
.Y(n_415)
);

INVx2_ASAP7_75t_SL g416 ( 
.A(n_39),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_69),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_147),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_214),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_26),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_28),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_97),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_23),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_219),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_217),
.Y(n_425)
);

BUFx10_ASAP7_75t_L g426 ( 
.A(n_111),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_68),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_183),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_54),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_9),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_215),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_131),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_12),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_133),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_43),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_216),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_29),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_117),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_61),
.Y(n_439)
);

BUFx3_ASAP7_75t_L g440 ( 
.A(n_80),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_83),
.Y(n_441)
);

INVx1_ASAP7_75t_SL g442 ( 
.A(n_212),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_0),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_31),
.Y(n_444)
);

BUFx10_ASAP7_75t_L g445 ( 
.A(n_64),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_35),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_6),
.Y(n_447)
);

BUFx2_ASAP7_75t_L g448 ( 
.A(n_152),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_66),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_51),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_222),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_42),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_130),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_29),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_83),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_179),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_96),
.Y(n_457)
);

INVx1_ASAP7_75t_SL g458 ( 
.A(n_90),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_37),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_129),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_49),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_93),
.Y(n_462)
);

BUFx10_ASAP7_75t_L g463 ( 
.A(n_145),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_92),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_21),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_27),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_231),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_107),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_12),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_87),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_44),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_20),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_3),
.Y(n_473)
);

CKINVDCx16_ASAP7_75t_R g474 ( 
.A(n_342),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_286),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_448),
.B(n_244),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_248),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_255),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_244),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_321),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_356),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_249),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_249),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_358),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_418),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_289),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_251),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_251),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_451),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_268),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_273),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_357),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_268),
.Y(n_493)
);

BUFx2_ASAP7_75t_L g494 ( 
.A(n_245),
.Y(n_494)
);

INVxp67_ASAP7_75t_L g495 ( 
.A(n_303),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_342),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_274),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_361),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_361),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_289),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_274),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_448),
.B(n_1),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_246),
.Y(n_503)
);

INVxp67_ASAP7_75t_L g504 ( 
.A(n_266),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_276),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_289),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_276),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_277),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_247),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_250),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_277),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_365),
.Y(n_512)
);

CKINVDCx14_ASAP7_75t_R g513 ( 
.A(n_414),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_279),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_279),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_252),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_253),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_281),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_281),
.Y(n_519)
);

NOR2xp67_ASAP7_75t_L g520 ( 
.A(n_303),
.B(n_1),
.Y(n_520)
);

INVxp67_ASAP7_75t_L g521 ( 
.A(n_266),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_300),
.B(n_4),
.Y(n_522)
);

NOR2xp67_ASAP7_75t_L g523 ( 
.A(n_416),
.B(n_299),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_258),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_289),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_386),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_447),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_289),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_260),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_263),
.Y(n_530)
);

INVxp67_ASAP7_75t_SL g531 ( 
.A(n_320),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_300),
.Y(n_532)
);

BUFx10_ASAP7_75t_L g533 ( 
.A(n_296),
.Y(n_533)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_455),
.Y(n_534)
);

CKINVDCx20_ASAP7_75t_R g535 ( 
.A(n_462),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_270),
.Y(n_536)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_348),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_280),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_289),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_315),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_348),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_282),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_315),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_324),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_324),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_325),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_325),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_284),
.Y(n_548)
);

CKINVDCx16_ASAP7_75t_R g549 ( 
.A(n_414),
.Y(n_549)
);

INVxp33_ASAP7_75t_L g550 ( 
.A(n_271),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_337),
.Y(n_551)
);

INVxp67_ASAP7_75t_SL g552 ( 
.A(n_320),
.Y(n_552)
);

CKINVDCx20_ASAP7_75t_R g553 ( 
.A(n_348),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_337),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_285),
.Y(n_555)
);

INVxp67_ASAP7_75t_L g556 ( 
.A(n_271),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_287),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_298),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_339),
.Y(n_559)
);

HB1xp67_ASAP7_75t_L g560 ( 
.A(n_306),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_309),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_311),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_311),
.Y(n_563)
);

BUFx2_ASAP7_75t_L g564 ( 
.A(n_320),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_312),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_339),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_314),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_340),
.B(n_4),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_340),
.Y(n_569)
);

INVxp67_ASAP7_75t_SL g570 ( 
.A(n_376),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_316),
.Y(n_571)
);

INVxp33_ASAP7_75t_SL g572 ( 
.A(n_318),
.Y(n_572)
);

CKINVDCx20_ASAP7_75t_R g573 ( 
.A(n_414),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_376),
.B(n_5),
.Y(n_574)
);

INVxp67_ASAP7_75t_L g575 ( 
.A(n_275),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_322),
.Y(n_576)
);

CKINVDCx20_ASAP7_75t_R g577 ( 
.A(n_414),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_353),
.Y(n_578)
);

CKINVDCx20_ASAP7_75t_R g579 ( 
.A(n_463),
.Y(n_579)
);

BUFx3_ASAP7_75t_L g580 ( 
.A(n_335),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_353),
.Y(n_581)
);

HB1xp67_ASAP7_75t_L g582 ( 
.A(n_326),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_362),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_328),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_331),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_338),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_362),
.B(n_7),
.Y(n_587)
);

INVxp67_ASAP7_75t_L g588 ( 
.A(n_275),
.Y(n_588)
);

CKINVDCx20_ASAP7_75t_R g589 ( 
.A(n_463),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_341),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_343),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_344),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_369),
.Y(n_593)
);

HB1xp67_ASAP7_75t_L g594 ( 
.A(n_345),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_369),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_375),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_311),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_375),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_379),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_379),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_383),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_383),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_347),
.Y(n_603)
);

CKINVDCx20_ASAP7_75t_R g604 ( 
.A(n_463),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_480),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_477),
.Y(n_606)
);

OAI21x1_ASAP7_75t_L g607 ( 
.A1(n_522),
.A2(n_396),
.B(n_393),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_478),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_479),
.B(n_393),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_479),
.Y(n_610)
);

CKINVDCx20_ASAP7_75t_R g611 ( 
.A(n_491),
.Y(n_611)
);

NAND2xp33_ASAP7_75t_L g612 ( 
.A(n_503),
.B(n_509),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_482),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_481),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_484),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g616 ( 
.A(n_564),
.B(n_376),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_485),
.Y(n_617)
);

CKINVDCx20_ASAP7_75t_R g618 ( 
.A(n_492),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_482),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_483),
.Y(n_620)
);

OAI21x1_ASAP7_75t_L g621 ( 
.A1(n_522),
.A2(n_408),
.B(n_396),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_489),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_549),
.B(n_311),
.Y(n_623)
);

CKINVDCx20_ASAP7_75t_R g624 ( 
.A(n_512),
.Y(n_624)
);

BUFx6f_ASAP7_75t_L g625 ( 
.A(n_486),
.Y(n_625)
);

INVx4_ASAP7_75t_L g626 ( 
.A(n_574),
.Y(n_626)
);

CKINVDCx20_ASAP7_75t_R g627 ( 
.A(n_526),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_486),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_475),
.Y(n_629)
);

HB1xp67_ASAP7_75t_L g630 ( 
.A(n_474),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g631 ( 
.A(n_486),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_483),
.B(n_408),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_487),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_R g634 ( 
.A(n_513),
.B(n_243),
.Y(n_634)
);

INVxp67_ASAP7_75t_L g635 ( 
.A(n_560),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_487),
.B(n_411),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_488),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_R g638 ( 
.A(n_510),
.B(n_256),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_488),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_500),
.Y(n_640)
);

INVx3_ASAP7_75t_L g641 ( 
.A(n_500),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_490),
.Y(n_642)
);

NAND3xp33_ASAP7_75t_L g643 ( 
.A(n_476),
.B(n_292),
.C(n_283),
.Y(n_643)
);

CKINVDCx16_ASAP7_75t_R g644 ( 
.A(n_549),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_R g645 ( 
.A(n_516),
.B(n_517),
.Y(n_645)
);

HB1xp67_ASAP7_75t_L g646 ( 
.A(n_474),
.Y(n_646)
);

HB1xp67_ASAP7_75t_L g647 ( 
.A(n_496),
.Y(n_647)
);

BUFx2_ASAP7_75t_L g648 ( 
.A(n_498),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_564),
.B(n_440),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_490),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_500),
.Y(n_651)
);

CKINVDCx20_ASAP7_75t_R g652 ( 
.A(n_527),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_493),
.B(n_440),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_493),
.Y(n_654)
);

BUFx6f_ASAP7_75t_L g655 ( 
.A(n_506),
.Y(n_655)
);

BUFx2_ASAP7_75t_L g656 ( 
.A(n_499),
.Y(n_656)
);

INVxp67_ASAP7_75t_SL g657 ( 
.A(n_497),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_497),
.Y(n_658)
);

INVx3_ASAP7_75t_L g659 ( 
.A(n_506),
.Y(n_659)
);

INVx3_ASAP7_75t_L g660 ( 
.A(n_506),
.Y(n_660)
);

INVx1_ASAP7_75t_SL g661 ( 
.A(n_537),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_501),
.B(n_411),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_524),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_525),
.Y(n_664)
);

BUFx3_ASAP7_75t_L g665 ( 
.A(n_580),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_529),
.Y(n_666)
);

CKINVDCx20_ASAP7_75t_R g667 ( 
.A(n_534),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_530),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_501),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_505),
.B(n_440),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_536),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_505),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_525),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_538),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_542),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_507),
.Y(n_676)
);

BUFx6f_ASAP7_75t_L g677 ( 
.A(n_525),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_548),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_507),
.B(n_301),
.Y(n_679)
);

BUFx6f_ASAP7_75t_L g680 ( 
.A(n_528),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_555),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_528),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_528),
.Y(n_683)
);

BUFx2_ASAP7_75t_L g684 ( 
.A(n_557),
.Y(n_684)
);

BUFx6f_ASAP7_75t_L g685 ( 
.A(n_539),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_539),
.Y(n_686)
);

BUFx6f_ASAP7_75t_L g687 ( 
.A(n_539),
.Y(n_687)
);

CKINVDCx20_ASAP7_75t_R g688 ( 
.A(n_535),
.Y(n_688)
);

NOR2xp67_ASAP7_75t_L g689 ( 
.A(n_508),
.B(n_296),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_558),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_R g691 ( 
.A(n_561),
.B(n_257),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_R g692 ( 
.A(n_565),
.B(n_259),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_508),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_567),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_511),
.B(n_412),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_562),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_571),
.Y(n_697)
);

BUFx2_ASAP7_75t_L g698 ( 
.A(n_576),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_511),
.B(n_301),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_562),
.Y(n_700)
);

CKINVDCx20_ASAP7_75t_R g701 ( 
.A(n_573),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_514),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_562),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_640),
.Y(n_704)
);

INVx5_ASAP7_75t_L g705 ( 
.A(n_625),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_623),
.B(n_572),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_623),
.B(n_584),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_SL g708 ( 
.A(n_644),
.B(n_577),
.Y(n_708)
);

AND2x6_ASAP7_75t_L g709 ( 
.A(n_610),
.B(n_574),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_657),
.B(n_533),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_629),
.Y(n_711)
);

AND2x4_ASAP7_75t_L g712 ( 
.A(n_657),
.B(n_531),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_626),
.B(n_533),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_640),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_610),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_626),
.B(n_533),
.Y(n_716)
);

INVx3_ASAP7_75t_L g717 ( 
.A(n_665),
.Y(n_717)
);

HB1xp67_ASAP7_75t_L g718 ( 
.A(n_630),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_665),
.B(n_585),
.Y(n_719)
);

INVx3_ASAP7_75t_L g720 ( 
.A(n_665),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_613),
.Y(n_721)
);

INVx5_ASAP7_75t_L g722 ( 
.A(n_625),
.Y(n_722)
);

INVxp33_ASAP7_75t_L g723 ( 
.A(n_630),
.Y(n_723)
);

BUFx6f_ASAP7_75t_L g724 ( 
.A(n_625),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_613),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_626),
.B(n_533),
.Y(n_726)
);

BUFx6f_ASAP7_75t_L g727 ( 
.A(n_625),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_619),
.Y(n_728)
);

BUFx6f_ASAP7_75t_L g729 ( 
.A(n_625),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_619),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_640),
.Y(n_731)
);

AOI22xp5_ASAP7_75t_L g732 ( 
.A1(n_635),
.A2(n_502),
.B1(n_590),
.B2(n_586),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_620),
.Y(n_733)
);

OR2x2_ASAP7_75t_L g734 ( 
.A(n_644),
.B(n_494),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_638),
.B(n_591),
.Y(n_735)
);

AOI22xp33_ASAP7_75t_L g736 ( 
.A1(n_643),
.A2(n_587),
.B1(n_568),
.B2(n_494),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_620),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_633),
.Y(n_738)
);

AND2x2_ASAP7_75t_L g739 ( 
.A(n_626),
.B(n_552),
.Y(n_739)
);

INVxp67_ASAP7_75t_SL g740 ( 
.A(n_689),
.Y(n_740)
);

INVx4_ASAP7_75t_L g741 ( 
.A(n_626),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_633),
.Y(n_742)
);

BUFx3_ASAP7_75t_L g743 ( 
.A(n_637),
.Y(n_743)
);

INVx2_ASAP7_75t_SL g744 ( 
.A(n_616),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_637),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_639),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_639),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_651),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_642),
.B(n_650),
.Y(n_749)
);

INVx1_ASAP7_75t_SL g750 ( 
.A(n_661),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_651),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_642),
.Y(n_752)
);

BUFx6f_ASAP7_75t_L g753 ( 
.A(n_625),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_651),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_664),
.Y(n_755)
);

BUFx2_ASAP7_75t_L g756 ( 
.A(n_646),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_635),
.B(n_592),
.Y(n_757)
);

INVx2_ASAP7_75t_SL g758 ( 
.A(n_616),
.Y(n_758)
);

AOI22x1_ASAP7_75t_L g759 ( 
.A1(n_650),
.A2(n_514),
.B1(n_518),
.B2(n_515),
.Y(n_759)
);

AND2x4_ASAP7_75t_L g760 ( 
.A(n_653),
.B(n_570),
.Y(n_760)
);

AO22x2_ASAP7_75t_L g761 ( 
.A1(n_643),
.A2(n_518),
.B1(n_519),
.B2(n_515),
.Y(n_761)
);

OR2x6_ASAP7_75t_L g762 ( 
.A(n_684),
.B(n_520),
.Y(n_762)
);

INVx4_ASAP7_75t_L g763 ( 
.A(n_625),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_664),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_638),
.B(n_603),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_616),
.B(n_541),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_691),
.B(n_692),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_654),
.Y(n_768)
);

BUFx3_ASAP7_75t_L g769 ( 
.A(n_654),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_679),
.B(n_699),
.Y(n_770)
);

CKINVDCx20_ASAP7_75t_R g771 ( 
.A(n_624),
.Y(n_771)
);

AO22x2_ASAP7_75t_L g772 ( 
.A1(n_661),
.A2(n_532),
.B1(n_540),
.B2(n_519),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_658),
.B(n_580),
.Y(n_773)
);

BUFx10_ASAP7_75t_L g774 ( 
.A(n_663),
.Y(n_774)
);

AOI22xp5_ASAP7_75t_L g775 ( 
.A1(n_612),
.A2(n_553),
.B1(n_520),
.B2(n_579),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_605),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_658),
.B(n_580),
.Y(n_777)
);

INVx4_ASAP7_75t_L g778 ( 
.A(n_628),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_649),
.B(n_582),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_669),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_669),
.Y(n_781)
);

AND2x4_ASAP7_75t_L g782 ( 
.A(n_653),
.B(n_504),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_672),
.Y(n_783)
);

AND2x2_ASAP7_75t_L g784 ( 
.A(n_679),
.B(n_550),
.Y(n_784)
);

AND2x6_ASAP7_75t_L g785 ( 
.A(n_672),
.B(n_412),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_645),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_664),
.Y(n_787)
);

CKINVDCx20_ASAP7_75t_R g788 ( 
.A(n_624),
.Y(n_788)
);

BUFx2_ASAP7_75t_L g789 ( 
.A(n_646),
.Y(n_789)
);

BUFx6f_ASAP7_75t_L g790 ( 
.A(n_628),
.Y(n_790)
);

BUFx6f_ASAP7_75t_L g791 ( 
.A(n_628),
.Y(n_791)
);

BUFx10_ASAP7_75t_L g792 ( 
.A(n_666),
.Y(n_792)
);

INVx4_ASAP7_75t_L g793 ( 
.A(n_628),
.Y(n_793)
);

BUFx10_ASAP7_75t_L g794 ( 
.A(n_668),
.Y(n_794)
);

AND2x6_ASAP7_75t_L g795 ( 
.A(n_676),
.B(n_419),
.Y(n_795)
);

INVxp67_ASAP7_75t_SL g796 ( 
.A(n_689),
.Y(n_796)
);

NAND3xp33_ASAP7_75t_L g797 ( 
.A(n_671),
.B(n_675),
.C(n_674),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_676),
.B(n_532),
.Y(n_798)
);

INVx2_ASAP7_75t_SL g799 ( 
.A(n_649),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_693),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_673),
.Y(n_801)
);

INVx1_ASAP7_75t_SL g802 ( 
.A(n_611),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_693),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_702),
.Y(n_804)
);

AOI22xp33_ASAP7_75t_L g805 ( 
.A1(n_607),
.A2(n_543),
.B1(n_544),
.B2(n_540),
.Y(n_805)
);

INVx6_ASAP7_75t_L g806 ( 
.A(n_653),
.Y(n_806)
);

BUFx3_ASAP7_75t_L g807 ( 
.A(n_702),
.Y(n_807)
);

OR2x2_ASAP7_75t_L g808 ( 
.A(n_684),
.B(n_594),
.Y(n_808)
);

NAND3xp33_ASAP7_75t_L g809 ( 
.A(n_678),
.B(n_495),
.C(n_521),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_SL g810 ( 
.A(n_691),
.B(n_692),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_645),
.B(n_589),
.Y(n_811)
);

AND2x6_ASAP7_75t_L g812 ( 
.A(n_670),
.B(n_419),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_673),
.Y(n_813)
);

AND2x2_ASAP7_75t_L g814 ( 
.A(n_679),
.B(n_543),
.Y(n_814)
);

AND2x4_ASAP7_75t_L g815 ( 
.A(n_670),
.B(n_556),
.Y(n_815)
);

AO21x2_ASAP7_75t_L g816 ( 
.A1(n_607),
.A2(n_621),
.B(n_609),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_673),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_703),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_682),
.Y(n_819)
);

INVx2_ASAP7_75t_SL g820 ( 
.A(n_649),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_699),
.B(n_544),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_682),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_670),
.B(n_545),
.Y(n_823)
);

BUFx6f_ASAP7_75t_L g824 ( 
.A(n_628),
.Y(n_824)
);

AND2x4_ASAP7_75t_L g825 ( 
.A(n_699),
.B(n_575),
.Y(n_825)
);

INVx4_ASAP7_75t_SL g826 ( 
.A(n_628),
.Y(n_826)
);

OAI22xp5_ASAP7_75t_L g827 ( 
.A1(n_698),
.A2(n_690),
.B1(n_694),
.B2(n_681),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_634),
.B(n_604),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_609),
.B(n_545),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_606),
.Y(n_830)
);

HB1xp67_ASAP7_75t_L g831 ( 
.A(n_698),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_682),
.Y(n_832)
);

CKINVDCx11_ASAP7_75t_R g833 ( 
.A(n_627),
.Y(n_833)
);

INVx4_ASAP7_75t_L g834 ( 
.A(n_628),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_683),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_683),
.Y(n_836)
);

BUFx6f_ASAP7_75t_L g837 ( 
.A(n_631),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_683),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_686),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_703),
.Y(n_840)
);

INVxp67_ASAP7_75t_SL g841 ( 
.A(n_632),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_632),
.B(n_546),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_636),
.B(n_662),
.Y(n_843)
);

AOI22xp33_ASAP7_75t_L g844 ( 
.A1(n_607),
.A2(n_547),
.B1(n_551),
.B2(n_546),
.Y(n_844)
);

AOI22xp33_ASAP7_75t_L g845 ( 
.A1(n_621),
.A2(n_551),
.B1(n_554),
.B2(n_547),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_703),
.Y(n_846)
);

INVx8_ASAP7_75t_L g847 ( 
.A(n_697),
.Y(n_847)
);

INVxp67_ASAP7_75t_SL g848 ( 
.A(n_636),
.Y(n_848)
);

BUFx3_ASAP7_75t_L g849 ( 
.A(n_631),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_686),
.Y(n_850)
);

CKINVDCx6p67_ASAP7_75t_R g851 ( 
.A(n_618),
.Y(n_851)
);

INVx1_ASAP7_75t_SL g852 ( 
.A(n_652),
.Y(n_852)
);

OR2x2_ASAP7_75t_L g853 ( 
.A(n_648),
.B(n_495),
.Y(n_853)
);

BUFx6f_ASAP7_75t_L g854 ( 
.A(n_631),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_662),
.Y(n_855)
);

INVx3_ASAP7_75t_L g856 ( 
.A(n_631),
.Y(n_856)
);

INVx6_ASAP7_75t_L g857 ( 
.A(n_631),
.Y(n_857)
);

INVx2_ASAP7_75t_SL g858 ( 
.A(n_634),
.Y(n_858)
);

INVx3_ASAP7_75t_L g859 ( 
.A(n_631),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_695),
.Y(n_860)
);

INVx2_ASAP7_75t_SL g861 ( 
.A(n_648),
.Y(n_861)
);

HB1xp67_ASAP7_75t_L g862 ( 
.A(n_656),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_695),
.Y(n_863)
);

INVx4_ASAP7_75t_L g864 ( 
.A(n_631),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_641),
.B(n_554),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_686),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_696),
.Y(n_867)
);

INVx3_ASAP7_75t_L g868 ( 
.A(n_741),
.Y(n_868)
);

AOI22xp5_ASAP7_75t_L g869 ( 
.A1(n_706),
.A2(n_656),
.B1(n_647),
.B2(n_428),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_861),
.B(n_647),
.Y(n_870)
);

OAI21xp5_ASAP7_75t_L g871 ( 
.A1(n_843),
.A2(n_621),
.B(n_432),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_704),
.Y(n_872)
);

OAI22xp5_ASAP7_75t_L g873 ( 
.A1(n_841),
.A2(n_351),
.B1(n_359),
.B2(n_349),
.Y(n_873)
);

HB1xp67_ASAP7_75t_L g874 ( 
.A(n_756),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_848),
.B(n_559),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_829),
.B(n_855),
.Y(n_876)
);

INVx4_ASAP7_75t_L g877 ( 
.A(n_741),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_829),
.B(n_559),
.Y(n_878)
);

INVx2_ASAP7_75t_SL g879 ( 
.A(n_750),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_743),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_860),
.B(n_566),
.Y(n_881)
);

BUFx3_ASAP7_75t_L g882 ( 
.A(n_847),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_743),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_863),
.B(n_566),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_739),
.B(n_569),
.Y(n_885)
);

NAND2x1_ASAP7_75t_L g886 ( 
.A(n_709),
.B(n_741),
.Y(n_886)
);

BUFx2_ASAP7_75t_L g887 ( 
.A(n_756),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_769),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_769),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_711),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_739),
.B(n_712),
.Y(n_891)
);

AOI22xp5_ASAP7_75t_L g892 ( 
.A1(n_707),
.A2(n_428),
.B1(n_438),
.B2(n_432),
.Y(n_892)
);

AOI22xp5_ASAP7_75t_L g893 ( 
.A1(n_812),
.A2(n_712),
.B1(n_709),
.B2(n_757),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_858),
.B(n_438),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_807),
.Y(n_895)
);

NOR2xp33_ASAP7_75t_SL g896 ( 
.A(n_786),
.B(n_608),
.Y(n_896)
);

OR2x6_ASAP7_75t_L g897 ( 
.A(n_847),
.B(n_588),
.Y(n_897)
);

AND2x4_ASAP7_75t_L g898 ( 
.A(n_770),
.B(n_569),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_807),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_858),
.B(n_456),
.Y(n_900)
);

NOR2x2_ASAP7_75t_L g901 ( 
.A(n_762),
.B(n_366),
.Y(n_901)
);

AOI22xp33_ASAP7_75t_L g902 ( 
.A1(n_812),
.A2(n_772),
.B1(n_761),
.B2(n_709),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_704),
.Y(n_903)
);

AOI22xp33_ASAP7_75t_L g904 ( 
.A1(n_812),
.A2(n_772),
.B1(n_761),
.B2(n_709),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_715),
.Y(n_905)
);

AOI22xp5_ASAP7_75t_L g906 ( 
.A1(n_812),
.A2(n_456),
.B1(n_330),
.B2(n_578),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_715),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_712),
.B(n_710),
.Y(n_908)
);

OAI21xp5_ASAP7_75t_L g909 ( 
.A1(n_725),
.A2(n_581),
.B(n_578),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_842),
.B(n_581),
.Y(n_910)
);

NOR2xp33_ASAP7_75t_L g911 ( 
.A(n_806),
.B(n_267),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_719),
.B(n_583),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_814),
.B(n_821),
.Y(n_913)
);

BUFx3_ASAP7_75t_L g914 ( 
.A(n_847),
.Y(n_914)
);

O2A1O1Ixp33_ASAP7_75t_L g915 ( 
.A1(n_823),
.A2(n_416),
.B(n_292),
.C(n_302),
.Y(n_915)
);

NOR2xp67_ASAP7_75t_L g916 ( 
.A(n_786),
.B(n_614),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_714),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_725),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_728),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_728),
.Y(n_920)
);

AND2x4_ASAP7_75t_SL g921 ( 
.A(n_774),
.B(n_688),
.Y(n_921)
);

NAND2xp33_ASAP7_75t_L g922 ( 
.A(n_709),
.B(n_311),
.Y(n_922)
);

INVxp33_ASAP7_75t_L g923 ( 
.A(n_766),
.Y(n_923)
);

OR2x6_ASAP7_75t_L g924 ( 
.A(n_847),
.B(n_523),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_SL g925 ( 
.A(n_861),
.B(n_583),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_814),
.B(n_593),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_730),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_821),
.B(n_593),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_760),
.B(n_595),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_SL g930 ( 
.A(n_713),
.B(n_716),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_SL g931 ( 
.A(n_726),
.B(n_595),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_730),
.Y(n_932)
);

INVx5_ASAP7_75t_L g933 ( 
.A(n_709),
.Y(n_933)
);

INVx2_ASAP7_75t_SL g934 ( 
.A(n_789),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_760),
.B(n_596),
.Y(n_935)
);

INVx2_ASAP7_75t_SL g936 ( 
.A(n_789),
.Y(n_936)
);

AND2x6_ASAP7_75t_SL g937 ( 
.A(n_762),
.B(n_283),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_SL g938 ( 
.A(n_767),
.B(n_596),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_L g939 ( 
.A(n_806),
.B(n_294),
.Y(n_939)
);

AOI22xp33_ASAP7_75t_L g940 ( 
.A1(n_812),
.A2(n_598),
.B1(n_600),
.B2(n_599),
.Y(n_940)
);

INVxp33_ASAP7_75t_SL g941 ( 
.A(n_711),
.Y(n_941)
);

AOI21x1_ASAP7_75t_L g942 ( 
.A1(n_817),
.A2(n_700),
.B(n_696),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_SL g943 ( 
.A(n_810),
.B(n_598),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_SL g944 ( 
.A(n_776),
.B(n_615),
.Y(n_944)
);

AOI22xp33_ASAP7_75t_L g945 ( 
.A1(n_812),
.A2(n_599),
.B1(n_601),
.B2(n_600),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_760),
.B(n_601),
.Y(n_946)
);

OR2x2_ASAP7_75t_L g947 ( 
.A(n_853),
.B(n_734),
.Y(n_947)
);

OR2x6_ASAP7_75t_L g948 ( 
.A(n_762),
.B(n_523),
.Y(n_948)
);

AOI22xp5_ASAP7_75t_L g949 ( 
.A1(n_812),
.A2(n_709),
.B1(n_758),
.B2(n_744),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_SL g950 ( 
.A(n_805),
.B(n_602),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_714),
.Y(n_951)
);

OR2x2_ASAP7_75t_L g952 ( 
.A(n_853),
.B(n_617),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_779),
.B(n_602),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_744),
.B(n_242),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_758),
.B(n_278),
.Y(n_955)
);

AOI22xp33_ASAP7_75t_L g956 ( 
.A1(n_772),
.A2(n_463),
.B1(n_458),
.B2(n_426),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_799),
.B(n_820),
.Y(n_957)
);

OR2x2_ASAP7_75t_L g958 ( 
.A(n_734),
.B(n_622),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_L g959 ( 
.A(n_806),
.B(n_374),
.Y(n_959)
);

NOR2xp33_ASAP7_75t_L g960 ( 
.A(n_806),
.B(n_380),
.Y(n_960)
);

BUFx6f_ASAP7_75t_L g961 ( 
.A(n_724),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_784),
.B(n_701),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_733),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_L g964 ( 
.A(n_799),
.B(n_384),
.Y(n_964)
);

BUFx3_ASAP7_75t_L g965 ( 
.A(n_774),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_820),
.B(n_385),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_784),
.B(n_313),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_770),
.B(n_323),
.Y(n_968)
);

NOR2xp67_ASAP7_75t_SL g969 ( 
.A(n_797),
.B(n_302),
.Y(n_969)
);

AOI22xp33_ASAP7_75t_L g970 ( 
.A1(n_772),
.A2(n_426),
.B1(n_445),
.B2(n_254),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_721),
.B(n_377),
.Y(n_971)
);

AOI22xp33_ASAP7_75t_L g972 ( 
.A1(n_761),
.A2(n_426),
.B1(n_445),
.B2(n_254),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_SL g973 ( 
.A(n_844),
.B(n_330),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_768),
.B(n_442),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_733),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_737),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_SL g977 ( 
.A(n_845),
.B(n_261),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_749),
.A2(n_700),
.B(n_696),
.Y(n_978)
);

BUFx6f_ASAP7_75t_L g979 ( 
.A(n_724),
.Y(n_979)
);

BUFx6f_ASAP7_75t_L g980 ( 
.A(n_724),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_737),
.Y(n_981)
);

BUFx3_ASAP7_75t_L g982 ( 
.A(n_774),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_738),
.Y(n_983)
);

INVxp67_ASAP7_75t_SL g984 ( 
.A(n_717),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_SL g985 ( 
.A(n_738),
.B(n_261),
.Y(n_985)
);

INVx4_ASAP7_75t_L g986 ( 
.A(n_785),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_SL g987 ( 
.A(n_742),
.B(n_295),
.Y(n_987)
);

NOR2xp33_ASAP7_75t_L g988 ( 
.A(n_740),
.B(n_388),
.Y(n_988)
);

AND2x2_ASAP7_75t_L g989 ( 
.A(n_831),
.B(n_627),
.Y(n_989)
);

A2O1A1Ixp33_ASAP7_75t_L g990 ( 
.A1(n_742),
.A2(n_307),
.B(n_329),
.C(n_319),
.Y(n_990)
);

INVx8_ASAP7_75t_L g991 ( 
.A(n_762),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_745),
.B(n_641),
.Y(n_992)
);

AOI22xp5_ASAP7_75t_L g993 ( 
.A1(n_782),
.A2(n_262),
.B1(n_265),
.B2(n_264),
.Y(n_993)
);

INVx4_ASAP7_75t_L g994 ( 
.A(n_717),
.Y(n_994)
);

NAND3xp33_ASAP7_75t_SL g995 ( 
.A(n_776),
.B(n_390),
.C(n_389),
.Y(n_995)
);

AOI22x1_ASAP7_75t_L g996 ( 
.A1(n_745),
.A2(n_307),
.B1(n_329),
.B2(n_319),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_796),
.B(n_395),
.Y(n_997)
);

NOR2x1p5_ASAP7_75t_L g998 ( 
.A(n_808),
.B(n_399),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_746),
.B(n_641),
.Y(n_999)
);

OR2x2_ASAP7_75t_L g1000 ( 
.A(n_808),
.B(n_667),
.Y(n_1000)
);

AOI22xp33_ASAP7_75t_L g1001 ( 
.A1(n_761),
.A2(n_426),
.B1(n_445),
.B2(n_254),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_746),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_747),
.Y(n_1003)
);

BUFx5_ASAP7_75t_L g1004 ( 
.A(n_785),
.Y(n_1004)
);

AOI22xp33_ASAP7_75t_L g1005 ( 
.A1(n_785),
.A2(n_445),
.B1(n_254),
.B2(n_350),
.Y(n_1005)
);

AOI22xp5_ASAP7_75t_L g1006 ( 
.A1(n_782),
.A2(n_815),
.B1(n_825),
.B2(n_785),
.Y(n_1006)
);

AOI22xp33_ASAP7_75t_L g1007 ( 
.A1(n_785),
.A2(n_795),
.B1(n_736),
.B2(n_782),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_830),
.Y(n_1008)
);

NOR2xp33_ASAP7_75t_L g1009 ( 
.A(n_735),
.B(n_400),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_747),
.B(n_641),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_731),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_752),
.B(n_780),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_L g1013 ( 
.A(n_765),
.B(n_404),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_731),
.Y(n_1014)
);

AND2x4_ASAP7_75t_L g1015 ( 
.A(n_815),
.B(n_332),
.Y(n_1015)
);

OR2x2_ASAP7_75t_L g1016 ( 
.A(n_802),
.B(n_852),
.Y(n_1016)
);

INVxp67_ASAP7_75t_L g1017 ( 
.A(n_862),
.Y(n_1017)
);

A2O1A1Ixp33_ASAP7_75t_L g1018 ( 
.A1(n_752),
.A2(n_334),
.B(n_336),
.C(n_332),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_780),
.B(n_641),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_L g1020 ( 
.A(n_815),
.B(n_406),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_SL g1021 ( 
.A(n_781),
.B(n_295),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_SL g1022 ( 
.A(n_781),
.B(n_333),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_L g1023 ( 
.A(n_825),
.B(n_732),
.Y(n_1023)
);

INVx2_ASAP7_75t_SL g1024 ( 
.A(n_718),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_SL g1025 ( 
.A(n_783),
.B(n_333),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_748),
.Y(n_1026)
);

AND3x1_ASAP7_75t_L g1027 ( 
.A(n_708),
.B(n_336),
.C(n_334),
.Y(n_1027)
);

NOR2xp33_ASAP7_75t_L g1028 ( 
.A(n_825),
.B(n_407),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_L g1029 ( 
.A(n_783),
.B(n_409),
.Y(n_1029)
);

OAI22xp5_ASAP7_75t_L g1030 ( 
.A1(n_800),
.A2(n_415),
.B1(n_410),
.B2(n_417),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_SL g1031 ( 
.A(n_800),
.B(n_367),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_748),
.Y(n_1032)
);

NOR3xp33_ASAP7_75t_L g1033 ( 
.A(n_827),
.B(n_355),
.C(n_352),
.Y(n_1033)
);

AND2x2_ASAP7_75t_L g1034 ( 
.A(n_792),
.B(n_667),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_803),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_803),
.B(n_659),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_804),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_804),
.B(n_659),
.Y(n_1038)
);

BUFx3_ASAP7_75t_L g1039 ( 
.A(n_792),
.Y(n_1039)
);

INVx3_ASAP7_75t_L g1040 ( 
.A(n_717),
.Y(n_1040)
);

INVx2_ASAP7_75t_SL g1041 ( 
.A(n_792),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_865),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_798),
.B(n_773),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_890),
.Y(n_1044)
);

INVx1_ASAP7_75t_SL g1045 ( 
.A(n_887),
.Y(n_1045)
);

BUFx6f_ASAP7_75t_L g1046 ( 
.A(n_933),
.Y(n_1046)
);

AOI22xp33_ASAP7_75t_L g1047 ( 
.A1(n_902),
.A2(n_795),
.B1(n_785),
.B2(n_775),
.Y(n_1047)
);

INVx3_ASAP7_75t_L g1048 ( 
.A(n_933),
.Y(n_1048)
);

AND2x4_ASAP7_75t_L g1049 ( 
.A(n_882),
.B(n_811),
.Y(n_1049)
);

AND2x4_ASAP7_75t_L g1050 ( 
.A(n_882),
.B(n_828),
.Y(n_1050)
);

INVx3_ASAP7_75t_L g1051 ( 
.A(n_933),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_905),
.Y(n_1052)
);

AND2x4_ASAP7_75t_L g1053 ( 
.A(n_914),
.B(n_830),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_872),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_L g1055 ( 
.A(n_923),
.B(n_941),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_953),
.B(n_908),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_912),
.B(n_777),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_872),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_903),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_907),
.Y(n_1060)
);

BUFx3_ASAP7_75t_L g1061 ( 
.A(n_914),
.Y(n_1061)
);

AND2x2_ASAP7_75t_L g1062 ( 
.A(n_898),
.B(n_794),
.Y(n_1062)
);

OAI22xp5_ASAP7_75t_SL g1063 ( 
.A1(n_1023),
.A2(n_771),
.B1(n_788),
.B2(n_723),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_930),
.A2(n_720),
.B(n_856),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_918),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_919),
.Y(n_1066)
);

NOR3xp33_ASAP7_75t_SL g1067 ( 
.A(n_1008),
.B(n_422),
.C(n_421),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_920),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_927),
.Y(n_1069)
);

AND2x4_ASAP7_75t_L g1070 ( 
.A(n_933),
.B(n_720),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_891),
.B(n_785),
.Y(n_1071)
);

HB1xp67_ASAP7_75t_L g1072 ( 
.A(n_874),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_903),
.Y(n_1073)
);

BUFx2_ASAP7_75t_L g1074 ( 
.A(n_934),
.Y(n_1074)
);

NOR2xp33_ASAP7_75t_R g1075 ( 
.A(n_944),
.B(n_771),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_876),
.B(n_795),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_932),
.Y(n_1077)
);

BUFx6f_ASAP7_75t_L g1078 ( 
.A(n_961),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_917),
.Y(n_1079)
);

BUFx6f_ASAP7_75t_L g1080 ( 
.A(n_961),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_898),
.B(n_795),
.Y(n_1081)
);

AND2x4_ASAP7_75t_L g1082 ( 
.A(n_965),
.B(n_982),
.Y(n_1082)
);

AND2x4_ASAP7_75t_L g1083 ( 
.A(n_965),
.B(n_720),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_898),
.B(n_878),
.Y(n_1084)
);

OR2x6_ASAP7_75t_L g1085 ( 
.A(n_991),
.B(n_809),
.Y(n_1085)
);

INVx4_ASAP7_75t_L g1086 ( 
.A(n_877),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_913),
.B(n_795),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_917),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_951),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_921),
.Y(n_1090)
);

AND2x2_ASAP7_75t_L g1091 ( 
.A(n_1023),
.B(n_794),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_885),
.B(n_795),
.Y(n_1092)
);

BUFx6f_ASAP7_75t_L g1093 ( 
.A(n_961),
.Y(n_1093)
);

AND2x4_ASAP7_75t_L g1094 ( 
.A(n_982),
.B(n_1039),
.Y(n_1094)
);

AOI22xp33_ASAP7_75t_L g1095 ( 
.A1(n_904),
.A2(n_956),
.B1(n_1007),
.B2(n_970),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_951),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_1011),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_963),
.Y(n_1098)
);

BUFx2_ASAP7_75t_L g1099 ( 
.A(n_936),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_929),
.B(n_795),
.Y(n_1100)
);

BUFx2_ASAP7_75t_L g1101 ( 
.A(n_962),
.Y(n_1101)
);

NOR3xp33_ASAP7_75t_L g1102 ( 
.A(n_952),
.B(n_833),
.C(n_355),
.Y(n_1102)
);

NOR3xp33_ASAP7_75t_SL g1103 ( 
.A(n_995),
.B(n_433),
.C(n_430),
.Y(n_1103)
);

BUFx4f_ASAP7_75t_L g1104 ( 
.A(n_991),
.Y(n_1104)
);

CKINVDCx11_ASAP7_75t_R g1105 ( 
.A(n_897),
.Y(n_1105)
);

BUFx3_ASAP7_75t_L g1106 ( 
.A(n_921),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_1011),
.Y(n_1107)
);

NOR2xp33_ASAP7_75t_L g1108 ( 
.A(n_923),
.B(n_794),
.Y(n_1108)
);

NOR2xp33_ASAP7_75t_L g1109 ( 
.A(n_1017),
.B(n_788),
.Y(n_1109)
);

BUFx2_ASAP7_75t_L g1110 ( 
.A(n_989),
.Y(n_1110)
);

BUFx2_ASAP7_75t_L g1111 ( 
.A(n_1016),
.Y(n_1111)
);

INVx4_ASAP7_75t_L g1112 ( 
.A(n_877),
.Y(n_1112)
);

INVx5_ASAP7_75t_L g1113 ( 
.A(n_986),
.Y(n_1113)
);

BUFx10_ASAP7_75t_L g1114 ( 
.A(n_1041),
.Y(n_1114)
);

AOI22xp33_ASAP7_75t_L g1115 ( 
.A1(n_972),
.A2(n_851),
.B1(n_754),
.B2(n_755),
.Y(n_1115)
);

NOR3xp33_ASAP7_75t_SL g1116 ( 
.A(n_1020),
.B(n_439),
.C(n_437),
.Y(n_1116)
);

AND3x1_ASAP7_75t_SL g1117 ( 
.A(n_998),
.B(n_360),
.C(n_352),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_975),
.Y(n_1118)
);

AND2x4_ASAP7_75t_L g1119 ( 
.A(n_1039),
.B(n_826),
.Y(n_1119)
);

BUFx6f_ASAP7_75t_L g1120 ( 
.A(n_961),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_935),
.B(n_817),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_946),
.B(n_818),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_976),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_897),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_981),
.Y(n_1125)
);

HB1xp67_ASAP7_75t_L g1126 ( 
.A(n_1024),
.Y(n_1126)
);

BUFx3_ASAP7_75t_L g1127 ( 
.A(n_879),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_1014),
.Y(n_1128)
);

AND2x4_ASAP7_75t_L g1129 ( 
.A(n_1006),
.B(n_826),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_968),
.B(n_818),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_1014),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_1029),
.B(n_822),
.Y(n_1132)
);

HB1xp67_ASAP7_75t_L g1133 ( 
.A(n_1000),
.Y(n_1133)
);

AOI22xp5_ASAP7_75t_L g1134 ( 
.A1(n_893),
.A2(n_857),
.B1(n_816),
.B2(n_778),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_983),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1002),
.Y(n_1136)
);

BUFx2_ASAP7_75t_L g1137 ( 
.A(n_870),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1003),
.Y(n_1138)
);

INVx2_ASAP7_75t_SL g1139 ( 
.A(n_886),
.Y(n_1139)
);

BUFx3_ASAP7_75t_L g1140 ( 
.A(n_991),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_897),
.Y(n_1141)
);

HB1xp67_ASAP7_75t_L g1142 ( 
.A(n_947),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1035),
.Y(n_1143)
);

INVx5_ASAP7_75t_L g1144 ( 
.A(n_986),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_1029),
.B(n_822),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1037),
.Y(n_1146)
);

NOR2xp33_ASAP7_75t_R g1147 ( 
.A(n_896),
.B(n_851),
.Y(n_1147)
);

INVx2_ASAP7_75t_SL g1148 ( 
.A(n_868),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_926),
.B(n_836),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_957),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_SL g1151 ( 
.A(n_986),
.B(n_724),
.Y(n_1151)
);

AND2x2_ASAP7_75t_L g1152 ( 
.A(n_928),
.B(n_816),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_910),
.B(n_836),
.Y(n_1153)
);

INVx2_ASAP7_75t_L g1154 ( 
.A(n_1026),
.Y(n_1154)
);

NAND3xp33_ASAP7_75t_SL g1155 ( 
.A(n_869),
.B(n_443),
.C(n_441),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_967),
.B(n_840),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_875),
.B(n_840),
.Y(n_1157)
);

NAND3xp33_ASAP7_75t_SL g1158 ( 
.A(n_1033),
.B(n_958),
.C(n_993),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_911),
.B(n_846),
.Y(n_1159)
);

BUFx2_ASAP7_75t_L g1160 ( 
.A(n_1034),
.Y(n_1160)
);

NOR2xp33_ASAP7_75t_L g1161 ( 
.A(n_925),
.B(n_938),
.Y(n_1161)
);

INVx3_ASAP7_75t_L g1162 ( 
.A(n_877),
.Y(n_1162)
);

BUFx4f_ASAP7_75t_L g1163 ( 
.A(n_868),
.Y(n_1163)
);

INVx4_ASAP7_75t_L g1164 ( 
.A(n_979),
.Y(n_1164)
);

NOR3xp33_ASAP7_75t_SL g1165 ( 
.A(n_1020),
.B(n_454),
.C(n_444),
.Y(n_1165)
);

INVx6_ASAP7_75t_L g1166 ( 
.A(n_979),
.Y(n_1166)
);

BUFx3_ASAP7_75t_L g1167 ( 
.A(n_979),
.Y(n_1167)
);

BUFx6f_ASAP7_75t_L g1168 ( 
.A(n_979),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1012),
.Y(n_1169)
);

INVx2_ASAP7_75t_SL g1170 ( 
.A(n_980),
.Y(n_1170)
);

A2O1A1Ixp33_ASAP7_75t_L g1171 ( 
.A1(n_922),
.A2(n_368),
.B(n_378),
.C(n_360),
.Y(n_1171)
);

AND2x2_ASAP7_75t_L g1172 ( 
.A(n_1015),
.B(n_816),
.Y(n_1172)
);

NOR2xp33_ASAP7_75t_R g1173 ( 
.A(n_937),
.B(n_1009),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_SL g1174 ( 
.A(n_1004),
.B(n_949),
.Y(n_1174)
);

AND2x4_ASAP7_75t_L g1175 ( 
.A(n_924),
.B(n_826),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_992),
.Y(n_1176)
);

AND2x2_ASAP7_75t_L g1177 ( 
.A(n_1015),
.B(n_846),
.Y(n_1177)
);

AOI22xp5_ASAP7_75t_L g1178 ( 
.A1(n_892),
.A2(n_857),
.B1(n_778),
.B2(n_793),
.Y(n_1178)
);

NAND2x1p5_ASAP7_75t_L g1179 ( 
.A(n_980),
.B(n_856),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_1026),
.Y(n_1180)
);

NAND2xp33_ASAP7_75t_SL g1181 ( 
.A(n_881),
.B(n_763),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_1032),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_999),
.Y(n_1183)
);

AOI22xp33_ASAP7_75t_SL g1184 ( 
.A1(n_948),
.A2(n_461),
.B1(n_465),
.B2(n_459),
.Y(n_1184)
);

BUFx6f_ASAP7_75t_L g1185 ( 
.A(n_980),
.Y(n_1185)
);

INVx3_ASAP7_75t_L g1186 ( 
.A(n_994),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1010),
.Y(n_1187)
);

BUFx4f_ASAP7_75t_L g1188 ( 
.A(n_924),
.Y(n_1188)
);

INVx2_ASAP7_75t_SL g1189 ( 
.A(n_980),
.Y(n_1189)
);

BUFx6f_ASAP7_75t_L g1190 ( 
.A(n_1040),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1019),
.Y(n_1191)
);

INVxp67_ASAP7_75t_SL g1192 ( 
.A(n_984),
.Y(n_1192)
);

HB1xp67_ASAP7_75t_L g1193 ( 
.A(n_1015),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_924),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_911),
.B(n_866),
.Y(n_1195)
);

AND2x6_ASAP7_75t_L g1196 ( 
.A(n_1004),
.B(n_856),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_939),
.B(n_866),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1036),
.Y(n_1198)
);

AND2x2_ASAP7_75t_L g1199 ( 
.A(n_909),
.B(n_867),
.Y(n_1199)
);

AND2x4_ASAP7_75t_SL g1200 ( 
.A(n_948),
.B(n_763),
.Y(n_1200)
);

OAI22xp5_ASAP7_75t_L g1201 ( 
.A1(n_884),
.A2(n_759),
.B1(n_778),
.B2(n_763),
.Y(n_1201)
);

BUFx8_ASAP7_75t_L g1202 ( 
.A(n_880),
.Y(n_1202)
);

BUFx4f_ASAP7_75t_L g1203 ( 
.A(n_883),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_1032),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_939),
.B(n_759),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1042),
.B(n_751),
.Y(n_1206)
);

BUFx6f_ASAP7_75t_L g1207 ( 
.A(n_1040),
.Y(n_1207)
);

HB1xp67_ASAP7_75t_L g1208 ( 
.A(n_916),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1038),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_888),
.Y(n_1210)
);

AO22x1_ASAP7_75t_L g1211 ( 
.A1(n_1009),
.A2(n_368),
.B1(n_382),
.B2(n_378),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_942),
.Y(n_1212)
);

BUFx3_ASAP7_75t_L g1213 ( 
.A(n_889),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_895),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_925),
.B(n_751),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_899),
.Y(n_1216)
);

BUFx4f_ASAP7_75t_L g1217 ( 
.A(n_948),
.Y(n_1217)
);

CKINVDCx8_ASAP7_75t_R g1218 ( 
.A(n_1028),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1043),
.B(n_754),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_959),
.B(n_755),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1031),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_994),
.Y(n_1222)
);

INVxp33_ASAP7_75t_L g1223 ( 
.A(n_1028),
.Y(n_1223)
);

INVx3_ASAP7_75t_L g1224 ( 
.A(n_1004),
.Y(n_1224)
);

AND2x6_ASAP7_75t_SL g1225 ( 
.A(n_1013),
.B(n_382),
.Y(n_1225)
);

NOR3xp33_ASAP7_75t_SL g1226 ( 
.A(n_1030),
.B(n_469),
.C(n_468),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_1004),
.Y(n_1227)
);

INVx3_ASAP7_75t_SL g1228 ( 
.A(n_901),
.Y(n_1228)
);

INVx2_ASAP7_75t_SL g1229 ( 
.A(n_1004),
.Y(n_1229)
);

AND2x6_ASAP7_75t_L g1230 ( 
.A(n_1004),
.B(n_859),
.Y(n_1230)
);

AND2x4_ASAP7_75t_L g1231 ( 
.A(n_938),
.B(n_826),
.Y(n_1231)
);

INVx2_ASAP7_75t_L g1232 ( 
.A(n_1004),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_985),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_985),
.Y(n_1234)
);

BUFx6f_ASAP7_75t_L g1235 ( 
.A(n_950),
.Y(n_1235)
);

INVx4_ASAP7_75t_L g1236 ( 
.A(n_940),
.Y(n_1236)
);

BUFx3_ASAP7_75t_L g1237 ( 
.A(n_959),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1031),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1056),
.B(n_964),
.Y(n_1239)
);

INVxp67_ASAP7_75t_SL g1240 ( 
.A(n_1078),
.Y(n_1240)
);

OAI21x1_ASAP7_75t_L g1241 ( 
.A1(n_1212),
.A2(n_871),
.B(n_978),
.Y(n_1241)
);

OAI21x1_ASAP7_75t_L g1242 ( 
.A1(n_1212),
.A2(n_977),
.B(n_987),
.Y(n_1242)
);

OAI21xp33_ASAP7_75t_SL g1243 ( 
.A1(n_1169),
.A2(n_943),
.B(n_900),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1084),
.B(n_1169),
.Y(n_1244)
);

NOR2xp33_ASAP7_75t_L g1245 ( 
.A(n_1223),
.B(n_894),
.Y(n_1245)
);

OAI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1205),
.A2(n_931),
.B(n_930),
.Y(n_1246)
);

BUFx2_ASAP7_75t_L g1247 ( 
.A(n_1075),
.Y(n_1247)
);

AOI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1132),
.A2(n_931),
.B(n_943),
.Y(n_1248)
);

AND2x2_ASAP7_75t_L g1249 ( 
.A(n_1137),
.B(n_1027),
.Y(n_1249)
);

AOI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1145),
.A2(n_973),
.B(n_950),
.Y(n_1250)
);

INVx3_ASAP7_75t_L g1251 ( 
.A(n_1086),
.Y(n_1251)
);

INVx5_ASAP7_75t_L g1252 ( 
.A(n_1046),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1052),
.Y(n_1253)
);

INVx1_ASAP7_75t_SL g1254 ( 
.A(n_1045),
.Y(n_1254)
);

BUFx2_ASAP7_75t_L g1255 ( 
.A(n_1074),
.Y(n_1255)
);

AOI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_1153),
.A2(n_973),
.B(n_900),
.Y(n_1256)
);

OAI21x1_ASAP7_75t_L g1257 ( 
.A1(n_1064),
.A2(n_977),
.B(n_987),
.Y(n_1257)
);

INVx3_ASAP7_75t_SL g1258 ( 
.A(n_1090),
.Y(n_1258)
);

A2O1A1Ixp33_ASAP7_75t_L g1259 ( 
.A1(n_1161),
.A2(n_1237),
.B(n_1223),
.C(n_1171),
.Y(n_1259)
);

BUFx6f_ASAP7_75t_L g1260 ( 
.A(n_1078),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1091),
.B(n_964),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_SL g1262 ( 
.A1(n_1229),
.A2(n_894),
.B(n_906),
.Y(n_1262)
);

INVx2_ASAP7_75t_L g1263 ( 
.A(n_1054),
.Y(n_1263)
);

AOI21x1_ASAP7_75t_L g1264 ( 
.A1(n_1220),
.A2(n_1022),
.B(n_1021),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_SL g1265 ( 
.A(n_1237),
.B(n_1113),
.Y(n_1265)
);

OAI21x1_ASAP7_75t_L g1266 ( 
.A1(n_1224),
.A2(n_1022),
.B(n_1021),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1060),
.Y(n_1267)
);

BUFx6f_ASAP7_75t_L g1268 ( 
.A(n_1078),
.Y(n_1268)
);

AND2x4_ASAP7_75t_L g1269 ( 
.A(n_1140),
.B(n_945),
.Y(n_1269)
);

AO31x2_ASAP7_75t_L g1270 ( 
.A1(n_1201),
.A2(n_1171),
.A3(n_1018),
.B(n_990),
.Y(n_1270)
);

INVx5_ASAP7_75t_L g1271 ( 
.A(n_1046),
.Y(n_1271)
);

OAI21x1_ASAP7_75t_L g1272 ( 
.A1(n_1174),
.A2(n_1025),
.B(n_996),
.Y(n_1272)
);

AOI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1057),
.A2(n_960),
.B(n_988),
.Y(n_1273)
);

NOR2xp33_ASAP7_75t_L g1274 ( 
.A(n_1091),
.B(n_988),
.Y(n_1274)
);

OA21x2_ASAP7_75t_L g1275 ( 
.A1(n_1152),
.A2(n_1025),
.B(n_1018),
.Y(n_1275)
);

NOR2xp33_ASAP7_75t_L g1276 ( 
.A(n_1218),
.B(n_997),
.Y(n_1276)
);

BUFx12f_ASAP7_75t_L g1277 ( 
.A(n_1105),
.Y(n_1277)
);

AO31x2_ASAP7_75t_L g1278 ( 
.A1(n_1159),
.A2(n_990),
.A3(n_966),
.B(n_960),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1065),
.Y(n_1279)
);

OA21x2_ASAP7_75t_L g1280 ( 
.A1(n_1152),
.A2(n_787),
.B(n_764),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1066),
.Y(n_1281)
);

OAI21xp33_ASAP7_75t_L g1282 ( 
.A1(n_1109),
.A2(n_966),
.B(n_873),
.Y(n_1282)
);

BUFx6f_ASAP7_75t_L g1283 ( 
.A(n_1078),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1137),
.B(n_1150),
.Y(n_1284)
);

OAI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1092),
.A2(n_1076),
.B(n_1087),
.Y(n_1285)
);

NOR2xp67_ASAP7_75t_L g1286 ( 
.A(n_1044),
.B(n_997),
.Y(n_1286)
);

BUFx6f_ASAP7_75t_L g1287 ( 
.A(n_1078),
.Y(n_1287)
);

AOI21xp33_ASAP7_75t_L g1288 ( 
.A1(n_1095),
.A2(n_1013),
.B(n_955),
.Y(n_1288)
);

AOI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1219),
.A2(n_1157),
.B(n_1163),
.Y(n_1289)
);

OAI21x1_ASAP7_75t_L g1290 ( 
.A1(n_1224),
.A2(n_859),
.B(n_787),
.Y(n_1290)
);

INVx4_ASAP7_75t_L g1291 ( 
.A(n_1119),
.Y(n_1291)
);

OAI21x1_ASAP7_75t_L g1292 ( 
.A1(n_1224),
.A2(n_859),
.B(n_801),
.Y(n_1292)
);

AOI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1163),
.A2(n_1149),
.B(n_1144),
.Y(n_1293)
);

OAI22xp5_ASAP7_75t_L g1294 ( 
.A1(n_1192),
.A2(n_954),
.B1(n_974),
.B2(n_971),
.Y(n_1294)
);

AOI221x1_ASAP7_75t_L g1295 ( 
.A1(n_1181),
.A2(n_420),
.B1(n_423),
.B2(n_427),
.C(n_394),
.Y(n_1295)
);

AOI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_1163),
.A2(n_834),
.B(n_793),
.Y(n_1296)
);

AOI22xp33_ASAP7_75t_L g1297 ( 
.A1(n_1236),
.A2(n_1001),
.B1(n_1005),
.B2(n_387),
.Y(n_1297)
);

OAI22xp5_ASAP7_75t_L g1298 ( 
.A1(n_1086),
.A2(n_915),
.B1(n_387),
.B2(n_398),
.Y(n_1298)
);

AO31x2_ASAP7_75t_L g1299 ( 
.A1(n_1195),
.A2(n_764),
.A3(n_813),
.B(n_801),
.Y(n_1299)
);

NOR2xp33_ASAP7_75t_L g1300 ( 
.A(n_1218),
.B(n_969),
.Y(n_1300)
);

NAND2x1_ASAP7_75t_L g1301 ( 
.A(n_1086),
.B(n_857),
.Y(n_1301)
);

AO31x2_ASAP7_75t_L g1302 ( 
.A1(n_1197),
.A2(n_819),
.A3(n_867),
.B(n_835),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1054),
.Y(n_1303)
);

AO31x2_ASAP7_75t_L g1304 ( 
.A1(n_1221),
.A2(n_838),
.A3(n_819),
.B(n_832),
.Y(n_1304)
);

OAI21x1_ASAP7_75t_L g1305 ( 
.A1(n_1227),
.A2(n_832),
.B(n_813),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1177),
.B(n_835),
.Y(n_1306)
);

HB1xp67_ASAP7_75t_L g1307 ( 
.A(n_1072),
.Y(n_1307)
);

AO31x2_ASAP7_75t_L g1308 ( 
.A1(n_1233),
.A2(n_850),
.A3(n_838),
.B(n_839),
.Y(n_1308)
);

INVx5_ASAP7_75t_L g1309 ( 
.A(n_1046),
.Y(n_1309)
);

AO31x2_ASAP7_75t_L g1310 ( 
.A1(n_1234),
.A2(n_850),
.A3(n_839),
.B(n_700),
.Y(n_1310)
);

AOI21xp5_ASAP7_75t_L g1311 ( 
.A1(n_1113),
.A2(n_1144),
.B(n_1181),
.Y(n_1311)
);

BUFx6f_ASAP7_75t_L g1312 ( 
.A(n_1080),
.Y(n_1312)
);

A2O1A1Ixp33_ASAP7_75t_L g1313 ( 
.A1(n_1130),
.A2(n_427),
.B(n_457),
.C(n_452),
.Y(n_1313)
);

OAI21xp5_ASAP7_75t_L g1314 ( 
.A1(n_1100),
.A2(n_834),
.B(n_793),
.Y(n_1314)
);

OAI21x1_ASAP7_75t_L g1315 ( 
.A1(n_1174),
.A2(n_660),
.B(n_659),
.Y(n_1315)
);

OAI21x1_ASAP7_75t_L g1316 ( 
.A1(n_1227),
.A2(n_660),
.B(n_659),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1177),
.B(n_834),
.Y(n_1317)
);

AO31x2_ASAP7_75t_L g1318 ( 
.A1(n_1238),
.A2(n_1058),
.A3(n_1073),
.B(n_1059),
.Y(n_1318)
);

AOI21xp5_ASAP7_75t_SL g1319 ( 
.A1(n_1229),
.A2(n_849),
.B(n_727),
.Y(n_1319)
);

AOI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1113),
.A2(n_864),
.B(n_727),
.Y(n_1320)
);

OAI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1134),
.A2(n_864),
.B(n_849),
.Y(n_1321)
);

BUFx12f_ASAP7_75t_L g1322 ( 
.A(n_1105),
.Y(n_1322)
);

AOI22xp5_ASAP7_75t_L g1323 ( 
.A1(n_1158),
.A2(n_472),
.B1(n_471),
.B2(n_857),
.Y(n_1323)
);

AND2x2_ASAP7_75t_SL g1324 ( 
.A(n_1188),
.B(n_901),
.Y(n_1324)
);

OA21x2_ASAP7_75t_L g1325 ( 
.A1(n_1172),
.A2(n_597),
.B(n_563),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1068),
.Y(n_1326)
);

BUFx3_ASAP7_75t_L g1327 ( 
.A(n_1140),
.Y(n_1327)
);

BUFx3_ASAP7_75t_L g1328 ( 
.A(n_1104),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1058),
.Y(n_1329)
);

INVx2_ASAP7_75t_SL g1330 ( 
.A(n_1106),
.Y(n_1330)
);

OAI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1071),
.A2(n_864),
.B(n_722),
.Y(n_1331)
);

OAI22xp5_ASAP7_75t_L g1332 ( 
.A1(n_1112),
.A2(n_423),
.B1(n_452),
.B2(n_457),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1062),
.B(n_394),
.Y(n_1333)
);

AO31x2_ASAP7_75t_L g1334 ( 
.A1(n_1059),
.A2(n_563),
.A3(n_597),
.B(n_367),
.Y(n_1334)
);

HB1xp67_ASAP7_75t_L g1335 ( 
.A(n_1193),
.Y(n_1335)
);

OAI22xp5_ASAP7_75t_L g1336 ( 
.A1(n_1112),
.A2(n_450),
.B1(n_449),
.B2(n_446),
.Y(n_1336)
);

AOI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1113),
.A2(n_727),
.B(n_724),
.Y(n_1337)
);

OAI21x1_ASAP7_75t_L g1338 ( 
.A1(n_1232),
.A2(n_660),
.B(n_659),
.Y(n_1338)
);

OAI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1215),
.A2(n_722),
.B(n_705),
.Y(n_1339)
);

AOI21xp5_ASAP7_75t_L g1340 ( 
.A1(n_1113),
.A2(n_729),
.B(n_727),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1069),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1062),
.B(n_398),
.Y(n_1342)
);

AOI21xp5_ASAP7_75t_L g1343 ( 
.A1(n_1144),
.A2(n_729),
.B(n_727),
.Y(n_1343)
);

AOI21x1_ASAP7_75t_L g1344 ( 
.A1(n_1151),
.A2(n_597),
.B(n_563),
.Y(n_1344)
);

OAI21x1_ASAP7_75t_L g1345 ( 
.A1(n_1232),
.A2(n_1179),
.B(n_1151),
.Y(n_1345)
);

OR2x2_ASAP7_75t_L g1346 ( 
.A(n_1142),
.B(n_420),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1108),
.B(n_435),
.Y(n_1347)
);

AO31x2_ASAP7_75t_L g1348 ( 
.A1(n_1073),
.A2(n_467),
.A3(n_464),
.B(n_470),
.Y(n_1348)
);

AOI21xp5_ASAP7_75t_L g1349 ( 
.A1(n_1144),
.A2(n_753),
.B(n_729),
.Y(n_1349)
);

OAI21x1_ASAP7_75t_L g1350 ( 
.A1(n_1179),
.A2(n_660),
.B(n_467),
.Y(n_1350)
);

OAI21x1_ASAP7_75t_L g1351 ( 
.A1(n_1179),
.A2(n_660),
.B(n_446),
.Y(n_1351)
);

HB1xp67_ASAP7_75t_L g1352 ( 
.A(n_1074),
.Y(n_1352)
);

OAI21x1_ASAP7_75t_L g1353 ( 
.A1(n_1206),
.A2(n_449),
.B(n_435),
.Y(n_1353)
);

AOI21xp33_ASAP7_75t_L g1354 ( 
.A1(n_1047),
.A2(n_464),
.B(n_450),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1098),
.B(n_470),
.Y(n_1355)
);

AND2x4_ASAP7_75t_L g1356 ( 
.A(n_1082),
.B(n_729),
.Y(n_1356)
);

BUFx6f_ASAP7_75t_L g1357 ( 
.A(n_1080),
.Y(n_1357)
);

O2A1O1Ixp5_ASAP7_75t_L g1358 ( 
.A1(n_1211),
.A2(n_1098),
.B(n_1183),
.C(n_1176),
.Y(n_1358)
);

CKINVDCx5p33_ASAP7_75t_R g1359 ( 
.A(n_1044),
.Y(n_1359)
);

OAI21x1_ASAP7_75t_L g1360 ( 
.A1(n_1079),
.A2(n_473),
.B(n_413),
.Y(n_1360)
);

AOI21xp5_ASAP7_75t_SL g1361 ( 
.A1(n_1112),
.A2(n_854),
.B(n_753),
.Y(n_1361)
);

A2O1A1Ixp33_ASAP7_75t_L g1362 ( 
.A1(n_1156),
.A2(n_473),
.B(n_413),
.C(n_366),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1101),
.B(n_311),
.Y(n_1363)
);

AO21x1_ASAP7_75t_L g1364 ( 
.A1(n_1172),
.A2(n_335),
.B(n_655),
.Y(n_1364)
);

OAI21x1_ASAP7_75t_L g1365 ( 
.A1(n_1079),
.A2(n_753),
.B(n_729),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1077),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1118),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1101),
.B(n_350),
.Y(n_1368)
);

OR2x6_ASAP7_75t_L g1369 ( 
.A(n_1106),
.B(n_753),
.Y(n_1369)
);

OAI22xp5_ASAP7_75t_L g1370 ( 
.A1(n_1236),
.A2(n_1081),
.B1(n_1125),
.B2(n_1123),
.Y(n_1370)
);

OAI21xp33_ASAP7_75t_L g1371 ( 
.A1(n_1055),
.A2(n_381),
.B(n_350),
.Y(n_1371)
);

AOI21xp5_ASAP7_75t_L g1372 ( 
.A1(n_1144),
.A2(n_790),
.B(n_753),
.Y(n_1372)
);

INVxp67_ASAP7_75t_SL g1373 ( 
.A(n_1080),
.Y(n_1373)
);

AO31x2_ASAP7_75t_L g1374 ( 
.A1(n_1088),
.A2(n_680),
.A3(n_655),
.B(n_677),
.Y(n_1374)
);

OAI21x1_ASAP7_75t_L g1375 ( 
.A1(n_1088),
.A2(n_791),
.B(n_790),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1089),
.Y(n_1376)
);

OAI21x1_ASAP7_75t_L g1377 ( 
.A1(n_1089),
.A2(n_1097),
.B(n_1096),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_SL g1378 ( 
.A(n_1235),
.B(n_790),
.Y(n_1378)
);

NOR2xp67_ASAP7_75t_SL g1379 ( 
.A(n_1090),
.B(n_350),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1211),
.B(n_790),
.Y(n_1380)
);

NAND2x1p5_ASAP7_75t_L g1381 ( 
.A(n_1104),
.B(n_705),
.Y(n_1381)
);

AND2x4_ASAP7_75t_L g1382 ( 
.A(n_1082),
.B(n_790),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1135),
.B(n_791),
.Y(n_1383)
);

OAI21x1_ASAP7_75t_L g1384 ( 
.A1(n_1096),
.A2(n_824),
.B(n_791),
.Y(n_1384)
);

OAI21x1_ASAP7_75t_SL g1385 ( 
.A1(n_1164),
.A2(n_8),
.B(n_9),
.Y(n_1385)
);

AND3x4_ASAP7_75t_L g1386 ( 
.A(n_1102),
.B(n_11),
.C(n_13),
.Y(n_1386)
);

INVx2_ASAP7_75t_L g1387 ( 
.A(n_1097),
.Y(n_1387)
);

OA21x2_ASAP7_75t_L g1388 ( 
.A1(n_1107),
.A2(n_288),
.B(n_272),
.Y(n_1388)
);

A2O1A1Ixp33_ASAP7_75t_L g1389 ( 
.A1(n_1199),
.A2(n_350),
.B(n_381),
.C(n_429),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1136),
.B(n_791),
.Y(n_1390)
);

AOI21xp5_ASAP7_75t_SL g1391 ( 
.A1(n_1046),
.A2(n_1129),
.B(n_1070),
.Y(n_1391)
);

AOI21xp5_ASAP7_75t_L g1392 ( 
.A1(n_1187),
.A2(n_824),
.B(n_791),
.Y(n_1392)
);

INVx3_ASAP7_75t_SL g1393 ( 
.A(n_1124),
.Y(n_1393)
);

BUFx6f_ASAP7_75t_L g1394 ( 
.A(n_1080),
.Y(n_1394)
);

OAI21xp5_ASAP7_75t_L g1395 ( 
.A1(n_1191),
.A2(n_722),
.B(n_705),
.Y(n_1395)
);

BUFx4f_ASAP7_75t_L g1396 ( 
.A(n_1053),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1138),
.B(n_824),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1111),
.B(n_350),
.Y(n_1398)
);

OAI21x1_ASAP7_75t_L g1399 ( 
.A1(n_1107),
.A2(n_837),
.B(n_824),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1143),
.Y(n_1400)
);

AO21x1_ASAP7_75t_L g1401 ( 
.A1(n_1199),
.A2(n_677),
.B(n_655),
.Y(n_1401)
);

OAI21x1_ASAP7_75t_L g1402 ( 
.A1(n_1128),
.A2(n_837),
.B(n_824),
.Y(n_1402)
);

OAI21xp5_ASAP7_75t_L g1403 ( 
.A1(n_1198),
.A2(n_1209),
.B(n_1122),
.Y(n_1403)
);

OAI21xp5_ASAP7_75t_L g1404 ( 
.A1(n_1121),
.A2(n_1178),
.B(n_1146),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1210),
.Y(n_1405)
);

A2O1A1Ixp33_ASAP7_75t_L g1406 ( 
.A1(n_1155),
.A2(n_381),
.B(n_429),
.C(n_466),
.Y(n_1406)
);

OAI21x1_ASAP7_75t_L g1407 ( 
.A1(n_1128),
.A2(n_854),
.B(n_837),
.Y(n_1407)
);

AOI21xp5_ASAP7_75t_L g1408 ( 
.A1(n_1162),
.A2(n_854),
.B(n_837),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1111),
.B(n_837),
.Y(n_1409)
);

AND2x4_ASAP7_75t_L g1410 ( 
.A(n_1291),
.B(n_1129),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1318),
.Y(n_1411)
);

CKINVDCx5p33_ASAP7_75t_R g1412 ( 
.A(n_1359),
.Y(n_1412)
);

AOI21xp5_ASAP7_75t_L g1413 ( 
.A1(n_1273),
.A2(n_1239),
.B(n_1289),
.Y(n_1413)
);

AOI22xp33_ASAP7_75t_SL g1414 ( 
.A1(n_1274),
.A2(n_1173),
.B1(n_1063),
.B2(n_1236),
.Y(n_1414)
);

OAI221xp5_ASAP7_75t_L g1415 ( 
.A1(n_1282),
.A2(n_1184),
.B1(n_1110),
.B2(n_1226),
.C(n_1160),
.Y(n_1415)
);

OAI21x1_ASAP7_75t_SL g1416 ( 
.A1(n_1246),
.A2(n_1285),
.B(n_1403),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1318),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_1318),
.Y(n_1418)
);

BUFx12f_ASAP7_75t_L g1419 ( 
.A(n_1277),
.Y(n_1419)
);

OR2x6_ASAP7_75t_L g1420 ( 
.A(n_1391),
.B(n_1129),
.Y(n_1420)
);

OAI21x1_ASAP7_75t_L g1421 ( 
.A1(n_1241),
.A2(n_1154),
.B(n_1131),
.Y(n_1421)
);

OA21x2_ASAP7_75t_L g1422 ( 
.A1(n_1401),
.A2(n_1154),
.B(n_1131),
.Y(n_1422)
);

AOI22xp5_ASAP7_75t_L g1423 ( 
.A1(n_1274),
.A2(n_1110),
.B1(n_1133),
.B2(n_1160),
.Y(n_1423)
);

AOI22xp33_ASAP7_75t_L g1424 ( 
.A1(n_1288),
.A2(n_1217),
.B1(n_1188),
.B2(n_1228),
.Y(n_1424)
);

OAI21x1_ASAP7_75t_L g1425 ( 
.A1(n_1375),
.A2(n_1182),
.B(n_1180),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1318),
.Y(n_1426)
);

A2O1A1Ixp33_ASAP7_75t_L g1427 ( 
.A1(n_1276),
.A2(n_1261),
.B(n_1243),
.C(n_1358),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1263),
.Y(n_1428)
);

AOI21xp5_ASAP7_75t_L g1429 ( 
.A1(n_1293),
.A2(n_1162),
.B(n_1186),
.Y(n_1429)
);

BUFx6f_ASAP7_75t_L g1430 ( 
.A(n_1260),
.Y(n_1430)
);

A2O1A1Ixp33_ASAP7_75t_L g1431 ( 
.A1(n_1276),
.A2(n_1203),
.B(n_1116),
.C(n_1165),
.Y(n_1431)
);

OAI21x1_ASAP7_75t_L g1432 ( 
.A1(n_1375),
.A2(n_1182),
.B(n_1180),
.Y(n_1432)
);

NAND2x1p5_ASAP7_75t_L g1433 ( 
.A(n_1252),
.B(n_1235),
.Y(n_1433)
);

INVx1_ASAP7_75t_SL g1434 ( 
.A(n_1254),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1244),
.B(n_1099),
.Y(n_1435)
);

OAI221xp5_ASAP7_75t_L g1436 ( 
.A1(n_1323),
.A2(n_1347),
.B1(n_1286),
.B2(n_1245),
.C(n_1313),
.Y(n_1436)
);

AND2x4_ASAP7_75t_L g1437 ( 
.A(n_1291),
.B(n_1356),
.Y(n_1437)
);

AOI21xp5_ASAP7_75t_L g1438 ( 
.A1(n_1361),
.A2(n_1162),
.B(n_1186),
.Y(n_1438)
);

OAI21x1_ASAP7_75t_L g1439 ( 
.A1(n_1399),
.A2(n_1204),
.B(n_1186),
.Y(n_1439)
);

BUFx4f_ASAP7_75t_SL g1440 ( 
.A(n_1277),
.Y(n_1440)
);

OAI21xp5_ASAP7_75t_L g1441 ( 
.A1(n_1250),
.A2(n_1070),
.B(n_1214),
.Y(n_1441)
);

OR2x6_ASAP7_75t_L g1442 ( 
.A(n_1319),
.B(n_1235),
.Y(n_1442)
);

OAI21x1_ASAP7_75t_L g1443 ( 
.A1(n_1399),
.A2(n_1204),
.B(n_1051),
.Y(n_1443)
);

OAI21xp5_ASAP7_75t_L g1444 ( 
.A1(n_1256),
.A2(n_1070),
.B(n_1216),
.Y(n_1444)
);

OAI21x1_ASAP7_75t_L g1445 ( 
.A1(n_1257),
.A2(n_1051),
.B(n_1048),
.Y(n_1445)
);

INVx2_ASAP7_75t_L g1446 ( 
.A(n_1263),
.Y(n_1446)
);

OAI21xp5_ASAP7_75t_L g1447 ( 
.A1(n_1358),
.A2(n_1203),
.B(n_1148),
.Y(n_1447)
);

AND2x4_ASAP7_75t_L g1448 ( 
.A(n_1356),
.B(n_1164),
.Y(n_1448)
);

OR2x6_ASAP7_75t_L g1449 ( 
.A(n_1265),
.B(n_1235),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1245),
.B(n_1099),
.Y(n_1450)
);

OAI22xp5_ASAP7_75t_L g1451 ( 
.A1(n_1396),
.A2(n_1053),
.B1(n_1203),
.B2(n_1124),
.Y(n_1451)
);

AO21x2_ASAP7_75t_L g1452 ( 
.A1(n_1364),
.A2(n_1222),
.B(n_1231),
.Y(n_1452)
);

OR2x6_ASAP7_75t_L g1453 ( 
.A(n_1265),
.B(n_1235),
.Y(n_1453)
);

OAI21xp5_ASAP7_75t_L g1454 ( 
.A1(n_1404),
.A2(n_1148),
.B(n_1083),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1304),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1284),
.B(n_1126),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1307),
.B(n_1053),
.Y(n_1457)
);

AO21x2_ASAP7_75t_L g1458 ( 
.A1(n_1389),
.A2(n_1222),
.B(n_1231),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1304),
.Y(n_1459)
);

OAI21x1_ASAP7_75t_L g1460 ( 
.A1(n_1315),
.A2(n_1051),
.B(n_1048),
.Y(n_1460)
);

NOR2xp33_ASAP7_75t_L g1461 ( 
.A(n_1300),
.B(n_1228),
.Y(n_1461)
);

AND2x4_ASAP7_75t_L g1462 ( 
.A(n_1356),
.B(n_1164),
.Y(n_1462)
);

O2A1O1Ixp33_ASAP7_75t_L g1463 ( 
.A1(n_1259),
.A2(n_1208),
.B(n_1103),
.C(n_1067),
.Y(n_1463)
);

AOI221xp5_ASAP7_75t_L g1464 ( 
.A1(n_1313),
.A2(n_1225),
.B1(n_1147),
.B2(n_1050),
.C(n_1049),
.Y(n_1464)
);

NAND2x1p5_ASAP7_75t_L g1465 ( 
.A(n_1252),
.B(n_1167),
.Y(n_1465)
);

OAI21x1_ASAP7_75t_L g1466 ( 
.A1(n_1315),
.A2(n_1048),
.B(n_1115),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1304),
.Y(n_1467)
);

AOI21xp5_ASAP7_75t_L g1468 ( 
.A1(n_1311),
.A2(n_1189),
.B(n_1170),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1304),
.Y(n_1469)
);

OAI21x1_ASAP7_75t_L g1470 ( 
.A1(n_1350),
.A2(n_1230),
.B(n_1196),
.Y(n_1470)
);

AOI21x1_ASAP7_75t_L g1471 ( 
.A1(n_1378),
.A2(n_1231),
.B(n_1189),
.Y(n_1471)
);

OAI22xp33_ASAP7_75t_L g1472 ( 
.A1(n_1396),
.A2(n_1141),
.B1(n_1188),
.B2(n_1085),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1308),
.Y(n_1473)
);

NOR2xp33_ASAP7_75t_L g1474 ( 
.A(n_1300),
.B(n_1255),
.Y(n_1474)
);

OA21x2_ASAP7_75t_L g1475 ( 
.A1(n_1389),
.A2(n_1242),
.B(n_1360),
.Y(n_1475)
);

OAI22xp33_ASAP7_75t_L g1476 ( 
.A1(n_1333),
.A2(n_1141),
.B1(n_1085),
.B2(n_1217),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1307),
.B(n_1127),
.Y(n_1477)
);

OAI21x1_ASAP7_75t_L g1478 ( 
.A1(n_1350),
.A2(n_1230),
.B(n_1196),
.Y(n_1478)
);

OA21x2_ASAP7_75t_L g1479 ( 
.A1(n_1272),
.A2(n_1139),
.B(n_1170),
.Y(n_1479)
);

BUFx3_ASAP7_75t_L g1480 ( 
.A(n_1328),
.Y(n_1480)
);

AND2x4_ASAP7_75t_L g1481 ( 
.A(n_1382),
.B(n_1167),
.Y(n_1481)
);

OAI21x1_ASAP7_75t_L g1482 ( 
.A1(n_1365),
.A2(n_1230),
.B(n_1196),
.Y(n_1482)
);

OAI21xp5_ASAP7_75t_L g1483 ( 
.A1(n_1248),
.A2(n_1083),
.B(n_1196),
.Y(n_1483)
);

CKINVDCx20_ASAP7_75t_R g1484 ( 
.A(n_1359),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1249),
.B(n_1213),
.Y(n_1485)
);

BUFx2_ASAP7_75t_L g1486 ( 
.A(n_1240),
.Y(n_1486)
);

AO21x2_ASAP7_75t_L g1487 ( 
.A1(n_1321),
.A2(n_1175),
.B(n_1049),
.Y(n_1487)
);

OAI21x1_ASAP7_75t_SL g1488 ( 
.A1(n_1395),
.A2(n_1139),
.B(n_1196),
.Y(n_1488)
);

OAI21xp5_ASAP7_75t_L g1489 ( 
.A1(n_1259),
.A2(n_1230),
.B(n_1196),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_1303),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1308),
.Y(n_1491)
);

INVx3_ASAP7_75t_L g1492 ( 
.A(n_1260),
.Y(n_1492)
);

NOR2xp33_ASAP7_75t_L g1493 ( 
.A(n_1352),
.B(n_1049),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1308),
.Y(n_1494)
);

INVx4_ASAP7_75t_L g1495 ( 
.A(n_1252),
.Y(n_1495)
);

OAI21x1_ASAP7_75t_L g1496 ( 
.A1(n_1384),
.A2(n_1230),
.B(n_1093),
.Y(n_1496)
);

AOI22xp5_ASAP7_75t_L g1497 ( 
.A1(n_1386),
.A2(n_1050),
.B1(n_1085),
.B2(n_1117),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_SL g1498 ( 
.A(n_1294),
.B(n_1082),
.Y(n_1498)
);

OAI21x1_ASAP7_75t_L g1499 ( 
.A1(n_1402),
.A2(n_1230),
.B(n_1093),
.Y(n_1499)
);

HB1xp67_ASAP7_75t_L g1500 ( 
.A(n_1352),
.Y(n_1500)
);

AOI22xp33_ASAP7_75t_L g1501 ( 
.A1(n_1354),
.A2(n_1217),
.B1(n_1050),
.B2(n_1213),
.Y(n_1501)
);

OAI22xp5_ASAP7_75t_L g1502 ( 
.A1(n_1297),
.A2(n_1083),
.B1(n_1094),
.B2(n_1061),
.Y(n_1502)
);

AO21x1_ASAP7_75t_L g1503 ( 
.A1(n_1370),
.A2(n_1200),
.B(n_1175),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1303),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1329),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_1329),
.Y(n_1506)
);

OAI21xp5_ASAP7_75t_L g1507 ( 
.A1(n_1272),
.A2(n_1094),
.B(n_1119),
.Y(n_1507)
);

BUFx3_ASAP7_75t_L g1508 ( 
.A(n_1328),
.Y(n_1508)
);

OAI21x1_ASAP7_75t_L g1509 ( 
.A1(n_1407),
.A2(n_1093),
.B(n_1080),
.Y(n_1509)
);

OAI21x1_ASAP7_75t_L g1510 ( 
.A1(n_1290),
.A2(n_1120),
.B(n_1093),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1308),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1335),
.B(n_1127),
.Y(n_1512)
);

OAI21x1_ASAP7_75t_L g1513 ( 
.A1(n_1292),
.A2(n_1345),
.B(n_1392),
.Y(n_1513)
);

OAI22xp5_ASAP7_75t_L g1514 ( 
.A1(n_1297),
.A2(n_1094),
.B1(n_1061),
.B2(n_1085),
.Y(n_1514)
);

AOI221x1_ASAP7_75t_L g1515 ( 
.A1(n_1371),
.A2(n_1185),
.B1(n_1093),
.B2(n_1168),
.C(n_1120),
.Y(n_1515)
);

AO21x2_ASAP7_75t_L g1516 ( 
.A1(n_1378),
.A2(n_1175),
.B(n_1119),
.Y(n_1516)
);

BUFx6f_ASAP7_75t_L g1517 ( 
.A(n_1260),
.Y(n_1517)
);

INVx2_ASAP7_75t_SL g1518 ( 
.A(n_1252),
.Y(n_1518)
);

NOR2xp33_ASAP7_75t_L g1519 ( 
.A(n_1335),
.B(n_1194),
.Y(n_1519)
);

AOI21x1_ASAP7_75t_L g1520 ( 
.A1(n_1344),
.A2(n_1168),
.B(n_1120),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1247),
.B(n_1194),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1376),
.Y(n_1522)
);

AOI22xp33_ASAP7_75t_L g1523 ( 
.A1(n_1324),
.A2(n_1202),
.B1(n_1200),
.B2(n_1104),
.Y(n_1523)
);

INVx3_ASAP7_75t_L g1524 ( 
.A(n_1260),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1376),
.Y(n_1525)
);

AOI22xp33_ASAP7_75t_L g1526 ( 
.A1(n_1324),
.A2(n_1202),
.B1(n_1207),
.B2(n_1190),
.Y(n_1526)
);

OAI21x1_ASAP7_75t_L g1527 ( 
.A1(n_1345),
.A2(n_1168),
.B(n_1120),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1387),
.Y(n_1528)
);

OAI21x1_ASAP7_75t_L g1529 ( 
.A1(n_1305),
.A2(n_1168),
.B(n_1120),
.Y(n_1529)
);

BUFx2_ASAP7_75t_L g1530 ( 
.A(n_1240),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1269),
.B(n_1190),
.Y(n_1531)
);

BUFx6f_ASAP7_75t_L g1532 ( 
.A(n_1268),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1387),
.Y(n_1533)
);

INVxp67_ASAP7_75t_SL g1534 ( 
.A(n_1409),
.Y(n_1534)
);

O2A1O1Ixp33_ASAP7_75t_L g1535 ( 
.A1(n_1406),
.A2(n_1114),
.B(n_1202),
.C(n_1190),
.Y(n_1535)
);

OAI21x1_ASAP7_75t_L g1536 ( 
.A1(n_1316),
.A2(n_1185),
.B(n_1168),
.Y(n_1536)
);

OAI21x1_ASAP7_75t_L g1537 ( 
.A1(n_1338),
.A2(n_1185),
.B(n_1166),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1269),
.B(n_1190),
.Y(n_1538)
);

BUFx2_ASAP7_75t_SL g1539 ( 
.A(n_1271),
.Y(n_1539)
);

AO21x2_ASAP7_75t_L g1540 ( 
.A1(n_1331),
.A2(n_1185),
.B(n_1190),
.Y(n_1540)
);

O2A1O1Ixp33_ASAP7_75t_SL g1541 ( 
.A1(n_1301),
.A2(n_1114),
.B(n_1166),
.C(n_1207),
.Y(n_1541)
);

OAI21x1_ASAP7_75t_L g1542 ( 
.A1(n_1266),
.A2(n_1264),
.B(n_1351),
.Y(n_1542)
);

OAI21x1_ASAP7_75t_L g1543 ( 
.A1(n_1351),
.A2(n_1185),
.B(n_1166),
.Y(n_1543)
);

OAI21x1_ASAP7_75t_L g1544 ( 
.A1(n_1377),
.A2(n_1166),
.B(n_1046),
.Y(n_1544)
);

AOI21x1_ASAP7_75t_L g1545 ( 
.A1(n_1380),
.A2(n_1275),
.B(n_1408),
.Y(n_1545)
);

OAI21xp5_ASAP7_75t_L g1546 ( 
.A1(n_1406),
.A2(n_722),
.B(n_705),
.Y(n_1546)
);

INVx3_ASAP7_75t_L g1547 ( 
.A(n_1268),
.Y(n_1547)
);

AO21x2_ASAP7_75t_L g1548 ( 
.A1(n_1339),
.A2(n_1207),
.B(n_854),
.Y(n_1548)
);

OAI22xp33_ASAP7_75t_SL g1549 ( 
.A1(n_1342),
.A2(n_297),
.B1(n_293),
.B2(n_291),
.Y(n_1549)
);

INVx2_ASAP7_75t_SL g1550 ( 
.A(n_1271),
.Y(n_1550)
);

BUFx2_ASAP7_75t_L g1551 ( 
.A(n_1373),
.Y(n_1551)
);

OAI21x1_ASAP7_75t_L g1552 ( 
.A1(n_1353),
.A2(n_1207),
.B(n_854),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1310),
.Y(n_1553)
);

HB1xp67_ASAP7_75t_L g1554 ( 
.A(n_1363),
.Y(n_1554)
);

OAI21x1_ASAP7_75t_L g1555 ( 
.A1(n_1337),
.A2(n_1207),
.B(n_722),
.Y(n_1555)
);

OAI21x1_ASAP7_75t_L g1556 ( 
.A1(n_1340),
.A2(n_705),
.B(n_677),
.Y(n_1556)
);

NOR2xp33_ASAP7_75t_L g1557 ( 
.A(n_1393),
.B(n_1114),
.Y(n_1557)
);

AOI21x1_ASAP7_75t_L g1558 ( 
.A1(n_1275),
.A2(n_677),
.B(n_655),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1310),
.Y(n_1559)
);

OAI21x1_ASAP7_75t_L g1560 ( 
.A1(n_1343),
.A2(n_677),
.B(n_655),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1310),
.Y(n_1561)
);

AOI22xp33_ASAP7_75t_L g1562 ( 
.A1(n_1386),
.A2(n_429),
.B1(n_381),
.B2(n_466),
.Y(n_1562)
);

INVx3_ASAP7_75t_L g1563 ( 
.A(n_1268),
.Y(n_1563)
);

CKINVDCx5p33_ASAP7_75t_R g1564 ( 
.A(n_1322),
.Y(n_1564)
);

NOR2xp33_ASAP7_75t_SL g1565 ( 
.A(n_1322),
.B(n_269),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1269),
.B(n_381),
.Y(n_1566)
);

OAI22xp5_ASAP7_75t_SL g1567 ( 
.A1(n_1393),
.A2(n_381),
.B1(n_429),
.B2(n_466),
.Y(n_1567)
);

OAI21x1_ASAP7_75t_L g1568 ( 
.A1(n_1349),
.A2(n_687),
.B(n_685),
.Y(n_1568)
);

OAI21x1_ASAP7_75t_L g1569 ( 
.A1(n_1372),
.A2(n_1314),
.B(n_1280),
.Y(n_1569)
);

AOI22xp33_ASAP7_75t_L g1570 ( 
.A1(n_1368),
.A2(n_466),
.B1(n_429),
.B2(n_680),
.Y(n_1570)
);

AO31x2_ASAP7_75t_L g1571 ( 
.A1(n_1295),
.A2(n_687),
.A3(n_685),
.B(n_680),
.Y(n_1571)
);

INVx2_ASAP7_75t_L g1572 ( 
.A(n_1310),
.Y(n_1572)
);

HB1xp67_ASAP7_75t_L g1573 ( 
.A(n_1398),
.Y(n_1573)
);

OAI21x1_ASAP7_75t_L g1574 ( 
.A1(n_1280),
.A2(n_1320),
.B(n_1325),
.Y(n_1574)
);

AOI22xp33_ASAP7_75t_L g1575 ( 
.A1(n_1346),
.A2(n_466),
.B1(n_429),
.B2(n_680),
.Y(n_1575)
);

OAI21xp5_ASAP7_75t_L g1576 ( 
.A1(n_1362),
.A2(n_397),
.B(n_304),
.Y(n_1576)
);

AND2x4_ASAP7_75t_L g1577 ( 
.A(n_1382),
.B(n_655),
.Y(n_1577)
);

OAI21x1_ASAP7_75t_L g1578 ( 
.A1(n_1280),
.A2(n_687),
.B(n_685),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1299),
.Y(n_1579)
);

OA21x2_ASAP7_75t_L g1580 ( 
.A1(n_1362),
.A2(n_392),
.B(n_290),
.Y(n_1580)
);

OA21x2_ASAP7_75t_L g1581 ( 
.A1(n_1383),
.A2(n_1397),
.B(n_1390),
.Y(n_1581)
);

INVx3_ASAP7_75t_L g1582 ( 
.A(n_1268),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1299),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1299),
.Y(n_1584)
);

OAI22xp5_ASAP7_75t_L g1585 ( 
.A1(n_1317),
.A2(n_466),
.B1(n_305),
.B2(n_308),
.Y(n_1585)
);

HB1xp67_ASAP7_75t_L g1586 ( 
.A(n_1327),
.Y(n_1586)
);

OAI21x1_ASAP7_75t_L g1587 ( 
.A1(n_1325),
.A2(n_687),
.B(n_685),
.Y(n_1587)
);

OAI21x1_ASAP7_75t_L g1588 ( 
.A1(n_1325),
.A2(n_687),
.B(n_685),
.Y(n_1588)
);

OAI21x1_ASAP7_75t_L g1589 ( 
.A1(n_1296),
.A2(n_687),
.B(n_685),
.Y(n_1589)
);

A2O1A1Ixp33_ASAP7_75t_L g1590 ( 
.A1(n_1253),
.A2(n_1367),
.B(n_1400),
.C(n_1366),
.Y(n_1590)
);

BUFx3_ASAP7_75t_L g1591 ( 
.A(n_1327),
.Y(n_1591)
);

AO21x2_ASAP7_75t_L g1592 ( 
.A1(n_1262),
.A2(n_687),
.B(n_685),
.Y(n_1592)
);

NOR2xp33_ASAP7_75t_L g1593 ( 
.A(n_1258),
.B(n_1330),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1299),
.Y(n_1594)
);

OAI21x1_ASAP7_75t_L g1595 ( 
.A1(n_1275),
.A2(n_680),
.B(n_677),
.Y(n_1595)
);

OR2x2_ASAP7_75t_L g1596 ( 
.A(n_1278),
.B(n_655),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1590),
.Y(n_1597)
);

AND2x4_ASAP7_75t_L g1598 ( 
.A(n_1531),
.B(n_1538),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1528),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1528),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1533),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1485),
.B(n_1267),
.Y(n_1602)
);

BUFx2_ASAP7_75t_L g1603 ( 
.A(n_1591),
.Y(n_1603)
);

AOI22xp33_ASAP7_75t_L g1604 ( 
.A1(n_1562),
.A2(n_1336),
.B1(n_1332),
.B2(n_1405),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_1418),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1418),
.Y(n_1606)
);

CKINVDCx8_ASAP7_75t_R g1607 ( 
.A(n_1564),
.Y(n_1607)
);

NAND2x1p5_ASAP7_75t_L g1608 ( 
.A(n_1410),
.B(n_1271),
.Y(n_1608)
);

OAI22xp33_ASAP7_75t_L g1609 ( 
.A1(n_1497),
.A2(n_1355),
.B1(n_1326),
.B2(n_1279),
.Y(n_1609)
);

INVx3_ASAP7_75t_L g1610 ( 
.A(n_1495),
.Y(n_1610)
);

NAND3xp33_ASAP7_75t_SL g1611 ( 
.A(n_1414),
.B(n_1341),
.C(n_1281),
.Y(n_1611)
);

AOI22xp5_ASAP7_75t_L g1612 ( 
.A1(n_1464),
.A2(n_1379),
.B1(n_1258),
.B2(n_1298),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1533),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1428),
.Y(n_1614)
);

CKINVDCx20_ASAP7_75t_R g1615 ( 
.A(n_1484),
.Y(n_1615)
);

AOI22xp33_ASAP7_75t_L g1616 ( 
.A1(n_1436),
.A2(n_1388),
.B1(n_1306),
.B2(n_1385),
.Y(n_1616)
);

CKINVDCx5p33_ASAP7_75t_R g1617 ( 
.A(n_1419),
.Y(n_1617)
);

AOI221xp5_ASAP7_75t_L g1618 ( 
.A1(n_1415),
.A2(n_1382),
.B1(n_1278),
.B2(n_391),
.C(n_310),
.Y(n_1618)
);

OAI22xp5_ASAP7_75t_L g1619 ( 
.A1(n_1423),
.A2(n_1497),
.B1(n_1457),
.B2(n_1450),
.Y(n_1619)
);

AOI22xp5_ASAP7_75t_SL g1620 ( 
.A1(n_1461),
.A2(n_1388),
.B1(n_1373),
.B2(n_317),
.Y(n_1620)
);

OAI22xp5_ASAP7_75t_L g1621 ( 
.A1(n_1423),
.A2(n_1369),
.B1(n_1251),
.B2(n_1309),
.Y(n_1621)
);

AO221x2_ASAP7_75t_L g1622 ( 
.A1(n_1567),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.C(n_16),
.Y(n_1622)
);

AOI22xp5_ASAP7_75t_L g1623 ( 
.A1(n_1514),
.A2(n_1369),
.B1(n_1251),
.B2(n_1388),
.Y(n_1623)
);

OAI211xp5_ASAP7_75t_L g1624 ( 
.A1(n_1463),
.A2(n_424),
.B(n_327),
.C(n_346),
.Y(n_1624)
);

AOI22xp33_ASAP7_75t_L g1625 ( 
.A1(n_1567),
.A2(n_1485),
.B1(n_1501),
.B2(n_1476),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1435),
.B(n_1369),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1428),
.Y(n_1627)
);

INVx2_ASAP7_75t_SL g1628 ( 
.A(n_1591),
.Y(n_1628)
);

AOI21xp33_ASAP7_75t_L g1629 ( 
.A1(n_1549),
.A2(n_1278),
.B(n_1394),
.Y(n_1629)
);

AOI221xp5_ASAP7_75t_L g1630 ( 
.A1(n_1549),
.A2(n_1278),
.B1(n_354),
.B2(n_363),
.C(n_370),
.Y(n_1630)
);

NAND3xp33_ASAP7_75t_SL g1631 ( 
.A(n_1565),
.B(n_425),
.C(n_460),
.Y(n_1631)
);

HB1xp67_ASAP7_75t_L g1632 ( 
.A(n_1486),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1474),
.B(n_14),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1446),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1500),
.B(n_15),
.Y(n_1635)
);

NOR2xp33_ASAP7_75t_L g1636 ( 
.A(n_1498),
.B(n_1283),
.Y(n_1636)
);

NAND3xp33_ASAP7_75t_SL g1637 ( 
.A(n_1565),
.B(n_405),
.C(n_453),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1493),
.B(n_1519),
.Y(n_1638)
);

OAI22xp5_ASAP7_75t_L g1639 ( 
.A1(n_1431),
.A2(n_1309),
.B1(n_1271),
.B2(n_1357),
.Y(n_1639)
);

OA21x2_ASAP7_75t_L g1640 ( 
.A1(n_1574),
.A2(n_1302),
.B(n_1334),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1456),
.B(n_16),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1446),
.Y(n_1642)
);

BUFx3_ASAP7_75t_L g1643 ( 
.A(n_1591),
.Y(n_1643)
);

INVx4_ASAP7_75t_L g1644 ( 
.A(n_1412),
.Y(n_1644)
);

OAI21x1_ASAP7_75t_L g1645 ( 
.A1(n_1574),
.A2(n_1381),
.B(n_1302),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1512),
.B(n_17),
.Y(n_1646)
);

INVx2_ASAP7_75t_SL g1647 ( 
.A(n_1586),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1477),
.B(n_1573),
.Y(n_1648)
);

CKINVDCx5p33_ASAP7_75t_R g1649 ( 
.A(n_1419),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1490),
.Y(n_1650)
);

OAI21x1_ASAP7_75t_L g1651 ( 
.A1(n_1513),
.A2(n_1381),
.B(n_1302),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1490),
.Y(n_1652)
);

AND2x2_ASAP7_75t_SL g1653 ( 
.A(n_1486),
.B(n_1283),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1566),
.B(n_1531),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1504),
.Y(n_1655)
);

INVx5_ASAP7_75t_L g1656 ( 
.A(n_1420),
.Y(n_1656)
);

AOI22xp33_ASAP7_75t_L g1657 ( 
.A1(n_1576),
.A2(n_677),
.B1(n_680),
.B2(n_1394),
.Y(n_1657)
);

BUFx6f_ASAP7_75t_L g1658 ( 
.A(n_1437),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_SL g1659 ( 
.A(n_1427),
.B(n_1283),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1566),
.B(n_17),
.Y(n_1660)
);

OAI22xp5_ASAP7_75t_L g1661 ( 
.A1(n_1424),
.A2(n_1309),
.B1(n_1357),
.B2(n_1312),
.Y(n_1661)
);

OAI22xp5_ASAP7_75t_L g1662 ( 
.A1(n_1489),
.A2(n_1309),
.B1(n_1357),
.B2(n_1312),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1538),
.B(n_1434),
.Y(n_1663)
);

OA21x2_ASAP7_75t_L g1664 ( 
.A1(n_1578),
.A2(n_1302),
.B(n_1334),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1434),
.B(n_1348),
.Y(n_1665)
);

INVx3_ASAP7_75t_SL g1666 ( 
.A(n_1412),
.Y(n_1666)
);

AOI21xp33_ASAP7_75t_L g1667 ( 
.A1(n_1576),
.A2(n_1394),
.B(n_1287),
.Y(n_1667)
);

HB1xp67_ASAP7_75t_L g1668 ( 
.A(n_1530),
.Y(n_1668)
);

BUFx10_ASAP7_75t_L g1669 ( 
.A(n_1564),
.Y(n_1669)
);

AO31x2_ASAP7_75t_L g1670 ( 
.A1(n_1583),
.A2(n_1334),
.A3(n_1348),
.B(n_1374),
.Y(n_1670)
);

OR2x4_ASAP7_75t_L g1671 ( 
.A(n_1557),
.B(n_1283),
.Y(n_1671)
);

NAND3xp33_ASAP7_75t_L g1672 ( 
.A(n_1580),
.B(n_1413),
.C(n_1535),
.Y(n_1672)
);

HB1xp67_ASAP7_75t_L g1673 ( 
.A(n_1530),
.Y(n_1673)
);

OAI22xp5_ASAP7_75t_L g1674 ( 
.A1(n_1489),
.A2(n_1357),
.B1(n_1312),
.B2(n_1287),
.Y(n_1674)
);

OAI22xp5_ASAP7_75t_L g1675 ( 
.A1(n_1526),
.A2(n_1394),
.B1(n_1312),
.B2(n_1287),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1554),
.B(n_1348),
.Y(n_1676)
);

AOI22xp33_ASAP7_75t_L g1677 ( 
.A1(n_1580),
.A2(n_680),
.B1(n_1287),
.B2(n_364),
.Y(n_1677)
);

INVx2_ASAP7_75t_L g1678 ( 
.A(n_1426),
.Y(n_1678)
);

BUFx2_ASAP7_75t_L g1679 ( 
.A(n_1480),
.Y(n_1679)
);

CKINVDCx11_ASAP7_75t_R g1680 ( 
.A(n_1440),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1504),
.Y(n_1681)
);

CKINVDCx5p33_ASAP7_75t_R g1682 ( 
.A(n_1593),
.Y(n_1682)
);

INVx4_ASAP7_75t_L g1683 ( 
.A(n_1437),
.Y(n_1683)
);

BUFx2_ASAP7_75t_SL g1684 ( 
.A(n_1480),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1505),
.Y(n_1685)
);

OR2x2_ASAP7_75t_L g1686 ( 
.A(n_1534),
.B(n_1348),
.Y(n_1686)
);

INVx2_ASAP7_75t_SL g1687 ( 
.A(n_1521),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1437),
.B(n_22),
.Y(n_1688)
);

INVx6_ASAP7_75t_L g1689 ( 
.A(n_1437),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1481),
.B(n_1270),
.Y(n_1690)
);

NOR2xp33_ASAP7_75t_R g1691 ( 
.A(n_1480),
.B(n_115),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1505),
.Y(n_1692)
);

AOI22xp33_ASAP7_75t_SL g1693 ( 
.A1(n_1580),
.A2(n_1270),
.B1(n_364),
.B2(n_269),
.Y(n_1693)
);

AOI221xp5_ASAP7_75t_L g1694 ( 
.A1(n_1416),
.A2(n_371),
.B1(n_436),
.B2(n_434),
.C(n_431),
.Y(n_1694)
);

AOI22xp33_ASAP7_75t_SL g1695 ( 
.A1(n_1580),
.A2(n_1270),
.B1(n_269),
.B2(n_401),
.Y(n_1695)
);

OAI22xp33_ASAP7_75t_L g1696 ( 
.A1(n_1420),
.A2(n_1270),
.B1(n_269),
.B2(n_401),
.Y(n_1696)
);

AND2x4_ASAP7_75t_L g1697 ( 
.A(n_1420),
.B(n_1374),
.Y(n_1697)
);

BUFx6f_ASAP7_75t_L g1698 ( 
.A(n_1448),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1481),
.B(n_1508),
.Y(n_1699)
);

INVx2_ASAP7_75t_L g1700 ( 
.A(n_1426),
.Y(n_1700)
);

AOI22xp33_ASAP7_75t_L g1701 ( 
.A1(n_1487),
.A2(n_269),
.B1(n_364),
.B2(n_401),
.Y(n_1701)
);

OAI221xp5_ASAP7_75t_L g1702 ( 
.A1(n_1451),
.A2(n_403),
.B1(n_402),
.B2(n_373),
.C(n_372),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1506),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1481),
.B(n_24),
.Y(n_1704)
);

OAI22xp5_ASAP7_75t_L g1705 ( 
.A1(n_1420),
.A2(n_401),
.B1(n_364),
.B2(n_269),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1506),
.Y(n_1706)
);

NAND2xp33_ASAP7_75t_R g1707 ( 
.A(n_1420),
.B(n_1374),
.Y(n_1707)
);

AOI22xp33_ASAP7_75t_L g1708 ( 
.A1(n_1487),
.A2(n_401),
.B1(n_364),
.B2(n_1334),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_SL g1709 ( 
.A(n_1447),
.B(n_1483),
.Y(n_1709)
);

AND2x4_ASAP7_75t_L g1710 ( 
.A(n_1448),
.B(n_1374),
.Y(n_1710)
);

A2O1A1Ixp33_ASAP7_75t_L g1711 ( 
.A1(n_1546),
.A2(n_364),
.B(n_401),
.C(n_30),
.Y(n_1711)
);

AOI22xp33_ASAP7_75t_SL g1712 ( 
.A1(n_1487),
.A2(n_24),
.B1(n_26),
.B2(n_30),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1522),
.Y(n_1713)
);

NAND2xp33_ASAP7_75t_L g1714 ( 
.A(n_1430),
.B(n_31),
.Y(n_1714)
);

HB1xp67_ASAP7_75t_L g1715 ( 
.A(n_1551),
.Y(n_1715)
);

OAI22xp5_ASAP7_75t_L g1716 ( 
.A1(n_1454),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_1716)
);

AOI22xp33_ASAP7_75t_L g1717 ( 
.A1(n_1416),
.A2(n_33),
.B1(n_37),
.B2(n_38),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1525),
.Y(n_1718)
);

INVx3_ASAP7_75t_L g1719 ( 
.A(n_1495),
.Y(n_1719)
);

OAI21x1_ASAP7_75t_L g1720 ( 
.A1(n_1513),
.A2(n_241),
.B(n_236),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1525),
.Y(n_1721)
);

AND2x6_ASAP7_75t_L g1722 ( 
.A(n_1410),
.B(n_122),
.Y(n_1722)
);

AND2x4_ASAP7_75t_L g1723 ( 
.A(n_1448),
.B(n_125),
.Y(n_1723)
);

OAI22xp5_ASAP7_75t_L g1724 ( 
.A1(n_1523),
.A2(n_38),
.B1(n_39),
.B2(n_41),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1481),
.B(n_41),
.Y(n_1725)
);

HB1xp67_ASAP7_75t_L g1726 ( 
.A(n_1551),
.Y(n_1726)
);

O2A1O1Ixp33_ASAP7_75t_SL g1727 ( 
.A1(n_1441),
.A2(n_46),
.B(n_49),
.C(n_50),
.Y(n_1727)
);

AOI22xp33_ASAP7_75t_L g1728 ( 
.A1(n_1410),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1411),
.Y(n_1729)
);

INVx4_ASAP7_75t_L g1730 ( 
.A(n_1430),
.Y(n_1730)
);

CKINVDCx5p33_ASAP7_75t_R g1731 ( 
.A(n_1508),
.Y(n_1731)
);

HB1xp67_ASAP7_75t_L g1732 ( 
.A(n_1479),
.Y(n_1732)
);

OR2x2_ASAP7_75t_L g1733 ( 
.A(n_1449),
.B(n_52),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1411),
.Y(n_1734)
);

INVx2_ASAP7_75t_L g1735 ( 
.A(n_1417),
.Y(n_1735)
);

BUFx2_ASAP7_75t_L g1736 ( 
.A(n_1508),
.Y(n_1736)
);

NAND2xp33_ASAP7_75t_L g1737 ( 
.A(n_1430),
.B(n_53),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1410),
.B(n_55),
.Y(n_1738)
);

OR2x6_ASAP7_75t_L g1739 ( 
.A(n_1442),
.B(n_230),
.Y(n_1739)
);

AOI22xp33_ASAP7_75t_L g1740 ( 
.A1(n_1458),
.A2(n_57),
.B1(n_59),
.B2(n_60),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1417),
.Y(n_1741)
);

BUFx2_ASAP7_75t_L g1742 ( 
.A(n_1448),
.Y(n_1742)
);

OR2x6_ASAP7_75t_L g1743 ( 
.A(n_1442),
.B(n_228),
.Y(n_1743)
);

INVx2_ASAP7_75t_L g1744 ( 
.A(n_1553),
.Y(n_1744)
);

AOI22xp33_ASAP7_75t_SL g1745 ( 
.A1(n_1502),
.A2(n_59),
.B1(n_60),
.B2(n_61),
.Y(n_1745)
);

OAI22xp33_ASAP7_75t_L g1746 ( 
.A1(n_1472),
.A2(n_62),
.B1(n_63),
.B2(n_65),
.Y(n_1746)
);

OR2x6_ASAP7_75t_L g1747 ( 
.A(n_1442),
.B(n_223),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1455),
.Y(n_1748)
);

BUFx6f_ASAP7_75t_L g1749 ( 
.A(n_1462),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1455),
.Y(n_1750)
);

INVx3_ASAP7_75t_L g1751 ( 
.A(n_1495),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1459),
.Y(n_1752)
);

NAND2x1_ASAP7_75t_L g1753 ( 
.A(n_1495),
.B(n_209),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1462),
.B(n_66),
.Y(n_1754)
);

AOI22xp33_ASAP7_75t_L g1755 ( 
.A1(n_1458),
.A2(n_1546),
.B1(n_1575),
.B2(n_1503),
.Y(n_1755)
);

AOI22xp33_ASAP7_75t_L g1756 ( 
.A1(n_1458),
.A2(n_67),
.B1(n_68),
.B2(n_69),
.Y(n_1756)
);

A2O1A1Ixp33_ASAP7_75t_L g1757 ( 
.A1(n_1444),
.A2(n_1441),
.B(n_1507),
.C(n_1478),
.Y(n_1757)
);

AOI21xp33_ASAP7_75t_L g1758 ( 
.A1(n_1452),
.A2(n_1596),
.B(n_1585),
.Y(n_1758)
);

INVx3_ASAP7_75t_L g1759 ( 
.A(n_1462),
.Y(n_1759)
);

AOI22xp33_ASAP7_75t_L g1760 ( 
.A1(n_1503),
.A2(n_1467),
.B1(n_1469),
.B2(n_1473),
.Y(n_1760)
);

BUFx3_ASAP7_75t_L g1761 ( 
.A(n_1430),
.Y(n_1761)
);

CKINVDCx16_ASAP7_75t_R g1762 ( 
.A(n_1539),
.Y(n_1762)
);

OAI21xp33_ASAP7_75t_L g1763 ( 
.A1(n_1444),
.A2(n_70),
.B(n_71),
.Y(n_1763)
);

OR2x6_ASAP7_75t_L g1764 ( 
.A(n_1442),
.B(n_205),
.Y(n_1764)
);

OAI21xp5_ASAP7_75t_L g1765 ( 
.A1(n_1438),
.A2(n_70),
.B(n_71),
.Y(n_1765)
);

INVx3_ASAP7_75t_L g1766 ( 
.A(n_1462),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1459),
.Y(n_1767)
);

AOI21xp5_ASAP7_75t_L g1768 ( 
.A1(n_1429),
.A2(n_72),
.B(n_74),
.Y(n_1768)
);

INVx4_ASAP7_75t_SL g1769 ( 
.A(n_1449),
.Y(n_1769)
);

AOI22xp33_ASAP7_75t_L g1770 ( 
.A1(n_1467),
.A2(n_74),
.B1(n_75),
.B2(n_76),
.Y(n_1770)
);

OAI22xp5_ASAP7_75t_L g1771 ( 
.A1(n_1449),
.A2(n_75),
.B1(n_76),
.B2(n_77),
.Y(n_1771)
);

AOI21xp33_ASAP7_75t_L g1772 ( 
.A1(n_1452),
.A2(n_77),
.B(n_81),
.Y(n_1772)
);

CKINVDCx5p33_ASAP7_75t_R g1773 ( 
.A(n_1539),
.Y(n_1773)
);

CKINVDCx20_ASAP7_75t_R g1774 ( 
.A(n_1518),
.Y(n_1774)
);

OAI22xp5_ASAP7_75t_L g1775 ( 
.A1(n_1449),
.A2(n_82),
.B1(n_84),
.B2(n_85),
.Y(n_1775)
);

BUFx6f_ASAP7_75t_L g1776 ( 
.A(n_1430),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1577),
.B(n_84),
.Y(n_1777)
);

BUFx2_ASAP7_75t_L g1778 ( 
.A(n_1517),
.Y(n_1778)
);

CKINVDCx20_ASAP7_75t_R g1779 ( 
.A(n_1518),
.Y(n_1779)
);

OAI221xp5_ASAP7_75t_L g1780 ( 
.A1(n_1570),
.A2(n_86),
.B1(n_87),
.B2(n_88),
.C(n_89),
.Y(n_1780)
);

AOI22xp33_ASAP7_75t_L g1781 ( 
.A1(n_1469),
.A2(n_86),
.B1(n_90),
.B2(n_93),
.Y(n_1781)
);

INVx4_ASAP7_75t_L g1782 ( 
.A(n_1517),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1473),
.Y(n_1783)
);

OR2x2_ASAP7_75t_L g1784 ( 
.A(n_1449),
.B(n_95),
.Y(n_1784)
);

A2O1A1Ixp33_ASAP7_75t_L g1785 ( 
.A1(n_1470),
.A2(n_103),
.B(n_104),
.C(n_106),
.Y(n_1785)
);

CKINVDCx12_ASAP7_75t_R g1786 ( 
.A(n_1453),
.Y(n_1786)
);

AND2x2_ASAP7_75t_L g1787 ( 
.A(n_1577),
.B(n_104),
.Y(n_1787)
);

CKINVDCx5p33_ASAP7_75t_R g1788 ( 
.A(n_1517),
.Y(n_1788)
);

BUFx2_ASAP7_75t_SL g1789 ( 
.A(n_1550),
.Y(n_1789)
);

BUFx4f_ASAP7_75t_SL g1790 ( 
.A(n_1517),
.Y(n_1790)
);

AND2x2_ASAP7_75t_L g1791 ( 
.A(n_1577),
.B(n_106),
.Y(n_1791)
);

AND2x4_ASAP7_75t_L g1792 ( 
.A(n_1453),
.B(n_164),
.Y(n_1792)
);

AOI22xp33_ASAP7_75t_L g1793 ( 
.A1(n_1491),
.A2(n_108),
.B1(n_109),
.B2(n_110),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1577),
.B(n_108),
.Y(n_1794)
);

INVx4_ASAP7_75t_L g1795 ( 
.A(n_1517),
.Y(n_1795)
);

AOI22xp33_ASAP7_75t_L g1796 ( 
.A1(n_1491),
.A2(n_112),
.B1(n_113),
.B2(n_126),
.Y(n_1796)
);

OR2x2_ASAP7_75t_L g1797 ( 
.A(n_1453),
.B(n_135),
.Y(n_1797)
);

INVx2_ASAP7_75t_L g1798 ( 
.A(n_1553),
.Y(n_1798)
);

CKINVDCx20_ASAP7_75t_R g1799 ( 
.A(n_1550),
.Y(n_1799)
);

AND2x4_ASAP7_75t_L g1800 ( 
.A(n_1516),
.B(n_138),
.Y(n_1800)
);

AOI22xp33_ASAP7_75t_L g1801 ( 
.A1(n_1494),
.A2(n_200),
.B1(n_141),
.B2(n_142),
.Y(n_1801)
);

INVx3_ASAP7_75t_L g1802 ( 
.A(n_1465),
.Y(n_1802)
);

CKINVDCx11_ASAP7_75t_R g1803 ( 
.A(n_1532),
.Y(n_1803)
);

NOR2xp33_ASAP7_75t_L g1804 ( 
.A(n_1453),
.B(n_140),
.Y(n_1804)
);

AOI221xp5_ASAP7_75t_L g1805 ( 
.A1(n_1609),
.A2(n_1561),
.B1(n_1584),
.B2(n_1579),
.C(n_1511),
.Y(n_1805)
);

AOI221xp5_ASAP7_75t_L g1806 ( 
.A1(n_1609),
.A2(n_1561),
.B1(n_1584),
.B2(n_1579),
.C(n_1511),
.Y(n_1806)
);

AOI22xp33_ASAP7_75t_L g1807 ( 
.A1(n_1622),
.A2(n_1494),
.B1(n_1572),
.B2(n_1559),
.Y(n_1807)
);

AOI22xp33_ASAP7_75t_L g1808 ( 
.A1(n_1622),
.A2(n_1572),
.B1(n_1559),
.B2(n_1594),
.Y(n_1808)
);

AOI22xp33_ASAP7_75t_L g1809 ( 
.A1(n_1622),
.A2(n_1583),
.B1(n_1594),
.B2(n_1596),
.Y(n_1809)
);

AOI22xp33_ASAP7_75t_L g1810 ( 
.A1(n_1611),
.A2(n_1516),
.B1(n_1453),
.B2(n_1452),
.Y(n_1810)
);

OR2x2_ASAP7_75t_L g1811 ( 
.A(n_1663),
.B(n_1516),
.Y(n_1811)
);

OAI22xp5_ASAP7_75t_L g1812 ( 
.A1(n_1612),
.A2(n_1492),
.B1(n_1524),
.B2(n_1582),
.Y(n_1812)
);

OAI211xp5_ASAP7_75t_SL g1813 ( 
.A1(n_1717),
.A2(n_1541),
.B(n_1547),
.C(n_1492),
.Y(n_1813)
);

AOI22xp33_ASAP7_75t_L g1814 ( 
.A1(n_1618),
.A2(n_1422),
.B1(n_1442),
.B2(n_1581),
.Y(n_1814)
);

NOR2xp33_ASAP7_75t_L g1815 ( 
.A(n_1619),
.B(n_1492),
.Y(n_1815)
);

AOI22xp33_ASAP7_75t_L g1816 ( 
.A1(n_1763),
.A2(n_1422),
.B1(n_1581),
.B2(n_1540),
.Y(n_1816)
);

OAI22xp5_ASAP7_75t_L g1817 ( 
.A1(n_1728),
.A2(n_1717),
.B1(n_1745),
.B2(n_1604),
.Y(n_1817)
);

OAI22xp33_ASAP7_75t_L g1818 ( 
.A1(n_1746),
.A2(n_1515),
.B1(n_1433),
.B2(n_1465),
.Y(n_1818)
);

OAI22xp5_ASAP7_75t_L g1819 ( 
.A1(n_1728),
.A2(n_1604),
.B1(n_1781),
.B2(n_1770),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1602),
.B(n_1492),
.Y(n_1820)
);

AOI22xp33_ASAP7_75t_L g1821 ( 
.A1(n_1696),
.A2(n_1422),
.B1(n_1581),
.B2(n_1540),
.Y(n_1821)
);

AOI22xp33_ASAP7_75t_L g1822 ( 
.A1(n_1696),
.A2(n_1625),
.B1(n_1630),
.B2(n_1746),
.Y(n_1822)
);

INVx4_ASAP7_75t_L g1823 ( 
.A(n_1773),
.Y(n_1823)
);

OR2x6_ASAP7_75t_L g1824 ( 
.A(n_1739),
.B(n_1743),
.Y(n_1824)
);

AOI211xp5_ASAP7_75t_SL g1825 ( 
.A1(n_1727),
.A2(n_1524),
.B(n_1563),
.C(n_1547),
.Y(n_1825)
);

OAI22xp5_ASAP7_75t_L g1826 ( 
.A1(n_1770),
.A2(n_1793),
.B1(n_1781),
.B2(n_1711),
.Y(n_1826)
);

INVx1_ASAP7_75t_SL g1827 ( 
.A(n_1682),
.Y(n_1827)
);

AOI22xp33_ASAP7_75t_L g1828 ( 
.A1(n_1625),
.A2(n_1422),
.B1(n_1581),
.B2(n_1540),
.Y(n_1828)
);

AOI222xp33_ASAP7_75t_L g1829 ( 
.A1(n_1793),
.A2(n_1421),
.B1(n_1488),
.B2(n_1524),
.C1(n_1582),
.C2(n_1547),
.Y(n_1829)
);

OAI22xp5_ASAP7_75t_L g1830 ( 
.A1(n_1711),
.A2(n_1582),
.B1(n_1524),
.B2(n_1547),
.Y(n_1830)
);

OAI221xp5_ASAP7_75t_SL g1831 ( 
.A1(n_1740),
.A2(n_1468),
.B1(n_1563),
.B2(n_1582),
.C(n_1515),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1638),
.B(n_1563),
.Y(n_1832)
);

AOI21xp5_ASAP7_75t_L g1833 ( 
.A1(n_1714),
.A2(n_1488),
.B(n_1482),
.Y(n_1833)
);

OAI22xp5_ASAP7_75t_L g1834 ( 
.A1(n_1796),
.A2(n_1563),
.B1(n_1433),
.B2(n_1532),
.Y(n_1834)
);

AOI22xp33_ASAP7_75t_L g1835 ( 
.A1(n_1740),
.A2(n_1548),
.B1(n_1592),
.B2(n_1475),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1599),
.Y(n_1836)
);

BUFx6f_ASAP7_75t_L g1837 ( 
.A(n_1803),
.Y(n_1837)
);

OAI22xp5_ASAP7_75t_L g1838 ( 
.A1(n_1796),
.A2(n_1433),
.B1(n_1532),
.B2(n_1465),
.Y(n_1838)
);

OAI221xp5_ASAP7_75t_L g1839 ( 
.A1(n_1756),
.A2(n_1545),
.B1(n_1471),
.B2(n_1479),
.C(n_1475),
.Y(n_1839)
);

OAI22xp5_ASAP7_75t_L g1840 ( 
.A1(n_1756),
.A2(n_1532),
.B1(n_1471),
.B2(n_1479),
.Y(n_1840)
);

AOI22xp33_ASAP7_75t_L g1841 ( 
.A1(n_1597),
.A2(n_1548),
.B1(n_1592),
.B2(n_1475),
.Y(n_1841)
);

AOI22xp33_ASAP7_75t_SL g1842 ( 
.A1(n_1620),
.A2(n_1691),
.B1(n_1765),
.B2(n_1737),
.Y(n_1842)
);

AND2x2_ASAP7_75t_L g1843 ( 
.A(n_1648),
.B(n_1532),
.Y(n_1843)
);

OAI22xp5_ASAP7_75t_L g1844 ( 
.A1(n_1716),
.A2(n_1479),
.B1(n_1545),
.B2(n_1475),
.Y(n_1844)
);

AOI21xp5_ASAP7_75t_L g1845 ( 
.A1(n_1659),
.A2(n_1757),
.B(n_1727),
.Y(n_1845)
);

OAI22xp33_ASAP7_75t_L g1846 ( 
.A1(n_1780),
.A2(n_1558),
.B1(n_1520),
.B2(n_1592),
.Y(n_1846)
);

OAI22xp33_ASAP7_75t_L g1847 ( 
.A1(n_1724),
.A2(n_1558),
.B1(n_1520),
.B2(n_1571),
.Y(n_1847)
);

AOI22xp33_ASAP7_75t_L g1848 ( 
.A1(n_1712),
.A2(n_1548),
.B1(n_1421),
.B2(n_1466),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1600),
.Y(n_1849)
);

BUFx4f_ASAP7_75t_L g1850 ( 
.A(n_1722),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1601),
.Y(n_1851)
);

AOI22xp33_ASAP7_75t_L g1852 ( 
.A1(n_1633),
.A2(n_1466),
.B1(n_1595),
.B2(n_1432),
.Y(n_1852)
);

AND2x2_ASAP7_75t_L g1853 ( 
.A(n_1598),
.B(n_1571),
.Y(n_1853)
);

OAI22xp5_ASAP7_75t_L g1854 ( 
.A1(n_1785),
.A2(n_1571),
.B1(n_1543),
.B2(n_1537),
.Y(n_1854)
);

AOI22xp33_ASAP7_75t_L g1855 ( 
.A1(n_1701),
.A2(n_1595),
.B1(n_1425),
.B2(n_1432),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1613),
.Y(n_1856)
);

OAI22xp5_ASAP7_75t_L g1857 ( 
.A1(n_1785),
.A2(n_1571),
.B1(n_1543),
.B2(n_1537),
.Y(n_1857)
);

AOI321xp33_ASAP7_75t_L g1858 ( 
.A1(n_1771),
.A2(n_1571),
.A3(n_1552),
.B1(n_1542),
.B2(n_1425),
.C(n_1569),
.Y(n_1858)
);

AOI22xp5_ASAP7_75t_L g1859 ( 
.A1(n_1775),
.A2(n_1544),
.B1(n_1460),
.B2(n_1527),
.Y(n_1859)
);

OR2x2_ASAP7_75t_L g1860 ( 
.A(n_1690),
.B(n_1527),
.Y(n_1860)
);

OAI22xp5_ASAP7_75t_L g1861 ( 
.A1(n_1733),
.A2(n_1460),
.B1(n_1536),
.B2(n_1552),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1614),
.Y(n_1862)
);

OAI221xp5_ASAP7_75t_L g1863 ( 
.A1(n_1616),
.A2(n_1542),
.B1(n_1569),
.B2(n_1445),
.C(n_1555),
.Y(n_1863)
);

AOI22xp33_ASAP7_75t_L g1864 ( 
.A1(n_1701),
.A2(n_1693),
.B1(n_1695),
.B2(n_1641),
.Y(n_1864)
);

OAI22xp5_ASAP7_75t_L g1865 ( 
.A1(n_1784),
.A2(n_1801),
.B1(n_1738),
.B2(n_1616),
.Y(n_1865)
);

AOI22xp33_ASAP7_75t_L g1866 ( 
.A1(n_1739),
.A2(n_1588),
.B1(n_1587),
.B2(n_1578),
.Y(n_1866)
);

OAI22xp5_ASAP7_75t_L g1867 ( 
.A1(n_1801),
.A2(n_1536),
.B1(n_1510),
.B2(n_1555),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1627),
.Y(n_1868)
);

OAI21x1_ASAP7_75t_L g1869 ( 
.A1(n_1651),
.A2(n_1589),
.B(n_1560),
.Y(n_1869)
);

AND2x2_ASAP7_75t_L g1870 ( 
.A(n_1598),
.B(n_1509),
.Y(n_1870)
);

AND2x2_ASAP7_75t_L g1871 ( 
.A(n_1598),
.B(n_1509),
.Y(n_1871)
);

AOI221xp5_ASAP7_75t_L g1872 ( 
.A1(n_1772),
.A2(n_153),
.B1(n_167),
.B2(n_173),
.C(n_174),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1634),
.Y(n_1873)
);

AOI22xp33_ASAP7_75t_L g1874 ( 
.A1(n_1739),
.A2(n_1588),
.B1(n_1587),
.B2(n_1544),
.Y(n_1874)
);

AOI22xp5_ASAP7_75t_L g1875 ( 
.A1(n_1621),
.A2(n_1445),
.B1(n_1478),
.B2(n_1470),
.Y(n_1875)
);

INVx2_ASAP7_75t_L g1876 ( 
.A(n_1735),
.Y(n_1876)
);

OAI22xp33_ASAP7_75t_L g1877 ( 
.A1(n_1743),
.A2(n_1482),
.B1(n_1499),
.B2(n_1496),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1654),
.B(n_1742),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1642),
.Y(n_1879)
);

OAI221xp5_ASAP7_75t_L g1880 ( 
.A1(n_1672),
.A2(n_1443),
.B1(n_1439),
.B2(n_1529),
.C(n_189),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1650),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1687),
.B(n_1443),
.Y(n_1882)
);

AOI22xp33_ASAP7_75t_L g1883 ( 
.A1(n_1743),
.A2(n_1439),
.B1(n_1529),
.B2(n_1499),
.Y(n_1883)
);

OAI22xp5_ASAP7_75t_L g1884 ( 
.A1(n_1657),
.A2(n_1510),
.B1(n_1496),
.B2(n_1556),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1647),
.B(n_1568),
.Y(n_1885)
);

AOI21xp5_ASAP7_75t_L g1886 ( 
.A1(n_1659),
.A2(n_1556),
.B(n_1589),
.Y(n_1886)
);

OAI22xp33_ASAP7_75t_L g1887 ( 
.A1(n_1747),
.A2(n_1568),
.B1(n_1560),
.B2(n_185),
.Y(n_1887)
);

AND2x2_ASAP7_75t_L g1888 ( 
.A(n_1704),
.B(n_180),
.Y(n_1888)
);

AOI221xp5_ASAP7_75t_SL g1889 ( 
.A1(n_1768),
.A2(n_182),
.B1(n_192),
.B2(n_195),
.C(n_196),
.Y(n_1889)
);

OAI211xp5_ASAP7_75t_SL g1890 ( 
.A1(n_1607),
.A2(n_1680),
.B(n_1694),
.C(n_1725),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1626),
.B(n_1731),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_L g1892 ( 
.A(n_1646),
.B(n_1635),
.Y(n_1892)
);

AO21x2_ASAP7_75t_L g1893 ( 
.A1(n_1629),
.A2(n_1758),
.B(n_1665),
.Y(n_1893)
);

AOI222xp33_ASAP7_75t_L g1894 ( 
.A1(n_1660),
.A2(n_1709),
.B1(n_1637),
.B2(n_1631),
.C1(n_1722),
.C2(n_1804),
.Y(n_1894)
);

OAI221xp5_ASAP7_75t_L g1895 ( 
.A1(n_1624),
.A2(n_1702),
.B1(n_1677),
.B2(n_1623),
.C(n_1667),
.Y(n_1895)
);

OAI211xp5_ASAP7_75t_SL g1896 ( 
.A1(n_1680),
.A2(n_1709),
.B(n_1757),
.C(n_1803),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1699),
.B(n_1754),
.Y(n_1897)
);

AOI22xp33_ASAP7_75t_L g1898 ( 
.A1(n_1747),
.A2(n_1764),
.B1(n_1755),
.B2(n_1722),
.Y(n_1898)
);

INVx2_ASAP7_75t_L g1899 ( 
.A(n_1735),
.Y(n_1899)
);

AO31x2_ASAP7_75t_L g1900 ( 
.A1(n_1744),
.A2(n_1798),
.A3(n_1605),
.B(n_1606),
.Y(n_1900)
);

OAI22xp5_ASAP7_75t_L g1901 ( 
.A1(n_1657),
.A2(n_1762),
.B1(n_1799),
.B2(n_1774),
.Y(n_1901)
);

AOI222xp33_ASAP7_75t_L g1902 ( 
.A1(n_1722),
.A2(n_1804),
.B1(n_1705),
.B2(n_1755),
.C1(n_1792),
.C2(n_1677),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1652),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1655),
.Y(n_1904)
);

AOI21xp5_ASAP7_75t_SL g1905 ( 
.A1(n_1723),
.A2(n_1764),
.B(n_1747),
.Y(n_1905)
);

AOI22xp33_ASAP7_75t_SL g1906 ( 
.A1(n_1691),
.A2(n_1722),
.B1(n_1764),
.B2(n_1656),
.Y(n_1906)
);

AND2x2_ASAP7_75t_L g1907 ( 
.A(n_1759),
.B(n_1766),
.Y(n_1907)
);

AOI221xp5_ASAP7_75t_L g1908 ( 
.A1(n_1676),
.A2(n_1760),
.B1(n_1767),
.B2(n_1752),
.C(n_1783),
.Y(n_1908)
);

AOI22xp33_ASAP7_75t_L g1909 ( 
.A1(n_1792),
.A2(n_1800),
.B1(n_1686),
.B2(n_1787),
.Y(n_1909)
);

OAI211xp5_ASAP7_75t_SL g1910 ( 
.A1(n_1632),
.A2(n_1668),
.B(n_1726),
.C(n_1715),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1681),
.Y(n_1911)
);

AOI221xp5_ASAP7_75t_L g1912 ( 
.A1(n_1760),
.A2(n_1750),
.B1(n_1748),
.B2(n_1741),
.C(n_1734),
.Y(n_1912)
);

BUFx2_ASAP7_75t_L g1913 ( 
.A(n_1643),
.Y(n_1913)
);

OAI22xp33_ASAP7_75t_L g1914 ( 
.A1(n_1671),
.A2(n_1797),
.B1(n_1656),
.B2(n_1689),
.Y(n_1914)
);

AOI22xp33_ASAP7_75t_L g1915 ( 
.A1(n_1792),
.A2(n_1800),
.B1(n_1794),
.B2(n_1777),
.Y(n_1915)
);

OAI22xp5_ASAP7_75t_L g1916 ( 
.A1(n_1779),
.A2(n_1688),
.B1(n_1683),
.B2(n_1636),
.Y(n_1916)
);

OR2x6_ASAP7_75t_L g1917 ( 
.A(n_1697),
.B(n_1684),
.Y(n_1917)
);

AOI22xp33_ASAP7_75t_L g1918 ( 
.A1(n_1791),
.A2(n_1708),
.B1(n_1710),
.B2(n_1697),
.Y(n_1918)
);

AND2x2_ASAP7_75t_L g1919 ( 
.A(n_1759),
.B(n_1766),
.Y(n_1919)
);

AOI21x1_ASAP7_75t_L g1920 ( 
.A1(n_1640),
.A2(n_1732),
.B(n_1675),
.Y(n_1920)
);

CKINVDCx5p33_ASAP7_75t_R g1921 ( 
.A(n_1617),
.Y(n_1921)
);

OAI22xp5_ASAP7_75t_L g1922 ( 
.A1(n_1683),
.A2(n_1636),
.B1(n_1653),
.B2(n_1666),
.Y(n_1922)
);

INVx2_ASAP7_75t_L g1923 ( 
.A(n_1703),
.Y(n_1923)
);

OAI22xp5_ASAP7_75t_L g1924 ( 
.A1(n_1653),
.A2(n_1666),
.B1(n_1644),
.B2(n_1671),
.Y(n_1924)
);

AOI22xp33_ASAP7_75t_SL g1925 ( 
.A1(n_1656),
.A2(n_1661),
.B1(n_1723),
.B2(n_1697),
.Y(n_1925)
);

AOI22xp33_ASAP7_75t_L g1926 ( 
.A1(n_1708),
.A2(n_1710),
.B1(n_1723),
.B2(n_1689),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1685),
.Y(n_1927)
);

INVx2_ASAP7_75t_L g1928 ( 
.A(n_1703),
.Y(n_1928)
);

AO21x2_ASAP7_75t_L g1929 ( 
.A1(n_1645),
.A2(n_1732),
.B(n_1692),
.Y(n_1929)
);

AOI22xp33_ASAP7_75t_SL g1930 ( 
.A1(n_1656),
.A2(n_1689),
.B1(n_1710),
.B2(n_1662),
.Y(n_1930)
);

AOI22xp33_ASAP7_75t_L g1931 ( 
.A1(n_1698),
.A2(n_1749),
.B1(n_1658),
.B2(n_1715),
.Y(n_1931)
);

A2O1A1Ixp33_ASAP7_75t_L g1932 ( 
.A1(n_1720),
.A2(n_1643),
.B(n_1753),
.C(n_1673),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1706),
.Y(n_1933)
);

AOI22xp33_ASAP7_75t_L g1934 ( 
.A1(n_1698),
.A2(n_1749),
.B1(n_1658),
.B2(n_1673),
.Y(n_1934)
);

NOR2xp33_ASAP7_75t_L g1935 ( 
.A(n_1679),
.B(n_1736),
.Y(n_1935)
);

AOI21xp5_ASAP7_75t_L g1936 ( 
.A1(n_1674),
.A2(n_1639),
.B(n_1726),
.Y(n_1936)
);

AND2x2_ASAP7_75t_L g1937 ( 
.A(n_1698),
.B(n_1749),
.Y(n_1937)
);

AOI22xp33_ASAP7_75t_L g1938 ( 
.A1(n_1698),
.A2(n_1749),
.B1(n_1658),
.B2(n_1668),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1632),
.Y(n_1939)
);

OAI22xp5_ASAP7_75t_L g1940 ( 
.A1(n_1644),
.A2(n_1790),
.B1(n_1788),
.B2(n_1603),
.Y(n_1940)
);

AOI22xp33_ASAP7_75t_L g1941 ( 
.A1(n_1658),
.A2(n_1721),
.B1(n_1713),
.B2(n_1718),
.Y(n_1941)
);

AOI21xp5_ASAP7_75t_L g1942 ( 
.A1(n_1628),
.A2(n_1608),
.B(n_1751),
.Y(n_1942)
);

AND2x6_ASAP7_75t_L g1943 ( 
.A(n_1802),
.B(n_1719),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1713),
.Y(n_1944)
);

OAI22xp33_ASAP7_75t_L g1945 ( 
.A1(n_1707),
.A2(n_1608),
.B1(n_1649),
.B2(n_1790),
.Y(n_1945)
);

BUFx2_ASAP7_75t_L g1946 ( 
.A(n_1761),
.Y(n_1946)
);

NAND2xp5_ASAP7_75t_L g1947 ( 
.A(n_1778),
.B(n_1789),
.Y(n_1947)
);

AOI22xp33_ASAP7_75t_SL g1948 ( 
.A1(n_1802),
.A2(n_1707),
.B1(n_1761),
.B2(n_1615),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_L g1949 ( 
.A(n_1776),
.B(n_1730),
.Y(n_1949)
);

BUFx3_ASAP7_75t_L g1950 ( 
.A(n_1776),
.Y(n_1950)
);

AOI22xp33_ASAP7_75t_L g1951 ( 
.A1(n_1718),
.A2(n_1721),
.B1(n_1769),
.B2(n_1669),
.Y(n_1951)
);

AOI221xp5_ASAP7_75t_L g1952 ( 
.A1(n_1744),
.A2(n_1798),
.B1(n_1606),
.B2(n_1700),
.C(n_1605),
.Y(n_1952)
);

INVx3_ASAP7_75t_L g1953 ( 
.A(n_1776),
.Y(n_1953)
);

AOI22xp33_ASAP7_75t_L g1954 ( 
.A1(n_1769),
.A2(n_1669),
.B1(n_1700),
.B2(n_1678),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1786),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1670),
.Y(n_1956)
);

AND2x2_ASAP7_75t_L g1957 ( 
.A(n_1730),
.B(n_1795),
.Y(n_1957)
);

AOI22xp33_ASAP7_75t_SL g1958 ( 
.A1(n_1640),
.A2(n_1664),
.B1(n_1678),
.B2(n_1776),
.Y(n_1958)
);

AND2x2_ASAP7_75t_L g1959 ( 
.A(n_1782),
.B(n_1795),
.Y(n_1959)
);

OAI21xp33_ASAP7_75t_L g1960 ( 
.A1(n_1610),
.A2(n_1751),
.B(n_1782),
.Y(n_1960)
);

AOI33xp33_ASAP7_75t_L g1961 ( 
.A1(n_1610),
.A2(n_736),
.A3(n_1728),
.B1(n_1717),
.B2(n_1781),
.B3(n_1770),
.Y(n_1961)
);

AO21x2_ASAP7_75t_L g1962 ( 
.A1(n_1640),
.A2(n_1670),
.B(n_1664),
.Y(n_1962)
);

AND2x2_ASAP7_75t_L g1963 ( 
.A(n_1670),
.B(n_1664),
.Y(n_1963)
);

AND2x2_ASAP7_75t_L g1964 ( 
.A(n_1670),
.B(n_1602),
.Y(n_1964)
);

AND2x4_ASAP7_75t_L g1965 ( 
.A(n_1769),
.B(n_1598),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1599),
.Y(n_1966)
);

AOI22xp33_ASAP7_75t_L g1967 ( 
.A1(n_1622),
.A2(n_1609),
.B1(n_1562),
.B2(n_1414),
.Y(n_1967)
);

OAI22xp5_ASAP7_75t_L g1968 ( 
.A1(n_1612),
.A2(n_1562),
.B1(n_1414),
.B2(n_1274),
.Y(n_1968)
);

OAI22xp5_ASAP7_75t_L g1969 ( 
.A1(n_1612),
.A2(n_1562),
.B1(n_1414),
.B2(n_1274),
.Y(n_1969)
);

INVx5_ASAP7_75t_SL g1970 ( 
.A(n_1739),
.Y(n_1970)
);

OAI22xp33_ASAP7_75t_L g1971 ( 
.A1(n_1609),
.A2(n_1497),
.B1(n_1612),
.B2(n_1611),
.Y(n_1971)
);

AOI21xp5_ASAP7_75t_L g1972 ( 
.A1(n_1711),
.A2(n_1489),
.B(n_1696),
.Y(n_1972)
);

OAI22xp33_ASAP7_75t_L g1973 ( 
.A1(n_1609),
.A2(n_1497),
.B1(n_1612),
.B2(n_1611),
.Y(n_1973)
);

AOI221xp5_ASAP7_75t_L g1974 ( 
.A1(n_1609),
.A2(n_1211),
.B1(n_1282),
.B2(n_736),
.C(n_502),
.Y(n_1974)
);

OAI22xp5_ASAP7_75t_L g1975 ( 
.A1(n_1612),
.A2(n_1562),
.B1(n_1414),
.B2(n_1274),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_L g1976 ( 
.A(n_1602),
.B(n_1500),
.Y(n_1976)
);

AOI22xp33_ASAP7_75t_L g1977 ( 
.A1(n_1622),
.A2(n_1609),
.B1(n_1562),
.B2(n_1414),
.Y(n_1977)
);

OAI211xp5_ASAP7_75t_SL g1978 ( 
.A1(n_1717),
.A2(n_1282),
.B(n_1067),
.C(n_1165),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1599),
.Y(n_1979)
);

INVx3_ASAP7_75t_L g1980 ( 
.A(n_1643),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_L g1981 ( 
.A(n_1602),
.B(n_1500),
.Y(n_1981)
);

NAND3xp33_ASAP7_75t_L g1982 ( 
.A(n_1622),
.B(n_1717),
.C(n_1630),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_L g1983 ( 
.A(n_1602),
.B(n_1500),
.Y(n_1983)
);

OAI221xp5_ASAP7_75t_L g1984 ( 
.A1(n_1630),
.A2(n_1414),
.B1(n_1282),
.B2(n_1562),
.C(n_869),
.Y(n_1984)
);

AOI22xp33_ASAP7_75t_L g1985 ( 
.A1(n_1622),
.A2(n_1609),
.B1(n_1562),
.B2(n_1414),
.Y(n_1985)
);

AOI22xp33_ASAP7_75t_L g1986 ( 
.A1(n_1622),
.A2(n_1609),
.B1(n_1562),
.B2(n_1414),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1599),
.Y(n_1987)
);

OAI221xp5_ASAP7_75t_L g1988 ( 
.A1(n_1630),
.A2(n_1414),
.B1(n_1282),
.B2(n_1562),
.C(n_869),
.Y(n_1988)
);

OAI22xp5_ASAP7_75t_L g1989 ( 
.A1(n_1612),
.A2(n_1562),
.B1(n_1414),
.B2(n_1274),
.Y(n_1989)
);

HB1xp67_ASAP7_75t_L g1990 ( 
.A(n_1632),
.Y(n_1990)
);

INVx2_ASAP7_75t_L g1991 ( 
.A(n_1729),
.Y(n_1991)
);

AOI22xp33_ASAP7_75t_SL g1992 ( 
.A1(n_1622),
.A2(n_1620),
.B1(n_477),
.B2(n_481),
.Y(n_1992)
);

OAI211xp5_ASAP7_75t_L g1993 ( 
.A1(n_1728),
.A2(n_1282),
.B(n_1414),
.C(n_1218),
.Y(n_1993)
);

AOI22xp33_ASAP7_75t_L g1994 ( 
.A1(n_1622),
.A2(n_1609),
.B1(n_1562),
.B2(n_1414),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_L g1995 ( 
.A(n_1602),
.B(n_1500),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1599),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_L g1997 ( 
.A(n_1976),
.B(n_1981),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1939),
.Y(n_1998)
);

AND2x4_ASAP7_75t_L g1999 ( 
.A(n_1917),
.B(n_1870),
.Y(n_1999)
);

AND2x2_ASAP7_75t_L g2000 ( 
.A(n_1853),
.B(n_1871),
.Y(n_2000)
);

AND2x2_ASAP7_75t_L g2001 ( 
.A(n_1964),
.B(n_1843),
.Y(n_2001)
);

HB1xp67_ASAP7_75t_L g2002 ( 
.A(n_1990),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1836),
.Y(n_2003)
);

AND2x2_ASAP7_75t_L g2004 ( 
.A(n_1832),
.B(n_1820),
.Y(n_2004)
);

OAI22xp33_ASAP7_75t_L g2005 ( 
.A1(n_1982),
.A2(n_1819),
.B1(n_1817),
.B2(n_1984),
.Y(n_2005)
);

OR2x2_ASAP7_75t_L g2006 ( 
.A(n_1811),
.B(n_1860),
.Y(n_2006)
);

BUFx3_ASAP7_75t_L g2007 ( 
.A(n_1837),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_L g2008 ( 
.A(n_1983),
.B(n_1995),
.Y(n_2008)
);

AND2x4_ASAP7_75t_L g2009 ( 
.A(n_1917),
.B(n_1824),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1849),
.Y(n_2010)
);

AND2x2_ASAP7_75t_L g2011 ( 
.A(n_1878),
.B(n_1851),
.Y(n_2011)
);

INVx2_ASAP7_75t_SL g2012 ( 
.A(n_1980),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1856),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1966),
.Y(n_2014)
);

AOI22xp33_ASAP7_75t_L g2015 ( 
.A1(n_1992),
.A2(n_1826),
.B1(n_1994),
.B2(n_1985),
.Y(n_2015)
);

INVxp67_ASAP7_75t_L g2016 ( 
.A(n_1935),
.Y(n_2016)
);

AO31x2_ASAP7_75t_L g2017 ( 
.A1(n_1840),
.A2(n_1844),
.A3(n_1857),
.B(n_1854),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_L g2018 ( 
.A(n_1935),
.B(n_1897),
.Y(n_2018)
);

AND2x2_ASAP7_75t_L g2019 ( 
.A(n_1979),
.B(n_1987),
.Y(n_2019)
);

BUFx6f_ASAP7_75t_SL g2020 ( 
.A(n_1824),
.Y(n_2020)
);

HB1xp67_ASAP7_75t_L g2021 ( 
.A(n_1913),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1996),
.Y(n_2022)
);

OR2x2_ASAP7_75t_L g2023 ( 
.A(n_1882),
.B(n_1917),
.Y(n_2023)
);

AND2x6_ASAP7_75t_L g2024 ( 
.A(n_1970),
.B(n_1965),
.Y(n_2024)
);

AND2x2_ASAP7_75t_L g2025 ( 
.A(n_1907),
.B(n_1919),
.Y(n_2025)
);

INVx1_ASAP7_75t_SL g2026 ( 
.A(n_1827),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1862),
.Y(n_2027)
);

OR2x2_ASAP7_75t_SL g2028 ( 
.A(n_1837),
.B(n_1891),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1868),
.Y(n_2029)
);

INVxp67_ASAP7_75t_R g2030 ( 
.A(n_1924),
.Y(n_2030)
);

AND2x2_ASAP7_75t_L g2031 ( 
.A(n_1885),
.B(n_1929),
.Y(n_2031)
);

AOI22xp33_ASAP7_75t_L g2032 ( 
.A1(n_1967),
.A2(n_1994),
.B1(n_1977),
.B2(n_1985),
.Y(n_2032)
);

INVx2_ASAP7_75t_SL g2033 ( 
.A(n_1980),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1873),
.Y(n_2034)
);

AO31x2_ASAP7_75t_L g2035 ( 
.A1(n_1845),
.A2(n_1972),
.A3(n_1956),
.B(n_1867),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_1879),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_L g2037 ( 
.A(n_1815),
.B(n_1946),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1881),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1903),
.Y(n_2039)
);

AOI22xp33_ASAP7_75t_L g2040 ( 
.A1(n_1967),
.A2(n_1977),
.B1(n_1986),
.B2(n_1973),
.Y(n_2040)
);

OR2x6_ASAP7_75t_L g2041 ( 
.A(n_1905),
.B(n_1824),
.Y(n_2041)
);

AND2x2_ASAP7_75t_L g2042 ( 
.A(n_1929),
.B(n_1815),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_1904),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_1911),
.Y(n_2044)
);

INVx3_ASAP7_75t_L g2045 ( 
.A(n_1943),
.Y(n_2045)
);

INVx6_ASAP7_75t_L g2046 ( 
.A(n_1837),
.Y(n_2046)
);

BUFx6f_ASAP7_75t_L g2047 ( 
.A(n_1850),
.Y(n_2047)
);

OR2x2_ASAP7_75t_L g2048 ( 
.A(n_1876),
.B(n_1899),
.Y(n_2048)
);

INVx4_ASAP7_75t_R g2049 ( 
.A(n_1937),
.Y(n_2049)
);

AND2x2_ASAP7_75t_L g2050 ( 
.A(n_1809),
.B(n_1828),
.Y(n_2050)
);

INVx3_ASAP7_75t_L g2051 ( 
.A(n_1943),
.Y(n_2051)
);

AND2x2_ASAP7_75t_L g2052 ( 
.A(n_1809),
.B(n_1828),
.Y(n_2052)
);

AOI22xp33_ASAP7_75t_L g2053 ( 
.A1(n_1986),
.A2(n_1971),
.B1(n_1822),
.B2(n_1974),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_1927),
.Y(n_2054)
);

HB1xp67_ASAP7_75t_L g2055 ( 
.A(n_1947),
.Y(n_2055)
);

OR2x2_ASAP7_75t_L g2056 ( 
.A(n_1991),
.B(n_1893),
.Y(n_2056)
);

AND2x2_ASAP7_75t_L g2057 ( 
.A(n_1963),
.B(n_1893),
.Y(n_2057)
);

AND2x2_ASAP7_75t_L g2058 ( 
.A(n_1920),
.B(n_1807),
.Y(n_2058)
);

AND2x2_ASAP7_75t_L g2059 ( 
.A(n_1807),
.B(n_1931),
.Y(n_2059)
);

BUFx2_ASAP7_75t_L g2060 ( 
.A(n_1943),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_1933),
.Y(n_2061)
);

INVx3_ASAP7_75t_L g2062 ( 
.A(n_1943),
.Y(n_2062)
);

AOI22xp5_ASAP7_75t_L g2063 ( 
.A1(n_1968),
.A2(n_1989),
.B1(n_1975),
.B2(n_1969),
.Y(n_2063)
);

INVx2_ASAP7_75t_L g2064 ( 
.A(n_1923),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_1944),
.Y(n_2065)
);

INVx3_ASAP7_75t_L g2066 ( 
.A(n_1943),
.Y(n_2066)
);

INVx2_ASAP7_75t_L g2067 ( 
.A(n_1928),
.Y(n_2067)
);

INVx2_ASAP7_75t_SL g2068 ( 
.A(n_1950),
.Y(n_2068)
);

AND2x2_ASAP7_75t_L g2069 ( 
.A(n_1931),
.B(n_1934),
.Y(n_2069)
);

AND2x4_ASAP7_75t_SL g2070 ( 
.A(n_1957),
.B(n_1959),
.Y(n_2070)
);

INVx1_ASAP7_75t_SL g2071 ( 
.A(n_1892),
.Y(n_2071)
);

BUFx2_ASAP7_75t_L g2072 ( 
.A(n_1950),
.Y(n_2072)
);

NOR2x1_ASAP7_75t_SL g2073 ( 
.A(n_1922),
.B(n_1940),
.Y(n_2073)
);

OR2x2_ASAP7_75t_L g2074 ( 
.A(n_1909),
.B(n_1934),
.Y(n_2074)
);

INVx2_ASAP7_75t_SL g2075 ( 
.A(n_1953),
.Y(n_2075)
);

AND2x2_ASAP7_75t_L g2076 ( 
.A(n_1938),
.B(n_1958),
.Y(n_2076)
);

OR2x2_ASAP7_75t_L g2077 ( 
.A(n_1909),
.B(n_1938),
.Y(n_2077)
);

BUFx2_ASAP7_75t_L g2078 ( 
.A(n_1953),
.Y(n_2078)
);

AND2x2_ASAP7_75t_L g2079 ( 
.A(n_1808),
.B(n_1835),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_1912),
.Y(n_2080)
);

INVx2_ASAP7_75t_L g2081 ( 
.A(n_1900),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_1910),
.Y(n_2082)
);

INVx3_ASAP7_75t_L g2083 ( 
.A(n_1869),
.Y(n_2083)
);

OR2x2_ASAP7_75t_L g2084 ( 
.A(n_1962),
.B(n_1808),
.Y(n_2084)
);

OR2x2_ASAP7_75t_L g2085 ( 
.A(n_1962),
.B(n_1916),
.Y(n_2085)
);

BUFx3_ASAP7_75t_L g2086 ( 
.A(n_1823),
.Y(n_2086)
);

OAI22xp33_ASAP7_75t_L g2087 ( 
.A1(n_1988),
.A2(n_1825),
.B1(n_1865),
.B2(n_1895),
.Y(n_2087)
);

OR2x2_ASAP7_75t_L g2088 ( 
.A(n_1970),
.B(n_1936),
.Y(n_2088)
);

OAI22xp5_ASAP7_75t_L g2089 ( 
.A1(n_1822),
.A2(n_1842),
.B1(n_1993),
.B2(n_1898),
.Y(n_2089)
);

INVx2_ASAP7_75t_SL g2090 ( 
.A(n_1949),
.Y(n_2090)
);

AND2x2_ASAP7_75t_L g2091 ( 
.A(n_1835),
.B(n_1918),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_1908),
.Y(n_2092)
);

OR2x2_ASAP7_75t_L g2093 ( 
.A(n_1970),
.B(n_1839),
.Y(n_2093)
);

INVx2_ASAP7_75t_SL g2094 ( 
.A(n_1955),
.Y(n_2094)
);

AND2x2_ASAP7_75t_L g2095 ( 
.A(n_1918),
.B(n_1841),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_1960),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_1805),
.Y(n_2097)
);

AND2x2_ASAP7_75t_L g2098 ( 
.A(n_1841),
.B(n_1915),
.Y(n_2098)
);

BUFx3_ASAP7_75t_L g2099 ( 
.A(n_1888),
.Y(n_2099)
);

NAND2xp5_ASAP7_75t_L g2100 ( 
.A(n_1915),
.B(n_1942),
.Y(n_2100)
);

AND2x2_ASAP7_75t_L g2101 ( 
.A(n_1829),
.B(n_1852),
.Y(n_2101)
);

OAI221xp5_ASAP7_75t_L g2102 ( 
.A1(n_1978),
.A2(n_1894),
.B1(n_1890),
.B2(n_1831),
.C(n_1889),
.Y(n_2102)
);

NAND2xp5_ASAP7_75t_L g2103 ( 
.A(n_1961),
.B(n_1812),
.Y(n_2103)
);

OR2x2_ASAP7_75t_L g2104 ( 
.A(n_1816),
.B(n_1861),
.Y(n_2104)
);

CKINVDCx11_ASAP7_75t_R g2105 ( 
.A(n_1901),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_L g2106 ( 
.A(n_1961),
.B(n_1902),
.Y(n_2106)
);

AND2x2_ASAP7_75t_L g2107 ( 
.A(n_1852),
.B(n_1883),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_1806),
.Y(n_2108)
);

AND2x4_ASAP7_75t_L g2109 ( 
.A(n_1954),
.B(n_1951),
.Y(n_2109)
);

BUFx3_ASAP7_75t_L g2110 ( 
.A(n_1921),
.Y(n_2110)
);

NAND3xp33_ASAP7_75t_L g2111 ( 
.A(n_1872),
.B(n_1858),
.C(n_1816),
.Y(n_2111)
);

OR2x2_ASAP7_75t_L g2112 ( 
.A(n_2006),
.B(n_1821),
.Y(n_2112)
);

OR2x2_ASAP7_75t_L g2113 ( 
.A(n_2006),
.B(n_1821),
.Y(n_2113)
);

INVx2_ASAP7_75t_L g2114 ( 
.A(n_2056),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_2013),
.Y(n_2115)
);

INVx2_ASAP7_75t_L g2116 ( 
.A(n_2056),
.Y(n_2116)
);

NAND2xp5_ASAP7_75t_L g2117 ( 
.A(n_2002),
.B(n_1810),
.Y(n_2117)
);

AND2x2_ASAP7_75t_SL g2118 ( 
.A(n_2009),
.B(n_1926),
.Y(n_2118)
);

OAI21xp5_ASAP7_75t_SL g2119 ( 
.A1(n_2063),
.A2(n_1896),
.B(n_1906),
.Y(n_2119)
);

OA222x2_ASAP7_75t_L g2120 ( 
.A1(n_2041),
.A2(n_1948),
.B1(n_1945),
.B2(n_1925),
.C1(n_1926),
.C2(n_1914),
.Y(n_2120)
);

OAI22xp33_ASAP7_75t_L g2121 ( 
.A1(n_2106),
.A2(n_1838),
.B1(n_1834),
.B2(n_1818),
.Y(n_2121)
);

BUFx2_ASAP7_75t_L g2122 ( 
.A(n_2099),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_2013),
.Y(n_2123)
);

INVx2_ASAP7_75t_L g2124 ( 
.A(n_2081),
.Y(n_2124)
);

INVxp67_ASAP7_75t_L g2125 ( 
.A(n_2021),
.Y(n_2125)
);

CKINVDCx8_ASAP7_75t_R g2126 ( 
.A(n_2024),
.Y(n_2126)
);

INVx2_ASAP7_75t_SL g2127 ( 
.A(n_2049),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_2014),
.Y(n_2128)
);

AND2x2_ASAP7_75t_L g2129 ( 
.A(n_2025),
.B(n_1875),
.Y(n_2129)
);

AND2x2_ASAP7_75t_L g2130 ( 
.A(n_2025),
.B(n_2000),
.Y(n_2130)
);

NAND2xp33_ASAP7_75t_SL g2131 ( 
.A(n_2060),
.B(n_1951),
.Y(n_2131)
);

NAND3xp33_ASAP7_75t_L g2132 ( 
.A(n_2082),
.B(n_1813),
.C(n_1814),
.Y(n_2132)
);

OAI33xp33_ASAP7_75t_L g2133 ( 
.A1(n_2005),
.A2(n_2087),
.A3(n_2089),
.B1(n_2092),
.B2(n_2080),
.B3(n_2097),
.Y(n_2133)
);

NAND4xp25_ASAP7_75t_L g2134 ( 
.A(n_2032),
.B(n_1932),
.C(n_1814),
.D(n_1859),
.Y(n_2134)
);

INVx2_ASAP7_75t_SL g2135 ( 
.A(n_2070),
.Y(n_2135)
);

NAND2xp5_ASAP7_75t_L g2136 ( 
.A(n_2018),
.B(n_2055),
.Y(n_2136)
);

OAI22xp33_ASAP7_75t_L g2137 ( 
.A1(n_2102),
.A2(n_1833),
.B1(n_1877),
.B2(n_1880),
.Y(n_2137)
);

AND2x2_ASAP7_75t_L g2138 ( 
.A(n_2000),
.B(n_2004),
.Y(n_2138)
);

AOI22xp5_ASAP7_75t_L g2139 ( 
.A1(n_2040),
.A2(n_1930),
.B1(n_1864),
.B2(n_1810),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_2014),
.Y(n_2140)
);

NOR2xp33_ASAP7_75t_L g2141 ( 
.A(n_2016),
.B(n_1932),
.Y(n_2141)
);

NOR2xp33_ASAP7_75t_L g2142 ( 
.A(n_2037),
.B(n_1830),
.Y(n_2142)
);

OAI22xp5_ASAP7_75t_L g2143 ( 
.A1(n_2053),
.A2(n_1864),
.B1(n_1954),
.B2(n_1883),
.Y(n_2143)
);

OAI211xp5_ASAP7_75t_L g2144 ( 
.A1(n_2015),
.A2(n_1863),
.B(n_1848),
.C(n_1886),
.Y(n_2144)
);

AO21x2_ASAP7_75t_L g2145 ( 
.A1(n_2111),
.A2(n_1846),
.B(n_1847),
.Y(n_2145)
);

CKINVDCx20_ASAP7_75t_R g2146 ( 
.A(n_2110),
.Y(n_2146)
);

OAI221xp5_ASAP7_75t_L g2147 ( 
.A1(n_2080),
.A2(n_2103),
.B1(n_2108),
.B2(n_2084),
.C(n_2058),
.Y(n_2147)
);

OAI322xp33_ASAP7_75t_L g2148 ( 
.A1(n_2085),
.A2(n_1887),
.A3(n_1884),
.B1(n_1848),
.B2(n_1941),
.C1(n_1874),
.C2(n_1866),
.Y(n_2148)
);

NAND3xp33_ASAP7_75t_L g2149 ( 
.A(n_2058),
.B(n_1874),
.C(n_1941),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_2022),
.Y(n_2150)
);

NAND3xp33_ASAP7_75t_L g2151 ( 
.A(n_2096),
.B(n_2042),
.C(n_2085),
.Y(n_2151)
);

HB1xp67_ASAP7_75t_L g2152 ( 
.A(n_2031),
.Y(n_2152)
);

OAI22xp5_ASAP7_75t_L g2153 ( 
.A1(n_2099),
.A2(n_1866),
.B1(n_1855),
.B2(n_1952),
.Y(n_2153)
);

INVx3_ASAP7_75t_L g2154 ( 
.A(n_2045),
.Y(n_2154)
);

OAI33xp33_ASAP7_75t_L g2155 ( 
.A1(n_2084),
.A2(n_1855),
.A3(n_1997),
.B1(n_2008),
.B2(n_2104),
.B3(n_2010),
.Y(n_2155)
);

A2O1A1Ixp33_ASAP7_75t_L g2156 ( 
.A1(n_2101),
.A2(n_2079),
.B(n_2107),
.C(n_2050),
.Y(n_2156)
);

CKINVDCx5p33_ASAP7_75t_R g2157 ( 
.A(n_2110),
.Y(n_2157)
);

CKINVDCx16_ASAP7_75t_R g2158 ( 
.A(n_2020),
.Y(n_2158)
);

AND2x2_ASAP7_75t_L g2159 ( 
.A(n_2004),
.B(n_2001),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_2022),
.Y(n_2160)
);

HB1xp67_ASAP7_75t_L g2161 ( 
.A(n_2031),
.Y(n_2161)
);

INVx3_ASAP7_75t_L g2162 ( 
.A(n_2045),
.Y(n_2162)
);

NOR4xp25_ASAP7_75t_SL g2163 ( 
.A(n_2060),
.B(n_2072),
.C(n_2078),
.D(n_2073),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_2034),
.Y(n_2164)
);

OAI33xp33_ASAP7_75t_L g2165 ( 
.A1(n_2104),
.A2(n_2003),
.A3(n_1998),
.B1(n_2100),
.B2(n_2036),
.B3(n_2054),
.Y(n_2165)
);

OR2x2_ASAP7_75t_L g2166 ( 
.A(n_2001),
.B(n_2011),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_2034),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_2039),
.Y(n_2168)
);

INVx2_ASAP7_75t_L g2169 ( 
.A(n_2064),
.Y(n_2169)
);

OAI221xp5_ASAP7_75t_L g2170 ( 
.A1(n_2101),
.A2(n_2052),
.B1(n_2050),
.B2(n_2079),
.C(n_2093),
.Y(n_2170)
);

OAI332xp33_ASAP7_75t_L g2171 ( 
.A1(n_2071),
.A2(n_2088),
.A3(n_2093),
.B1(n_2077),
.B2(n_2074),
.B3(n_2029),
.C1(n_2038),
.C2(n_2027),
.Y(n_2171)
);

OAI21xp33_ASAP7_75t_L g2172 ( 
.A1(n_2042),
.A2(n_2107),
.B(n_2052),
.Y(n_2172)
);

BUFx6f_ASAP7_75t_L g2173 ( 
.A(n_2007),
.Y(n_2173)
);

BUFx3_ASAP7_75t_L g2174 ( 
.A(n_2046),
.Y(n_2174)
);

OAI31xp33_ASAP7_75t_L g2175 ( 
.A1(n_2091),
.A2(n_2098),
.A3(n_2095),
.B(n_2076),
.Y(n_2175)
);

OAI33xp33_ASAP7_75t_L g2176 ( 
.A1(n_2061),
.A2(n_2039),
.A3(n_2043),
.B1(n_2044),
.B2(n_2065),
.B3(n_2074),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_2043),
.Y(n_2177)
);

NAND2xp5_ASAP7_75t_L g2178 ( 
.A(n_2011),
.B(n_2090),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_2044),
.Y(n_2179)
);

AOI22xp33_ASAP7_75t_L g2180 ( 
.A1(n_2091),
.A2(n_2095),
.B1(n_2098),
.B2(n_2059),
.Y(n_2180)
);

AND2x2_ASAP7_75t_L g2181 ( 
.A(n_1999),
.B(n_2019),
.Y(n_2181)
);

NAND2xp33_ASAP7_75t_R g2182 ( 
.A(n_2041),
.B(n_2062),
.Y(n_2182)
);

BUFx10_ASAP7_75t_L g2183 ( 
.A(n_2046),
.Y(n_2183)
);

HB1xp67_ASAP7_75t_L g2184 ( 
.A(n_2019),
.Y(n_2184)
);

INVx2_ASAP7_75t_L g2185 ( 
.A(n_2067),
.Y(n_2185)
);

OAI211xp5_ASAP7_75t_L g2186 ( 
.A1(n_2105),
.A2(n_2076),
.B(n_2057),
.C(n_2023),
.Y(n_2186)
);

AND4x1_ASAP7_75t_L g2187 ( 
.A(n_2073),
.B(n_2028),
.C(n_2030),
.D(n_2059),
.Y(n_2187)
);

OAI211xp5_ASAP7_75t_L g2188 ( 
.A1(n_2105),
.A2(n_2057),
.B(n_2023),
.C(n_2088),
.Y(n_2188)
);

AND2x2_ASAP7_75t_L g2189 ( 
.A(n_1999),
.B(n_2017),
.Y(n_2189)
);

NOR2xp33_ASAP7_75t_L g2190 ( 
.A(n_2026),
.B(n_2086),
.Y(n_2190)
);

AND2x4_ASAP7_75t_L g2191 ( 
.A(n_2009),
.B(n_2062),
.Y(n_2191)
);

NAND4xp25_ASAP7_75t_L g2192 ( 
.A(n_2086),
.B(n_2078),
.C(n_2083),
.D(n_2072),
.Y(n_2192)
);

NAND2xp5_ASAP7_75t_L g2193 ( 
.A(n_2141),
.B(n_2035),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_2115),
.Y(n_2194)
);

AND2x2_ASAP7_75t_L g2195 ( 
.A(n_2189),
.B(n_2017),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_2123),
.Y(n_2196)
);

AND2x2_ASAP7_75t_L g2197 ( 
.A(n_2189),
.B(n_2017),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_2128),
.Y(n_2198)
);

AND2x2_ASAP7_75t_L g2199 ( 
.A(n_2159),
.B(n_2017),
.Y(n_2199)
);

AND2x2_ASAP7_75t_L g2200 ( 
.A(n_2159),
.B(n_2138),
.Y(n_2200)
);

NOR2x1_ASAP7_75t_L g2201 ( 
.A(n_2192),
.B(n_2062),
.Y(n_2201)
);

INVx2_ASAP7_75t_L g2202 ( 
.A(n_2114),
.Y(n_2202)
);

AND2x2_ASAP7_75t_L g2203 ( 
.A(n_2138),
.B(n_2017),
.Y(n_2203)
);

OR2x2_ASAP7_75t_L g2204 ( 
.A(n_2184),
.B(n_2035),
.Y(n_2204)
);

INVx2_ASAP7_75t_L g2205 ( 
.A(n_2114),
.Y(n_2205)
);

OR2x2_ASAP7_75t_L g2206 ( 
.A(n_2166),
.B(n_2035),
.Y(n_2206)
);

INVx2_ASAP7_75t_L g2207 ( 
.A(n_2116),
.Y(n_2207)
);

OR2x2_ASAP7_75t_L g2208 ( 
.A(n_2136),
.B(n_2035),
.Y(n_2208)
);

OR2x2_ASAP7_75t_L g2209 ( 
.A(n_2152),
.B(n_2161),
.Y(n_2209)
);

AND2x2_ASAP7_75t_L g2210 ( 
.A(n_2130),
.B(n_2035),
.Y(n_2210)
);

AND2x2_ASAP7_75t_L g2211 ( 
.A(n_2130),
.B(n_2129),
.Y(n_2211)
);

INVx2_ASAP7_75t_L g2212 ( 
.A(n_2124),
.Y(n_2212)
);

AND2x2_ASAP7_75t_L g2213 ( 
.A(n_2129),
.B(n_1999),
.Y(n_2213)
);

NAND4xp75_ASAP7_75t_L g2214 ( 
.A(n_2120),
.B(n_2094),
.C(n_2069),
.D(n_2090),
.Y(n_2214)
);

NOR2xp67_ASAP7_75t_L g2215 ( 
.A(n_2151),
.B(n_2051),
.Y(n_2215)
);

AND2x4_ASAP7_75t_L g2216 ( 
.A(n_2154),
.B(n_2051),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_2140),
.Y(n_2217)
);

NAND2xp5_ASAP7_75t_L g2218 ( 
.A(n_2141),
.B(n_2033),
.Y(n_2218)
);

NAND2xp5_ASAP7_75t_L g2219 ( 
.A(n_2142),
.B(n_2012),
.Y(n_2219)
);

INVx1_ASAP7_75t_SL g2220 ( 
.A(n_2122),
.Y(n_2220)
);

NAND2xp5_ASAP7_75t_L g2221 ( 
.A(n_2142),
.B(n_2150),
.Y(n_2221)
);

AND2x2_ASAP7_75t_L g2222 ( 
.A(n_2181),
.B(n_2154),
.Y(n_2222)
);

HB1xp67_ASAP7_75t_L g2223 ( 
.A(n_2160),
.Y(n_2223)
);

INVxp67_ASAP7_75t_L g2224 ( 
.A(n_2145),
.Y(n_2224)
);

NOR2xp33_ASAP7_75t_L g2225 ( 
.A(n_2157),
.B(n_2070),
.Y(n_2225)
);

NAND2xp5_ASAP7_75t_SL g2226 ( 
.A(n_2187),
.B(n_2045),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_2164),
.Y(n_2227)
);

OR2x2_ASAP7_75t_L g2228 ( 
.A(n_2112),
.B(n_2012),
.Y(n_2228)
);

INVxp67_ASAP7_75t_L g2229 ( 
.A(n_2145),
.Y(n_2229)
);

AOI22xp33_ASAP7_75t_L g2230 ( 
.A1(n_2147),
.A2(n_2109),
.B1(n_2069),
.B2(n_2077),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_2167),
.Y(n_2231)
);

AND2x2_ASAP7_75t_L g2232 ( 
.A(n_2162),
.B(n_2083),
.Y(n_2232)
);

BUFx2_ASAP7_75t_L g2233 ( 
.A(n_2162),
.Y(n_2233)
);

BUFx2_ASAP7_75t_L g2234 ( 
.A(n_2162),
.Y(n_2234)
);

INVxp67_ASAP7_75t_SL g2235 ( 
.A(n_2117),
.Y(n_2235)
);

AND2x4_ASAP7_75t_L g2236 ( 
.A(n_2191),
.B(n_2066),
.Y(n_2236)
);

OR2x2_ASAP7_75t_L g2237 ( 
.A(n_2113),
.B(n_2094),
.Y(n_2237)
);

AND2x2_ASAP7_75t_L g2238 ( 
.A(n_2178),
.B(n_2083),
.Y(n_2238)
);

HB1xp67_ASAP7_75t_L g2239 ( 
.A(n_2168),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_2177),
.Y(n_2240)
);

INVxp67_ASAP7_75t_L g2241 ( 
.A(n_2145),
.Y(n_2241)
);

AND2x2_ASAP7_75t_L g2242 ( 
.A(n_2191),
.B(n_2030),
.Y(n_2242)
);

AND2x2_ASAP7_75t_L g2243 ( 
.A(n_2191),
.B(n_2009),
.Y(n_2243)
);

INVx1_ASAP7_75t_L g2244 ( 
.A(n_2179),
.Y(n_2244)
);

AND2x2_ASAP7_75t_L g2245 ( 
.A(n_2163),
.B(n_2066),
.Y(n_2245)
);

AND2x4_ASAP7_75t_L g2246 ( 
.A(n_2135),
.B(n_2066),
.Y(n_2246)
);

AND2x2_ASAP7_75t_L g2247 ( 
.A(n_2135),
.B(n_2068),
.Y(n_2247)
);

OR2x2_ASAP7_75t_L g2248 ( 
.A(n_2125),
.B(n_2172),
.Y(n_2248)
);

NAND2xp5_ASAP7_75t_L g2249 ( 
.A(n_2156),
.B(n_2068),
.Y(n_2249)
);

OR2x2_ASAP7_75t_L g2250 ( 
.A(n_2149),
.B(n_2028),
.Y(n_2250)
);

NAND2xp5_ASAP7_75t_L g2251 ( 
.A(n_2156),
.B(n_2075),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_2169),
.Y(n_2252)
);

NAND2xp5_ASAP7_75t_L g2253 ( 
.A(n_2180),
.B(n_2075),
.Y(n_2253)
);

OR2x2_ASAP7_75t_L g2254 ( 
.A(n_2153),
.B(n_2048),
.Y(n_2254)
);

NAND2xp5_ASAP7_75t_L g2255 ( 
.A(n_2199),
.B(n_2171),
.Y(n_2255)
);

OAI21xp5_ASAP7_75t_L g2256 ( 
.A1(n_2214),
.A2(n_2229),
.B(n_2224),
.Y(n_2256)
);

AND2x2_ASAP7_75t_L g2257 ( 
.A(n_2199),
.B(n_2127),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_2223),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_2223),
.Y(n_2259)
);

NAND2xp5_ASAP7_75t_L g2260 ( 
.A(n_2199),
.B(n_2137),
.Y(n_2260)
);

NAND2xp5_ASAP7_75t_L g2261 ( 
.A(n_2203),
.B(n_2193),
.Y(n_2261)
);

NAND2xp5_ASAP7_75t_L g2262 ( 
.A(n_2203),
.B(n_2144),
.Y(n_2262)
);

NAND2xp5_ASAP7_75t_L g2263 ( 
.A(n_2203),
.B(n_2175),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_2239),
.Y(n_2264)
);

OR2x2_ASAP7_75t_L g2265 ( 
.A(n_2208),
.B(n_2134),
.Y(n_2265)
);

OR2x2_ASAP7_75t_SL g2266 ( 
.A(n_2193),
.B(n_2158),
.Y(n_2266)
);

HB1xp67_ASAP7_75t_L g2267 ( 
.A(n_2239),
.Y(n_2267)
);

INVx2_ASAP7_75t_L g2268 ( 
.A(n_2195),
.Y(n_2268)
);

NAND2xp5_ASAP7_75t_L g2269 ( 
.A(n_2195),
.B(n_2132),
.Y(n_2269)
);

INVx1_ASAP7_75t_SL g2270 ( 
.A(n_2220),
.Y(n_2270)
);

NAND2xp5_ASAP7_75t_L g2271 ( 
.A(n_2195),
.B(n_2121),
.Y(n_2271)
);

NAND2xp5_ASAP7_75t_L g2272 ( 
.A(n_2197),
.B(n_2190),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_2194),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_2194),
.Y(n_2274)
);

INVx2_ASAP7_75t_L g2275 ( 
.A(n_2197),
.Y(n_2275)
);

INVx2_ASAP7_75t_L g2276 ( 
.A(n_2197),
.Y(n_2276)
);

OAI21xp5_ASAP7_75t_L g2277 ( 
.A1(n_2214),
.A2(n_2119),
.B(n_2170),
.Y(n_2277)
);

INVxp67_ASAP7_75t_L g2278 ( 
.A(n_2253),
.Y(n_2278)
);

INVxp67_ASAP7_75t_SL g2279 ( 
.A(n_2215),
.Y(n_2279)
);

AND2x2_ASAP7_75t_L g2280 ( 
.A(n_2210),
.B(n_2127),
.Y(n_2280)
);

AND2x4_ASAP7_75t_L g2281 ( 
.A(n_2201),
.B(n_2174),
.Y(n_2281)
);

OR2x2_ASAP7_75t_L g2282 ( 
.A(n_2208),
.B(n_2186),
.Y(n_2282)
);

AND2x2_ASAP7_75t_L g2283 ( 
.A(n_2210),
.B(n_2174),
.Y(n_2283)
);

INVx2_ASAP7_75t_L g2284 ( 
.A(n_2204),
.Y(n_2284)
);

NAND2xp5_ASAP7_75t_L g2285 ( 
.A(n_2221),
.B(n_2190),
.Y(n_2285)
);

INVx2_ASAP7_75t_L g2286 ( 
.A(n_2204),
.Y(n_2286)
);

OR2x2_ASAP7_75t_L g2287 ( 
.A(n_2221),
.B(n_2188),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_2196),
.Y(n_2288)
);

AND2x2_ASAP7_75t_L g2289 ( 
.A(n_2210),
.B(n_2173),
.Y(n_2289)
);

INVx2_ASAP7_75t_L g2290 ( 
.A(n_2209),
.Y(n_2290)
);

INVx2_ASAP7_75t_SL g2291 ( 
.A(n_2236),
.Y(n_2291)
);

HB1xp67_ASAP7_75t_L g2292 ( 
.A(n_2248),
.Y(n_2292)
);

NAND2xp5_ASAP7_75t_L g2293 ( 
.A(n_2235),
.B(n_2211),
.Y(n_2293)
);

INVx1_ASAP7_75t_L g2294 ( 
.A(n_2196),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_2198),
.Y(n_2295)
);

OR2x2_ASAP7_75t_L g2296 ( 
.A(n_2206),
.B(n_2173),
.Y(n_2296)
);

INVx2_ASAP7_75t_SL g2297 ( 
.A(n_2236),
.Y(n_2297)
);

OR2x2_ASAP7_75t_L g2298 ( 
.A(n_2206),
.B(n_2173),
.Y(n_2298)
);

OR2x6_ASAP7_75t_L g2299 ( 
.A(n_2224),
.B(n_2041),
.Y(n_2299)
);

NAND2xp5_ASAP7_75t_L g2300 ( 
.A(n_2235),
.B(n_2185),
.Y(n_2300)
);

AND2x2_ASAP7_75t_L g2301 ( 
.A(n_2211),
.B(n_2173),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_2198),
.Y(n_2302)
);

AND2x2_ASAP7_75t_L g2303 ( 
.A(n_2211),
.B(n_2183),
.Y(n_2303)
);

INVxp67_ASAP7_75t_L g2304 ( 
.A(n_2253),
.Y(n_2304)
);

AND2x2_ASAP7_75t_L g2305 ( 
.A(n_2200),
.B(n_2183),
.Y(n_2305)
);

INVx2_ASAP7_75t_L g2306 ( 
.A(n_2209),
.Y(n_2306)
);

INVx2_ASAP7_75t_L g2307 ( 
.A(n_2212),
.Y(n_2307)
);

NAND2xp5_ASAP7_75t_L g2308 ( 
.A(n_2229),
.B(n_2185),
.Y(n_2308)
);

OR2x2_ASAP7_75t_L g2309 ( 
.A(n_2293),
.B(n_2248),
.Y(n_2309)
);

OR2x2_ASAP7_75t_L g2310 ( 
.A(n_2293),
.B(n_2251),
.Y(n_2310)
);

NAND2xp5_ASAP7_75t_L g2311 ( 
.A(n_2269),
.B(n_2241),
.Y(n_2311)
);

NAND2xp5_ASAP7_75t_L g2312 ( 
.A(n_2269),
.B(n_2241),
.Y(n_2312)
);

INVx2_ASAP7_75t_L g2313 ( 
.A(n_2268),
.Y(n_2313)
);

AND2x2_ASAP7_75t_L g2314 ( 
.A(n_2279),
.B(n_2200),
.Y(n_2314)
);

INVxp33_ASAP7_75t_SL g2315 ( 
.A(n_2270),
.Y(n_2315)
);

AO21x2_ASAP7_75t_L g2316 ( 
.A1(n_2256),
.A2(n_2249),
.B(n_2251),
.Y(n_2316)
);

OR2x2_ASAP7_75t_L g2317 ( 
.A(n_2261),
.B(n_2200),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_2273),
.Y(n_2318)
);

NAND2x1_ASAP7_75t_L g2319 ( 
.A(n_2281),
.B(n_2201),
.Y(n_2319)
);

BUFx3_ASAP7_75t_L g2320 ( 
.A(n_2270),
.Y(n_2320)
);

NAND2xp5_ASAP7_75t_L g2321 ( 
.A(n_2285),
.B(n_2219),
.Y(n_2321)
);

INVx1_ASAP7_75t_L g2322 ( 
.A(n_2273),
.Y(n_2322)
);

OR2x2_ASAP7_75t_L g2323 ( 
.A(n_2261),
.B(n_2249),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_2274),
.Y(n_2324)
);

AND2x4_ASAP7_75t_L g2325 ( 
.A(n_2291),
.B(n_2242),
.Y(n_2325)
);

INVx1_ASAP7_75t_L g2326 ( 
.A(n_2274),
.Y(n_2326)
);

NAND2xp5_ASAP7_75t_L g2327 ( 
.A(n_2285),
.B(n_2219),
.Y(n_2327)
);

INVx2_ASAP7_75t_L g2328 ( 
.A(n_2268),
.Y(n_2328)
);

OR2x2_ASAP7_75t_L g2329 ( 
.A(n_2290),
.B(n_2218),
.Y(n_2329)
);

NOR2xp33_ASAP7_75t_L g2330 ( 
.A(n_2260),
.B(n_2146),
.Y(n_2330)
);

INVx1_ASAP7_75t_L g2331 ( 
.A(n_2288),
.Y(n_2331)
);

NAND2xp5_ASAP7_75t_L g2332 ( 
.A(n_2262),
.B(n_2218),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_2288),
.Y(n_2333)
);

NOR3xp33_ASAP7_75t_L g2334 ( 
.A(n_2256),
.B(n_2133),
.C(n_2165),
.Y(n_2334)
);

NOR4xp25_ASAP7_75t_SL g2335 ( 
.A(n_2258),
.B(n_2226),
.C(n_2157),
.D(n_2182),
.Y(n_2335)
);

AND2x2_ASAP7_75t_L g2336 ( 
.A(n_2257),
.B(n_2242),
.Y(n_2336)
);

NAND2xp5_ASAP7_75t_L g2337 ( 
.A(n_2262),
.B(n_2220),
.Y(n_2337)
);

INVx1_ASAP7_75t_L g2338 ( 
.A(n_2294),
.Y(n_2338)
);

NAND2xp5_ASAP7_75t_L g2339 ( 
.A(n_2260),
.B(n_2217),
.Y(n_2339)
);

BUFx2_ASAP7_75t_L g2340 ( 
.A(n_2292),
.Y(n_2340)
);

AND2x2_ASAP7_75t_L g2341 ( 
.A(n_2257),
.B(n_2242),
.Y(n_2341)
);

NAND2xp5_ASAP7_75t_L g2342 ( 
.A(n_2278),
.B(n_2217),
.Y(n_2342)
);

BUFx3_ASAP7_75t_L g2343 ( 
.A(n_2266),
.Y(n_2343)
);

INVx2_ASAP7_75t_L g2344 ( 
.A(n_2268),
.Y(n_2344)
);

NAND2xp5_ASAP7_75t_L g2345 ( 
.A(n_2304),
.B(n_2227),
.Y(n_2345)
);

INVx1_ASAP7_75t_L g2346 ( 
.A(n_2294),
.Y(n_2346)
);

INVxp67_ASAP7_75t_SL g2347 ( 
.A(n_2267),
.Y(n_2347)
);

INVxp67_ASAP7_75t_L g2348 ( 
.A(n_2265),
.Y(n_2348)
);

NOR2xp33_ASAP7_75t_L g2349 ( 
.A(n_2287),
.B(n_2146),
.Y(n_2349)
);

HB1xp67_ASAP7_75t_L g2350 ( 
.A(n_2258),
.Y(n_2350)
);

NOR2x1_ASAP7_75t_L g2351 ( 
.A(n_2287),
.B(n_2245),
.Y(n_2351)
);

INVx2_ASAP7_75t_L g2352 ( 
.A(n_2275),
.Y(n_2352)
);

HB1xp67_ASAP7_75t_L g2353 ( 
.A(n_2259),
.Y(n_2353)
);

INVx4_ASAP7_75t_L g2354 ( 
.A(n_2281),
.Y(n_2354)
);

AND2x4_ASAP7_75t_L g2355 ( 
.A(n_2291),
.B(n_2215),
.Y(n_2355)
);

INVx1_ASAP7_75t_L g2356 ( 
.A(n_2295),
.Y(n_2356)
);

OR2x2_ASAP7_75t_L g2357 ( 
.A(n_2290),
.B(n_2227),
.Y(n_2357)
);

AND2x2_ASAP7_75t_L g2358 ( 
.A(n_2280),
.B(n_2222),
.Y(n_2358)
);

INVx2_ASAP7_75t_L g2359 ( 
.A(n_2275),
.Y(n_2359)
);

INVx1_ASAP7_75t_L g2360 ( 
.A(n_2350),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_2353),
.Y(n_2361)
);

AND2x2_ASAP7_75t_L g2362 ( 
.A(n_2314),
.B(n_2291),
.Y(n_2362)
);

OAI21xp5_ASAP7_75t_SL g2363 ( 
.A1(n_2351),
.A2(n_2277),
.B(n_2255),
.Y(n_2363)
);

AOI221xp5_ASAP7_75t_L g2364 ( 
.A1(n_2334),
.A2(n_2255),
.B1(n_2271),
.B2(n_2277),
.C(n_2265),
.Y(n_2364)
);

NAND2xp5_ASAP7_75t_L g2365 ( 
.A(n_2320),
.B(n_2271),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_2318),
.Y(n_2366)
);

INVx2_ASAP7_75t_L g2367 ( 
.A(n_2320),
.Y(n_2367)
);

AOI31xp33_ASAP7_75t_L g2368 ( 
.A1(n_2351),
.A2(n_2349),
.A3(n_2348),
.B(n_2337),
.Y(n_2368)
);

NAND2xp5_ASAP7_75t_L g2369 ( 
.A(n_2320),
.B(n_2272),
.Y(n_2369)
);

NAND2xp5_ASAP7_75t_L g2370 ( 
.A(n_2340),
.B(n_2272),
.Y(n_2370)
);

AOI22xp5_ASAP7_75t_L g2371 ( 
.A1(n_2316),
.A2(n_2263),
.B1(n_2330),
.B2(n_2155),
.Y(n_2371)
);

INVx1_ASAP7_75t_L g2372 ( 
.A(n_2318),
.Y(n_2372)
);

INVxp67_ASAP7_75t_SL g2373 ( 
.A(n_2315),
.Y(n_2373)
);

OAI22xp5_ASAP7_75t_L g2374 ( 
.A1(n_2343),
.A2(n_2266),
.B1(n_2263),
.B2(n_2282),
.Y(n_2374)
);

NAND2xp5_ASAP7_75t_L g2375 ( 
.A(n_2340),
.B(n_2290),
.Y(n_2375)
);

NAND2xp5_ASAP7_75t_L g2376 ( 
.A(n_2332),
.B(n_2306),
.Y(n_2376)
);

INVx1_ASAP7_75t_L g2377 ( 
.A(n_2322),
.Y(n_2377)
);

INVx1_ASAP7_75t_L g2378 ( 
.A(n_2322),
.Y(n_2378)
);

AOI21xp5_ASAP7_75t_L g2379 ( 
.A1(n_2316),
.A2(n_2282),
.B(n_2250),
.Y(n_2379)
);

OAI322xp33_ASAP7_75t_L g2380 ( 
.A1(n_2309),
.A2(n_2275),
.A3(n_2276),
.B1(n_2284),
.B2(n_2286),
.C1(n_2306),
.C2(n_2250),
.Y(n_2380)
);

AOI22xp33_ASAP7_75t_L g2381 ( 
.A1(n_2316),
.A2(n_2276),
.B1(n_2143),
.B2(n_2230),
.Y(n_2381)
);

AND2x2_ASAP7_75t_L g2382 ( 
.A(n_2314),
.B(n_2297),
.Y(n_2382)
);

INVx1_ASAP7_75t_SL g2383 ( 
.A(n_2343),
.Y(n_2383)
);

OAI22xp5_ASAP7_75t_L g2384 ( 
.A1(n_2323),
.A2(n_2276),
.B1(n_2297),
.B2(n_2280),
.Y(n_2384)
);

AOI22xp33_ASAP7_75t_SL g2385 ( 
.A1(n_2311),
.A2(n_2286),
.B1(n_2284),
.B2(n_2245),
.Y(n_2385)
);

INVx1_ASAP7_75t_L g2386 ( 
.A(n_2324),
.Y(n_2386)
);

OAI21xp5_ASAP7_75t_L g2387 ( 
.A1(n_2312),
.A2(n_2259),
.B(n_2264),
.Y(n_2387)
);

AOI21xp5_ASAP7_75t_L g2388 ( 
.A1(n_2319),
.A2(n_2281),
.B(n_2300),
.Y(n_2388)
);

NAND4xp25_ASAP7_75t_L g2389 ( 
.A(n_2354),
.B(n_2264),
.C(n_2306),
.D(n_2281),
.Y(n_2389)
);

OAI32xp33_ASAP7_75t_L g2390 ( 
.A1(n_2323),
.A2(n_2284),
.A3(n_2286),
.B1(n_2296),
.B2(n_2298),
.Y(n_2390)
);

AOI22xp5_ASAP7_75t_L g2391 ( 
.A1(n_2339),
.A2(n_2131),
.B1(n_2139),
.B2(n_2254),
.Y(n_2391)
);

NAND2xp5_ASAP7_75t_L g2392 ( 
.A(n_2321),
.B(n_2295),
.Y(n_2392)
);

NAND2xp5_ASAP7_75t_L g2393 ( 
.A(n_2327),
.B(n_2302),
.Y(n_2393)
);

NOR2xp33_ASAP7_75t_L g2394 ( 
.A(n_2354),
.B(n_2297),
.Y(n_2394)
);

INVx1_ASAP7_75t_L g2395 ( 
.A(n_2324),
.Y(n_2395)
);

AOI32xp33_ASAP7_75t_L g2396 ( 
.A1(n_2355),
.A2(n_2289),
.A3(n_2245),
.B1(n_2131),
.B2(n_2283),
.Y(n_2396)
);

OAI322xp33_ASAP7_75t_L g2397 ( 
.A1(n_2309),
.A2(n_2254),
.A3(n_2296),
.B1(n_2298),
.B2(n_2302),
.C1(n_2300),
.C2(n_2237),
.Y(n_2397)
);

NAND2xp5_ASAP7_75t_L g2398 ( 
.A(n_2347),
.B(n_2283),
.Y(n_2398)
);

INVx1_ASAP7_75t_L g2399 ( 
.A(n_2326),
.Y(n_2399)
);

AOI22xp5_ASAP7_75t_L g2400 ( 
.A1(n_2355),
.A2(n_2176),
.B1(n_2289),
.B2(n_2299),
.Y(n_2400)
);

NAND2xp5_ASAP7_75t_SL g2401 ( 
.A(n_2368),
.B(n_2355),
.Y(n_2401)
);

NOR4xp25_ASAP7_75t_SL g2402 ( 
.A(n_2363),
.B(n_2326),
.C(n_2333),
.D(n_2338),
.Y(n_2402)
);

INVx1_ASAP7_75t_L g2403 ( 
.A(n_2366),
.Y(n_2403)
);

OAI22xp5_ASAP7_75t_L g2404 ( 
.A1(n_2381),
.A2(n_2319),
.B1(n_2317),
.B2(n_2335),
.Y(n_2404)
);

INVx1_ASAP7_75t_L g2405 ( 
.A(n_2372),
.Y(n_2405)
);

NAND2xp5_ASAP7_75t_L g2406 ( 
.A(n_2373),
.B(n_2310),
.Y(n_2406)
);

INVx1_ASAP7_75t_SL g2407 ( 
.A(n_2383),
.Y(n_2407)
);

AOI21xp33_ASAP7_75t_L g2408 ( 
.A1(n_2364),
.A2(n_2310),
.B(n_2357),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_2377),
.Y(n_2409)
);

INVxp67_ASAP7_75t_L g2410 ( 
.A(n_2373),
.Y(n_2410)
);

OAI32xp33_ASAP7_75t_L g2411 ( 
.A1(n_2374),
.A2(n_2365),
.A3(n_2389),
.B1(n_2369),
.B2(n_2381),
.Y(n_2411)
);

NAND2xp5_ASAP7_75t_L g2412 ( 
.A(n_2367),
.B(n_2342),
.Y(n_2412)
);

OR2x2_ASAP7_75t_L g2413 ( 
.A(n_2376),
.B(n_2317),
.Y(n_2413)
);

OR2x2_ASAP7_75t_L g2414 ( 
.A(n_2392),
.B(n_2345),
.Y(n_2414)
);

NAND2xp5_ASAP7_75t_L g2415 ( 
.A(n_2367),
.B(n_2329),
.Y(n_2415)
);

NAND3xp33_ASAP7_75t_L g2416 ( 
.A(n_2379),
.B(n_2354),
.C(n_2331),
.Y(n_2416)
);

NAND2xp5_ASAP7_75t_L g2417 ( 
.A(n_2371),
.B(n_2329),
.Y(n_2417)
);

INVxp67_ASAP7_75t_L g2418 ( 
.A(n_2375),
.Y(n_2418)
);

AOI222xp33_ASAP7_75t_L g2419 ( 
.A1(n_2387),
.A2(n_2359),
.B1(n_2328),
.B2(n_2313),
.C1(n_2344),
.C2(n_2352),
.Y(n_2419)
);

INVx1_ASAP7_75t_SL g2420 ( 
.A(n_2362),
.Y(n_2420)
);

NAND2xp5_ASAP7_75t_L g2421 ( 
.A(n_2360),
.B(n_2361),
.Y(n_2421)
);

OAI211xp5_ASAP7_75t_SL g2422 ( 
.A1(n_2396),
.A2(n_2346),
.B(n_2333),
.C(n_2338),
.Y(n_2422)
);

INVxp67_ASAP7_75t_L g2423 ( 
.A(n_2394),
.Y(n_2423)
);

INVx1_ASAP7_75t_L g2424 ( 
.A(n_2378),
.Y(n_2424)
);

OAI21xp33_ASAP7_75t_L g2425 ( 
.A1(n_2400),
.A2(n_2325),
.B(n_2356),
.Y(n_2425)
);

INVx1_ASAP7_75t_L g2426 ( 
.A(n_2386),
.Y(n_2426)
);

HB1xp67_ASAP7_75t_L g2427 ( 
.A(n_2398),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_2395),
.Y(n_2428)
);

AND2x2_ASAP7_75t_L g2429 ( 
.A(n_2362),
.B(n_2336),
.Y(n_2429)
);

OAI221xp5_ASAP7_75t_L g2430 ( 
.A1(n_2385),
.A2(n_2359),
.B1(n_2344),
.B2(n_2313),
.C(n_2352),
.Y(n_2430)
);

OAI221xp5_ASAP7_75t_SL g2431 ( 
.A1(n_2391),
.A2(n_2388),
.B1(n_2370),
.B2(n_2382),
.C(n_2393),
.Y(n_2431)
);

NAND5xp2_ASAP7_75t_L g2432 ( 
.A(n_2431),
.B(n_2394),
.C(n_2382),
.D(n_2399),
.E(n_2341),
.Y(n_2432)
);

INVx1_ASAP7_75t_L g2433 ( 
.A(n_2410),
.Y(n_2433)
);

INVx1_ASAP7_75t_L g2434 ( 
.A(n_2415),
.Y(n_2434)
);

HB1xp67_ASAP7_75t_L g2435 ( 
.A(n_2407),
.Y(n_2435)
);

NAND2xp5_ASAP7_75t_L g2436 ( 
.A(n_2420),
.B(n_2384),
.Y(n_2436)
);

NOR2x1_ASAP7_75t_L g2437 ( 
.A(n_2416),
.B(n_2401),
.Y(n_2437)
);

NAND2xp5_ASAP7_75t_SL g2438 ( 
.A(n_2401),
.B(n_2404),
.Y(n_2438)
);

INVx1_ASAP7_75t_L g2439 ( 
.A(n_2426),
.Y(n_2439)
);

NAND2xp5_ASAP7_75t_L g2440 ( 
.A(n_2427),
.B(n_2358),
.Y(n_2440)
);

CKINVDCx5p33_ASAP7_75t_R g2441 ( 
.A(n_2406),
.Y(n_2441)
);

INVx1_ASAP7_75t_L g2442 ( 
.A(n_2426),
.Y(n_2442)
);

OAI22xp5_ASAP7_75t_L g2443 ( 
.A1(n_2402),
.A2(n_2355),
.B1(n_2335),
.B2(n_2354),
.Y(n_2443)
);

INVx1_ASAP7_75t_L g2444 ( 
.A(n_2403),
.Y(n_2444)
);

AND2x4_ASAP7_75t_L g2445 ( 
.A(n_2429),
.B(n_2325),
.Y(n_2445)
);

AND2x2_ASAP7_75t_L g2446 ( 
.A(n_2429),
.B(n_2336),
.Y(n_2446)
);

INVx1_ASAP7_75t_L g2447 ( 
.A(n_2405),
.Y(n_2447)
);

INVx1_ASAP7_75t_L g2448 ( 
.A(n_2409),
.Y(n_2448)
);

INVx1_ASAP7_75t_L g2449 ( 
.A(n_2424),
.Y(n_2449)
);

OAI22x1_ASAP7_75t_L g2450 ( 
.A1(n_2417),
.A2(n_2325),
.B1(n_2331),
.B2(n_2356),
.Y(n_2450)
);

NAND3xp33_ASAP7_75t_SL g2451 ( 
.A(n_2419),
.B(n_2328),
.C(n_2380),
.Y(n_2451)
);

INVxp67_ASAP7_75t_L g2452 ( 
.A(n_2421),
.Y(n_2452)
);

INVx1_ASAP7_75t_L g2453 ( 
.A(n_2428),
.Y(n_2453)
);

NOR4xp25_ASAP7_75t_SL g2454 ( 
.A(n_2422),
.B(n_2390),
.C(n_2346),
.D(n_2397),
.Y(n_2454)
);

HB1xp67_ASAP7_75t_L g2455 ( 
.A(n_2423),
.Y(n_2455)
);

INVx1_ASAP7_75t_L g2456 ( 
.A(n_2413),
.Y(n_2456)
);

NAND2xp5_ASAP7_75t_L g2457 ( 
.A(n_2435),
.B(n_2418),
.Y(n_2457)
);

NOR2xp33_ASAP7_75t_L g2458 ( 
.A(n_2441),
.B(n_2452),
.Y(n_2458)
);

NAND4xp25_ASAP7_75t_L g2459 ( 
.A(n_2432),
.B(n_2411),
.C(n_2425),
.D(n_2412),
.Y(n_2459)
);

INVx1_ASAP7_75t_L g2460 ( 
.A(n_2455),
.Y(n_2460)
);

NOR2xp33_ASAP7_75t_L g2461 ( 
.A(n_2441),
.B(n_2411),
.Y(n_2461)
);

INVx1_ASAP7_75t_L g2462 ( 
.A(n_2456),
.Y(n_2462)
);

INVx1_ASAP7_75t_L g2463 ( 
.A(n_2456),
.Y(n_2463)
);

NAND4xp25_ASAP7_75t_L g2464 ( 
.A(n_2437),
.B(n_2408),
.C(n_2413),
.D(n_2414),
.Y(n_2464)
);

INVx2_ASAP7_75t_L g2465 ( 
.A(n_2445),
.Y(n_2465)
);

OAI22xp33_ASAP7_75t_L g2466 ( 
.A1(n_2454),
.A2(n_2451),
.B1(n_2450),
.B2(n_2438),
.Y(n_2466)
);

INVx1_ASAP7_75t_L g2467 ( 
.A(n_2439),
.Y(n_2467)
);

INVx1_ASAP7_75t_L g2468 ( 
.A(n_2442),
.Y(n_2468)
);

INVx2_ASAP7_75t_L g2469 ( 
.A(n_2445),
.Y(n_2469)
);

NAND2xp5_ASAP7_75t_L g2470 ( 
.A(n_2446),
.B(n_2414),
.Y(n_2470)
);

NOR2xp33_ASAP7_75t_L g2471 ( 
.A(n_2438),
.B(n_2430),
.Y(n_2471)
);

AOI322xp5_ASAP7_75t_L g2472 ( 
.A1(n_2466),
.A2(n_2434),
.A3(n_2433),
.B1(n_2447),
.B2(n_2436),
.C1(n_2448),
.C2(n_2449),
.Y(n_2472)
);

AOI211xp5_ASAP7_75t_L g2473 ( 
.A1(n_2466),
.A2(n_2443),
.B(n_2447),
.C(n_2453),
.Y(n_2473)
);

INVx1_ASAP7_75t_L g2474 ( 
.A(n_2470),
.Y(n_2474)
);

NAND2xp5_ASAP7_75t_SL g2475 ( 
.A(n_2461),
.B(n_2445),
.Y(n_2475)
);

NAND2xp5_ASAP7_75t_L g2476 ( 
.A(n_2471),
.B(n_2446),
.Y(n_2476)
);

NAND3xp33_ASAP7_75t_L g2477 ( 
.A(n_2471),
.B(n_2444),
.C(n_2440),
.Y(n_2477)
);

INVx1_ASAP7_75t_L g2478 ( 
.A(n_2457),
.Y(n_2478)
);

NOR2x1_ASAP7_75t_L g2479 ( 
.A(n_2458),
.B(n_2450),
.Y(n_2479)
);

NOR2xp33_ASAP7_75t_L g2480 ( 
.A(n_2464),
.B(n_2325),
.Y(n_2480)
);

AOI221xp5_ASAP7_75t_L g2481 ( 
.A1(n_2459),
.A2(n_2148),
.B1(n_2308),
.B2(n_2357),
.C(n_2307),
.Y(n_2481)
);

OR2x2_ASAP7_75t_L g2482 ( 
.A(n_2460),
.B(n_2465),
.Y(n_2482)
);

CKINVDCx5p33_ASAP7_75t_R g2483 ( 
.A(n_2478),
.Y(n_2483)
);

INVx1_ASAP7_75t_L g2484 ( 
.A(n_2482),
.Y(n_2484)
);

AOI221x1_ASAP7_75t_L g2485 ( 
.A1(n_2474),
.A2(n_2463),
.B1(n_2462),
.B2(n_2467),
.C(n_2468),
.Y(n_2485)
);

INVx1_ASAP7_75t_L g2486 ( 
.A(n_2476),
.Y(n_2486)
);

AOI221xp5_ASAP7_75t_L g2487 ( 
.A1(n_2473),
.A2(n_2469),
.B1(n_2308),
.B2(n_2307),
.C(n_2341),
.Y(n_2487)
);

NAND3xp33_ASAP7_75t_SL g2488 ( 
.A(n_2472),
.B(n_2358),
.C(n_2301),
.Y(n_2488)
);

NAND2xp5_ASAP7_75t_L g2489 ( 
.A(n_2479),
.B(n_2301),
.Y(n_2489)
);

NOR3x2_ASAP7_75t_L g2490 ( 
.A(n_2483),
.B(n_2475),
.C(n_2477),
.Y(n_2490)
);

NAND2x1p5_ASAP7_75t_L g2491 ( 
.A(n_2484),
.B(n_2486),
.Y(n_2491)
);

CKINVDCx20_ASAP7_75t_R g2492 ( 
.A(n_2489),
.Y(n_2492)
);

BUFx2_ASAP7_75t_L g2493 ( 
.A(n_2487),
.Y(n_2493)
);

HB1xp67_ASAP7_75t_L g2494 ( 
.A(n_2485),
.Y(n_2494)
);

NOR2xp33_ASAP7_75t_L g2495 ( 
.A(n_2488),
.B(n_2480),
.Y(n_2495)
);

NAND2xp5_ASAP7_75t_L g2496 ( 
.A(n_2484),
.B(n_2481),
.Y(n_2496)
);

OAI211xp5_ASAP7_75t_L g2497 ( 
.A1(n_2485),
.A2(n_2234),
.B(n_2233),
.C(n_2225),
.Y(n_2497)
);

NOR4xp25_ASAP7_75t_L g2498 ( 
.A(n_2496),
.B(n_2303),
.C(n_2307),
.D(n_2238),
.Y(n_2498)
);

NAND4xp25_ASAP7_75t_L g2499 ( 
.A(n_2495),
.B(n_2007),
.C(n_2303),
.D(n_2305),
.Y(n_2499)
);

A2O1A1Ixp33_ASAP7_75t_L g2500 ( 
.A1(n_2494),
.A2(n_2237),
.B(n_2228),
.C(n_2305),
.Y(n_2500)
);

NAND4xp25_ASAP7_75t_L g2501 ( 
.A(n_2493),
.B(n_2234),
.C(n_2233),
.D(n_2216),
.Y(n_2501)
);

AO22x2_ASAP7_75t_L g2502 ( 
.A1(n_2497),
.A2(n_2228),
.B1(n_2240),
.B2(n_2231),
.Y(n_2502)
);

NAND5xp2_ASAP7_75t_L g2503 ( 
.A(n_2491),
.B(n_2213),
.C(n_2247),
.D(n_2243),
.E(n_2222),
.Y(n_2503)
);

OAI221xp5_ASAP7_75t_L g2504 ( 
.A1(n_2491),
.A2(n_2299),
.B1(n_2041),
.B2(n_2126),
.C(n_2046),
.Y(n_2504)
);

HB1xp67_ASAP7_75t_L g2505 ( 
.A(n_2500),
.Y(n_2505)
);

INVx1_ASAP7_75t_L g2506 ( 
.A(n_2502),
.Y(n_2506)
);

AOI221xp5_ASAP7_75t_L g2507 ( 
.A1(n_2498),
.A2(n_2492),
.B1(n_2490),
.B2(n_2231),
.C(n_2240),
.Y(n_2507)
);

NOR2x2_ASAP7_75t_L g2508 ( 
.A(n_2499),
.B(n_2299),
.Y(n_2508)
);

XNOR2xp5_ASAP7_75t_L g2509 ( 
.A(n_2505),
.B(n_2501),
.Y(n_2509)
);

INVx2_ASAP7_75t_L g2510 ( 
.A(n_2508),
.Y(n_2510)
);

NAND2x1_ASAP7_75t_L g2511 ( 
.A(n_2510),
.B(n_2506),
.Y(n_2511)
);

AOI22xp5_ASAP7_75t_L g2512 ( 
.A1(n_2509),
.A2(n_2507),
.B1(n_2504),
.B2(n_2503),
.Y(n_2512)
);

XNOR2xp5_ASAP7_75t_L g2513 ( 
.A(n_2512),
.B(n_2299),
.Y(n_2513)
);

HB1xp67_ASAP7_75t_L g2514 ( 
.A(n_2511),
.Y(n_2514)
);

AND2x2_ASAP7_75t_L g2515 ( 
.A(n_2512),
.B(n_2222),
.Y(n_2515)
);

AOI21xp33_ASAP7_75t_L g2516 ( 
.A1(n_2514),
.A2(n_2299),
.B(n_2252),
.Y(n_2516)
);

AOI22xp33_ASAP7_75t_L g2517 ( 
.A1(n_2513),
.A2(n_2515),
.B1(n_2244),
.B2(n_2202),
.Y(n_2517)
);

OAI21xp5_ASAP7_75t_L g2518 ( 
.A1(n_2517),
.A2(n_2238),
.B(n_2213),
.Y(n_2518)
);

AOI22xp33_ASAP7_75t_R g2519 ( 
.A1(n_2516),
.A2(n_2244),
.B1(n_2202),
.B2(n_2205),
.Y(n_2519)
);

AOI322xp5_ASAP7_75t_L g2520 ( 
.A1(n_2519),
.A2(n_2213),
.A3(n_2238),
.B1(n_2109),
.B2(n_2118),
.C1(n_2232),
.C2(n_2207),
.Y(n_2520)
);

OAI221xp5_ASAP7_75t_R g2521 ( 
.A1(n_2520),
.A2(n_2518),
.B1(n_2182),
.B2(n_2232),
.C(n_2046),
.Y(n_2521)
);

AOI211xp5_ASAP7_75t_L g2522 ( 
.A1(n_2521),
.A2(n_2232),
.B(n_2246),
.C(n_2047),
.Y(n_2522)
);


endmodule