module fake_jpeg_8587_n_331 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_331);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_331;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_38),
.Y(n_53)
);

NAND2x1_ASAP7_75t_L g37 ( 
.A(n_32),
.B(n_0),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_37),
.A2(n_25),
.B1(n_24),
.B2(n_19),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_33),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_39),
.B(n_41),
.Y(n_66)
);

BUFx10_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_25),
.Y(n_43)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_46),
.B(n_48),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_47),
.A2(n_59),
.B(n_24),
.Y(n_95)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_37),
.A2(n_28),
.B1(n_33),
.B2(n_26),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_50),
.A2(n_48),
.B1(n_32),
.B2(n_55),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_42),
.A2(n_28),
.B1(n_26),
.B2(n_19),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_51),
.A2(n_57),
.B1(n_20),
.B2(n_27),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_55),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_39),
.A2(n_28),
.B1(n_34),
.B2(n_20),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_58),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_42),
.A2(n_28),
.B1(n_27),
.B2(n_19),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_63),
.B(n_65),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_67),
.B(n_68),
.Y(n_92)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_70),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_71),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_38),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_72),
.B(n_87),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_46),
.B(n_36),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_73),
.B(n_79),
.Y(n_105)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_74),
.B(n_76),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_75),
.A2(n_88),
.B1(n_95),
.B2(n_77),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_66),
.Y(n_76)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_78),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_50),
.B(n_32),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_52),
.A2(n_32),
.B1(n_34),
.B2(n_21),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_84),
.A2(n_25),
.B1(n_24),
.B2(n_21),
.Y(n_98)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_53),
.Y(n_86)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_86),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_62),
.B(n_20),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_89),
.Y(n_118)
);

NAND3xp33_ASAP7_75t_SL g90 ( 
.A(n_65),
.B(n_32),
.C(n_40),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_18),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_54),
.B(n_27),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_90),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_95),
.A2(n_23),
.B(n_21),
.Y(n_103)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_96),
.B(n_101),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_98),
.A2(n_100),
.B1(n_111),
.B2(n_83),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_72),
.A2(n_49),
.B1(n_56),
.B2(n_63),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_93),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_76),
.A2(n_49),
.B1(n_56),
.B2(n_58),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_102),
.A2(n_104),
.B1(n_109),
.B2(n_112),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_103),
.A2(n_17),
.B(n_22),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_92),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_107),
.B(n_108),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_87),
.B(n_23),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_80),
.A2(n_23),
.B1(n_18),
.B2(n_31),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_74),
.A2(n_69),
.B1(n_14),
.B2(n_9),
.Y(n_112)
);

NAND2xp67_ASAP7_75t_SL g151 ( 
.A(n_113),
.B(n_40),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_77),
.B(n_13),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_114),
.B(n_120),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_73),
.B(n_0),
.Y(n_115)
);

AOI21xp33_ASAP7_75t_L g133 ( 
.A1(n_115),
.A2(n_93),
.B(n_79),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_116),
.A2(n_121),
.B1(n_78),
.B2(n_81),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_80),
.B(n_40),
.C(n_70),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_117),
.B(n_91),
.C(n_71),
.Y(n_146)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_85),
.Y(n_119)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_119),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_73),
.B(n_18),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_88),
.A2(n_64),
.B1(n_61),
.B2(n_18),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_85),
.Y(n_122)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_122),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_123),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_125),
.B(n_127),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_100),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_110),
.Y(n_129)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_129),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_99),
.B(n_75),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_131),
.B(n_137),
.Y(n_155)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_121),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_132),
.B(n_134),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_133),
.A2(n_149),
.B(n_151),
.Y(n_166)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_111),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_117),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_135),
.B(n_139),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_136),
.A2(n_140),
.B1(n_97),
.B2(n_71),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_99),
.B(n_79),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_98),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_138),
.B(n_142),
.Y(n_158)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_104),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_101),
.A2(n_81),
.B1(n_83),
.B2(n_86),
.Y(n_140)
);

A2O1A1Ixp33_ASAP7_75t_L g141 ( 
.A1(n_120),
.A2(n_84),
.B(n_40),
.C(n_17),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_141),
.B(n_147),
.Y(n_168)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_110),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_107),
.B(n_91),
.Y(n_143)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_143),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_144),
.A2(n_122),
.B(n_114),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_146),
.B(n_105),
.C(n_113),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_119),
.B(n_91),
.Y(n_148)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_148),
.Y(n_169)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_109),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_132),
.A2(n_103),
.B1(n_113),
.B2(n_105),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_153),
.A2(n_162),
.B1(n_130),
.B2(n_126),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_154),
.B(n_124),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_156),
.B(n_157),
.C(n_29),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_137),
.B(n_105),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_143),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_159),
.B(n_163),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_151),
.A2(n_115),
.B(n_118),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_160),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_127),
.A2(n_115),
.B1(n_118),
.B2(n_106),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_148),
.Y(n_163)
);

XNOR2x1_ASAP7_75t_L g165 ( 
.A(n_133),
.B(n_108),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_165),
.B(n_176),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_134),
.A2(n_96),
.B1(n_97),
.B2(n_106),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_167),
.A2(n_171),
.B1(n_141),
.B2(n_149),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_140),
.Y(n_172)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_172),
.Y(n_182)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_129),
.Y(n_174)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_174),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_128),
.Y(n_175)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_175),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_128),
.A2(n_17),
.B(n_22),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_145),
.Y(n_177)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_177),
.Y(n_199)
);

OA21x2_ASAP7_75t_SL g178 ( 
.A1(n_131),
.A2(n_40),
.B(n_22),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_178),
.B(n_179),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_139),
.A2(n_110),
.B(n_82),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_144),
.A2(n_17),
.B(n_22),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_180),
.B(n_31),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_183),
.B(n_200),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_158),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_184),
.B(n_189),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_166),
.B(n_146),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_185),
.B(n_193),
.C(n_197),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_172),
.A2(n_138),
.B1(n_147),
.B2(n_136),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_187),
.A2(n_171),
.B1(n_164),
.B2(n_170),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_188),
.A2(n_192),
.B1(n_201),
.B2(n_162),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_167),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_152),
.A2(n_141),
.B1(n_150),
.B2(n_124),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_166),
.B(n_145),
.Y(n_193)
);

OA22x2_ASAP7_75t_L g194 ( 
.A1(n_178),
.A2(n_142),
.B1(n_130),
.B2(n_126),
.Y(n_194)
);

OAI22x1_ASAP7_75t_L g227 ( 
.A1(n_194),
.A2(n_154),
.B1(n_29),
.B2(n_94),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_195),
.A2(n_155),
.B(n_94),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_156),
.B(n_125),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_152),
.A2(n_142),
.B1(n_31),
.B2(n_29),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_179),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_202),
.B(n_204),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_157),
.B(n_129),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_203),
.B(n_205),
.C(n_176),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_170),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_168),
.A2(n_94),
.B1(n_31),
.B2(n_29),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_206),
.A2(n_173),
.B1(n_169),
.B2(n_180),
.Y(n_225)
);

OR2x2_ASAP7_75t_L g207 ( 
.A(n_159),
.B(n_10),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_207),
.B(n_13),
.Y(n_226)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_186),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_L g239 ( 
.A1(n_209),
.A2(n_213),
.B1(n_215),
.B2(n_217),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_193),
.B(n_165),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_211),
.B(n_212),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_185),
.B(n_153),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_181),
.A2(n_168),
.B(n_164),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_184),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_216),
.Y(n_237)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_194),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_196),
.B(n_160),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_219),
.B(n_222),
.C(n_232),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_182),
.A2(n_177),
.B1(n_163),
.B2(n_161),
.Y(n_220)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_220),
.Y(n_249)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_191),
.Y(n_221)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_221),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_181),
.A2(n_161),
.B(n_169),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_223),
.A2(n_224),
.B1(n_228),
.B2(n_206),
.Y(n_236)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_225),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_226),
.B(n_229),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_SL g244 ( 
.A(n_227),
.B(n_194),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_195),
.A2(n_155),
.B1(n_173),
.B2(n_174),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_207),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_190),
.Y(n_230)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_230),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_231),
.B(n_200),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_196),
.B(n_7),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_203),
.B(n_1),
.C(n_2),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_233),
.B(n_205),
.C(n_198),
.Y(n_240)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_236),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_215),
.B(n_199),
.Y(n_238)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_238),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_240),
.B(n_243),
.C(n_9),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_214),
.B(n_194),
.Y(n_241)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_241),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_210),
.B(n_197),
.C(n_183),
.Y(n_243)
);

OAI321xp33_ASAP7_75t_L g259 ( 
.A1(n_244),
.A2(n_227),
.A3(n_219),
.B1(n_208),
.B2(n_211),
.C(n_233),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_218),
.B(n_221),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_247),
.Y(n_261)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_223),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_248),
.B(n_251),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_250),
.B(n_255),
.Y(n_271)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_225),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_213),
.B(n_198),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g274 ( 
.A(n_253),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_210),
.B(n_208),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_254),
.B(n_9),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_232),
.B(n_7),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_224),
.B(n_7),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_256),
.A2(n_239),
.B1(n_246),
.B2(n_251),
.Y(n_257)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_257),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_259),
.B(n_265),
.Y(n_280)
);

NOR3xp33_ASAP7_75t_SL g263 ( 
.A(n_244),
.B(n_212),
.C(n_222),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_263),
.B(n_264),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_248),
.A2(n_1),
.B(n_2),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_266),
.B(n_267),
.C(n_269),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_243),
.B(n_1),
.C(n_2),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_254),
.B(n_11),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_237),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_270)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_270),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_246),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_272)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_272),
.Y(n_283)
);

AOI321xp33_ASAP7_75t_L g273 ( 
.A1(n_242),
.A2(n_253),
.A3(n_249),
.B1(n_241),
.B2(n_234),
.C(n_240),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_273),
.B(n_235),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_261),
.B(n_238),
.Y(n_276)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_276),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_265),
.B(n_242),
.C(n_234),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_278),
.B(n_266),
.C(n_267),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_260),
.B(n_247),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_279),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_268),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_281),
.B(n_284),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_262),
.B(n_252),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_268),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_285),
.B(n_272),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_274),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_286),
.B(n_288),
.Y(n_292)
);

MAJx2_ASAP7_75t_L g295 ( 
.A(n_287),
.B(n_263),
.C(n_273),
.Y(n_295)
);

INVxp67_ASAP7_75t_SL g288 ( 
.A(n_270),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_282),
.A2(n_258),
.B1(n_277),
.B2(n_283),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_290),
.B(n_299),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_294),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_295),
.B(n_11),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_296),
.B(n_298),
.C(n_300),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_289),
.A2(n_235),
.B1(n_245),
.B2(n_271),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_297),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_287),
.B(n_269),
.C(n_264),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_280),
.B(n_245),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_276),
.A2(n_279),
.B1(n_280),
.B2(n_275),
.Y(n_300)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_275),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_302),
.B(n_12),
.Y(n_306)
);

AO21x1_ASAP7_75t_L g305 ( 
.A1(n_301),
.A2(n_278),
.B(n_12),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_305),
.B(n_307),
.Y(n_313)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_306),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_302),
.B(n_300),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_296),
.B(n_298),
.C(n_293),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_310),
.B(n_11),
.C(n_14),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_292),
.B(n_12),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_311),
.A2(n_299),
.B(n_291),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_312),
.B(n_304),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_314),
.B(n_315),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_305),
.A2(n_295),
.B(n_14),
.Y(n_316)
);

NOR3xp33_ASAP7_75t_L g323 ( 
.A(n_316),
.B(n_313),
.C(n_320),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_317),
.B(n_4),
.C(n_5),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_309),
.B(n_15),
.Y(n_318)
);

AO21x1_ASAP7_75t_L g321 ( 
.A1(n_318),
.A2(n_319),
.B(n_16),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_303),
.A2(n_16),
.B(n_5),
.Y(n_319)
);

AOI31xp33_ASAP7_75t_L g326 ( 
.A1(n_321),
.A2(n_322),
.A3(n_323),
.B(n_325),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_313),
.Y(n_325)
);

NAND2xp33_ASAP7_75t_SL g327 ( 
.A(n_324),
.B(n_308),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_308),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_328),
.B(n_326),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_6),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_6),
.Y(n_331)
);


endmodule