module fake_jpeg_31249_n_162 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_162);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_162;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_48),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

BUFx16f_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

BUFx16f_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_39),
.B(n_49),
.Y(n_55)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_5),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_34),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_7),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_33),
.B(n_41),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_10),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_21),
.Y(n_63)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_16),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_13),
.B(n_9),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_5),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_6),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_40),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_26),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_15),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_19),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_2),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_0),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_73),
.B(n_76),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_62),
.B(n_0),
.Y(n_74)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_74),
.Y(n_84)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_77),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_78),
.Y(n_85)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_79),
.Y(n_87)
);

CKINVDCx14_ASAP7_75t_R g80 ( 
.A(n_53),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_80),
.B(n_58),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_23),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_81),
.B(n_67),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_75),
.B(n_62),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_86),
.B(n_91),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_78),
.A2(n_71),
.B1(n_61),
.B2(n_54),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_88),
.A2(n_69),
.B1(n_52),
.B2(n_63),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_90),
.B(n_57),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_74),
.B(n_65),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_60),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_95),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_81),
.B(n_72),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_93),
.B(n_96),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_94),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_59),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_84),
.A2(n_70),
.B1(n_61),
.B2(n_71),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_97),
.A2(n_105),
.B1(n_106),
.B2(n_115),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_86),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_100),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_89),
.B(n_96),
.C(n_83),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_99),
.B(n_103),
.C(n_102),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_53),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_101),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_93),
.B(n_57),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_103),
.A2(n_111),
.B(n_11),
.Y(n_130)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_82),
.Y(n_104)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_104),
.Y(n_135)
);

OAI22xp33_ASAP7_75t_L g105 ( 
.A1(n_85),
.A2(n_79),
.B1(n_64),
.B2(n_66),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_91),
.A2(n_56),
.B1(n_66),
.B2(n_52),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_82),
.B(n_51),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_108),
.B(n_110),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_87),
.B(n_50),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_87),
.A2(n_76),
.B(n_50),
.Y(n_111)
);

NAND2x1p5_ASAP7_75t_L g112 ( 
.A(n_85),
.B(n_56),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_112),
.A2(n_114),
.B(n_107),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_113),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_94),
.A2(n_69),
.B1(n_68),
.B2(n_25),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_89),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_116),
.B(n_12),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_86),
.B(n_55),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_117),
.B(n_14),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_118),
.A2(n_127),
.B1(n_132),
.B2(n_18),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_101),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_119),
.B(n_130),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_112),
.A2(n_20),
.B(n_45),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_122),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_123),
.B(n_131),
.C(n_136),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_113),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_125),
.A2(n_15),
.B1(n_47),
.B2(n_24),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_99),
.B(n_6),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_126),
.B(n_133),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_105),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_100),
.A2(n_10),
.B(n_11),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_129),
.B(n_134),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_109),
.B(n_31),
.C(n_44),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_114),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_35),
.C(n_43),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_137),
.B(n_28),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_138),
.A2(n_139),
.B1(n_147),
.B2(n_30),
.Y(n_154)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_135),
.Y(n_140)
);

INVx1_ASAP7_75t_SL g151 ( 
.A(n_140),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_123),
.B(n_42),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_141),
.B(n_129),
.C(n_131),
.Y(n_150)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_134),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_144),
.A2(n_149),
.B(n_120),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_128),
.A2(n_122),
.B1(n_121),
.B2(n_124),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_150),
.B(n_152),
.Y(n_156)
);

AOI322xp5_ASAP7_75t_L g153 ( 
.A1(n_142),
.A2(n_124),
.A3(n_128),
.B1(n_136),
.B2(n_37),
.C1(n_29),
.C2(n_36),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_153),
.A2(n_154),
.B1(n_142),
.B2(n_143),
.Y(n_155)
);

AOI321xp33_ASAP7_75t_L g158 ( 
.A1(n_155),
.A2(n_157),
.A3(n_153),
.B1(n_141),
.B2(n_146),
.C(n_38),
.Y(n_158)
);

OAI22xp33_ASAP7_75t_L g157 ( 
.A1(n_151),
.A2(n_143),
.B1(n_148),
.B2(n_145),
.Y(n_157)
);

BUFx24_ASAP7_75t_SL g159 ( 
.A(n_158),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_159),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_160),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_156),
.Y(n_162)
);


endmodule