module fake_jpeg_17031_n_302 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_302);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_302;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_288;
wire n_272;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_241;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

INVx4_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx1_ASAP7_75t_SL g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx24_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_26),
.B(n_28),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_16),
.B(n_22),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_16),
.B(n_11),
.Y(n_29)
);

BUFx24_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_16),
.B(n_11),
.Y(n_32)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx16f_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx16f_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_43),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_26),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_44),
.A2(n_13),
.B1(n_30),
.B2(n_34),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_48),
.A2(n_65),
.B1(n_43),
.B2(n_39),
.Y(n_85)
);

CKINVDCx14_ASAP7_75t_R g49 ( 
.A(n_36),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_49),
.B(n_55),
.Y(n_84)
);

OA22x2_ASAP7_75t_L g50 ( 
.A1(n_36),
.A2(n_46),
.B1(n_34),
.B2(n_30),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_50),
.B(n_51),
.Y(n_82)
);

OA22x2_ASAP7_75t_L g51 ( 
.A1(n_36),
.A2(n_46),
.B1(n_19),
.B2(n_31),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_28),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_53),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_38),
.Y(n_53)
);

CKINVDCx14_ASAP7_75t_R g55 ( 
.A(n_36),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_41),
.A2(n_13),
.B1(n_19),
.B2(n_22),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_56),
.A2(n_57),
.B1(n_61),
.B2(n_67),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_45),
.A2(n_35),
.B1(n_33),
.B2(n_19),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_40),
.B(n_29),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_59),
.B(n_32),
.Y(n_69)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_41),
.A2(n_19),
.B1(n_20),
.B2(n_14),
.Y(n_61)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_62),
.Y(n_88)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_64),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_42),
.A2(n_35),
.B1(n_33),
.B2(n_15),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_42),
.A2(n_14),
.B1(n_20),
.B2(n_26),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_68),
.B(n_70),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_69),
.B(n_86),
.Y(n_89)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

O2A1O1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_50),
.A2(n_42),
.B(n_31),
.C(n_23),
.Y(n_71)
);

CKINVDCx14_ASAP7_75t_R g101 ( 
.A(n_71),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_52),
.A2(n_53),
.B1(n_59),
.B2(n_38),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_51),
.Y(n_93)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g78 ( 
.A(n_51),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_78),
.B(n_81),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_67),
.A2(n_47),
.B1(n_43),
.B2(n_39),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_79),
.A2(n_85),
.B1(n_63),
.B2(n_65),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_62),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_49),
.B(n_38),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_50),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_50),
.Y(n_105)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_90),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_77),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_91),
.B(n_103),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_93),
.A2(n_95),
.B1(n_105),
.B2(n_107),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_72),
.B(n_50),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_94),
.B(n_82),
.Y(n_109)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_96),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_72),
.B(n_50),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_98),
.A2(n_106),
.B(n_108),
.Y(n_128)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_99),
.Y(n_127)
);

AOI21xp33_ASAP7_75t_L g102 ( 
.A1(n_86),
.A2(n_38),
.B(n_55),
.Y(n_102)
);

OAI21xp33_ASAP7_75t_L g113 ( 
.A1(n_102),
.A2(n_88),
.B(n_84),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_80),
.Y(n_103)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_68),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_104),
.B(n_92),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_73),
.B(n_75),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_87),
.A2(n_67),
.B1(n_56),
.B2(n_63),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_73),
.B(n_51),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_109),
.B(n_126),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_94),
.B(n_81),
.C(n_88),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_110),
.B(n_112),
.C(n_114),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_107),
.B(n_51),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_111),
.A2(n_82),
.B(n_78),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_106),
.B(n_69),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_113),
.A2(n_93),
.B(n_101),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_89),
.B(n_64),
.C(n_60),
.Y(n_114)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_90),
.Y(n_116)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_116),
.Y(n_135)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_96),
.Y(n_118)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_118),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_89),
.B(n_84),
.Y(n_119)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_119),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_106),
.C(n_98),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_120),
.B(n_57),
.C(n_83),
.Y(n_159)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_99),
.Y(n_121)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_121),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_92),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_122),
.B(n_124),
.Y(n_139)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_123),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_100),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_98),
.B(n_82),
.Y(n_126)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_126),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_103),
.B(n_83),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_129),
.B(n_132),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_104),
.B(n_70),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_131),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_97),
.Y(n_132)
);

BUFx5_ASAP7_75t_L g133 ( 
.A(n_124),
.Y(n_133)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_133),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_112),
.B(n_93),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_134),
.B(n_159),
.C(n_57),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g136 ( 
.A(n_111),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_136),
.B(n_145),
.Y(n_160)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_137),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_138),
.A2(n_128),
.B1(n_110),
.B2(n_114),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_130),
.A2(n_95),
.B1(n_108),
.B2(n_78),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_140),
.A2(n_111),
.B1(n_109),
.B2(n_130),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_115),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_141),
.B(n_146),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_119),
.B(n_91),
.Y(n_142)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_142),
.Y(n_176)
);

INVx13_ASAP7_75t_L g145 ( 
.A(n_116),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_118),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_148),
.A2(n_127),
.B1(n_71),
.B2(n_61),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_115),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_150),
.B(n_151),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_117),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_132),
.B(n_108),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_152),
.B(n_128),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_125),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_155),
.B(n_157),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_125),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_133),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_161),
.B(n_163),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_152),
.B(n_120),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_162),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_155),
.Y(n_163)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_164),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_165),
.A2(n_170),
.B1(n_181),
.B2(n_186),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_157),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_166),
.B(n_173),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_168),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_140),
.A2(n_82),
.B1(n_127),
.B2(n_121),
.Y(n_170)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_171),
.Y(n_194)
);

BUFx12f_ASAP7_75t_L g172 ( 
.A(n_145),
.Y(n_172)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_172),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_135),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_142),
.B(n_71),
.Y(n_174)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_174),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_179),
.B(n_184),
.C(n_143),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_149),
.Y(n_180)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_180),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_151),
.A2(n_136),
.B1(n_154),
.B2(n_138),
.Y(n_181)
);

OA21x2_ASAP7_75t_L g182 ( 
.A1(n_137),
.A2(n_79),
.B(n_51),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_182),
.B(n_183),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_156),
.A2(n_74),
.B(n_70),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_143),
.B(n_68),
.C(n_37),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_135),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_185),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_156),
.A2(n_148),
.B1(n_159),
.B2(n_147),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_188),
.B(n_189),
.C(n_198),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_184),
.B(n_134),
.C(n_147),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_179),
.B(n_139),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_191),
.B(n_199),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_186),
.B(n_150),
.C(n_141),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_164),
.B(n_158),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_168),
.B(n_153),
.C(n_149),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_201),
.B(n_204),
.C(n_207),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_177),
.A2(n_153),
.B(n_146),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_202),
.B(n_174),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_170),
.B(n_144),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_178),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_205),
.B(n_172),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_183),
.B(n_144),
.C(n_37),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_162),
.B(n_48),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_209),
.B(n_171),
.C(n_163),
.Y(n_216)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_210),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_200),
.B(n_176),
.Y(n_211)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_211),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_193),
.B(n_175),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_213),
.A2(n_209),
.B(n_23),
.Y(n_230)
);

AOI21xp33_ASAP7_75t_L g214 ( 
.A1(n_206),
.A2(n_162),
.B(n_160),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_214),
.B(n_217),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_216),
.B(n_31),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_194),
.A2(n_190),
.B1(n_187),
.B2(n_196),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_198),
.A2(n_195),
.B1(n_201),
.B2(n_166),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_218),
.B(n_222),
.Y(n_240)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_219),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_191),
.B(n_169),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_220),
.B(n_228),
.C(n_21),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_199),
.A2(n_169),
.B1(n_167),
.B2(n_182),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_192),
.B(n_172),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_223),
.Y(n_239)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_197),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_224),
.B(n_227),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_208),
.B(n_161),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_225),
.B(n_11),
.Y(n_232)
);

INVx2_ASAP7_75t_SL g226 ( 
.A(n_203),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_226),
.B(n_0),
.Y(n_242)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_204),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_188),
.B(n_189),
.C(n_207),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_195),
.A2(n_182),
.B1(n_92),
.B2(n_47),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_229),
.A2(n_25),
.B1(n_24),
.B2(n_15),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_230),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_231),
.B(n_241),
.C(n_243),
.Y(n_252)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_232),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_213),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_238),
.B(n_219),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_212),
.B(n_37),
.C(n_39),
.Y(n_241)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_242),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_212),
.B(n_21),
.C(n_18),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_244),
.B(n_215),
.C(n_228),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_245),
.A2(n_229),
.B1(n_226),
.B2(n_216),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_247),
.B(n_249),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_248),
.B(n_250),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_238),
.B(n_220),
.Y(n_249)
);

INVx6_ASAP7_75t_L g250 ( 
.A(n_233),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_234),
.A2(n_221),
.B(n_215),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_251),
.A2(n_235),
.B(n_243),
.Y(n_260)
);

OAI21xp33_ASAP7_75t_L g253 ( 
.A1(n_237),
.A2(n_236),
.B(n_240),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_253),
.B(n_254),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_231),
.B(n_221),
.C(n_25),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_255),
.B(n_256),
.C(n_259),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_241),
.B(n_25),
.C(n_24),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_239),
.B(n_242),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_258),
.B(n_230),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_260),
.A2(n_270),
.B(n_1),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_261),
.B(n_265),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_264),
.A2(n_257),
.B1(n_250),
.B2(n_246),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_254),
.B(n_244),
.C(n_245),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_252),
.B(n_25),
.C(n_24),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_266),
.B(n_267),
.C(n_269),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_252),
.B(n_24),
.C(n_15),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_255),
.B(n_21),
.C(n_18),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_248),
.B(n_21),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_256),
.B(n_21),
.C(n_18),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_271),
.B(n_17),
.C(n_18),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_272),
.A2(n_274),
.B(n_2),
.Y(n_282)
);

OR2x2_ASAP7_75t_L g273 ( 
.A(n_263),
.B(n_253),
.Y(n_273)
);

OR2x2_ASAP7_75t_L g287 ( 
.A(n_273),
.B(n_278),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_268),
.A2(n_0),
.B(n_1),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_275),
.B(n_279),
.C(n_280),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_262),
.B(n_21),
.C(n_18),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_264),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_268),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_281),
.B(n_17),
.C(n_12),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_282),
.B(n_283),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_277),
.A2(n_3),
.B(n_5),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_276),
.B(n_18),
.C(n_12),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_285),
.B(n_279),
.C(n_276),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_273),
.A2(n_5),
.B(n_6),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_286),
.B(n_278),
.C(n_17),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_288),
.B(n_5),
.Y(n_290)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_289),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_290),
.A2(n_291),
.B(n_287),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_294),
.B(n_284),
.C(n_292),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_295),
.B(n_293),
.C(n_17),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_296),
.B(n_7),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_297),
.B(n_17),
.C(n_8),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_298),
.B(n_7),
.C(n_8),
.Y(n_299)
);

AOI322xp5_ASAP7_75t_L g300 ( 
.A1(n_299),
.A2(n_7),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.C1(n_294),
.C2(n_280),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_300),
.B(n_7),
.Y(n_301)
);

OA21x2_ASAP7_75t_L g302 ( 
.A1(n_301),
.A2(n_10),
.B(n_8),
.Y(n_302)
);


endmodule