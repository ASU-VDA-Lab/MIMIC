module fake_jpeg_29808_n_548 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_548);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_548;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx8_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx14_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_14),
.Y(n_36)
);

INVx8_ASAP7_75t_SL g37 ( 
.A(n_0),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_12),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_17),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_7),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_3),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

BUFx16f_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_13),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_5),
.Y(n_55)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_56),
.Y(n_141)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_17),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_57),
.B(n_84),
.Y(n_118)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_58),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_59),
.Y(n_143)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_60),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_61),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_62),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_63),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_64),
.Y(n_134)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_65),
.Y(n_128)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_66),
.Y(n_164)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_67),
.Y(n_116)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_68),
.Y(n_114)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_69),
.Y(n_120)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_70),
.Y(n_166)
);

INVx3_ASAP7_75t_SL g71 ( 
.A(n_31),
.Y(n_71)
);

INVx2_ASAP7_75t_SL g115 ( 
.A(n_71),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_39),
.B(n_15),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_72),
.B(n_79),
.Y(n_132)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_73),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_74),
.Y(n_150)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_30),
.Y(n_75)
);

INVx2_ASAP7_75t_SL g174 ( 
.A(n_75),
.Y(n_174)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_30),
.Y(n_76)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_76),
.Y(n_159)
);

HB1xp67_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_77),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_78),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_20),
.B(n_15),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

BUFx4f_ASAP7_75t_SL g177 ( 
.A(n_80),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

INVx8_ASAP7_75t_L g148 ( 
.A(n_81),
.Y(n_148)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_23),
.Y(n_82)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_82),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_37),
.Y(n_83)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_83),
.Y(n_163)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_37),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_85),
.B(n_101),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_20),
.B(n_1),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_86),
.B(n_110),
.Y(n_139)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_31),
.Y(n_87)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_87),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

INVx11_ASAP7_75t_L g122 ( 
.A(n_88),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

INVx11_ASAP7_75t_L g135 ( 
.A(n_89),
.Y(n_135)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_43),
.Y(n_90)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_90),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_91),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_51),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_92),
.Y(n_119)
);

BUFx8_ASAP7_75t_L g93 ( 
.A(n_30),
.Y(n_93)
);

CKINVDCx9p33_ASAP7_75t_R g131 ( 
.A(n_93),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_51),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g145 ( 
.A(n_94),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_18),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_95),
.Y(n_146)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_23),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g125 ( 
.A(n_96),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_51),
.Y(n_97)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_97),
.Y(n_142)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_30),
.Y(n_98)
);

BUFx16f_ASAP7_75t_L g124 ( 
.A(n_98),
.Y(n_124)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_42),
.Y(n_99)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_99),
.Y(n_149)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_30),
.Y(n_100)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_100),
.Y(n_162)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_26),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_42),
.Y(n_102)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_102),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_18),
.Y(n_103)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_103),
.Y(n_170)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_42),
.Y(n_104)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_104),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_18),
.Y(n_105)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_105),
.Y(n_175)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_23),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_106),
.B(n_107),
.Y(n_137)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_33),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_26),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_108),
.B(n_113),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_33),
.Y(n_109)
);

INVx6_ASAP7_75t_SL g165 ( 
.A(n_109),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_19),
.B(n_15),
.Y(n_110)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_47),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_111),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_33),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_112),
.A2(n_48),
.B1(n_47),
.B2(n_53),
.Y(n_152)
);

BUFx12f_ASAP7_75t_L g113 ( 
.A(n_47),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_86),
.B(n_53),
.C(n_52),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_117),
.B(n_32),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g123 ( 
.A(n_80),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_123),
.B(n_160),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_57),
.B(n_27),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_144),
.B(n_156),
.Y(n_203)
);

OA22x2_ASAP7_75t_L g189 ( 
.A1(n_152),
.A2(n_78),
.B1(n_59),
.B2(n_61),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_71),
.A2(n_48),
.B1(n_47),
.B2(n_29),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_153),
.A2(n_154),
.B1(n_171),
.B2(n_63),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_109),
.A2(n_25),
.B1(n_45),
.B2(n_40),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_110),
.B(n_25),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_79),
.B(n_36),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_157),
.B(n_158),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_77),
.B(n_27),
.Y(n_158)
);

AOI21xp33_ASAP7_75t_L g160 ( 
.A1(n_83),
.A2(n_52),
.B(n_46),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_93),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_167),
.B(n_169),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_113),
.B(n_24),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_112),
.A2(n_48),
.B1(n_47),
.B2(n_46),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_99),
.B(n_21),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_178),
.B(n_48),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_179),
.B(n_191),
.Y(n_268)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_116),
.Y(n_180)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_180),
.Y(n_264)
);

INVx6_ASAP7_75t_L g181 ( 
.A(n_122),
.Y(n_181)
);

BUFx2_ASAP7_75t_L g262 ( 
.A(n_181),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_127),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_182),
.B(n_187),
.Y(n_243)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_126),
.Y(n_183)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_183),
.Y(n_259)
);

BUFx12f_ASAP7_75t_L g184 ( 
.A(n_124),
.Y(n_184)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_184),
.Y(n_269)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_128),
.Y(n_185)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_185),
.Y(n_245)
);

INVx4_ASAP7_75t_SL g186 ( 
.A(n_131),
.Y(n_186)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_186),
.Y(n_246)
);

A2O1A1Ixp33_ASAP7_75t_L g187 ( 
.A1(n_139),
.A2(n_32),
.B(n_29),
.C(n_45),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_165),
.A2(n_105),
.B1(n_103),
.B2(n_56),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_188),
.A2(n_234),
.B1(n_115),
.B2(n_140),
.Y(n_237)
);

AO22x2_ASAP7_75t_L g255 ( 
.A1(n_189),
.A2(n_233),
.B1(n_140),
.B2(n_176),
.Y(n_255)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_166),
.Y(n_190)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_190),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_118),
.B(n_97),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_192),
.A2(n_193),
.B1(n_208),
.B2(n_224),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_132),
.A2(n_88),
.B1(n_64),
.B2(n_91),
.Y(n_193)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_126),
.Y(n_194)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_194),
.Y(n_277)
);

HB1xp67_ASAP7_75t_L g195 ( 
.A(n_159),
.Y(n_195)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_195),
.Y(n_280)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_120),
.Y(n_196)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_196),
.Y(n_241)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_138),
.Y(n_197)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_197),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_147),
.B(n_24),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_199),
.B(n_221),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_124),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_200),
.B(n_206),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_133),
.A2(n_89),
.B1(n_62),
.B2(n_74),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_201),
.A2(n_155),
.B1(n_150),
.B2(n_134),
.Y(n_238)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_142),
.Y(n_202)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_202),
.Y(n_257)
);

INVx6_ASAP7_75t_L g205 ( 
.A(n_122),
.Y(n_205)
);

INVx6_ASAP7_75t_L g263 ( 
.A(n_205),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_129),
.B(n_19),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_207),
.B(n_211),
.Y(n_244)
);

OAI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_170),
.A2(n_175),
.B1(n_155),
.B2(n_150),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_153),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_209),
.B(n_217),
.Y(n_251)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_159),
.Y(n_210)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_210),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_168),
.B(n_172),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_162),
.Y(n_212)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_212),
.Y(n_273)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_130),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_213),
.Y(n_252)
);

INVx3_ASAP7_75t_SL g214 ( 
.A(n_114),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_214),
.Y(n_258)
);

AND2x2_ASAP7_75t_SL g215 ( 
.A(n_149),
.B(n_94),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_215),
.B(n_121),
.C(n_148),
.Y(n_250)
);

BUFx12f_ASAP7_75t_L g216 ( 
.A(n_130),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_216),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_137),
.B(n_40),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_164),
.B(n_54),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_218),
.B(n_219),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_119),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_134),
.B(n_38),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_136),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_222),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_164),
.B(n_54),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_223),
.B(n_227),
.Y(n_270)
);

OAI22xp33_ASAP7_75t_L g224 ( 
.A1(n_135),
.A2(n_81),
.B1(n_92),
.B2(n_38),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_143),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_225),
.A2(n_228),
.B1(n_230),
.B2(n_232),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_115),
.A2(n_2),
.B(n_3),
.Y(n_226)
);

OAI21xp33_ASAP7_75t_SL g266 ( 
.A1(n_226),
.A2(n_235),
.B(n_236),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_174),
.B(n_36),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_119),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_114),
.B(n_151),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_229),
.B(n_2),
.Y(n_278)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_136),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_152),
.A2(n_28),
.B1(n_21),
.B2(n_48),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_231),
.A2(n_161),
.B1(n_28),
.B2(n_135),
.Y(n_275)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_125),
.Y(n_232)
);

OA22x2_ASAP7_75t_L g233 ( 
.A1(n_171),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_163),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_141),
.Y(n_235)
);

CKINVDCx12_ASAP7_75t_R g236 ( 
.A(n_177),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g303 ( 
.A1(n_237),
.A2(n_184),
.B1(n_216),
.B2(n_213),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_238),
.A2(n_248),
.B1(n_255),
.B2(n_274),
.Y(n_312)
);

AO22x1_ASAP7_75t_L g240 ( 
.A1(n_198),
.A2(n_177),
.B1(n_145),
.B2(n_141),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_240),
.B(n_247),
.Y(n_306)
);

AOI22x1_ASAP7_75t_SL g247 ( 
.A1(n_209),
.A2(n_146),
.B1(n_145),
.B2(n_125),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_221),
.A2(n_176),
.B1(n_143),
.B2(n_173),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_250),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_179),
.B(n_121),
.C(n_146),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_254),
.B(n_256),
.C(n_272),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_179),
.B(n_174),
.C(n_163),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_191),
.B(n_148),
.C(n_173),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_191),
.A2(n_233),
.B1(n_189),
.B2(n_215),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_275),
.A2(n_267),
.B1(n_246),
.B2(n_186),
.Y(n_288)
);

AOI32xp33_ASAP7_75t_L g276 ( 
.A1(n_204),
.A2(n_125),
.A3(n_177),
.B1(n_161),
.B2(n_6),
.Y(n_276)
);

AOI32xp33_ASAP7_75t_L g301 ( 
.A1(n_276),
.A2(n_215),
.A3(n_214),
.B1(n_232),
.B2(n_189),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_278),
.Y(n_294)
);

AND2x2_ASAP7_75t_SL g281 ( 
.A(n_240),
.B(n_226),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_281),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_244),
.B(n_220),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_282),
.B(n_287),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_249),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_283),
.B(n_285),
.Y(n_324)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_269),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_284),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_249),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_279),
.B(n_233),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_288),
.A2(n_238),
.B1(n_224),
.B2(n_235),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_270),
.B(n_199),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_289),
.B(n_291),
.Y(n_326)
);

BUFx3_ASAP7_75t_L g290 ( 
.A(n_269),
.Y(n_290)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_290),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_260),
.B(n_203),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_263),
.Y(n_292)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_292),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_247),
.A2(n_233),
.B(n_189),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_293),
.A2(n_255),
.B(n_265),
.Y(n_323)
);

INVx13_ASAP7_75t_L g295 ( 
.A(n_259),
.Y(n_295)
);

INVxp33_ASAP7_75t_L g316 ( 
.A(n_295),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_279),
.B(n_196),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_296),
.B(n_299),
.Y(n_342)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_257),
.Y(n_297)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_297),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_243),
.B(n_187),
.Y(n_298)
);

NAND3xp33_ASAP7_75t_L g339 ( 
.A(n_298),
.B(n_280),
.C(n_253),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_268),
.B(n_197),
.Y(n_299)
);

INVx13_ASAP7_75t_L g300 ( 
.A(n_259),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_300),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_301),
.A2(n_255),
.B1(n_272),
.B2(n_250),
.Y(n_317)
);

INVx13_ASAP7_75t_L g302 ( 
.A(n_239),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_302),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_303),
.A2(n_267),
.B1(n_275),
.B2(n_262),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_268),
.B(n_180),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_304),
.B(n_305),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_242),
.B(n_210),
.Y(n_305)
);

INVxp67_ASAP7_75t_SL g307 ( 
.A(n_258),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_307),
.B(n_314),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_268),
.B(n_229),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_309),
.B(n_313),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_266),
.A2(n_229),
.B(n_183),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_310),
.A2(n_252),
.B(n_277),
.Y(n_340)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_257),
.Y(n_311)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_311),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_278),
.B(n_202),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_251),
.B(n_230),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_241),
.Y(n_315)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_315),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_317),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_306),
.B(n_293),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g358 ( 
.A1(n_320),
.A2(n_323),
.B(n_325),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_312),
.A2(n_255),
.B1(n_256),
.B2(n_254),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_328),
.A2(n_338),
.B1(n_306),
.B2(n_286),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_329),
.A2(n_337),
.B1(n_343),
.B2(n_293),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_306),
.B(n_273),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g368 ( 
.A1(n_332),
.A2(n_340),
.B(n_310),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_288),
.A2(n_273),
.B1(n_261),
.B2(n_245),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_312),
.A2(n_225),
.B1(n_241),
.B2(n_253),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_339),
.B(n_298),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_288),
.A2(n_306),
.B1(n_281),
.B2(n_312),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_308),
.B(n_271),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_344),
.B(n_345),
.C(n_313),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_308),
.B(n_271),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_297),
.Y(n_346)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_346),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_348),
.A2(n_371),
.B1(n_337),
.B2(n_360),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_319),
.B(n_342),
.Y(n_350)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_350),
.Y(n_393)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_330),
.Y(n_352)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_352),
.Y(n_396)
);

CKINVDCx12_ASAP7_75t_R g353 ( 
.A(n_335),
.Y(n_353)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_353),
.Y(n_380)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_330),
.Y(n_354)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_354),
.Y(n_404)
);

CKINVDCx16_ASAP7_75t_R g355 ( 
.A(n_324),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_355),
.B(n_359),
.Y(n_385)
);

XOR2x2_ASAP7_75t_L g356 ( 
.A(n_345),
.B(n_281),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_356),
.B(n_332),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_344),
.B(n_308),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_357),
.B(n_375),
.C(n_327),
.Y(n_378)
);

OR2x2_ASAP7_75t_L g360 ( 
.A(n_322),
.B(n_287),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_360),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_361),
.A2(n_323),
.B1(n_340),
.B2(n_329),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_321),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_362),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_321),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_363),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_343),
.A2(n_281),
.B1(n_301),
.B2(n_310),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_364),
.B(n_365),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_319),
.B(n_296),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_326),
.B(n_291),
.Y(n_366)
);

INVxp33_ASAP7_75t_L g407 ( 
.A(n_366),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_326),
.B(n_299),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_367),
.B(n_369),
.Y(n_400)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_368),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_317),
.A2(n_281),
.B1(n_304),
.B2(n_303),
.Y(n_369)
);

CKINVDCx10_ASAP7_75t_R g370 ( 
.A(n_335),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_370),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_338),
.A2(n_314),
.B1(n_305),
.B2(n_294),
.Y(n_371)
);

AND2x6_ASAP7_75t_L g372 ( 
.A(n_322),
.B(n_300),
.Y(n_372)
);

NOR3xp33_ASAP7_75t_L g399 ( 
.A(n_372),
.B(n_334),
.C(n_309),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_SL g373 ( 
.A(n_331),
.B(n_282),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_373),
.Y(n_406)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_336),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_374),
.B(n_377),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_334),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_376),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_342),
.B(n_315),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_378),
.B(n_379),
.C(n_386),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_357),
.B(n_327),
.C(n_320),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_375),
.B(n_320),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_383),
.B(n_384),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_356),
.B(n_347),
.C(n_332),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_348),
.B(n_347),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_388),
.B(n_401),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_390),
.A2(n_389),
.B1(n_387),
.B2(n_393),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_391),
.A2(n_351),
.B1(n_360),
.B2(n_358),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_373),
.B(n_355),
.Y(n_392)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_392),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_366),
.B(n_289),
.Y(n_394)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_394),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_371),
.B(n_284),
.Y(n_397)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_397),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_399),
.B(n_283),
.Y(n_429)
);

XNOR2x1_ASAP7_75t_L g401 ( 
.A(n_364),
.B(n_346),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_350),
.B(n_290),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_402),
.B(n_277),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_SL g405 ( 
.A(n_356),
.B(n_341),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_405),
.B(n_311),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g444 ( 
.A(n_412),
.B(n_432),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_406),
.A2(n_376),
.B1(n_367),
.B2(n_365),
.Y(n_413)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_413),
.Y(n_443)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_396),
.Y(n_414)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_414),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_406),
.A2(n_377),
.B1(n_353),
.B2(n_370),
.Y(n_416)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_416),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_391),
.A2(n_361),
.B1(n_358),
.B2(n_369),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_417),
.B(n_419),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_381),
.A2(n_372),
.B1(n_368),
.B2(n_374),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_378),
.B(n_354),
.C(n_352),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_420),
.B(n_421),
.C(n_422),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_383),
.B(n_379),
.C(n_405),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_386),
.B(n_349),
.C(n_341),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_388),
.B(n_349),
.C(n_336),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_423),
.B(n_408),
.C(n_400),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_SL g447 ( 
.A(n_424),
.B(n_380),
.Y(n_447)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_396),
.Y(n_426)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_426),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_L g427 ( 
.A1(n_385),
.A2(n_363),
.B1(n_362),
.B2(n_318),
.Y(n_427)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_427),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_381),
.A2(n_318),
.B1(n_333),
.B2(n_292),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_428),
.B(n_429),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_407),
.B(n_290),
.Y(n_430)
);

CKINVDCx16_ASAP7_75t_R g457 ( 
.A(n_430),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_L g431 ( 
.A1(n_382),
.A2(n_333),
.B(n_284),
.Y(n_431)
);

AOI21xp5_ASAP7_75t_L g442 ( 
.A1(n_431),
.A2(n_437),
.B(n_380),
.Y(n_442)
);

HB1xp67_ASAP7_75t_L g433 ( 
.A(n_393),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g460 ( 
.A(n_433),
.Y(n_460)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_404),
.Y(n_434)
);

CKINVDCx16_ASAP7_75t_R g461 ( 
.A(n_434),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_389),
.A2(n_292),
.B1(n_285),
.B2(n_263),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_435),
.B(n_404),
.Y(n_448)
);

XNOR2x2_ASAP7_75t_L g436 ( 
.A(n_382),
.B(n_316),
.Y(n_436)
);

FAx1_ASAP7_75t_L g439 ( 
.A(n_436),
.B(n_429),
.CI(n_432),
.CON(n_439),
.SN(n_439)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_415),
.B(n_401),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_438),
.B(n_445),
.C(n_450),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_SL g463 ( 
.A(n_439),
.B(n_436),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_409),
.B(n_384),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_440),
.B(n_446),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_442),
.B(n_447),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_415),
.B(n_400),
.Y(n_445)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_448),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_421),
.B(n_409),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_418),
.B(n_408),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_453),
.B(n_455),
.C(n_458),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_420),
.B(n_422),
.C(n_423),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_418),
.B(n_398),
.C(n_395),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_449),
.B(n_395),
.Y(n_462)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_462),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_463),
.A2(n_472),
.B1(n_471),
.B2(n_479),
.Y(n_498)
);

INVxp67_ASAP7_75t_SL g464 ( 
.A(n_452),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_464),
.B(n_465),
.Y(n_482)
);

INVxp33_ASAP7_75t_L g465 ( 
.A(n_451),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g469 ( 
.A1(n_454),
.A2(n_443),
.B1(n_459),
.B2(n_444),
.Y(n_469)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_469),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_456),
.B(n_398),
.Y(n_470)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_470),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_444),
.A2(n_417),
.B1(n_412),
.B2(n_419),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_472),
.A2(n_479),
.B1(n_453),
.B2(n_438),
.Y(n_497)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_458),
.Y(n_473)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_473),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_461),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_474),
.B(n_476),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_460),
.B(n_410),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_SL g477 ( 
.A1(n_439),
.A2(n_425),
.B(n_411),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_477),
.B(n_431),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_455),
.B(n_424),
.C(n_428),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_478),
.B(n_441),
.C(n_445),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_448),
.A2(n_435),
.B1(n_434),
.B2(n_414),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_446),
.B(n_403),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_480),
.B(n_474),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_483),
.B(n_484),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_SL g484 ( 
.A(n_475),
.B(n_439),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_485),
.B(n_467),
.Y(n_505)
);

OAI21xp5_ASAP7_75t_L g503 ( 
.A1(n_487),
.A2(n_470),
.B(n_463),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_476),
.B(n_473),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_488),
.B(n_490),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_468),
.B(n_441),
.Y(n_490)
);

NOR2xp67_ASAP7_75t_SL g491 ( 
.A(n_468),
.B(n_447),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_SL g510 ( 
.A(n_491),
.B(n_184),
.Y(n_510)
);

OAI21xp5_ASAP7_75t_SL g493 ( 
.A1(n_469),
.A2(n_460),
.B(n_426),
.Y(n_493)
);

AOI21xp5_ASAP7_75t_L g507 ( 
.A1(n_493),
.A2(n_302),
.B(n_300),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_462),
.B(n_457),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_494),
.B(n_495),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_SL g495 ( 
.A(n_466),
.B(n_477),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_497),
.A2(n_295),
.B1(n_194),
.B2(n_222),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_498),
.B(n_497),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_490),
.B(n_467),
.C(n_450),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_499),
.B(n_504),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_SL g518 ( 
.A(n_500),
.B(n_507),
.Y(n_518)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_503),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_L g504 ( 
.A1(n_486),
.A2(n_471),
.B1(n_478),
.B2(n_403),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_505),
.B(n_506),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_485),
.B(n_239),
.C(n_264),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_483),
.B(n_307),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_SL g524 ( 
.A(n_508),
.B(n_512),
.Y(n_524)
);

AOI22xp33_ASAP7_75t_SL g509 ( 
.A1(n_489),
.A2(n_262),
.B1(n_302),
.B2(n_181),
.Y(n_509)
);

AOI21xp5_ASAP7_75t_SL g525 ( 
.A1(n_509),
.A2(n_295),
.B(n_216),
.Y(n_525)
);

AOI21xp5_ASAP7_75t_L g516 ( 
.A1(n_510),
.A2(n_494),
.B(n_482),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_492),
.B(n_264),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_L g523 ( 
.A(n_511),
.B(n_514),
.Y(n_523)
);

XOR2xp5_ASAP7_75t_L g517 ( 
.A(n_513),
.B(n_481),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_481),
.B(n_205),
.Y(n_514)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_516),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_L g533 ( 
.A1(n_517),
.A2(n_524),
.B1(n_5),
.B2(n_8),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_499),
.B(n_496),
.C(n_498),
.Y(n_519)
);

INVxp67_ASAP7_75t_L g529 ( 
.A(n_519),
.Y(n_529)
);

MAJx2_ASAP7_75t_L g520 ( 
.A(n_501),
.B(n_496),
.C(n_493),
.Y(n_520)
);

OAI21xp5_ASAP7_75t_L g530 ( 
.A1(n_520),
.A2(n_506),
.B(n_8),
.Y(n_530)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_525),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_502),
.B(n_2),
.C(n_3),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_SL g527 ( 
.A(n_526),
.B(n_5),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_527),
.B(n_528),
.Y(n_536)
);

AOI31xp33_ASAP7_75t_SL g528 ( 
.A1(n_515),
.A2(n_503),
.A3(n_509),
.B(n_513),
.Y(n_528)
);

HB1xp67_ASAP7_75t_L g539 ( 
.A(n_530),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_SL g532 ( 
.A(n_521),
.B(n_5),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_532),
.B(n_533),
.Y(n_537)
);

OAI21xp5_ASAP7_75t_SL g535 ( 
.A1(n_529),
.A2(n_522),
.B(n_525),
.Y(n_535)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_535),
.Y(n_541)
);

OAI21xp5_ASAP7_75t_SL g538 ( 
.A1(n_529),
.A2(n_520),
.B(n_518),
.Y(n_538)
);

AOI322xp5_ASAP7_75t_L g540 ( 
.A1(n_538),
.A2(n_534),
.A3(n_518),
.B1(n_531),
.B2(n_523),
.C1(n_8),
.C2(n_13),
.Y(n_540)
);

OAI21xp5_ASAP7_75t_L g544 ( 
.A1(n_540),
.A2(n_542),
.B(n_9),
.Y(n_544)
);

AOI322xp5_ASAP7_75t_L g542 ( 
.A1(n_536),
.A2(n_539),
.A3(n_537),
.B1(n_13),
.B2(n_14),
.C1(n_10),
.C2(n_9),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_541),
.B(n_9),
.C(n_10),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_543),
.B(n_544),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_545),
.B(n_9),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_546),
.Y(n_547)
);

AOI21xp5_ASAP7_75t_L g548 ( 
.A1(n_547),
.A2(n_14),
.B(n_541),
.Y(n_548)
);


endmodule