module fake_jpeg_14078_n_521 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_521);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_521;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_479;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx24_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_6),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_0),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_7),
.Y(n_50)
);

BUFx12_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_5),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_13),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_3),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_11),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_58),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_59),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_60),
.Y(n_143)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_61),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_62),
.Y(n_166)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

BUFx10_ASAP7_75t_L g191 ( 
.A(n_63),
.Y(n_191)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_64),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_65),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_21),
.B(n_17),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_66),
.B(n_70),
.Y(n_149)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_67),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_68),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

INVx6_ASAP7_75t_L g188 ( 
.A(n_69),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_21),
.B(n_15),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_23),
.Y(n_71)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_71),
.Y(n_194)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g163 ( 
.A(n_72),
.Y(n_163)
);

INVx3_ASAP7_75t_SL g73 ( 
.A(n_35),
.Y(n_73)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_73),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_49),
.B(n_1),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_74),
.B(n_78),
.Y(n_151)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_34),
.Y(n_75)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_75),
.Y(n_179)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_34),
.Y(n_76)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_76),
.Y(n_129)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_77),
.Y(n_193)
);

CKINVDCx6p67_ASAP7_75t_R g78 ( 
.A(n_35),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_23),
.Y(n_79)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_79),
.Y(n_122)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_80),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_23),
.Y(n_81)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_81),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_27),
.Y(n_82)
);

INVx8_ASAP7_75t_L g170 ( 
.A(n_82),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_27),
.Y(n_83)
);

INVx8_ASAP7_75t_L g197 ( 
.A(n_83),
.Y(n_197)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_22),
.Y(n_84)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_84),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_27),
.Y(n_85)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_85),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_36),
.Y(n_86)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_86),
.Y(n_152)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_40),
.Y(n_87)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_87),
.Y(n_148)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_35),
.Y(n_88)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_88),
.Y(n_156)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

INVx2_ASAP7_75t_SL g123 ( 
.A(n_89),
.Y(n_123)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_90),
.Y(n_158)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_18),
.Y(n_91)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_91),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_35),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_92),
.B(n_99),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_36),
.Y(n_93)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_93),
.Y(n_199)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_18),
.Y(n_94)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_94),
.Y(n_150)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_18),
.Y(n_95)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_95),
.Y(n_155)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_43),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_96),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_36),
.Y(n_97)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_97),
.Y(n_157)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_18),
.Y(n_98)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_98),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_24),
.B(n_1),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_24),
.Y(n_100)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_100),
.Y(n_124)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_30),
.Y(n_101)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_101),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_22),
.Y(n_102)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_102),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_18),
.B(n_15),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_103),
.B(n_109),
.Y(n_175)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_29),
.Y(n_104)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_104),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_40),
.A2(n_15),
.B1(n_2),
.B2(n_3),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_105),
.A2(n_48),
.B1(n_37),
.B2(n_57),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_42),
.Y(n_106)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_106),
.Y(n_177)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_30),
.Y(n_107)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_107),
.Y(n_128)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_42),
.Y(n_108)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_108),
.Y(n_180)
);

INVx13_ASAP7_75t_L g109 ( 
.A(n_43),
.Y(n_109)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_40),
.Y(n_110)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_110),
.Y(n_184)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_22),
.Y(n_111)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_111),
.Y(n_186)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_29),
.Y(n_112)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_112),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_33),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_113),
.B(n_119),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_42),
.Y(n_114)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_114),
.Y(n_132)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_33),
.Y(n_115)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_115),
.Y(n_154)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_33),
.Y(n_116)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_116),
.Y(n_159)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_46),
.Y(n_117)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_117),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_46),
.Y(n_118)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_118),
.Y(n_176)
);

BUFx12f_ASAP7_75t_L g119 ( 
.A(n_46),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_25),
.B(n_1),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_120),
.B(n_57),
.Y(n_171)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_28),
.Y(n_121)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_121),
.Y(n_185)
);

AO22x1_ASAP7_75t_SL g131 ( 
.A1(n_74),
.A2(n_37),
.B1(n_55),
.B2(n_54),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_131),
.A2(n_133),
.B1(n_153),
.B2(n_162),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_73),
.A2(n_28),
.B1(n_41),
.B2(n_38),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_99),
.B(n_66),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_134),
.B(n_137),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_135),
.A2(n_174),
.B1(n_169),
.B2(n_187),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_70),
.B(n_25),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_103),
.B(n_50),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_139),
.B(n_4),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_84),
.B(n_31),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_141),
.B(n_1),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_109),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_146),
.B(n_171),
.Y(n_215)
);

HAxp5_ASAP7_75t_SL g147 ( 
.A(n_78),
.B(n_48),
.CON(n_147),
.SN(n_147)
);

CKINVDCx14_ASAP7_75t_R g244 ( 
.A(n_147),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_75),
.A2(n_28),
.B1(n_38),
.B2(n_52),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_59),
.A2(n_38),
.B1(n_52),
.B2(n_54),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_61),
.A2(n_52),
.B1(n_55),
.B2(n_47),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_165),
.B(n_51),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_108),
.A2(n_44),
.B1(n_31),
.B2(n_47),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_167),
.A2(n_173),
.B1(n_181),
.B2(n_195),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_60),
.A2(n_50),
.B1(n_26),
.B2(n_45),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_62),
.A2(n_26),
.B1(n_45),
.B2(n_44),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_65),
.A2(n_39),
.B1(n_32),
.B2(n_3),
.Y(n_181)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_117),
.Y(n_189)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_189),
.Y(n_202)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_68),
.Y(n_190)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_190),
.Y(n_211)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_69),
.Y(n_192)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_192),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_78),
.A2(n_39),
.B1(n_32),
.B2(n_4),
.Y(n_195)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_180),
.Y(n_200)
);

BUFx2_ASAP7_75t_L g270 ( 
.A(n_200),
.Y(n_270)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_179),
.Y(n_201)
);

BUFx2_ASAP7_75t_L g290 ( 
.A(n_201),
.Y(n_290)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_157),
.Y(n_203)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_203),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_204),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_205),
.A2(n_240),
.B1(n_265),
.B2(n_140),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_175),
.B(n_119),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_206),
.B(n_207),
.C(n_222),
.Y(n_278)
);

AND2x2_ASAP7_75t_SL g207 ( 
.A(n_125),
.B(n_118),
.Y(n_207)
);

BUFx4f_ASAP7_75t_SL g210 ( 
.A(n_191),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_210),
.Y(n_291)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_196),
.Y(n_212)
);

INVx3_ASAP7_75t_L g308 ( 
.A(n_212),
.Y(n_308)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_177),
.Y(n_213)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_213),
.Y(n_286)
);

CKINVDCx14_ASAP7_75t_R g306 ( 
.A(n_216),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_141),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_217),
.B(n_223),
.Y(n_266)
);

INVx5_ASAP7_75t_L g218 ( 
.A(n_122),
.Y(n_218)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_218),
.Y(n_289)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_132),
.Y(n_219)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_219),
.Y(n_295)
);

INVx6_ASAP7_75t_L g220 ( 
.A(n_138),
.Y(n_220)
);

INVx6_ASAP7_75t_L g281 ( 
.A(n_220),
.Y(n_281)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_176),
.Y(n_221)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_221),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_175),
.B(n_2),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_172),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_224),
.B(n_226),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_172),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_225),
.B(n_228),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_149),
.B(n_5),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_124),
.Y(n_227)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_227),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_178),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_127),
.Y(n_229)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_229),
.Y(n_273)
);

BUFx12_ASAP7_75t_L g231 ( 
.A(n_191),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g277 ( 
.A(n_231),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_128),
.B(n_5),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_232),
.B(n_245),
.Y(n_316)
);

BUFx2_ASAP7_75t_SL g233 ( 
.A(n_136),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_233),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_149),
.A2(n_79),
.B1(n_106),
.B2(n_97),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_234),
.A2(n_235),
.B1(n_264),
.B2(n_207),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_168),
.A2(n_71),
.B1(n_93),
.B2(n_86),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_195),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_236),
.B(n_241),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_168),
.B(n_5),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_237),
.B(n_247),
.Y(n_283)
);

AND2x2_ASAP7_75t_SL g238 ( 
.A(n_126),
.B(n_114),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_238),
.B(n_206),
.C(n_222),
.Y(n_311)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_185),
.Y(n_239)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_239),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_L g240 ( 
.A1(n_162),
.A2(n_85),
.B1(n_83),
.B2(n_82),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_178),
.Y(n_241)
);

AO22x2_ASAP7_75t_L g242 ( 
.A1(n_147),
.A2(n_81),
.B1(n_51),
.B2(n_10),
.Y(n_242)
);

AO21x2_ASAP7_75t_SL g279 ( 
.A1(n_242),
.A2(n_194),
.B(n_188),
.Y(n_279)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_154),
.Y(n_243)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_243),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_191),
.Y(n_245)
);

BUFx2_ASAP7_75t_L g246 ( 
.A(n_122),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g305 ( 
.A(n_246),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_131),
.B(n_8),
.Y(n_247)
);

BUFx12_ASAP7_75t_L g248 ( 
.A(n_142),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_248),
.Y(n_293)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_148),
.Y(n_249)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_249),
.Y(n_304)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_159),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_250),
.B(n_251),
.Y(n_288)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_150),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_184),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_252),
.Y(n_300)
);

BUFx2_ASAP7_75t_L g253 ( 
.A(n_140),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_253),
.Y(n_298)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_155),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_254),
.A2(n_256),
.B1(n_257),
.B2(n_259),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_167),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_255),
.B(n_258),
.Y(n_294)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_163),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_163),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_181),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_164),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_160),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_260),
.B(n_261),
.Y(n_309)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_130),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_151),
.B(n_9),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_262),
.B(n_263),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_151),
.B(n_9),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_153),
.A2(n_51),
.B1(n_11),
.B2(n_12),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_L g265 ( 
.A1(n_198),
.A2(n_51),
.B1(n_12),
.B2(n_13),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_267),
.A2(n_276),
.B1(n_257),
.B2(n_225),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_236),
.A2(n_133),
.B(n_156),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_268),
.A2(n_269),
.B(n_282),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_204),
.A2(n_161),
.B(n_129),
.Y(n_269)
);

OAI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_241),
.A2(n_205),
.B1(n_209),
.B2(n_230),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_271),
.A2(n_314),
.B1(n_289),
.B2(n_273),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_272),
.A2(n_296),
.B1(n_310),
.B2(n_312),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_L g276 ( 
.A1(n_206),
.A2(n_197),
.B1(n_170),
.B2(n_199),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_279),
.A2(n_253),
.B1(n_246),
.B2(n_218),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_244),
.A2(n_186),
.B(n_123),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_208),
.B(n_144),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_287),
.B(n_260),
.Y(n_329)
);

AND2x2_ASAP7_75t_SL g292 ( 
.A(n_242),
.B(n_123),
.Y(n_292)
);

CKINVDCx14_ASAP7_75t_R g322 ( 
.A(n_292),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_242),
.A2(n_238),
.B1(n_207),
.B2(n_145),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_242),
.A2(n_183),
.B1(n_166),
.B2(n_138),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_311),
.B(n_256),
.Y(n_336)
);

OA21x2_ASAP7_75t_L g312 ( 
.A1(n_238),
.A2(n_193),
.B(n_182),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_249),
.A2(n_152),
.B1(n_183),
.B2(n_143),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_314),
.A2(n_220),
.B1(n_219),
.B2(n_221),
.Y(n_325)
);

O2A1O1Ixp33_ASAP7_75t_L g315 ( 
.A1(n_222),
.A2(n_158),
.B(n_143),
.C(n_166),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_315),
.A2(n_210),
.B(n_231),
.Y(n_341)
);

OAI32xp33_ASAP7_75t_L g318 ( 
.A1(n_292),
.A2(n_215),
.A3(n_261),
.B1(n_252),
.B2(n_201),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_318),
.B(n_324),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_319),
.A2(n_323),
.B1(n_328),
.B2(n_335),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_316),
.B(n_202),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g387 ( 
.A(n_320),
.B(n_334),
.Y(n_387)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_309),
.Y(n_321)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_321),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_287),
.B(n_216),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_325),
.B(n_341),
.Y(n_375)
);

CKINVDCx16_ASAP7_75t_R g326 ( 
.A(n_282),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_326),
.B(n_327),
.Y(n_361)
);

CKINVDCx14_ASAP7_75t_R g327 ( 
.A(n_288),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_279),
.A2(n_203),
.B1(n_213),
.B2(n_259),
.Y(n_328)
);

XNOR2x1_ASAP7_75t_L g379 ( 
.A(n_329),
.B(n_302),
.Y(n_379)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_291),
.Y(n_330)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_330),
.Y(n_369)
);

BUFx24_ASAP7_75t_L g331 ( 
.A(n_291),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g378 ( 
.A(n_331),
.Y(n_378)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_300),
.Y(n_332)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_332),
.Y(n_366)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_309),
.Y(n_333)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_333),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_266),
.B(n_211),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_279),
.A2(n_214),
.B1(n_200),
.B2(n_212),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_336),
.B(n_304),
.C(n_285),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_283),
.B(n_10),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_337),
.B(n_338),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_279),
.A2(n_210),
.B1(n_231),
.B2(n_51),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_280),
.B(n_10),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_340),
.B(n_342),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_267),
.A2(n_12),
.B1(n_248),
.B2(n_294),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_295),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_343),
.B(n_344),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_307),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_280),
.B(n_248),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_345),
.B(n_351),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_296),
.A2(n_292),
.B1(n_294),
.B2(n_301),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_346),
.A2(n_347),
.B1(n_348),
.B2(n_349),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_301),
.A2(n_269),
.B1(n_268),
.B2(n_311),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_278),
.A2(n_303),
.B1(n_312),
.B2(n_274),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_312),
.A2(n_278),
.B1(n_315),
.B2(n_306),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_350),
.A2(n_354),
.B1(n_325),
.B2(n_317),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_273),
.B(n_299),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_299),
.B(n_275),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_352),
.Y(n_376)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_295),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_353),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_275),
.A2(n_313),
.B1(n_289),
.B2(n_281),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_308),
.B(n_270),
.Y(n_355)
);

CKINVDCx16_ASAP7_75t_R g381 ( 
.A(n_355),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_356),
.A2(n_341),
.B1(n_330),
.B2(n_331),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_SL g357 ( 
.A1(n_326),
.A2(n_293),
.B(n_284),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g399 ( 
.A1(n_357),
.A2(n_358),
.B(n_360),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_339),
.A2(n_297),
.B(n_290),
.Y(n_358)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_339),
.A2(n_290),
.B(n_270),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_347),
.B(n_329),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_362),
.B(n_379),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_317),
.A2(n_281),
.B1(n_298),
.B2(n_308),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_368),
.A2(n_370),
.B1(n_384),
.B2(n_319),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_346),
.A2(n_302),
.B1(n_304),
.B2(n_286),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_351),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_380),
.B(n_321),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_382),
.B(n_385),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_SL g383 ( 
.A1(n_322),
.A2(n_285),
.B(n_286),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_L g404 ( 
.A1(n_383),
.A2(n_355),
.B(n_343),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_350),
.A2(n_300),
.B1(n_305),
.B2(n_277),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_336),
.B(n_277),
.C(n_305),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_324),
.B(n_345),
.Y(n_386)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_386),
.B(n_340),
.Y(n_395)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_388),
.Y(n_421)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_389),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_356),
.A2(n_342),
.B1(n_328),
.B2(n_335),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_390),
.B(n_393),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_365),
.A2(n_349),
.B1(n_333),
.B2(n_318),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_391),
.A2(n_408),
.B1(n_409),
.B2(n_411),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_374),
.A2(n_323),
.B1(n_338),
.B2(n_348),
.Y(n_393)
);

OAI21xp5_ASAP7_75t_SL g417 ( 
.A1(n_394),
.A2(n_406),
.B(n_413),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_SL g425 ( 
.A(n_395),
.B(n_379),
.Y(n_425)
);

INVx2_ASAP7_75t_SL g396 ( 
.A(n_366),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_396),
.B(n_401),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g397 ( 
.A1(n_373),
.A2(n_337),
.B1(n_352),
.B2(n_354),
.Y(n_397)
);

AOI22xp33_ASAP7_75t_L g432 ( 
.A1(n_397),
.A2(n_407),
.B1(n_381),
.B2(n_376),
.Y(n_432)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_359),
.Y(n_398)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_398),
.Y(n_424)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_359),
.Y(n_400)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_400),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_378),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_377),
.Y(n_402)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_402),
.Y(n_438)
);

INVxp33_ASAP7_75t_SL g403 ( 
.A(n_371),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_403),
.B(n_405),
.Y(n_427)
);

AOI21xp5_ASAP7_75t_SL g418 ( 
.A1(n_404),
.A2(n_357),
.B(n_361),
.Y(n_418)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_377),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_375),
.B(n_353),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_366),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_365),
.A2(n_331),
.B1(n_332),
.B2(n_373),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_367),
.A2(n_331),
.B1(n_361),
.B2(n_374),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_378),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_410),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_375),
.A2(n_368),
.B1(n_367),
.B2(n_384),
.Y(n_411)
);

OA22x2_ASAP7_75t_L g413 ( 
.A1(n_380),
.A2(n_375),
.B1(n_364),
.B2(n_383),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_375),
.A2(n_362),
.B1(n_370),
.B2(n_381),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_SL g426 ( 
.A1(n_414),
.A2(n_360),
.B(n_358),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_SL g458 ( 
.A1(n_418),
.A2(n_435),
.B(n_363),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_392),
.B(n_386),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_419),
.B(n_423),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_391),
.B(n_387),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_420),
.B(n_426),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_392),
.B(n_379),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_SL g443 ( 
.A(n_425),
.B(n_409),
.Y(n_443)
);

CKINVDCx16_ASAP7_75t_R g428 ( 
.A(n_406),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_428),
.B(n_429),
.Y(n_450)
);

CKINVDCx16_ASAP7_75t_R g429 ( 
.A(n_406),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_412),
.B(n_372),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_430),
.B(n_434),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_412),
.B(n_385),
.C(n_382),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_431),
.B(n_393),
.C(n_399),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_L g446 ( 
.A1(n_432),
.A2(n_411),
.B1(n_388),
.B2(n_394),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_395),
.B(n_372),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_SL g435 ( 
.A(n_395),
.B(n_371),
.C(n_387),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_430),
.B(n_414),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_439),
.B(n_445),
.Y(n_467)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_427),
.Y(n_441)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_441),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_SL g460 ( 
.A(n_443),
.B(n_425),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_444),
.B(n_437),
.C(n_421),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_431),
.B(n_408),
.Y(n_445)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_446),
.Y(n_470)
);

AND2x2_ASAP7_75t_L g447 ( 
.A(n_416),
.B(n_404),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_447),
.B(n_452),
.Y(n_459)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_427),
.Y(n_448)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_448),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_419),
.B(n_399),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_451),
.B(n_456),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_421),
.A2(n_389),
.B1(n_413),
.B2(n_400),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_422),
.B(n_402),
.Y(n_453)
);

NOR2xp67_ASAP7_75t_SL g474 ( 
.A(n_453),
.B(n_455),
.Y(n_474)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_424),
.Y(n_454)
);

INVx3_ASAP7_75t_L g472 ( 
.A(n_454),
.Y(n_472)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_424),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_423),
.B(n_398),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_436),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_457),
.B(n_458),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_SL g484 ( 
.A(n_460),
.B(n_443),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_440),
.B(n_426),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_462),
.B(n_463),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_SL g463 ( 
.A1(n_444),
.A2(n_418),
.B(n_416),
.Y(n_463)
);

FAx1_ASAP7_75t_SL g464 ( 
.A(n_442),
.B(n_434),
.CI(n_435),
.CON(n_464),
.SN(n_464)
);

AOI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_464),
.A2(n_447),
.B1(n_451),
.B2(n_450),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_440),
.B(n_417),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_465),
.B(n_468),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_445),
.B(n_417),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_471),
.B(n_467),
.C(n_439),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_475),
.B(n_483),
.C(n_485),
.Y(n_487)
);

AOI21xp5_ASAP7_75t_L g493 ( 
.A1(n_476),
.A2(n_482),
.B(n_461),
.Y(n_493)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_472),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_477),
.B(n_478),
.Y(n_494)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_472),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_474),
.Y(n_479)
);

OR2x2_ASAP7_75t_L g488 ( 
.A(n_479),
.B(n_480),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_467),
.B(n_449),
.C(n_456),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_462),
.B(n_449),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_484),
.B(n_486),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_465),
.B(n_452),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_466),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_475),
.B(n_471),
.C(n_470),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_489),
.B(n_490),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_481),
.B(n_469),
.C(n_468),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_480),
.B(n_485),
.C(n_483),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_491),
.B(n_461),
.C(n_469),
.Y(n_498)
);

AOI22xp33_ASAP7_75t_SL g492 ( 
.A1(n_484),
.A2(n_473),
.B1(n_459),
.B2(n_415),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_SL g504 ( 
.A1(n_492),
.A2(n_410),
.B1(n_390),
.B2(n_396),
.Y(n_504)
);

OAI21x1_ASAP7_75t_L g499 ( 
.A1(n_493),
.A2(n_413),
.B(n_458),
.Y(n_499)
);

OAI21xp5_ASAP7_75t_SL g496 ( 
.A1(n_479),
.A2(n_447),
.B(n_464),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g503 ( 
.A(n_496),
.B(n_460),
.Y(n_503)
);

AOI22xp5_ASAP7_75t_L g497 ( 
.A1(n_494),
.A2(n_415),
.B1(n_433),
.B2(n_405),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_497),
.B(n_503),
.Y(n_507)
);

OR2x2_ASAP7_75t_L g506 ( 
.A(n_498),
.B(n_501),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_499),
.B(n_500),
.Y(n_510)
);

O2A1O1Ixp33_ASAP7_75t_L g500 ( 
.A1(n_492),
.A2(n_413),
.B(n_437),
.C(n_438),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_488),
.A2(n_438),
.B1(n_436),
.B2(n_401),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_504),
.B(n_495),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_502),
.B(n_487),
.C(n_495),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_505),
.B(n_508),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_SL g509 ( 
.A(n_498),
.B(n_364),
.Y(n_509)
);

AOI21xp5_ASAP7_75t_L g514 ( 
.A1(n_509),
.A2(n_363),
.B(n_407),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_L g512 ( 
.A(n_507),
.B(n_503),
.Y(n_512)
);

OR2x2_ASAP7_75t_L g516 ( 
.A(n_512),
.B(n_510),
.Y(n_516)
);

AOI21xp5_ASAP7_75t_L g513 ( 
.A1(n_506),
.A2(n_501),
.B(n_500),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_513),
.B(n_514),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_516),
.B(n_511),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_517),
.Y(n_518)
);

OAI21xp5_ASAP7_75t_L g519 ( 
.A1(n_518),
.A2(n_515),
.B(n_508),
.Y(n_519)
);

NOR2xp67_ASAP7_75t_L g520 ( 
.A(n_519),
.B(n_396),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_520),
.B(n_369),
.Y(n_521)
);


endmodule