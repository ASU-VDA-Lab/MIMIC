module real_jpeg_27707_n_17 (n_8, n_0, n_2, n_338, n_10, n_9, n_12, n_6, n_337, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_17);

input n_8;
input n_0;
input n_2;
input n_338;
input n_10;
input n_9;
input n_12;
input n_6;
input n_337;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_332;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx5_ASAP7_75t_L g82 ( 
.A(n_0),
.Y(n_82)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_0),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_1),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_L g26 ( 
.A1(n_1),
.A2(n_22),
.B1(n_27),
.B2(n_28),
.Y(n_26)
);

O2A1O1Ixp33_ASAP7_75t_SL g169 ( 
.A1(n_1),
.A2(n_10),
.B(n_28),
.C(n_170),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_3),
.A2(n_53),
.B1(n_55),
.B2(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_3),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_3),
.A2(n_49),
.B1(n_50),
.B2(n_64),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_3),
.A2(n_23),
.B1(n_24),
.B2(n_64),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_3),
.A2(n_27),
.B1(n_28),
.B2(n_64),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_4),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_4),
.A2(n_30),
.B1(n_49),
.B2(n_50),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_4),
.A2(n_30),
.B1(n_53),
.B2(n_55),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g312 ( 
.A1(n_4),
.A2(n_23),
.B1(n_24),
.B2(n_30),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_5),
.A2(n_53),
.B1(n_55),
.B2(n_77),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_5),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_5),
.A2(n_49),
.B1(n_50),
.B2(n_77),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_5),
.A2(n_23),
.B1(n_24),
.B2(n_77),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_5),
.A2(n_27),
.B1(n_28),
.B2(n_77),
.Y(n_201)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_7),
.A2(n_49),
.B1(n_50),
.B2(n_168),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_7),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g227 ( 
.A1(n_7),
.A2(n_53),
.B1(n_55),
.B2(n_168),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_7),
.A2(n_23),
.B1(n_24),
.B2(n_168),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g307 ( 
.A1(n_7),
.A2(n_27),
.B1(n_28),
.B2(n_168),
.Y(n_307)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_8),
.A2(n_49),
.B1(n_50),
.B2(n_151),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_8),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_8),
.A2(n_53),
.B1(n_55),
.B2(n_151),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_8),
.A2(n_23),
.B1(n_24),
.B2(n_151),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_8),
.A2(n_27),
.B1(n_28),
.B2(n_151),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_9),
.A2(n_27),
.B1(n_28),
.B2(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_9),
.A2(n_34),
.B1(n_49),
.B2(n_50),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_9),
.A2(n_34),
.B1(n_53),
.B2(n_55),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_9),
.A2(n_23),
.B1(n_24),
.B2(n_34),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_10),
.B(n_55),
.Y(n_54)
);

A2O1A1O1Ixp25_ASAP7_75t_L g58 ( 
.A1(n_10),
.A2(n_54),
.B(n_55),
.C(n_59),
.D(n_62),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_10),
.B(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_10),
.Y(n_103)
);

OAI21xp33_ASAP7_75t_L g108 ( 
.A1(n_10),
.A2(n_81),
.B(n_85),
.Y(n_108)
);

A2O1A1O1Ixp25_ASAP7_75t_L g118 ( 
.A1(n_10),
.A2(n_24),
.B(n_119),
.C(n_120),
.D(n_122),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_10),
.B(n_24),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_10),
.B(n_21),
.Y(n_147)
);

OAI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_10),
.A2(n_27),
.B1(n_28),
.B2(n_103),
.Y(n_175)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

O2A1O1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_11),
.A2(n_55),
.B(n_60),
.C(n_61),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_11),
.A2(n_49),
.B1(n_50),
.B2(n_52),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_12),
.A2(n_49),
.B1(n_50),
.B2(n_84),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_12),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_12),
.A2(n_53),
.B1(n_55),
.B2(n_84),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_12),
.A2(n_23),
.B1(n_24),
.B2(n_84),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_12),
.A2(n_27),
.B1(n_28),
.B2(n_84),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_13),
.A2(n_49),
.B1(n_50),
.B2(n_132),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_13),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_13),
.A2(n_53),
.B1(n_55),
.B2(n_132),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_13),
.A2(n_23),
.B1(n_24),
.B2(n_132),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_13),
.A2(n_27),
.B1(n_28),
.B2(n_132),
.Y(n_270)
);

BUFx24_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_15),
.Y(n_71)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_15),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_15),
.A2(n_23),
.B1(n_24),
.B2(n_73),
.Y(n_121)
);

INVx11_ASAP7_75t_SL g51 ( 
.A(n_16),
.Y(n_51)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_37),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_35),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_31),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_20),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_25),
.B(n_29),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_21),
.B(n_26),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_21),
.A2(n_25),
.B1(n_29),
.B2(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_21),
.B(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_21),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_21),
.A2(n_25),
.B1(n_201),
.B2(n_219),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_21),
.A2(n_25),
.B1(n_33),
.B2(n_328),
.Y(n_327)
);

OAI21xp33_ASAP7_75t_L g170 ( 
.A1(n_22),
.A2(n_24),
.B(n_103),
.Y(n_170)
);

INVx5_ASAP7_75t_SL g24 ( 
.A(n_23),
.Y(n_24)
);

AOI32xp33_ASAP7_75t_L g133 ( 
.A1(n_23),
.A2(n_55),
.A3(n_119),
.B1(n_134),
.B2(n_135),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_25),
.A2(n_175),
.B(n_176),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_25),
.B(n_178),
.Y(n_203)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_25),
.Y(n_242)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_27),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_32),
.B(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_32),
.B(n_334),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_32),
.B(n_334),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_SL g37 ( 
.A1(n_38),
.A2(n_333),
.B(n_335),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_321),
.B(n_332),
.Y(n_38)
);

OAI321xp33_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_285),
.A3(n_314),
.B1(n_319),
.B2(n_320),
.C(n_337),
.Y(n_39)
);

AOI321xp33_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_235),
.A3(n_274),
.B1(n_279),
.B2(n_284),
.C(n_338),
.Y(n_40)
);

NOR3xp33_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_188),
.C(n_231),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_159),
.B(n_187),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_SL g43 ( 
.A1(n_44),
.A2(n_137),
.B(n_158),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_114),
.B(n_136),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_SL g45 ( 
.A1(n_46),
.A2(n_90),
.B(n_113),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_66),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_47),
.B(n_66),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_58),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_48),
.B(n_58),
.Y(n_99)
);

AOI32xp33_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_52),
.A3(n_53),
.B1(n_54),
.B2(n_56),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_49),
.B(n_110),
.Y(n_109)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_50),
.B(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_50),
.B(n_82),
.Y(n_81)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_52),
.Y(n_57)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_53),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_53),
.A2(n_55),
.B1(n_71),
.B2(n_72),
.Y(n_70)
);

NAND2xp33_ASAP7_75t_SL g135 ( 
.A(n_53),
.B(n_72),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_55),
.B(n_57),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_59),
.B(n_79),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_59),
.A2(n_61),
.B1(n_126),
.B2(n_127),
.Y(n_125)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_59),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_59),
.A2(n_61),
.B1(n_250),
.B2(n_251),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_59),
.A2(n_61),
.B1(n_251),
.B2(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_62),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_65),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g75 ( 
.A1(n_65),
.A2(n_76),
.B(n_78),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_65),
.B(n_103),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_65),
.A2(n_78),
.B(n_186),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_65),
.A2(n_155),
.B1(n_186),
.B2(n_210),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_65),
.A2(n_155),
.B1(n_210),
.B2(n_227),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_65),
.A2(n_155),
.B(n_260),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_80),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_69),
.B1(n_74),
.B2(n_75),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_68),
.B(n_75),
.C(n_80),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_70),
.B(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_70),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_70),
.A2(n_120),
.B1(n_182),
.B2(n_183),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_70),
.A2(n_120),
.B1(n_262),
.B2(n_263),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_70),
.A2(n_120),
.B1(n_263),
.B2(n_292),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_70),
.A2(n_120),
.B(n_326),
.Y(n_325)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_72),
.Y(n_134)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_76),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_83),
.B(n_85),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_81),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_81),
.B(n_87),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_81),
.A2(n_98),
.B1(n_131),
.B2(n_150),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_81),
.A2(n_89),
.B1(n_207),
.B2(n_208),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_81),
.A2(n_98),
.B1(n_208),
.B2(n_225),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_81),
.A2(n_98),
.B(n_225),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_83),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_86),
.B(n_88),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_88),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_88),
.A2(n_95),
.B1(n_166),
.B2(n_167),
.Y(n_165)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_103),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_100),
.B(n_112),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_99),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_92),
.B(n_99),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_93),
.A2(n_95),
.B1(n_96),
.B2(n_97),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_94),
.A2(n_98),
.B(n_105),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_97),
.A2(n_106),
.B(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_101),
.A2(n_107),
.B(n_111),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_104),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_102),
.B(n_104),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_108),
.B(n_109),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_116),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_115),
.B(n_116),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_128),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_125),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_125),
.C(n_128),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_120),
.B(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_120),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_122),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_124),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_123),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_124),
.A2(n_142),
.B(n_143),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_124),
.A2(n_143),
.B(n_222),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_124),
.A2(n_196),
.B1(n_222),
.B2(n_245),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_124),
.A2(n_196),
.B1(n_311),
.B2(n_312),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_127),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g128 ( 
.A(n_129),
.B(n_133),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_133),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_139),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_138),
.B(n_139),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_152),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_140),
.B(n_153),
.C(n_154),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_141),
.B(n_145),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_141),
.B(n_146),
.C(n_149),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_142),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_147),
.B1(n_148),
.B2(n_149),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_150),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_154),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_156),
.B(n_157),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_161),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_160),
.B(n_161),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_173),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_163),
.B(n_164),
.C(n_173),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_165),
.A2(n_169),
.B1(n_171),
.B2(n_172),
.Y(n_164)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_165),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_167),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_169),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_169),
.B(n_171),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_174),
.B(n_179),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_174),
.B(n_181),
.C(n_184),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_177),
.A2(n_242),
.B(n_243),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_181),
.B1(n_184),
.B2(n_185),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_183),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_189),
.A2(n_281),
.B(n_282),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_212),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_190),
.B(n_212),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_205),
.C(n_211),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_191),
.B(n_234),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_192),
.B(n_194),
.C(n_204),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_195),
.B1(n_199),
.B2(n_204),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_195),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_196),
.A2(n_197),
.B(n_198),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_199),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_202),
.B(n_203),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_201),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_202),
.A2(n_203),
.B(n_270),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_202),
.A2(n_242),
.B1(n_270),
.B2(n_297),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_202),
.A2(n_242),
.B1(n_297),
.B2(n_307),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_205),
.B(n_211),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_209),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_206),
.B(n_209),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_213),
.A2(n_228),
.B1(n_229),
.B2(n_230),
.Y(n_212)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_213),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_214),
.B(n_223),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_214),
.B(n_223),
.C(n_230),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_SL g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_215),
.B(n_218),
.C(n_220),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_218),
.B1(n_220),
.B2(n_221),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_219),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_221),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_226),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_224),
.B(n_226),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_227),
.Y(n_250)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_228),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_232),
.B(n_233),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_255),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_236),
.B(n_255),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_247),
.C(n_254),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_237),
.B(n_247),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_239),
.B1(n_240),
.B2(n_246),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_238),
.Y(n_246)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_SL g240 ( 
.A(n_241),
.B(n_244),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_241),
.B(n_244),
.C(n_246),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_245),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_248),
.A2(n_249),
.B1(n_252),
.B2(n_253),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_248),
.B(n_253),
.Y(n_271)
);

CKINVDCx14_ASAP7_75t_R g248 ( 
.A(n_249),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_252),
.A2(n_253),
.B1(n_268),
.B2(n_269),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_253),
.Y(n_252)
);

AOI21xp33_ASAP7_75t_L g301 ( 
.A1(n_253),
.A2(n_268),
.B(n_271),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_254),
.B(n_278),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_273),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_265),
.B1(n_266),
.B2(n_272),
.Y(n_256)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_257),
.Y(n_272)
);

OAI21xp33_ASAP7_75t_L g257 ( 
.A1(n_258),
.A2(n_261),
.B(n_264),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_258),
.B(n_261),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_260),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_264),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_264),
.A2(n_287),
.B1(n_288),
.B2(n_299),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_265),
.B(n_272),
.C(n_273),
.Y(n_315)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_271),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_275),
.A2(n_280),
.B(n_283),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_276),
.B(n_277),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_302),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_286),
.B(n_302),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_299),
.C(n_300),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_289),
.A2(n_290),
.B1(n_296),
.B2(n_298),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_291),
.A2(n_293),
.B1(n_294),
.B2(n_295),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_291),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_291),
.B(n_295),
.C(n_296),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_292),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_293),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_293),
.A2(n_295),
.B1(n_309),
.B2(n_310),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_295),
.B(n_306),
.C(n_310),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_296),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_296),
.A2(n_298),
.B1(n_304),
.B2(n_305),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_296),
.B(n_305),
.C(n_313),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_300),
.A2(n_301),
.B1(n_317),
.B2(n_318),
.Y(n_316)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_313),
.Y(n_302)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_308),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_307),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_310),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_312),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_315),
.B(n_316),
.Y(n_319)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_322),
.B(n_323),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_322),
.B(n_323),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_331),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_325),
.A2(n_327),
.B1(n_329),
.B2(n_330),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_325),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_327),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_327),
.B(n_330),
.C(n_331),
.Y(n_334)
);


endmodule