module real_aes_9897_n_376 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_374, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_376);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_374;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_376;
wire n_2043;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_2003;
wire n_2014;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_1797;
wire n_933;
wire n_485;
wire n_822;
wire n_1641;
wire n_750;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_1903;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1929;
wire n_1737;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_1888;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_1972;
wire n_593;
wire n_2029;
wire n_989;
wire n_431;
wire n_1044;
wire n_1730;
wire n_1744;
wire n_963;
wire n_2006;
wire n_551;
wire n_884;
wire n_2035;
wire n_814;
wire n_944;
wire n_1936;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1873;
wire n_1835;
wire n_1871;
wire n_1468;
wire n_1713;
wire n_1967;
wire n_1920;
wire n_870;
wire n_1248;
wire n_2021;
wire n_1602;
wire n_548;
wire n_1859;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1845;
wire n_1415;
wire n_2031;
wire n_1160;
wire n_1849;
wire n_2040;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1805;
wire n_1367;
wire n_744;
wire n_1994;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_2049;
wire n_1833;
wire n_1477;
wire n_1944;
wire n_595;
wire n_1893;
wire n_1960;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_2016;
wire n_962;
wire n_1599;
wire n_1959;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_1809;
wire n_682;
wire n_1745;
wire n_1820;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_1883;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_2022;
wire n_885;
wire n_950;
wire n_381;
wire n_1981;
wire n_1196;
wire n_1013;
wire n_1905;
wire n_808;
wire n_1639;
wire n_1224;
wire n_1694;
wire n_1872;
wire n_688;
wire n_1042;
wire n_1588;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_527;
wire n_1676;
wire n_1342;
wire n_2018;
wire n_1440;
wire n_1966;
wire n_552;
wire n_1346;
wire n_1383;
wire n_1890;
wire n_1675;
wire n_1954;
wire n_590;
wire n_1293;
wire n_1880;
wire n_432;
wire n_1882;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_1865;
wire n_1600;
wire n_805;
wire n_619;
wire n_1284;
wire n_1250;
wire n_1095;
wire n_1583;
wire n_1987;
wire n_859;
wire n_1465;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_1658;
wire n_1866;
wire n_954;
wire n_702;
wire n_1874;
wire n_1007;
wire n_1906;
wire n_898;
wire n_1926;
wire n_562;
wire n_1897;
wire n_1022;
wire n_1502;
wire n_1073;
wire n_404;
wire n_1632;
wire n_1301;
wire n_728;
wire n_1201;
wire n_2004;
wire n_997;
wire n_2000;
wire n_1105;
wire n_1768;
wire n_1243;
wire n_1846;
wire n_1003;
wire n_749;
wire n_1870;
wire n_914;
wire n_1837;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_1351;
wire n_972;
wire n_1813;
wire n_1978;
wire n_1628;
wire n_1587;
wire n_1821;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1825;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_2024;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1956;
wire n_1048;
wire n_1422;
wire n_787;
wire n_2038;
wire n_1214;
wire n_806;
wire n_715;
wire n_1714;
wire n_1940;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_1814;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1510;
wire n_1495;
wire n_1727;
wire n_712;
wire n_1921;
wire n_2041;
wire n_422;
wire n_861;
wire n_2007;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_724;
wire n_1648;
wire n_1914;
wire n_440;
wire n_1945;
wire n_1231;
wire n_2058;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_1793;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_1538;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_1787;
wire n_877;
wire n_424;
wire n_802;
wire n_1876;
wire n_2057;
wire n_1488;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1999;
wire n_1652;
wire n_684;
wire n_2050;
wire n_1178;
wire n_1979;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1828;
wire n_1860;
wire n_2012;
wire n_1018;
wire n_1563;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_1973;
wire n_635;
wire n_792;
wire n_1542;
wire n_1392;
wire n_665;
wire n_991;
wire n_667;
wire n_1712;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_1951;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_1260;
wire n_1606;
wire n_1129;
wire n_1760;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_1852;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1830;
wire n_1594;
wire n_2020;
wire n_1864;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1991;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_948;
wire n_399;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1839;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_1881;
wire n_1568;
wire n_1368;
wire n_994;
wire n_2059;
wire n_384;
wire n_1612;
wire n_1479;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1884;
wire n_1182;
wire n_872;
wire n_1401;
wire n_2045;
wire n_2017;
wire n_1946;
wire n_1086;
wire n_1189;
wire n_1070;
wire n_2036;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1741;
wire n_1456;
wire n_1879;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_1853;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_2009;
wire n_925;
wire n_1389;
wire n_1393;
wire n_1977;
wire n_1930;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_2005;
wire n_508;
wire n_1141;
wire n_2033;
wire n_1985;
wire n_1769;
wire n_1812;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_1971;
wire n_600;
wire n_964;
wire n_731;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_1854;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_658;
wire n_676;
wire n_1856;
wire n_531;
wire n_1848;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_1569;
wire n_895;
wire n_799;
wire n_490;
wire n_391;
wire n_1993;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_1145;
wire n_645;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_777;
wire n_985;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_2039;
wire n_2002;
wire n_734;
wire n_1623;
wire n_1907;
wire n_735;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_1857;
wire n_1984;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_1234;
wire n_1915;
wire n_622;
wire n_1634;
wire n_1353;
wire n_1002;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_1862;
wire n_1965;
wire n_850;
wire n_720;
wire n_2023;
wire n_1026;
wire n_1756;
wire n_1803;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_1699;
wire n_1794;
wire n_1748;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_1970;
wire n_526;
wire n_1513;
wire n_2015;
wire n_1983;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_1934;
wire n_809;
wire n_1532;
wire n_679;
wire n_520;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1784;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_1431;
wire n_721;
wire n_1806;
wire n_1829;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_1976;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1807;
wire n_459;
wire n_1172;
wire n_1689;
wire n_998;
wire n_1625;
wire n_1910;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1957;
wire n_1184;
wire n_583;
wire n_1998;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_2052;
wire n_1961;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_1904;
wire n_450;
wire n_1578;
wire n_1779;
wire n_473;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1908;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_1840;
wire n_968;
wire n_710;
wire n_1040;
wire n_1185;
wire n_661;
wire n_1102;
wire n_447;
wire n_1795;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_1788;
wire n_1938;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_2019;
wire n_869;
wire n_1816;
wire n_1952;
wire n_1811;
wire n_2042;
wire n_1066;
wire n_2046;
wire n_1917;
wire n_1377;
wire n_800;
wire n_1175;
wire n_1170;
wire n_778;
wire n_522;
wire n_1475;
wire n_1928;
wire n_977;
wire n_943;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1995;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_1980;
wire n_2013;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1932;
wire n_1707;
wire n_856;
wire n_594;
wire n_1146;
wire n_1685;
wire n_1810;
wire n_1435;
wire n_1800;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_1990;
wire n_427;
wire n_1540;
wire n_519;
wire n_1878;
wire n_1116;
wire n_709;
wire n_1834;
wire n_388;
wire n_1913;
wire n_1470;
wire n_816;
wire n_1899;
wire n_625;
wire n_953;
wire n_1565;
wire n_1953;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_584;
wire n_896;
wire n_1817;
wire n_2008;
wire n_1722;
wire n_528;
wire n_1638;
wire n_495;
wire n_1072;
wire n_1078;
wire n_1663;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1923;
wire n_2025;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1850;
wire n_1332;
wire n_1927;
wire n_1263;
wire n_1411;
wire n_1922;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1726;
wire n_1827;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1949;
wire n_1029;
wire n_1989;
wire n_1207;
wire n_1555;
wire n_1962;
wire n_664;
wire n_1017;
wire n_1942;
wire n_581;
wire n_2048;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_1608;
wire n_1167;
wire n_1939;
wire n_1327;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1792;
wire n_1006;
wire n_1869;
wire n_1259;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1414;
wire n_1241;
wire n_1671;
wire n_502;
wire n_434;
wire n_769;
wire n_1455;
wire n_1212;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1895;
wire n_1670;
wire n_1941;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_1986;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_632;
wire n_1344;
wire n_1603;
wire n_1450;
wire n_1720;
wire n_1331;
wire n_714;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_1948;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1886;
wire n_2032;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_1832;
wire n_727;
wire n_1083;
wire n_397;
wire n_1605;
wire n_1056;
wire n_1592;
wire n_1802;
wire n_1855;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1785;
wire n_1774;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1798;
wire n_1038;
wire n_1085;
wire n_2027;
wire n_845;
wire n_1838;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_1863;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_2053;
wire n_826;
wire n_628;
wire n_487;
wire n_831;
wire n_1772;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_2034;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_2028;
wire n_1693;
wire n_1791;
wire n_418;
wire n_771;
wire n_524;
wire n_1496;
wire n_1378;
wire n_1191;
wire n_705;
wire n_1206;
wire n_1824;
wire n_1933;
wire n_1270;
wire n_1988;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_1761;
wire n_863;
wire n_1226;
wire n_525;
wire n_1617;
wire n_1790;
wire n_644;
wire n_1150;
wire n_1861;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_929;
wire n_1143;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_1343;
wire n_719;
wire n_465;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_2011;
wire n_1757;
wire n_2055;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1799;
wire n_640;
wire n_1176;
wire n_1691;
wire n_1721;
wire n_1931;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1804;
wire n_1480;
wire n_1101;
wire n_1251;
wire n_1076;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_1964;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1844;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1937;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_1841;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_1596;
wire n_987;
wire n_2037;
wire n_1982;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_1822;
wire n_2030;
wire n_718;
wire n_1955;
wire n_669;
wire n_1091;
wire n_423;
wire n_1969;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_1777;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1819;
wire n_1887;
wire n_1674;
wire n_491;
wire n_1294;
wire n_1902;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_1889;
wire n_2044;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_1896;
wire n_767;
wire n_889;
wire n_1398;
wire n_1911;
wire n_379;
wire n_1847;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1912;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_1919;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1541;
wire n_1272;
wire n_408;
wire n_1754;
wire n_578;
wire n_892;
wire n_938;
wire n_774;
wire n_466;
wire n_1049;
wire n_559;
wire n_1277;
wire n_1584;
wire n_1950;
wire n_984;
wire n_726;
wire n_517;
wire n_931;
wire n_780;
wire n_1851;
wire n_530;
wire n_2047;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_1916;
wire n_532;
wire n_1025;
wire n_1875;
wire n_1826;
wire n_1836;
wire n_1909;
wire n_924;
wire n_1264;
wire n_1858;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1901;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1943;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1318;
wire n_1290;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_1818;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1974;
wire n_1547;
wire n_1823;
wire n_1867;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1891;
wire n_1267;
wire n_790;
wire n_1262;
wire n_1843;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1885;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1416;
wire n_1249;
wire n_387;
wire n_1239;
wire n_2056;
wire n_1796;
wire n_1662;
wire n_1992;
wire n_1963;
wire n_1958;
wire n_969;
wire n_1535;
wire n_2010;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1925;
wire n_1801;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_1968;
wire n_430;
wire n_1252;
wire n_1647;
wire n_1132;
wire n_1947;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_1996;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_2001;
wire n_965;
wire n_1894;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1808;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_1481;
wire n_1430;
wire n_907;
wire n_1758;
wire n_1005;
wire n_2051;
wire n_1312;
wire n_1697;
wire n_1877;
wire n_1900;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1842;
wire n_1536;
wire n_1746;
wire n_1898;
wire n_1711;
wire n_482;
wire n_633;
wire n_1892;
wire n_971;
wire n_1052;
wire n_1071;
wire n_2026;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_1573;
wire n_1130;
wire n_1918;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_1831;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_1300;
wire n_575;
wire n_1372;
wire n_698;
wire n_1997;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1815;
wire n_1924;
wire n_1412;
wire n_1868;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1975;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_1630;
wire n_1280;
wire n_729;
wire n_394;
wire n_1352;
wire n_1323;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_2054;
wire n_1236;
wire n_1523;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1935;
wire n_1645;
wire n_429;
OAI221xp5_ASAP7_75t_L g990 ( .A1(n_0), .A2(n_653), .B1(n_991), .B2(n_993), .C(n_1000), .Y(n_990) );
AOI21xp33_ASAP7_75t_L g1023 ( .A1(n_0), .A2(n_820), .B(n_1024), .Y(n_1023) );
AOI221xp5_ASAP7_75t_L g1283 ( .A1(n_1), .A2(n_71), .B1(n_555), .B2(n_898), .C(n_1284), .Y(n_1283) );
AOI22xp33_ASAP7_75t_SL g1306 ( .A1(n_1), .A2(n_203), .B1(n_452), .B2(n_1307), .Y(n_1306) );
CKINVDCx5p33_ASAP7_75t_R g1384 ( .A(n_2), .Y(n_1384) );
INVx1_ASAP7_75t_L g2000 ( .A(n_3), .Y(n_2000) );
INVx1_ASAP7_75t_L g951 ( .A(n_4), .Y(n_951) );
OAI22xp5_ASAP7_75t_L g1595 ( .A1(n_5), .A2(n_81), .B1(n_1175), .B2(n_1596), .Y(n_1595) );
INVx1_ASAP7_75t_L g1606 ( .A(n_5), .Y(n_1606) );
AOI22xp5_ASAP7_75t_L g1676 ( .A1(n_6), .A2(n_362), .B1(n_1677), .B2(n_1685), .Y(n_1676) );
CKINVDCx5p33_ASAP7_75t_R g1546 ( .A(n_7), .Y(n_1546) );
OAI221xp5_ASAP7_75t_L g1003 ( .A1(n_8), .A2(n_208), .B1(n_643), .B2(n_647), .C(n_651), .Y(n_1003) );
CKINVDCx5p33_ASAP7_75t_R g1030 ( .A(n_8), .Y(n_1030) );
AOI221xp5_ASAP7_75t_L g1054 ( .A1(n_9), .A2(n_347), .B1(n_471), .B2(n_1055), .C(n_1057), .Y(n_1054) );
INVx1_ASAP7_75t_L g1066 ( .A(n_9), .Y(n_1066) );
INVx1_ASAP7_75t_L g1439 ( .A(n_10), .Y(n_1439) );
AOI22xp33_ASAP7_75t_SL g475 ( .A1(n_11), .A2(n_336), .B1(n_470), .B2(n_476), .Y(n_475) );
INVxp33_ASAP7_75t_SL g574 ( .A(n_11), .Y(n_574) );
OAI22xp33_ASAP7_75t_L g1172 ( .A1(n_12), .A2(n_339), .B1(n_1173), .B2(n_1175), .Y(n_1172) );
INVx1_ASAP7_75t_L g1204 ( .A(n_12), .Y(n_1204) );
INVx1_ASAP7_75t_L g1602 ( .A(n_13), .Y(n_1602) );
OAI22xp5_ASAP7_75t_L g1619 ( .A1(n_13), .A2(n_93), .B1(n_979), .B2(n_984), .Y(n_1619) );
INVx1_ASAP7_75t_L g1039 ( .A(n_14), .Y(n_1039) );
INVxp33_ASAP7_75t_SL g450 ( .A(n_15), .Y(n_450) );
AOI221xp5_ASAP7_75t_L g526 ( .A1(n_15), .A2(n_180), .B1(n_527), .B2(n_532), .C(n_534), .Y(n_526) );
AOI22xp33_ASAP7_75t_L g1275 ( .A1(n_16), .A2(n_292), .B1(n_1233), .B2(n_1276), .Y(n_1275) );
INVxp33_ASAP7_75t_SL g1296 ( .A(n_16), .Y(n_1296) );
AOI22xp33_ASAP7_75t_SL g1103 ( .A1(n_17), .A2(n_172), .B1(n_465), .B2(n_856), .Y(n_1103) );
AOI221xp5_ASAP7_75t_L g1121 ( .A1(n_17), .A2(n_276), .B1(n_532), .B2(n_1122), .C(n_1124), .Y(n_1121) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_18), .A2(n_178), .B1(n_603), .B2(n_605), .Y(n_602) );
INVx1_ASAP7_75t_L g659 ( .A(n_18), .Y(n_659) );
INVx1_ASAP7_75t_L g1592 ( .A(n_19), .Y(n_1592) );
OAI221xp5_ASAP7_75t_L g1608 ( .A1(n_19), .A2(n_968), .B1(n_1189), .B2(n_1609), .C(n_1611), .Y(n_1608) );
CKINVDCx5p33_ASAP7_75t_R g914 ( .A(n_20), .Y(n_914) );
OAI22xp5_ASAP7_75t_L g751 ( .A1(n_21), .A2(n_752), .B1(n_826), .B2(n_827), .Y(n_751) );
INVx1_ASAP7_75t_L g827 ( .A(n_21), .Y(n_827) );
AOI22xp33_ASAP7_75t_L g1168 ( .A1(n_22), .A2(n_221), .B1(n_528), .B2(n_1169), .Y(n_1168) );
OAI22xp5_ASAP7_75t_L g1177 ( .A1(n_22), .A2(n_221), .B1(n_1178), .B2(n_1179), .Y(n_1177) );
AOI22xp5_ASAP7_75t_L g1688 ( .A1(n_23), .A2(n_316), .B1(n_1689), .B2(n_1693), .Y(n_1688) );
AOI22xp33_ASAP7_75t_L g1157 ( .A1(n_24), .A2(n_247), .B1(n_1158), .B2(n_1160), .Y(n_1157) );
INVxp67_ASAP7_75t_SL g1187 ( .A(n_24), .Y(n_1187) );
OAI22xp5_ASAP7_75t_L g1365 ( .A1(n_25), .A2(n_348), .B1(n_1178), .B2(n_1179), .Y(n_1365) );
AOI22xp33_ASAP7_75t_SL g1406 ( .A1(n_25), .A2(n_348), .B1(n_1232), .B2(n_1407), .Y(n_1406) );
INVx1_ASAP7_75t_L g788 ( .A(n_26), .Y(n_788) );
OAI22xp5_ASAP7_75t_L g825 ( .A1(n_26), .A2(n_364), .B1(n_573), .B2(n_576), .Y(n_825) );
AOI221xp5_ASAP7_75t_L g1041 ( .A1(n_27), .A2(n_52), .B1(n_948), .B2(n_1042), .C(n_1043), .Y(n_1041) );
AOI22xp33_ASAP7_75t_L g1072 ( .A1(n_27), .A2(n_319), .B1(n_1073), .B2(n_1074), .Y(n_1072) );
CKINVDCx16_ASAP7_75t_R g1725 ( .A(n_28), .Y(n_1725) );
CKINVDCx5p33_ASAP7_75t_R g997 ( .A(n_29), .Y(n_997) );
INVx1_ASAP7_75t_L g1045 ( .A(n_30), .Y(n_1045) );
AOI221xp5_ASAP7_75t_L g1068 ( .A1(n_30), .A2(n_52), .B1(n_549), .B2(n_1069), .C(n_1071), .Y(n_1068) );
AOI22xp33_ASAP7_75t_L g1485 ( .A1(n_31), .A2(n_104), .B1(n_603), .B2(n_1486), .Y(n_1485) );
INVx1_ASAP7_75t_L g1508 ( .A(n_31), .Y(n_1508) );
OAI22xp5_ASAP7_75t_L g1005 ( .A1(n_32), .A2(n_83), .B1(n_747), .B2(n_1006), .Y(n_1005) );
INVx1_ASAP7_75t_L g1020 ( .A(n_32), .Y(n_1020) );
AOI22xp33_ASAP7_75t_SL g1484 ( .A1(n_33), .A2(n_63), .B1(n_823), .B2(n_1467), .Y(n_1484) );
AOI21xp33_ASAP7_75t_L g1500 ( .A1(n_33), .A2(n_654), .B(n_963), .Y(n_1500) );
INVx1_ASAP7_75t_L g1059 ( .A(n_34), .Y(n_1059) );
INVxp33_ASAP7_75t_L g1525 ( .A(n_35), .Y(n_1525) );
AOI221xp5_ASAP7_75t_L g1552 ( .A1(n_35), .A2(n_103), .B1(n_1226), .B2(n_1483), .C(n_1553), .Y(n_1552) );
OAI221xp5_ASAP7_75t_L g1930 ( .A1(n_36), .A2(n_109), .B1(n_641), .B2(n_646), .C(n_1653), .Y(n_1930) );
OAI22xp5_ASAP7_75t_L g1951 ( .A1(n_36), .A2(n_109), .B1(n_624), .B2(n_1448), .Y(n_1951) );
AOI22xp33_ASAP7_75t_SL g1534 ( .A1(n_37), .A2(n_191), .B1(n_1535), .B2(n_1536), .Y(n_1534) );
AOI22xp33_ASAP7_75t_L g1566 ( .A1(n_37), .A2(n_191), .B1(n_1567), .B2(n_1569), .Y(n_1566) );
INVx1_ASAP7_75t_L g794 ( .A(n_38), .Y(n_794) );
OAI211xp5_ASAP7_75t_SL g798 ( .A1(n_38), .A2(n_799), .B(n_800), .C(n_807), .Y(n_798) );
AOI221xp5_ASAP7_75t_L g1196 ( .A1(n_39), .A2(n_141), .B1(n_854), .B2(n_856), .C(n_1197), .Y(n_1196) );
OAI22xp5_ASAP7_75t_L g1207 ( .A1(n_39), .A2(n_176), .B1(n_1208), .B2(n_1210), .Y(n_1207) );
AOI22xp33_ASAP7_75t_L g853 ( .A1(n_40), .A2(n_254), .B1(n_854), .B2(n_856), .Y(n_853) );
INVxp33_ASAP7_75t_SL g884 ( .A(n_40), .Y(n_884) );
AOI22xp33_ASAP7_75t_SL g478 ( .A1(n_41), .A2(n_328), .B1(n_465), .B2(n_479), .Y(n_478) );
INVxp33_ASAP7_75t_L g571 ( .A(n_41), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g848 ( .A1(n_42), .A2(n_332), .B1(n_849), .B2(n_850), .Y(n_848) );
AOI22xp33_ASAP7_75t_L g880 ( .A1(n_42), .A2(n_138), .B1(n_527), .B2(n_881), .Y(n_880) );
INVx1_ASAP7_75t_L g382 ( .A(n_43), .Y(n_382) );
INVx1_ASAP7_75t_L g1328 ( .A(n_44), .Y(n_1328) );
AOI22xp33_ASAP7_75t_L g1356 ( .A1(n_44), .A2(n_308), .B1(n_881), .B2(n_1357), .Y(n_1356) );
AOI22xp33_ASAP7_75t_L g852 ( .A1(n_45), .A2(n_258), .B1(n_849), .B2(n_850), .Y(n_852) );
INVxp67_ASAP7_75t_SL g862 ( .A(n_45), .Y(n_862) );
INVx1_ASAP7_75t_L g1229 ( .A(n_46), .Y(n_1229) );
OAI221xp5_ASAP7_75t_L g1250 ( .A1(n_46), .A2(n_968), .B1(n_1189), .B2(n_1251), .C(n_1255), .Y(n_1250) );
INVx1_ASAP7_75t_L g1319 ( .A(n_47), .Y(n_1319) );
AOI22xp33_ASAP7_75t_L g1589 ( .A1(n_48), .A2(n_210), .B1(n_1483), .B2(n_1590), .Y(n_1589) );
INVx1_ASAP7_75t_L g1613 ( .A(n_48), .Y(n_1613) );
AOI22xp5_ASAP7_75t_L g1712 ( .A1(n_49), .A2(n_187), .B1(n_1677), .B2(n_1685), .Y(n_1712) );
AOI22xp33_ASAP7_75t_L g1964 ( .A1(n_49), .A2(n_1965), .B1(n_1968), .B2(n_2056), .Y(n_1964) );
XNOR2xp5_ASAP7_75t_L g1970 ( .A(n_49), .B(n_1971), .Y(n_1970) );
INVx1_ASAP7_75t_L g760 ( .A(n_50), .Y(n_760) );
AOI221xp5_ASAP7_75t_L g817 ( .A1(n_50), .A2(n_307), .B1(n_818), .B2(n_821), .C(n_824), .Y(n_817) );
AOI22xp33_ASAP7_75t_L g1744 ( .A1(n_51), .A2(n_243), .B1(n_1714), .B2(n_1745), .Y(n_1744) );
INVx1_ASAP7_75t_L g441 ( .A(n_53), .Y(n_441) );
INVx1_ASAP7_75t_L g1240 ( .A(n_54), .Y(n_1240) );
OAI22xp5_ASAP7_75t_L g1264 ( .A1(n_54), .A2(n_261), .B1(n_1208), .B2(n_1210), .Y(n_1264) );
AOI22xp33_ASAP7_75t_SL g1539 ( .A1(n_55), .A2(n_334), .B1(n_470), .B2(n_1540), .Y(n_1539) );
AOI221xp5_ASAP7_75t_L g1560 ( .A1(n_55), .A2(n_334), .B1(n_1561), .B2(n_1562), .C(n_1564), .Y(n_1560) );
INVx1_ASAP7_75t_L g1941 ( .A(n_56), .Y(n_1941) );
INVxp33_ASAP7_75t_L g1322 ( .A(n_57), .Y(n_1322) );
AOI221xp5_ASAP7_75t_L g1349 ( .A1(n_57), .A2(n_324), .B1(n_1233), .B2(n_1350), .C(n_1351), .Y(n_1349) );
INVx1_ASAP7_75t_L g1167 ( .A(n_58), .Y(n_1167) );
OAI211xp5_ASAP7_75t_SL g1190 ( .A1(n_58), .A2(n_928), .B(n_1191), .C(n_1198), .Y(n_1190) );
OAI22xp5_ASAP7_75t_L g1973 ( .A1(n_59), .A2(n_356), .B1(n_1974), .B2(n_1978), .Y(n_1973) );
AOI22xp33_ASAP7_75t_L g2012 ( .A1(n_59), .A2(n_274), .B1(n_849), .B2(n_1538), .Y(n_2012) );
CKINVDCx5p33_ASAP7_75t_R g1108 ( .A(n_60), .Y(n_1108) );
INVx1_ASAP7_75t_L g697 ( .A(n_61), .Y(n_697) );
AOI22xp33_ASAP7_75t_L g724 ( .A1(n_61), .A2(n_317), .B1(n_467), .B2(n_725), .Y(n_724) );
XOR2x2_ASAP7_75t_L g1086 ( .A(n_62), .B(n_1087), .Y(n_1086) );
AOI22xp5_ASAP7_75t_L g1696 ( .A1(n_62), .A2(n_152), .B1(n_1677), .B2(n_1685), .Y(n_1696) );
INVx1_ASAP7_75t_L g1499 ( .A(n_63), .Y(n_1499) );
AOI22xp33_ASAP7_75t_L g903 ( .A1(n_64), .A2(n_372), .B1(n_900), .B2(n_901), .Y(n_903) );
OAI22xp33_ASAP7_75t_L g967 ( .A1(n_64), .A2(n_352), .B1(n_968), .B2(n_970), .Y(n_967) );
INVx1_ASAP7_75t_L g1464 ( .A(n_65), .Y(n_1464) );
OAI221xp5_ASAP7_75t_L g1470 ( .A1(n_65), .A2(n_314), .B1(n_1471), .B2(n_1472), .C(n_1473), .Y(n_1470) );
AOI22xp33_ASAP7_75t_SL g1541 ( .A1(n_66), .A2(n_148), .B1(n_470), .B2(n_1536), .Y(n_1541) );
INVxp67_ASAP7_75t_SL g1549 ( .A(n_66), .Y(n_1549) );
AO221x2_ASAP7_75t_L g1702 ( .A1(n_67), .A2(n_278), .B1(n_1689), .B2(n_1693), .C(n_1703), .Y(n_1702) );
CKINVDCx16_ASAP7_75t_R g1727 ( .A(n_68), .Y(n_1727) );
INVx1_ASAP7_75t_L g1959 ( .A(n_69), .Y(n_1959) );
AOI22xp5_ASAP7_75t_SL g1731 ( .A1(n_70), .A2(n_260), .B1(n_1693), .B2(n_1714), .Y(n_1731) );
AOI22xp33_ASAP7_75t_SL g1303 ( .A1(n_71), .A2(n_183), .B1(n_1304), .B2(n_1305), .Y(n_1303) );
INVx1_ASAP7_75t_L g1340 ( .A(n_72), .Y(n_1340) );
CKINVDCx5p33_ASAP7_75t_R g1100 ( .A(n_73), .Y(n_1100) );
INVx1_ASAP7_75t_L g1038 ( .A(n_74), .Y(n_1038) );
INVxp33_ASAP7_75t_SL g1101 ( .A(n_75), .Y(n_1101) );
AOI221xp5_ASAP7_75t_L g1113 ( .A1(n_75), .A2(n_269), .B1(n_561), .B2(n_1114), .C(n_1116), .Y(n_1113) );
AOI22xp33_ASAP7_75t_L g1002 ( .A1(n_76), .A2(n_200), .B1(n_963), .B2(n_999), .Y(n_1002) );
OAI22xp5_ASAP7_75t_L g1010 ( .A1(n_76), .A2(n_200), .B1(n_573), .B2(n_594), .Y(n_1010) );
INVx1_ASAP7_75t_L g1339 ( .A(n_77), .Y(n_1339) );
CKINVDCx14_ASAP7_75t_R g1783 ( .A(n_78), .Y(n_1783) );
INVxp67_ASAP7_75t_SL g1277 ( .A(n_79), .Y(n_1277) );
AOI22xp33_ASAP7_75t_SL g1308 ( .A1(n_79), .A2(n_224), .B1(n_452), .B2(n_472), .Y(n_1308) );
AOI22xp33_ASAP7_75t_SL g1104 ( .A1(n_80), .A2(n_276), .B1(n_470), .B2(n_476), .Y(n_1104) );
AOI22xp33_ASAP7_75t_L g1126 ( .A1(n_80), .A2(n_172), .B1(n_1079), .B2(n_1127), .Y(n_1126) );
INVx1_ASAP7_75t_L g1607 ( .A(n_81), .Y(n_1607) );
OAI221xp5_ASAP7_75t_L g765 ( .A1(n_82), .A2(n_110), .B1(n_641), .B2(n_766), .C(n_767), .Y(n_765) );
INVx1_ASAP7_75t_L g813 ( .A(n_82), .Y(n_813) );
AOI22xp33_ASAP7_75t_L g1022 ( .A1(n_83), .A2(n_133), .B1(n_511), .B2(n_1018), .Y(n_1022) );
INVxp67_ASAP7_75t_SL g1094 ( .A(n_84), .Y(n_1094) );
OAI22xp33_ASAP7_75t_L g1112 ( .A1(n_84), .A2(n_320), .B1(n_516), .B2(n_521), .Y(n_1112) );
XOR2xp5_ASAP7_75t_L g890 ( .A(n_85), .B(n_891), .Y(n_890) );
AOI22xp33_ASAP7_75t_SL g1542 ( .A1(n_86), .A2(n_128), .B1(n_1535), .B2(n_1540), .Y(n_1542) );
INVxp67_ASAP7_75t_L g1559 ( .A(n_86), .Y(n_1559) );
INVx1_ASAP7_75t_L g1098 ( .A(n_87), .Y(n_1098) );
INVx1_ASAP7_75t_L g949 ( .A(n_88), .Y(n_949) );
INVx1_ASAP7_75t_L g1370 ( .A(n_89), .Y(n_1370) );
AOI22xp33_ASAP7_75t_L g1400 ( .A1(n_89), .A2(n_106), .B1(n_898), .B2(n_1233), .Y(n_1400) );
CKINVDCx5p33_ASAP7_75t_R g1345 ( .A(n_90), .Y(n_1345) );
AOI22xp33_ASAP7_75t_L g1742 ( .A1(n_91), .A2(n_233), .B1(n_1677), .B2(n_1743), .Y(n_1742) );
AOI22xp33_ASAP7_75t_L g897 ( .A1(n_92), .A2(n_333), .B1(n_527), .B2(n_898), .Y(n_897) );
INVx1_ASAP7_75t_L g932 ( .A(n_92), .Y(n_932) );
AOI221xp5_ASAP7_75t_L g1603 ( .A1(n_93), .A2(n_369), .B1(n_845), .B2(n_1197), .C(n_1604), .Y(n_1603) );
INVx1_ASAP7_75t_L g1593 ( .A(n_94), .Y(n_1593) );
OAI211xp5_ASAP7_75t_L g1598 ( .A1(n_94), .A2(n_928), .B(n_1599), .C(n_1605), .Y(n_1598) );
INVx1_ASAP7_75t_L g1926 ( .A(n_95), .Y(n_1926) );
OAI222xp33_ASAP7_75t_L g1424 ( .A1(n_96), .A2(n_166), .B1(n_331), .B2(n_490), .C1(n_766), .C2(n_1425), .Y(n_1424) );
INVx1_ASAP7_75t_L g1450 ( .A(n_96), .Y(n_1450) );
OAI211xp5_ASAP7_75t_SL g707 ( .A1(n_97), .A2(n_708), .B(n_709), .C(n_712), .Y(n_707) );
AOI22xp33_ASAP7_75t_L g731 ( .A1(n_97), .A2(n_213), .B1(n_727), .B2(n_732), .Y(n_731) );
AOI22xp33_ASAP7_75t_L g1594 ( .A1(n_98), .A2(n_253), .B1(n_528), .B2(n_1169), .Y(n_1594) );
OAI22xp5_ASAP7_75t_L g1614 ( .A1(n_98), .A2(n_253), .B1(n_1178), .B2(n_1179), .Y(n_1614) );
CKINVDCx5p33_ASAP7_75t_R g763 ( .A(n_99), .Y(n_763) );
CKINVDCx5p33_ASAP7_75t_R g777 ( .A(n_100), .Y(n_777) );
AOI221xp5_ASAP7_75t_L g1633 ( .A1(n_101), .A2(n_259), .B1(n_816), .B2(n_1233), .C(n_1634), .Y(n_1633) );
INVx1_ASAP7_75t_L g1651 ( .A(n_101), .Y(n_1651) );
INVx1_ASAP7_75t_L g1342 ( .A(n_102), .Y(n_1342) );
INVxp33_ASAP7_75t_SL g1531 ( .A(n_103), .Y(n_1531) );
OAI22xp5_ASAP7_75t_L g1513 ( .A1(n_104), .A2(n_112), .B1(n_927), .B2(n_961), .Y(n_1513) );
CKINVDCx14_ASAP7_75t_R g1704 ( .A(n_105), .Y(n_1704) );
INVx1_ASAP7_75t_L g1368 ( .A(n_106), .Y(n_1368) );
OAI22xp5_ASAP7_75t_L g621 ( .A1(n_107), .A2(n_367), .B1(n_622), .B2(n_624), .Y(n_621) );
OAI221xp5_ASAP7_75t_L g640 ( .A1(n_107), .A2(n_367), .B1(n_641), .B2(n_646), .C(n_650), .Y(n_640) );
AOI22xp33_ASAP7_75t_L g1482 ( .A1(n_108), .A2(n_124), .B1(n_804), .B2(n_1483), .Y(n_1482) );
INVx1_ASAP7_75t_L g1503 ( .A(n_108), .Y(n_1503) );
INVx1_ASAP7_75t_L g811 ( .A(n_110), .Y(n_811) );
OR2x2_ASAP7_75t_L g417 ( .A(n_111), .B(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g438 ( .A(n_111), .Y(n_438) );
BUFx2_ASAP7_75t_L g462 ( .A(n_111), .Y(n_462) );
BUFx2_ASAP7_75t_L g493 ( .A(n_111), .Y(n_493) );
OAI222xp33_ASAP7_75t_L g1515 ( .A1(n_112), .A2(n_157), .B1(n_252), .B2(n_491), .C1(n_1208), .C2(n_1210), .Y(n_1515) );
AOI22xp33_ASAP7_75t_SL g2007 ( .A1(n_113), .A2(n_266), .B1(n_1535), .B2(n_2008), .Y(n_2007) );
AOI22xp33_ASAP7_75t_SL g2015 ( .A1(n_113), .A2(n_266), .B1(n_1274), .B2(n_1405), .Y(n_2015) );
AOI22xp33_ASAP7_75t_SL g998 ( .A1(n_114), .A2(n_162), .B1(n_963), .B2(n_999), .Y(n_998) );
INVx1_ASAP7_75t_L g1016 ( .A(n_114), .Y(n_1016) );
INVx1_ASAP7_75t_L g1223 ( .A(n_115), .Y(n_1223) );
INVx1_ASAP7_75t_L g1343 ( .A(n_116), .Y(n_1343) );
INVx1_ASAP7_75t_L g1492 ( .A(n_117), .Y(n_1492) );
OAI221xp5_ASAP7_75t_L g1509 ( .A1(n_117), .A2(n_225), .B1(n_1203), .B2(n_1510), .C(n_1512), .Y(n_1509) );
AOI22xp33_ASAP7_75t_SL g1105 ( .A1(n_118), .A2(n_229), .B1(n_470), .B2(n_476), .Y(n_1105) );
INVxp33_ASAP7_75t_SL g1130 ( .A(n_118), .Y(n_1130) );
CKINVDCx5p33_ASAP7_75t_R g1636 ( .A(n_119), .Y(n_1636) );
CKINVDCx5p33_ASAP7_75t_R g1260 ( .A(n_120), .Y(n_1260) );
INVx1_ASAP7_75t_L g1321 ( .A(n_121), .Y(n_1321) );
OAI221xp5_ASAP7_75t_L g1323 ( .A1(n_122), .A2(n_357), .B1(n_766), .B2(n_767), .C(n_1324), .Y(n_1323) );
OAI22xp5_ASAP7_75t_L g1348 ( .A1(n_122), .A2(n_357), .B1(n_865), .B2(n_1279), .Y(n_1348) );
CKINVDCx5p33_ASAP7_75t_R g1387 ( .A(n_123), .Y(n_1387) );
INVx1_ASAP7_75t_L g1502 ( .A(n_124), .Y(n_1502) );
AOI221xp5_ASAP7_75t_L g596 ( .A1(n_125), .A2(n_216), .B1(n_597), .B2(n_598), .C(n_600), .Y(n_596) );
INVxp67_ASAP7_75t_SL g671 ( .A(n_125), .Y(n_671) );
AOI22xp33_ASAP7_75t_SL g1106 ( .A1(n_126), .A2(n_287), .B1(n_465), .B2(n_856), .Y(n_1106) );
INVxp33_ASAP7_75t_L g1129 ( .A(n_126), .Y(n_1129) );
INVxp33_ASAP7_75t_L g1925 ( .A(n_127), .Y(n_1925) );
AOI221xp5_ASAP7_75t_L g1952 ( .A1(n_127), .A2(n_374), .B1(n_549), .B2(n_1233), .C(n_1953), .Y(n_1952) );
INVxp33_ASAP7_75t_L g1571 ( .A(n_128), .Y(n_1571) );
INVx1_ASAP7_75t_L g1164 ( .A(n_129), .Y(n_1164) );
OAI221xp5_ASAP7_75t_L g1180 ( .A1(n_129), .A2(n_968), .B1(n_1181), .B2(n_1185), .C(n_1189), .Y(n_1180) );
INVx1_ASAP7_75t_L g1058 ( .A(n_130), .Y(n_1058) );
OAI221xp5_ASAP7_75t_L g1062 ( .A1(n_130), .A2(n_347), .B1(n_620), .B2(n_1063), .C(n_1065), .Y(n_1062) );
AOI22xp33_ASAP7_75t_L g1231 ( .A1(n_131), .A2(n_151), .B1(n_1232), .B2(n_1233), .Y(n_1231) );
OAI22xp5_ASAP7_75t_L g1258 ( .A1(n_131), .A2(n_151), .B1(n_924), .B2(n_970), .Y(n_1258) );
OAI221xp5_ASAP7_75t_L g1376 ( .A1(n_132), .A2(n_928), .B1(n_1377), .B2(n_1381), .C(n_1386), .Y(n_1376) );
AOI22xp33_ASAP7_75t_SL g1404 ( .A1(n_132), .A2(n_240), .B1(n_818), .B2(n_1405), .Y(n_1404) );
OAI22xp33_ASAP7_75t_L g1007 ( .A1(n_133), .A2(n_158), .B1(n_490), .B2(n_746), .Y(n_1007) );
OAI22xp5_ASAP7_75t_L g1278 ( .A1(n_134), .A2(n_194), .B1(n_1279), .B2(n_1280), .Y(n_1278) );
INVxp67_ASAP7_75t_SL g1293 ( .A(n_134), .Y(n_1293) );
INVx1_ASAP7_75t_L g1529 ( .A(n_135), .Y(n_1529) );
INVx1_ASAP7_75t_L g445 ( .A(n_136), .Y(n_445) );
XNOR2xp5_ASAP7_75t_L g1920 ( .A(n_137), .B(n_1921), .Y(n_1920) );
AOI22xp33_ASAP7_75t_SL g843 ( .A1(n_138), .A2(n_304), .B1(n_844), .B2(n_846), .Y(n_843) );
AOI221xp5_ASAP7_75t_L g613 ( .A1(n_139), .A2(n_182), .B1(n_598), .B2(n_614), .C(n_616), .Y(n_613) );
INVx1_ASAP7_75t_L g637 ( .A(n_139), .Y(n_637) );
INVx1_ASAP7_75t_L g1580 ( .A(n_140), .Y(n_1580) );
OAI22xp5_ASAP7_75t_L g1206 ( .A1(n_141), .A2(n_227), .B1(n_979), .B2(n_984), .Y(n_1206) );
INVx1_ASAP7_75t_L g1374 ( .A(n_142), .Y(n_1374) );
AOI22xp33_ASAP7_75t_L g1401 ( .A1(n_142), .A2(n_150), .B1(n_1402), .B2(n_1403), .Y(n_1401) );
INVx1_ASAP7_75t_L g886 ( .A(n_143), .Y(n_886) );
INVxp67_ASAP7_75t_L g1332 ( .A(n_144), .Y(n_1332) );
AOI221xp5_ASAP7_75t_L g1353 ( .A1(n_144), .A2(n_231), .B1(n_705), .B2(n_1354), .C(n_1355), .Y(n_1353) );
CKINVDCx5p33_ASAP7_75t_R g1643 ( .A(n_145), .Y(n_1643) );
AOI22xp33_ASAP7_75t_L g2027 ( .A1(n_146), .A2(n_257), .B1(n_1350), .B2(n_2028), .Y(n_2027) );
OAI22xp5_ASAP7_75t_L g2047 ( .A1(n_146), .A2(n_257), .B1(n_2048), .B2(n_2050), .Y(n_2047) );
XOR2x2_ASAP7_75t_L g1214 ( .A(n_147), .B(n_1215), .Y(n_1214) );
INVxp33_ASAP7_75t_L g1572 ( .A(n_148), .Y(n_1572) );
CKINVDCx5p33_ASAP7_75t_R g1270 ( .A(n_149), .Y(n_1270) );
INVx1_ASAP7_75t_L g1373 ( .A(n_150), .Y(n_1373) );
CKINVDCx5p33_ASAP7_75t_R g711 ( .A(n_153), .Y(n_711) );
AOI221xp5_ASAP7_75t_L g1639 ( .A1(n_154), .A2(n_282), .B1(n_597), .B2(n_1071), .C(n_1640), .Y(n_1639) );
INVx1_ASAP7_75t_L g1660 ( .A(n_154), .Y(n_1660) );
OAI22xp5_ASAP7_75t_L g1980 ( .A1(n_155), .A2(n_274), .B1(n_1981), .B2(n_1985), .Y(n_1980) );
INVxp33_ASAP7_75t_SL g2040 ( .A(n_155), .Y(n_2040) );
CKINVDCx5p33_ASAP7_75t_R g1630 ( .A(n_156), .Y(n_1630) );
AOI221xp5_ASAP7_75t_L g1506 ( .A1(n_157), .A2(n_296), .B1(n_467), .B2(n_956), .C(n_1507), .Y(n_1506) );
INVx1_ASAP7_75t_L g1026 ( .A(n_158), .Y(n_1026) );
INVxp67_ASAP7_75t_SL g1522 ( .A(n_159), .Y(n_1522) );
OAI22xp33_ASAP7_75t_L g1550 ( .A1(n_159), .A2(n_197), .B1(n_865), .B2(n_1551), .Y(n_1550) );
INVx1_ASAP7_75t_L g595 ( .A(n_160), .Y(n_595) );
XNOR2xp5_ASAP7_75t_L g1625 ( .A(n_161), .B(n_1626), .Y(n_1625) );
INVx1_ASAP7_75t_L g1013 ( .A(n_162), .Y(n_1013) );
CKINVDCx5p33_ASAP7_75t_R g1143 ( .A(n_163), .Y(n_1143) );
AOI21xp33_ASAP7_75t_L g704 ( .A1(n_164), .A2(n_533), .B(n_705), .Y(n_704) );
AOI22xp33_ASAP7_75t_L g726 ( .A1(n_164), .A2(n_196), .B1(n_727), .B2(n_729), .Y(n_726) );
INVxp33_ASAP7_75t_L g1933 ( .A(n_165), .Y(n_1933) );
AOI22xp33_ASAP7_75t_L g1957 ( .A1(n_165), .A2(n_175), .B1(n_1073), .B2(n_1074), .Y(n_1957) );
INVx1_ASAP7_75t_L g1460 ( .A(n_166), .Y(n_1460) );
INVx1_ASAP7_75t_L g1242 ( .A(n_167), .Y(n_1242) );
OAI22xp5_ASAP7_75t_L g1262 ( .A1(n_167), .A2(n_242), .B1(n_984), .B2(n_1263), .Y(n_1262) );
AOI22xp5_ASAP7_75t_SL g1730 ( .A1(n_168), .A2(n_193), .B1(n_1677), .B2(n_1685), .Y(n_1730) );
OAI22xp33_ASAP7_75t_L g717 ( .A1(n_169), .A2(n_213), .B1(n_573), .B2(n_576), .Y(n_717) );
AOI22xp33_ASAP7_75t_L g735 ( .A1(n_169), .A2(n_295), .B1(n_467), .B2(n_736), .Y(n_735) );
OAI22xp33_ASAP7_75t_SL g1631 ( .A1(n_170), .A2(n_343), .B1(n_1448), .B2(n_1632), .Y(n_1631) );
OAI221xp5_ASAP7_75t_L g1652 ( .A1(n_170), .A2(n_343), .B1(n_641), .B2(n_646), .C(n_1653), .Y(n_1652) );
CKINVDCx5p33_ASAP7_75t_R g710 ( .A(n_171), .Y(n_710) );
INVx1_ASAP7_75t_L g1681 ( .A(n_173), .Y(n_1681) );
INVxp67_ASAP7_75t_SL g773 ( .A(n_174), .Y(n_773) );
AOI221xp5_ASAP7_75t_L g805 ( .A1(n_174), .A2(n_338), .B1(n_549), .B2(n_551), .C(n_806), .Y(n_805) );
INVxp67_ASAP7_75t_SL g1938 ( .A(n_175), .Y(n_1938) );
INVx1_ASAP7_75t_L g1194 ( .A(n_176), .Y(n_1194) );
AOI22xp33_ASAP7_75t_SL g469 ( .A1(n_177), .A2(n_226), .B1(n_470), .B2(n_472), .Y(n_469) );
AOI22xp33_ASAP7_75t_L g557 ( .A1(n_177), .A2(n_291), .B1(n_558), .B2(n_561), .Y(n_557) );
INVx1_ASAP7_75t_L g673 ( .A(n_178), .Y(n_673) );
OAI22xp5_ASAP7_75t_L g585 ( .A1(n_179), .A2(n_586), .B1(n_687), .B2(n_688), .Y(n_585) );
INVx1_ASAP7_75t_L g688 ( .A(n_179), .Y(n_688) );
INVxp33_ASAP7_75t_SL g431 ( .A(n_180), .Y(n_431) );
INVx1_ASAP7_75t_L g1944 ( .A(n_181), .Y(n_1944) );
INVx1_ASAP7_75t_L g634 ( .A(n_182), .Y(n_634) );
AOI22xp33_ASAP7_75t_L g1286 ( .A1(n_183), .A2(n_203), .B1(n_818), .B2(n_1160), .Y(n_1286) );
CKINVDCx5p33_ASAP7_75t_R g1638 ( .A(n_184), .Y(n_1638) );
INVx1_ASAP7_75t_L g1220 ( .A(n_185), .Y(n_1220) );
CKINVDCx16_ASAP7_75t_R g1722 ( .A(n_186), .Y(n_1722) );
AOI22xp33_ASAP7_75t_L g617 ( .A1(n_188), .A2(n_238), .B1(n_618), .B2(n_619), .Y(n_617) );
INVx1_ASAP7_75t_L g631 ( .A(n_188), .Y(n_631) );
INVx1_ASAP7_75t_L g1682 ( .A(n_189), .Y(n_1682) );
NAND2xp5_ASAP7_75t_L g1687 ( .A(n_189), .B(n_1680), .Y(n_1687) );
INVx1_ASAP7_75t_L g1433 ( .A(n_190), .Y(n_1433) );
CKINVDCx5p33_ASAP7_75t_R g1635 ( .A(n_192), .Y(n_1635) );
INVx1_ASAP7_75t_L g1360 ( .A(n_193), .Y(n_1360) );
INVxp67_ASAP7_75t_SL g1294 ( .A(n_194), .Y(n_1294) );
INVx2_ASAP7_75t_L g394 ( .A(n_195), .Y(n_394) );
INVx1_ASAP7_75t_L g699 ( .A(n_196), .Y(n_699) );
INVxp67_ASAP7_75t_SL g1523 ( .A(n_197), .Y(n_1523) );
INVxp67_ASAP7_75t_L g1435 ( .A(n_198), .Y(n_1435) );
OAI222xp33_ASAP7_75t_L g1452 ( .A1(n_198), .A2(n_206), .B1(n_301), .B2(n_906), .C1(n_1063), .C2(n_1211), .Y(n_1452) );
INVx1_ASAP7_75t_L g1645 ( .A(n_199), .Y(n_1645) );
BUFx3_ASAP7_75t_L g502 ( .A(n_201), .Y(n_502) );
INVx1_ASAP7_75t_L g531 ( .A(n_201), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g2024 ( .A1(n_202), .A2(n_207), .B1(n_1405), .B2(n_2025), .Y(n_2024) );
INVx1_ASAP7_75t_L g2038 ( .A(n_202), .Y(n_2038) );
OAI211xp5_ASAP7_75t_L g752 ( .A1(n_204), .A2(n_753), .B(n_755), .C(n_797), .Y(n_752) );
INVx1_ASAP7_75t_L g946 ( .A(n_205), .Y(n_946) );
INVxp67_ASAP7_75t_L g1438 ( .A(n_206), .Y(n_1438) );
INVx1_ASAP7_75t_L g2032 ( .A(n_207), .Y(n_2032) );
CKINVDCx5p33_ASAP7_75t_R g1031 ( .A(n_208), .Y(n_1031) );
AOI22xp33_ASAP7_75t_L g464 ( .A1(n_209), .A2(n_291), .B1(n_465), .B2(n_466), .Y(n_464) );
AOI221xp5_ASAP7_75t_L g548 ( .A1(n_209), .A2(n_226), .B1(n_549), .B2(n_551), .C(n_555), .Y(n_548) );
INVx1_ASAP7_75t_L g1612 ( .A(n_210), .Y(n_1612) );
CKINVDCx5p33_ASAP7_75t_R g1380 ( .A(n_211), .Y(n_1380) );
INVx1_ASAP7_75t_L g1046 ( .A(n_212), .Y(n_1046) );
AOI22xp33_ASAP7_75t_L g2005 ( .A1(n_214), .A2(n_346), .B1(n_849), .B2(n_2006), .Y(n_2005) );
AOI22xp33_ASAP7_75t_L g2016 ( .A1(n_214), .A2(n_346), .B1(n_2017), .B2(n_2019), .Y(n_2016) );
AOI22xp33_ASAP7_75t_L g1224 ( .A1(n_215), .A2(n_350), .B1(n_1225), .B2(n_1226), .Y(n_1224) );
INVxp67_ASAP7_75t_SL g1257 ( .A(n_215), .Y(n_1257) );
INVxp67_ASAP7_75t_SL g665 ( .A(n_216), .Y(n_665) );
AOI22xp33_ASAP7_75t_L g904 ( .A1(n_217), .A2(n_352), .B1(n_532), .B2(n_905), .Y(n_904) );
OAI22xp33_ASAP7_75t_L g923 ( .A1(n_217), .A2(n_372), .B1(n_924), .B2(n_928), .Y(n_923) );
CKINVDCx5p33_ASAP7_75t_R g919 ( .A(n_218), .Y(n_919) );
INVxp33_ASAP7_75t_SL g836 ( .A(n_219), .Y(n_836) );
AOI22xp33_ASAP7_75t_SL g869 ( .A1(n_219), .A2(n_264), .B1(n_533), .B2(n_562), .Y(n_869) );
INVxp67_ASAP7_75t_SL g834 ( .A(n_220), .Y(n_834) );
OAI221xp5_ASAP7_75t_L g863 ( .A1(n_220), .A2(n_265), .B1(n_864), .B2(n_865), .C(n_867), .Y(n_863) );
INVx1_ASAP7_75t_L g497 ( .A(n_222), .Y(n_497) );
INVx1_ASAP7_75t_L g546 ( .A(n_222), .Y(n_546) );
INVx1_ASAP7_75t_L g591 ( .A(n_223), .Y(n_591) );
INVxp33_ASAP7_75t_L g1290 ( .A(n_224), .Y(n_1290) );
INVx1_ASAP7_75t_L g1491 ( .A(n_225), .Y(n_1491) );
INVx1_ASAP7_75t_L g1195 ( .A(n_227), .Y(n_1195) );
INVx1_ASAP7_75t_L g1526 ( .A(n_228), .Y(n_1526) );
INVxp67_ASAP7_75t_SL g1111 ( .A(n_229), .Y(n_1111) );
XNOR2xp5_ASAP7_75t_L g1421 ( .A(n_230), .B(n_1422), .Y(n_1421) );
INVxp67_ASAP7_75t_L g1330 ( .A(n_231), .Y(n_1330) );
INVxp67_ASAP7_75t_SL g1937 ( .A(n_232), .Y(n_1937) );
AOI221xp5_ASAP7_75t_L g1956 ( .A1(n_232), .A2(n_310), .B1(n_1069), .B2(n_1071), .C(n_1561), .Y(n_1956) );
OAI22xp5_ASAP7_75t_L g405 ( .A1(n_233), .A2(n_406), .B1(n_407), .B2(n_581), .Y(n_405) );
INVx1_ASAP7_75t_L g581 ( .A(n_233), .Y(n_581) );
INVxp67_ASAP7_75t_L g1428 ( .A(n_234), .Y(n_1428) );
AOI221xp5_ASAP7_75t_L g1455 ( .A1(n_234), .A2(n_340), .B1(n_597), .B2(n_600), .C(n_1456), .Y(n_1455) );
OAI21xp33_ASAP7_75t_L g1035 ( .A1(n_235), .A2(n_1036), .B(n_1060), .Y(n_1035) );
INVx1_ASAP7_75t_L g1085 ( .A(n_235), .Y(n_1085) );
CKINVDCx20_ASAP7_75t_R g1781 ( .A(n_236), .Y(n_1781) );
CKINVDCx5p33_ASAP7_75t_R g505 ( .A(n_237), .Y(n_505) );
INVx1_ASAP7_75t_L g638 ( .A(n_238), .Y(n_638) );
INVxp67_ASAP7_75t_SL g1287 ( .A(n_239), .Y(n_1287) );
AOI22xp33_ASAP7_75t_SL g1309 ( .A1(n_239), .A2(n_312), .B1(n_465), .B2(n_1305), .Y(n_1309) );
OAI221xp5_ASAP7_75t_L g1366 ( .A1(n_240), .A2(n_968), .B1(n_1367), .B2(n_1371), .C(n_1375), .Y(n_1366) );
XOR2xp5_ASAP7_75t_L g987 ( .A(n_241), .B(n_988), .Y(n_987) );
AOI221xp5_ASAP7_75t_L g1243 ( .A1(n_242), .A2(n_261), .B1(n_1244), .B2(n_1245), .C(n_1246), .Y(n_1243) );
CKINVDCx14_ASAP7_75t_R g1706 ( .A(n_244), .Y(n_1706) );
AOI22xp33_ASAP7_75t_L g715 ( .A1(n_245), .A2(n_298), .B1(n_510), .B2(n_562), .Y(n_715) );
OAI22xp5_ASAP7_75t_L g745 ( .A1(n_245), .A2(n_370), .B1(n_746), .B2(n_747), .Y(n_745) );
XNOR2xp5_ASAP7_75t_L g1475 ( .A(n_246), .B(n_1476), .Y(n_1475) );
INVxp67_ASAP7_75t_SL g1188 ( .A(n_247), .Y(n_1188) );
INVx1_ASAP7_75t_L g1053 ( .A(n_248), .Y(n_1053) );
AOI221xp5_ASAP7_75t_L g1076 ( .A1(n_248), .A2(n_321), .B1(n_882), .B2(n_1024), .C(n_1077), .Y(n_1076) );
INVx1_ASAP7_75t_L g1601 ( .A(n_249), .Y(n_1601) );
OAI22xp5_ASAP7_75t_L g1620 ( .A1(n_249), .A2(n_369), .B1(n_1208), .B2(n_1210), .Y(n_1620) );
CKINVDCx5p33_ASAP7_75t_R g954 ( .A(n_250), .Y(n_954) );
CKINVDCx5p33_ASAP7_75t_R g1391 ( .A(n_251), .Y(n_1391) );
AOI22xp33_ASAP7_75t_L g1505 ( .A1(n_252), .A2(n_360), .B1(n_1042), .B2(n_1335), .Y(n_1505) );
INVxp67_ASAP7_75t_SL g873 ( .A(n_254), .Y(n_873) );
AOI221xp5_ASAP7_75t_L g1273 ( .A1(n_255), .A2(n_273), .B1(n_824), .B2(n_901), .C(n_1274), .Y(n_1273) );
INVxp33_ASAP7_75t_SL g1297 ( .A(n_255), .Y(n_1297) );
INVx1_ASAP7_75t_L g626 ( .A(n_256), .Y(n_626) );
INVxp33_ASAP7_75t_SL g885 ( .A(n_258), .Y(n_885) );
INVx1_ASAP7_75t_L g1649 ( .A(n_259), .Y(n_1649) );
AOI22xp33_ASAP7_75t_L g899 ( .A1(n_262), .A2(n_272), .B1(n_900), .B2(n_901), .Y(n_899) );
INVx1_ASAP7_75t_L g941 ( .A(n_262), .Y(n_941) );
CKINVDCx20_ASAP7_75t_R g1267 ( .A(n_263), .Y(n_1267) );
INVxp33_ASAP7_75t_SL g841 ( .A(n_264), .Y(n_841) );
INVxp67_ASAP7_75t_SL g833 ( .A(n_265), .Y(n_833) );
INVx1_ASAP7_75t_L g779 ( .A(n_267), .Y(n_779) );
CKINVDCx5p33_ASAP7_75t_R g1644 ( .A(n_268), .Y(n_1644) );
INVxp33_ASAP7_75t_SL g1096 ( .A(n_269), .Y(n_1096) );
INVx1_ASAP7_75t_L g784 ( .A(n_270), .Y(n_784) );
OAI211xp5_ASAP7_75t_L g808 ( .A1(n_270), .A2(n_809), .B(n_810), .C(n_814), .Y(n_808) );
INVx1_ASAP7_75t_L g1449 ( .A(n_271), .Y(n_1449) );
INVx1_ASAP7_75t_L g937 ( .A(n_272), .Y(n_937) );
INVxp33_ASAP7_75t_L g1299 ( .A(n_273), .Y(n_1299) );
AOI22xp33_ASAP7_75t_L g1641 ( .A1(n_275), .A2(n_293), .B1(n_603), .B2(n_1462), .Y(n_1641) );
INVx1_ASAP7_75t_L g1656 ( .A(n_275), .Y(n_1656) );
INVx1_ASAP7_75t_L g1230 ( .A(n_277), .Y(n_1230) );
OAI211xp5_ASAP7_75t_SL g1237 ( .A1(n_277), .A2(n_928), .B(n_1238), .C(n_1247), .Y(n_1237) );
CKINVDCx5p33_ASAP7_75t_R g758 ( .A(n_279), .Y(n_758) );
INVx1_ASAP7_75t_L g1156 ( .A(n_280), .Y(n_1156) );
CKINVDCx20_ASAP7_75t_R g1573 ( .A(n_281), .Y(n_1573) );
INVx1_ASAP7_75t_L g1658 ( .A(n_282), .Y(n_1658) );
BUFx3_ASAP7_75t_L g504 ( .A(n_283), .Y(n_504) );
INVx1_ASAP7_75t_L g512 ( .A(n_283), .Y(n_512) );
INVx1_ASAP7_75t_L g859 ( .A(n_284), .Y(n_859) );
AO221x2_ASAP7_75t_L g1778 ( .A1(n_285), .A2(n_351), .B1(n_1745), .B2(n_1779), .C(n_1780), .Y(n_1778) );
AOI21xp33_ASAP7_75t_L g716 ( .A1(n_286), .A2(n_614), .B(n_616), .Y(n_716) );
INVx1_ASAP7_75t_L g743 ( .A(n_286), .Y(n_743) );
INVxp67_ASAP7_75t_SL g1120 ( .A(n_287), .Y(n_1120) );
AOI22xp5_ASAP7_75t_L g1697 ( .A1(n_288), .A2(n_289), .B1(n_1689), .B2(n_1693), .Y(n_1697) );
HB1xp67_ASAP7_75t_L g390 ( .A(n_290), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_290), .B(n_353), .Y(n_418) );
AND2x2_ASAP7_75t_L g439 ( .A(n_290), .B(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g486 ( .A(n_290), .Y(n_486) );
INVxp33_ASAP7_75t_SL g1300 ( .A(n_292), .Y(n_1300) );
INVx1_ASAP7_75t_L g1663 ( .A(n_293), .Y(n_1663) );
CKINVDCx5p33_ASAP7_75t_R g1385 ( .A(n_294), .Y(n_1385) );
OAI221xp5_ASAP7_75t_L g693 ( .A1(n_295), .A2(n_594), .B1(n_694), .B2(n_700), .C(n_706), .Y(n_693) );
OAI22xp5_ASAP7_75t_L g1516 ( .A1(n_296), .A2(n_360), .B1(n_984), .B2(n_1263), .Y(n_1516) );
INVx2_ASAP7_75t_L g499 ( .A(n_297), .Y(n_499) );
OR2x2_ASAP7_75t_L g514 ( .A(n_297), .B(n_497), .Y(n_514) );
INVx1_ASAP7_75t_L g744 ( .A(n_298), .Y(n_744) );
AOI22xp33_ASAP7_75t_L g1001 ( .A1(n_299), .A2(n_318), .B1(n_453), .B2(n_679), .Y(n_1001) );
OAI22xp5_ASAP7_75t_L g1009 ( .A1(n_299), .A2(n_318), .B1(n_576), .B2(n_708), .Y(n_1009) );
INVx1_ASAP7_75t_L g1430 ( .A(n_300), .Y(n_1430) );
INVxp67_ASAP7_75t_L g1436 ( .A(n_301), .Y(n_1436) );
OAI211xp5_ASAP7_75t_L g1989 ( .A1(n_302), .A2(n_1990), .B(n_1991), .C(n_1994), .Y(n_1989) );
AOI22xp33_ASAP7_75t_SL g2013 ( .A1(n_302), .A2(n_356), .B1(n_1514), .B2(n_2008), .Y(n_2013) );
INVx1_ASAP7_75t_L g995 ( .A(n_303), .Y(n_995) );
AOI21xp33_ASAP7_75t_L g1014 ( .A1(n_303), .A2(n_597), .B(n_705), .Y(n_1014) );
AOI221xp5_ASAP7_75t_L g874 ( .A1(n_304), .A2(n_332), .B1(n_705), .B2(n_875), .C(n_877), .Y(n_874) );
INVx1_ASAP7_75t_L g1946 ( .A(n_305), .Y(n_1946) );
AO22x2_ASAP7_75t_L g1361 ( .A1(n_306), .A2(n_1362), .B1(n_1363), .B2(n_1412), .Y(n_1361) );
INVx1_ASAP7_75t_L g1412 ( .A(n_306), .Y(n_1412) );
INVx1_ASAP7_75t_L g762 ( .A(n_307), .Y(n_762) );
INVxp67_ASAP7_75t_L g1336 ( .A(n_308), .Y(n_1336) );
AOI22xp5_ASAP7_75t_SL g1713 ( .A1(n_309), .A2(n_313), .B1(n_1693), .B2(n_1714), .Y(n_1713) );
INVxp33_ASAP7_75t_SL g1934 ( .A(n_310), .Y(n_1934) );
CKINVDCx5p33_ASAP7_75t_R g1378 ( .A(n_311), .Y(n_1378) );
INVxp33_ASAP7_75t_SL g1289 ( .A(n_312), .Y(n_1289) );
AOI221xp5_ASAP7_75t_L g1465 ( .A1(n_314), .A2(n_335), .B1(n_1466), .B2(n_1467), .C(n_1468), .Y(n_1465) );
CKINVDCx5p33_ASAP7_75t_R g1389 ( .A(n_315), .Y(n_1389) );
INVx1_ASAP7_75t_L g701 ( .A(n_317), .Y(n_701) );
INVxp67_ASAP7_75t_SL g1044 ( .A(n_319), .Y(n_1044) );
INVxp67_ASAP7_75t_SL g1091 ( .A(n_320), .Y(n_1091) );
INVx1_ASAP7_75t_L g1052 ( .A(n_321), .Y(n_1052) );
INVxp33_ASAP7_75t_SL g840 ( .A(n_322), .Y(n_840) );
AOI21xp33_ASAP7_75t_L g870 ( .A1(n_322), .A2(n_544), .B(n_871), .Y(n_870) );
OAI22xp5_ASAP7_75t_L g689 ( .A1(n_323), .A2(n_690), .B1(n_748), .B2(n_749), .Y(n_689) );
INVxp67_ASAP7_75t_SL g748 ( .A(n_323), .Y(n_748) );
INVxp33_ASAP7_75t_L g1318 ( .A(n_324), .Y(n_1318) );
OAI22xp33_ASAP7_75t_L g1234 ( .A1(n_325), .A2(n_368), .B1(n_912), .B2(n_1235), .Y(n_1234) );
INVx1_ASAP7_75t_L g1249 ( .A(n_325), .Y(n_1249) );
INVxp67_ASAP7_75t_SL g419 ( .A(n_326), .Y(n_419) );
OAI22xp5_ASAP7_75t_L g515 ( .A1(n_326), .A2(n_375), .B1(n_516), .B2(n_521), .Y(n_515) );
OAI221xp5_ASAP7_75t_SL g1049 ( .A1(n_327), .A2(n_365), .B1(n_672), .B2(n_1050), .C(n_1051), .Y(n_1049) );
AOI22xp33_ASAP7_75t_L g1078 ( .A1(n_327), .A2(n_365), .B1(n_533), .B2(n_1079), .Y(n_1078) );
INVxp67_ASAP7_75t_SL g565 ( .A(n_328), .Y(n_565) );
INVx1_ASAP7_75t_L g838 ( .A(n_329), .Y(n_838) );
INVx1_ASAP7_75t_L g1947 ( .A(n_330), .Y(n_1947) );
INVx1_ASAP7_75t_L g1446 ( .A(n_331), .Y(n_1446) );
INVx1_ASAP7_75t_L g933 ( .A(n_333), .Y(n_933) );
OAI332xp33_ASAP7_75t_L g1426 ( .A1(n_335), .A2(n_653), .A3(n_686), .B1(n_1427), .B2(n_1431), .B3(n_1434), .C1(n_1437), .C2(n_1442), .Y(n_1426) );
INVxp67_ASAP7_75t_SL g508 ( .A(n_336), .Y(n_508) );
AOI22xp33_ASAP7_75t_SL g1487 ( .A1(n_337), .A2(n_341), .B1(n_528), .B2(n_1170), .Y(n_1487) );
INVx1_ASAP7_75t_L g1495 ( .A(n_337), .Y(n_1495) );
INVxp67_ASAP7_75t_SL g782 ( .A(n_338), .Y(n_782) );
INVx1_ASAP7_75t_L g1201 ( .A(n_339), .Y(n_1201) );
INVx1_ASAP7_75t_L g1432 ( .A(n_340), .Y(n_1432) );
INVx1_ASAP7_75t_L g1496 ( .A(n_341), .Y(n_1496) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_342), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g1684 ( .A(n_342), .B(n_382), .Y(n_1684) );
AND3x2_ASAP7_75t_L g1690 ( .A(n_342), .B(n_382), .C(n_1681), .Y(n_1690) );
CKINVDCx5p33_ASAP7_75t_R g1583 ( .A(n_344), .Y(n_1583) );
INVx2_ASAP7_75t_L g395 ( .A(n_345), .Y(n_395) );
CKINVDCx5p33_ASAP7_75t_R g1588 ( .A(n_349), .Y(n_1588) );
INVxp67_ASAP7_75t_SL g1256 ( .A(n_350), .Y(n_1256) );
INVx1_ASAP7_75t_L g397 ( .A(n_353), .Y(n_397) );
INVx2_ASAP7_75t_L g440 ( .A(n_353), .Y(n_440) );
OR2x2_ASAP7_75t_L g691 ( .A(n_354), .B(n_489), .Y(n_691) );
CKINVDCx5p33_ASAP7_75t_R g1587 ( .A(n_355), .Y(n_1587) );
INVx1_ASAP7_75t_L g1928 ( .A(n_358), .Y(n_1928) );
INVx1_ASAP7_75t_L g964 ( .A(n_359), .Y(n_964) );
INVx1_ASAP7_75t_L g1998 ( .A(n_361), .Y(n_1998) );
INVx1_ASAP7_75t_L g612 ( .A(n_363), .Y(n_612) );
INVx1_ASAP7_75t_L g790 ( .A(n_364), .Y(n_790) );
INVx1_ASAP7_75t_L g1140 ( .A(n_366), .Y(n_1140) );
INVx1_ASAP7_75t_L g1248 ( .A(n_368), .Y(n_1248) );
INVx1_ASAP7_75t_L g713 ( .A(n_370), .Y(n_713) );
INVx1_ASAP7_75t_L g1152 ( .A(n_371), .Y(n_1152) );
INVx1_ASAP7_75t_L g590 ( .A(n_373), .Y(n_590) );
INVxp33_ASAP7_75t_L g1929 ( .A(n_374), .Y(n_1929) );
INVxp67_ASAP7_75t_SL g423 ( .A(n_375), .Y(n_423) );
AOI21xp5_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_398), .B(n_1668), .Y(n_376) );
BUFx3_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
BUFx3_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
AND2x4_ASAP7_75t_L g379 ( .A(n_380), .B(n_385), .Y(n_379) );
AND2x4_ASAP7_75t_L g1967 ( .A(n_380), .B(n_386), .Y(n_1967) );
NOR2xp33_ASAP7_75t_SL g380 ( .A(n_381), .B(n_383), .Y(n_380) );
INVx1_ASAP7_75t_SL g1963 ( .A(n_381), .Y(n_1963) );
NAND2xp5_ASAP7_75t_L g2059 ( .A(n_381), .B(n_383), .Y(n_2059) );
HB1xp67_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_L g1962 ( .A(n_383), .B(n_1963), .Y(n_1962) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
NOR2xp33_ASAP7_75t_L g386 ( .A(n_387), .B(n_391), .Y(n_386) );
INVxp67_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
OR2x6_ASAP7_75t_L g2055 ( .A(n_388), .B(n_493), .Y(n_2055) );
HB1xp67_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
AND2x2_ASAP7_75t_L g463 ( .A(n_389), .B(n_397), .Y(n_463) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
OR2x2_ASAP7_75t_L g654 ( .A(n_390), .B(n_655), .Y(n_654) );
INVx8_ASAP7_75t_L g2039 ( .A(n_391), .Y(n_2039) );
OR2x6_ASAP7_75t_L g391 ( .A(n_392), .B(n_396), .Y(n_391) );
OR2x2_ASAP7_75t_L g490 ( .A(n_392), .B(n_417), .Y(n_490) );
INVx2_ASAP7_75t_SL g658 ( .A(n_392), .Y(n_658) );
BUFx6f_ASAP7_75t_L g682 ( .A(n_392), .Y(n_682) );
BUFx2_ASAP7_75t_L g940 ( .A(n_392), .Y(n_940) );
INVx1_ASAP7_75t_L g953 ( .A(n_392), .Y(n_953) );
OAI22xp33_ASAP7_75t_L g1043 ( .A1(n_392), .A2(n_684), .B1(n_1044), .B2(n_1045), .Y(n_1043) );
OAI22xp33_ASAP7_75t_L g1057 ( .A1(n_392), .A2(n_684), .B1(n_1058), .B2(n_1059), .Y(n_1057) );
INVx2_ASAP7_75t_SL g1184 ( .A(n_392), .Y(n_1184) );
OR2x6_ASAP7_75t_L g2042 ( .A(n_392), .B(n_2043), .Y(n_2042) );
BUFx6f_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_394), .B(n_395), .Y(n_393) );
INVx1_ASAP7_75t_L g415 ( .A(n_394), .Y(n_415) );
INVx1_ASAP7_75t_L g428 ( .A(n_394), .Y(n_428) );
AND2x4_ASAP7_75t_L g436 ( .A(n_394), .B(n_429), .Y(n_436) );
AND2x2_ASAP7_75t_L g449 ( .A(n_394), .B(n_395), .Y(n_449) );
INVx2_ASAP7_75t_L g454 ( .A(n_394), .Y(n_454) );
INVx1_ASAP7_75t_L g422 ( .A(n_395), .Y(n_422) );
INVx2_ASAP7_75t_L g429 ( .A(n_395), .Y(n_429) );
INVx1_ASAP7_75t_L g456 ( .A(n_395), .Y(n_456) );
INVx1_ASAP7_75t_L g664 ( .A(n_395), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_395), .B(n_454), .Y(n_670) );
AND2x4_ASAP7_75t_L g2033 ( .A(n_396), .B(n_422), .Y(n_2033) );
INVx2_ASAP7_75t_SL g396 ( .A(n_397), .Y(n_396) );
OAI21xp33_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_1416), .B(n_1667), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g1667 ( .A(n_399), .B(n_1416), .Y(n_1667) );
AOI22x1_ASAP7_75t_L g399 ( .A1(n_400), .A2(n_401), .B1(n_1135), .B2(n_1415), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
XNOR2x1_ASAP7_75t_L g401 ( .A(n_402), .B(n_582), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx2_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_408), .B(n_487), .Y(n_407) );
AND4x1_ASAP7_75t_L g408 ( .A(n_409), .B(n_430), .C(n_444), .D(n_457), .Y(n_408) );
AOI221xp5_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_419), .B1(n_420), .B2(n_423), .C(n_424), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
AOI221xp5_ASAP7_75t_L g741 ( .A1(n_412), .A2(n_420), .B1(n_425), .B2(n_710), .C(n_711), .Y(n_741) );
AOI221xp5_ASAP7_75t_L g832 ( .A1(n_412), .A2(n_420), .B1(n_425), .B2(n_833), .C(n_834), .Y(n_832) );
AOI221xp5_ASAP7_75t_L g1037 ( .A1(n_412), .A2(n_420), .B1(n_425), .B2(n_1038), .C(n_1039), .Y(n_1037) );
HB1xp67_ASAP7_75t_L g1090 ( .A(n_412), .Y(n_1090) );
AOI221xp5_ASAP7_75t_L g1292 ( .A1(n_412), .A2(n_420), .B1(n_425), .B2(n_1293), .C(n_1294), .Y(n_1292) );
AOI221xp5_ASAP7_75t_L g1521 ( .A1(n_412), .A2(n_420), .B1(n_425), .B2(n_1522), .C(n_1523), .Y(n_1521) );
AND2x4_ASAP7_75t_L g412 ( .A(n_413), .B(n_416), .Y(n_412) );
AND2x4_ASAP7_75t_L g2034 ( .A(n_413), .B(n_2035), .Y(n_2034) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
AND2x2_ASAP7_75t_L g663 ( .A(n_415), .B(n_664), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_415), .B(n_664), .Y(n_685) );
AND2x4_ASAP7_75t_L g420 ( .A(n_416), .B(n_421), .Y(n_420) );
AND2x4_ASAP7_75t_L g425 ( .A(n_416), .B(n_426), .Y(n_425) );
NAND2x1_ASAP7_75t_SL g643 ( .A(n_416), .B(n_644), .Y(n_643) );
NAND2x1p5_ASAP7_75t_L g647 ( .A(n_416), .B(n_648), .Y(n_647) );
NAND2x1p5_ASAP7_75t_L g651 ( .A(n_416), .B(n_443), .Y(n_651) );
INVx3_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g962 ( .A(n_418), .Y(n_962) );
INVx1_ASAP7_75t_L g1093 ( .A(n_420), .Y(n_1093) );
AOI21xp5_ASAP7_75t_L g1473 ( .A1(n_420), .A2(n_425), .B(n_1449), .Y(n_1473) );
AND2x2_ASAP7_75t_L g1200 ( .A(n_421), .B(n_960), .Y(n_1200) );
AND2x2_ASAP7_75t_L g1388 ( .A(n_421), .B(n_960), .Y(n_1388) );
HB1xp67_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g645 ( .A(n_422), .Y(n_645) );
HB1xp67_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
AOI221xp5_ASAP7_75t_L g1089 ( .A1(n_425), .A2(n_1090), .B1(n_1091), .B2(n_1092), .C(n_1094), .Y(n_1089) );
INVx1_ASAP7_75t_L g847 ( .A(n_426), .Y(n_847) );
AOI22xp33_ASAP7_75t_L g1051 ( .A1(n_426), .A2(n_447), .B1(n_1052), .B2(n_1053), .Y(n_1051) );
HB1xp67_ASAP7_75t_L g1540 ( .A(n_426), .Y(n_1540) );
BUFx2_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
BUFx3_ASAP7_75t_L g443 ( .A(n_427), .Y(n_443) );
BUFx3_ASAP7_75t_L g468 ( .A(n_427), .Y(n_468) );
BUFx6f_ASAP7_75t_L g480 ( .A(n_427), .Y(n_480) );
BUFx6f_ASAP7_75t_L g999 ( .A(n_427), .Y(n_999) );
AND2x4_ASAP7_75t_L g2045 ( .A(n_427), .B(n_2046), .Y(n_2045) );
AND2x4_ASAP7_75t_L g427 ( .A(n_428), .B(n_429), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g430 ( .A1(n_431), .A2(n_432), .B1(n_441), .B2(n_442), .Y(n_430) );
AOI22xp33_ASAP7_75t_L g1317 ( .A1(n_432), .A2(n_442), .B1(n_1318), .B2(n_1319), .Y(n_1317) );
BUFx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
BUFx2_ASAP7_75t_L g759 ( .A(n_433), .Y(n_759) );
BUFx2_ASAP7_75t_L g837 ( .A(n_433), .Y(n_837) );
BUFx2_ASAP7_75t_L g1097 ( .A(n_433), .Y(n_1097) );
BUFx2_ASAP7_75t_L g1532 ( .A(n_433), .Y(n_1532) );
AND2x4_ASAP7_75t_L g433 ( .A(n_434), .B(n_437), .Y(n_433) );
INVx2_ASAP7_75t_L g672 ( .A(n_434), .Y(n_672) );
INVx1_ASAP7_75t_SL g996 ( .A(n_434), .Y(n_996) );
BUFx3_ASAP7_75t_L g1538 ( .A(n_434), .Y(n_1538) );
INVx3_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx3_ASAP7_75t_L g633 ( .A(n_435), .Y(n_633) );
BUFx6f_ASAP7_75t_L g787 ( .A(n_435), .Y(n_787) );
INVx3_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
BUFx6f_ASAP7_75t_L g474 ( .A(n_436), .Y(n_474) );
INVx1_ASAP7_75t_L g680 ( .A(n_436), .Y(n_680) );
INVx1_ASAP7_75t_L g2053 ( .A(n_436), .Y(n_2053) );
AND2x6_ASAP7_75t_L g442 ( .A(n_437), .B(n_443), .Y(n_442) );
AND2x4_ASAP7_75t_L g446 ( .A(n_437), .B(n_447), .Y(n_446) );
AND2x2_ASAP7_75t_L g451 ( .A(n_437), .B(n_452), .Y(n_451) );
AND2x2_ASAP7_75t_L g632 ( .A(n_437), .B(n_633), .Y(n_632) );
AND2x2_ASAP7_75t_L g635 ( .A(n_437), .B(n_480), .Y(n_635) );
AND2x2_ASAP7_75t_L g639 ( .A(n_437), .B(n_452), .Y(n_639) );
AND2x2_ASAP7_75t_L g764 ( .A(n_437), .B(n_452), .Y(n_764) );
AND2x2_ASAP7_75t_L g992 ( .A(n_437), .B(n_963), .Y(n_992) );
AOI22xp5_ASAP7_75t_L g1048 ( .A1(n_437), .A2(n_739), .B1(n_1049), .B2(n_1054), .Y(n_1048) );
AND2x2_ASAP7_75t_L g1301 ( .A(n_437), .B(n_452), .Y(n_1301) );
AND2x4_ASAP7_75t_L g437 ( .A(n_438), .B(n_439), .Y(n_437) );
INVx1_ASAP7_75t_L g483 ( .A(n_438), .Y(n_483) );
OR2x2_ASAP7_75t_L g977 ( .A(n_438), .B(n_514), .Y(n_977) );
INVx2_ASAP7_75t_L g927 ( .A(n_439), .Y(n_927) );
AND2x4_ASAP7_75t_L g969 ( .A(n_439), .B(n_738), .Y(n_969) );
AND2x2_ASAP7_75t_L g971 ( .A(n_439), .B(n_453), .Y(n_971) );
INVx1_ASAP7_75t_L g485 ( .A(n_440), .Y(n_485) );
INVx1_ASAP7_75t_L g655 ( .A(n_440), .Y(n_655) );
OAI221xp5_ASAP7_75t_L g534 ( .A1(n_441), .A2(n_445), .B1(n_535), .B2(n_540), .C(n_543), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g757 ( .A1(n_442), .A2(n_758), .B1(n_759), .B2(n_760), .Y(n_757) );
AOI22xp33_ASAP7_75t_L g835 ( .A1(n_442), .A2(n_836), .B1(n_837), .B2(n_838), .Y(n_835) );
AOI22xp33_ASAP7_75t_L g1095 ( .A1(n_442), .A2(n_1096), .B1(n_1097), .B2(n_1098), .Y(n_1095) );
AOI22xp33_ASAP7_75t_L g1295 ( .A1(n_442), .A2(n_837), .B1(n_1296), .B2(n_1297), .Y(n_1295) );
BUFx2_ASAP7_75t_L g1527 ( .A(n_442), .Y(n_1527) );
AOI22xp33_ASAP7_75t_L g1648 ( .A1(n_442), .A2(n_1097), .B1(n_1635), .B2(n_1649), .Y(n_1648) );
AOI22xp33_ASAP7_75t_L g1924 ( .A1(n_442), .A2(n_1532), .B1(n_1925), .B2(n_1926), .Y(n_1924) );
BUFx2_ASAP7_75t_L g1604 ( .A(n_443), .Y(n_1604) );
AOI22xp33_ASAP7_75t_L g444 ( .A1(n_445), .A2(n_446), .B1(n_450), .B2(n_451), .Y(n_444) );
AOI22xp33_ASAP7_75t_L g636 ( .A1(n_446), .A2(n_637), .B1(n_638), .B2(n_639), .Y(n_636) );
AOI221xp5_ASAP7_75t_L g742 ( .A1(n_446), .A2(n_451), .B1(n_743), .B2(n_744), .C(n_745), .Y(n_742) );
AOI22xp33_ASAP7_75t_L g761 ( .A1(n_446), .A2(n_762), .B1(n_763), .B2(n_764), .Y(n_761) );
AOI22xp33_ASAP7_75t_L g839 ( .A1(n_446), .A2(n_764), .B1(n_840), .B2(n_841), .Y(n_839) );
AOI22xp33_ASAP7_75t_L g1099 ( .A1(n_446), .A2(n_764), .B1(n_1100), .B2(n_1101), .Y(n_1099) );
AOI22xp33_ASAP7_75t_L g1298 ( .A1(n_446), .A2(n_1299), .B1(n_1300), .B2(n_1301), .Y(n_1298) );
AOI22xp33_ASAP7_75t_L g1320 ( .A1(n_446), .A2(n_451), .B1(n_1321), .B2(n_1322), .Y(n_1320) );
INVx1_ASAP7_75t_L g1471 ( .A(n_446), .Y(n_1471) );
BUFx2_ASAP7_75t_L g1530 ( .A(n_446), .Y(n_1530) );
AOI22xp33_ASAP7_75t_L g1650 ( .A1(n_446), .A2(n_764), .B1(n_1636), .B2(n_1651), .Y(n_1650) );
AOI22xp33_ASAP7_75t_L g1927 ( .A1(n_446), .A2(n_1301), .B1(n_1928), .B2(n_1929), .Y(n_1927) );
BUFx3_ASAP7_75t_L g465 ( .A(n_447), .Y(n_465) );
BUFx2_ASAP7_75t_L g725 ( .A(n_447), .Y(n_725) );
INVx2_ASAP7_75t_SL g447 ( .A(n_448), .Y(n_447) );
INVx2_ASAP7_75t_SL g963 ( .A(n_448), .Y(n_963) );
INVx2_ASAP7_75t_L g1514 ( .A(n_448), .Y(n_1514) );
INVx3_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
BUFx6f_ASAP7_75t_L g738 ( .A(n_449), .Y(n_738) );
BUFx6f_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
BUFx6f_ASAP7_75t_L g471 ( .A(n_453), .Y(n_471) );
INVx1_ASAP7_75t_L g728 ( .A(n_453), .Y(n_728) );
BUFx2_ASAP7_75t_L g849 ( .A(n_453), .Y(n_849) );
BUFx6f_ASAP7_75t_L g1042 ( .A(n_453), .Y(n_1042) );
AND2x4_ASAP7_75t_L g453 ( .A(n_454), .B(n_455), .Y(n_453) );
INVx1_ASAP7_75t_L g649 ( .A(n_454), .Y(n_649) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
AOI33xp33_ASAP7_75t_L g457 ( .A1(n_458), .A2(n_464), .A3(n_469), .B1(n_475), .B2(n_478), .B3(n_481), .Y(n_457) );
AOI33xp33_ASAP7_75t_L g1102 ( .A1(n_458), .A2(n_481), .A3(n_1103), .B1(n_1104), .B2(n_1105), .B3(n_1106), .Y(n_1102) );
AOI33xp33_ASAP7_75t_L g1302 ( .A1(n_458), .A2(n_481), .A3(n_1303), .B1(n_1306), .B2(n_1308), .B3(n_1309), .Y(n_1302) );
AOI33xp33_ASAP7_75t_L g1533 ( .A1(n_458), .A2(n_1534), .A3(n_1539), .B1(n_1541), .B2(n_1542), .B3(n_1543), .Y(n_1533) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
AND2x4_ASAP7_75t_L g460 ( .A(n_461), .B(n_463), .Y(n_460) );
BUFx2_ASAP7_75t_L g580 ( .A(n_461), .Y(n_580) );
INVx2_ASAP7_75t_L g720 ( .A(n_461), .Y(n_720) );
AND2x4_ASAP7_75t_L g723 ( .A(n_461), .B(n_463), .Y(n_723) );
AND2x2_ASAP7_75t_L g739 ( .A(n_461), .B(n_740), .Y(n_739) );
OR2x6_ASAP7_75t_L g895 ( .A(n_461), .B(n_896), .Y(n_895) );
OR2x2_ASAP7_75t_L g1480 ( .A(n_461), .B(n_1481), .Y(n_1480) );
OR2x2_ASAP7_75t_L g2022 ( .A(n_461), .B(n_896), .Y(n_2022) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
OR2x6_ASAP7_75t_L g653 ( .A(n_462), .B(n_654), .Y(n_653) );
BUFx2_ASAP7_75t_L g973 ( .A(n_462), .Y(n_973) );
INVx1_ASAP7_75t_L g943 ( .A(n_463), .Y(n_943) );
BUFx2_ASAP7_75t_SL g1254 ( .A(n_463), .Y(n_1254) );
HB1xp67_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
BUFx6f_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
AND2x4_ASAP7_75t_L g929 ( .A(n_468), .B(n_926), .Y(n_929) );
BUFx3_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx2_ASAP7_75t_SL g472 ( .A(n_473), .Y(n_472) );
OAI22xp5_ASAP7_75t_L g1341 ( .A1(n_473), .A2(n_952), .B1(n_1342), .B2(n_1343), .Y(n_1341) );
OAI22xp33_ASAP7_75t_L g1427 ( .A1(n_473), .A2(n_1428), .B1(n_1429), .B2(n_1430), .Y(n_1427) );
OAI221xp5_ASAP7_75t_L g1599 ( .A1(n_473), .A2(n_1600), .B1(n_1601), .B2(n_1602), .C(n_1603), .Y(n_1599) );
OAI22xp5_ASAP7_75t_L g1664 ( .A1(n_473), .A2(n_1630), .B1(n_1644), .B2(n_1665), .Y(n_1664) );
INVx2_ASAP7_75t_L g2006 ( .A(n_473), .Y(n_2006) );
INVx4_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx2_ASAP7_75t_SL g477 ( .A(n_474), .Y(n_477) );
INVx2_ASAP7_75t_SL g851 ( .A(n_474), .Y(n_851) );
INVx2_ASAP7_75t_SL g934 ( .A(n_474), .Y(n_934) );
BUFx3_ASAP7_75t_L g1307 ( .A(n_474), .Y(n_1307) );
INVx2_ASAP7_75t_SL g1369 ( .A(n_474), .Y(n_1369) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
OAI22xp5_ASAP7_75t_SL g1255 ( .A1(n_477), .A2(n_1192), .B1(n_1256), .B2(n_1257), .Y(n_1255) );
OAI22xp5_ASAP7_75t_L g1381 ( .A1(n_477), .A2(n_1382), .B1(n_1384), .B2(n_1385), .Y(n_1381) );
BUFx6f_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx2_ASAP7_75t_SL g857 ( .A(n_480), .Y(n_857) );
INVx2_ASAP7_75t_L g686 ( .A(n_481), .Y(n_686) );
AOI33xp33_ASAP7_75t_L g842 ( .A1(n_481), .A2(n_723), .A3(n_843), .B1(n_848), .B2(n_852), .B3(n_853), .Y(n_842) );
INVx6_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx5_ASAP7_75t_L g796 ( .A(n_482), .Y(n_796) );
OR2x6_ASAP7_75t_L g482 ( .A(n_483), .B(n_484), .Y(n_482) );
NAND2x1p5_ASAP7_75t_L g913 ( .A(n_483), .B(n_495), .Y(n_913) );
INVx2_ASAP7_75t_L g740 ( .A(n_484), .Y(n_740) );
BUFx2_ASAP7_75t_L g1246 ( .A(n_484), .Y(n_1246) );
NAND2x1p5_ASAP7_75t_L g484 ( .A(n_485), .B(n_486), .Y(n_484) );
INVx1_ASAP7_75t_L g2036 ( .A(n_485), .Y(n_2036) );
AOI21xp33_ASAP7_75t_SL g487 ( .A1(n_488), .A2(n_505), .B(n_506), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx2_ASAP7_75t_SL g627 ( .A(n_489), .Y(n_627) );
INVx5_ASAP7_75t_L g754 ( .A(n_489), .Y(n_754) );
INVx2_ASAP7_75t_L g1545 ( .A(n_489), .Y(n_1545) );
AND2x4_ASAP7_75t_L g489 ( .A(n_490), .B(n_491), .Y(n_489) );
INVx2_ASAP7_75t_L g1047 ( .A(n_490), .Y(n_1047) );
INVx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
AOI222xp33_ASAP7_75t_L g974 ( .A1(n_492), .A2(n_949), .B1(n_954), .B2(n_964), .C1(n_975), .C2(n_978), .Y(n_974) );
OR2x6_ASAP7_75t_L g1144 ( .A(n_492), .B(n_1145), .Y(n_1144) );
AND2x4_ASAP7_75t_L g492 ( .A(n_493), .B(n_494), .Y(n_492) );
AND2x4_ASAP7_75t_L g909 ( .A(n_493), .B(n_545), .Y(n_909) );
AND2x4_ASAP7_75t_L g1488 ( .A(n_493), .B(n_545), .Y(n_1488) );
INVx2_ASAP7_75t_L g1081 ( .A(n_494), .Y(n_1081) );
AND2x2_ASAP7_75t_L g494 ( .A(n_495), .B(n_500), .Y(n_494) );
AND2x4_ASAP7_75t_L g517 ( .A(n_495), .B(n_518), .Y(n_517) );
INVx1_ASAP7_75t_L g522 ( .A(n_495), .Y(n_522) );
BUFx2_ASAP7_75t_L g608 ( .A(n_495), .Y(n_608) );
AND2x4_ASAP7_75t_L g623 ( .A(n_495), .B(n_518), .Y(n_623) );
AND2x4_ASAP7_75t_L g625 ( .A(n_495), .B(n_524), .Y(n_625) );
AND2x2_ASAP7_75t_L g866 ( .A(n_495), .B(n_524), .Y(n_866) );
AND2x2_ASAP7_75t_L g1281 ( .A(n_495), .B(n_524), .Y(n_1281) );
AND2x4_ASAP7_75t_L g495 ( .A(n_496), .B(n_498), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
AND2x4_ASAP7_75t_L g545 ( .A(n_498), .B(n_546), .Y(n_545) );
INVx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
AND2x2_ASAP7_75t_L g556 ( .A(n_499), .B(n_546), .Y(n_556) );
INVx1_ASAP7_75t_L g1977 ( .A(n_499), .Y(n_1977) );
HB1xp67_ASAP7_75t_L g1984 ( .A(n_499), .Y(n_1984) );
INVx1_ASAP7_75t_L g1988 ( .A(n_499), .Y(n_1988) );
INVx6_ASAP7_75t_L g560 ( .A(n_500), .Y(n_560) );
INVx2_ASAP7_75t_L g615 ( .A(n_500), .Y(n_615) );
BUFx2_ASAP7_75t_L g1568 ( .A(n_500), .Y(n_1568) );
AND2x4_ASAP7_75t_L g1982 ( .A(n_500), .B(n_1983), .Y(n_1982) );
AND2x4_ASAP7_75t_L g500 ( .A(n_501), .B(n_503), .Y(n_500) );
INVx1_ASAP7_75t_L g525 ( .A(n_501), .Y(n_525) );
INVx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
AND2x4_ASAP7_75t_L g511 ( .A(n_502), .B(n_512), .Y(n_511) );
AND2x2_ASAP7_75t_L g554 ( .A(n_502), .B(n_504), .Y(n_554) );
INVx1_ASAP7_75t_L g520 ( .A(n_503), .Y(n_520) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
AND2x4_ASAP7_75t_L g530 ( .A(n_504), .B(n_531), .Y(n_530) );
AOI31xp33_ASAP7_75t_L g506 ( .A1(n_507), .A2(n_547), .A3(n_570), .B(n_578), .Y(n_506) );
AOI211xp5_ASAP7_75t_L g507 ( .A1(n_508), .A2(n_509), .B(n_515), .C(n_526), .Y(n_507) );
INVx1_ASAP7_75t_L g809 ( .A(n_509), .Y(n_809) );
AOI21xp33_ASAP7_75t_SL g861 ( .A1(n_509), .A2(n_862), .B(n_863), .Y(n_861) );
AOI211xp5_ASAP7_75t_L g1110 ( .A1(n_509), .A2(n_1111), .B(n_1112), .C(n_1113), .Y(n_1110) );
AOI221xp5_ASAP7_75t_L g1272 ( .A1(n_509), .A2(n_1273), .B1(n_1275), .B2(n_1277), .C(n_1278), .Y(n_1272) );
AOI211xp5_ASAP7_75t_L g1347 ( .A1(n_509), .A2(n_1339), .B(n_1348), .C(n_1349), .Y(n_1347) );
AOI211xp5_ASAP7_75t_L g1548 ( .A1(n_509), .A2(n_1549), .B(n_1550), .C(n_1552), .Y(n_1548) );
AOI211xp5_ASAP7_75t_SL g1629 ( .A1(n_509), .A2(n_1630), .B(n_1631), .C(n_1633), .Y(n_1629) );
AOI211xp5_ASAP7_75t_SL g1950 ( .A1(n_509), .A2(n_1941), .B(n_1951), .C(n_1952), .Y(n_1950) );
AND2x4_ASAP7_75t_L g509 ( .A(n_510), .B(n_513), .Y(n_509) );
INVx2_ASAP7_75t_SL g1159 ( .A(n_510), .Y(n_1159) );
BUFx3_ASAP7_75t_L g1232 ( .A(n_510), .Y(n_1232) );
BUFx6f_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
BUFx6f_ASAP7_75t_L g533 ( .A(n_511), .Y(n_533) );
INVx2_ASAP7_75t_SL g550 ( .A(n_511), .Y(n_550) );
BUFx6f_ASAP7_75t_L g597 ( .A(n_511), .Y(n_597) );
BUFx6f_ASAP7_75t_L g611 ( .A(n_511), .Y(n_611) );
HB1xp67_ASAP7_75t_L g618 ( .A(n_511), .Y(n_618) );
HB1xp67_ASAP7_75t_L g816 ( .A(n_511), .Y(n_816) );
BUFx3_ASAP7_75t_L g1170 ( .A(n_511), .Y(n_1170) );
BUFx2_ASAP7_75t_L g1561 ( .A(n_511), .Y(n_1561) );
AND2x6_ASAP7_75t_L g1979 ( .A(n_511), .B(n_1976), .Y(n_1979) );
INVx1_ASAP7_75t_L g539 ( .A(n_512), .Y(n_539) );
AND2x4_ASAP7_75t_L g564 ( .A(n_513), .B(n_553), .Y(n_564) );
AND2x2_ASAP7_75t_L g610 ( .A(n_513), .B(n_611), .Y(n_610) );
AOI222xp33_ASAP7_75t_L g1061 ( .A1(n_513), .A2(n_623), .B1(n_625), .B2(n_1038), .C1(n_1039), .C2(n_1062), .Y(n_1061) );
AOI221xp5_ASAP7_75t_L g1451 ( .A1(n_513), .A2(n_564), .B1(n_607), .B2(n_1439), .C(n_1452), .Y(n_1451) );
INVx2_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
OR2x2_ASAP7_75t_L g573 ( .A(n_514), .B(n_542), .Y(n_573) );
OR2x2_ASAP7_75t_L g576 ( .A(n_514), .B(n_577), .Y(n_576) );
INVx2_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g810 ( .A1(n_517), .A2(n_811), .B1(n_812), .B2(n_813), .Y(n_810) );
INVx1_ASAP7_75t_L g1279 ( .A(n_517), .Y(n_1279) );
INVx2_ASAP7_75t_SL g1551 ( .A(n_517), .Y(n_1551) );
AOI22xp5_ASAP7_75t_L g1029 ( .A1(n_518), .A2(n_524), .B1(n_1030), .B2(n_1031), .Y(n_1029) );
INVx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g917 ( .A(n_519), .Y(n_917) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g1997 ( .A(n_520), .Y(n_1997) );
INVx1_ASAP7_75t_L g812 ( .A(n_521), .Y(n_812) );
OR2x2_ASAP7_75t_L g521 ( .A(n_522), .B(n_523), .Y(n_521) );
INVx1_ASAP7_75t_SL g567 ( .A(n_522), .Y(n_567) );
OR2x6_ASAP7_75t_L g912 ( .A(n_523), .B(n_913), .Y(n_912) );
OR2x2_ASAP7_75t_L g1175 ( .A(n_523), .B(n_913), .Y(n_1175) );
INVx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
BUFx3_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
AND2x6_ASAP7_75t_L g1999 ( .A(n_525), .B(n_1977), .Y(n_1999) );
BUFx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
OR2x6_ASAP7_75t_L g979 ( .A(n_529), .B(n_977), .Y(n_979) );
OR2x2_ASAP7_75t_L g1263 ( .A(n_529), .B(n_977), .Y(n_1263) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
BUFx6f_ASAP7_75t_L g562 ( .A(n_530), .Y(n_562) );
INVx2_ASAP7_75t_L g577 ( .A(n_530), .Y(n_577) );
BUFx6f_ASAP7_75t_L g606 ( .A(n_530), .Y(n_606) );
INVx1_ASAP7_75t_L g1227 ( .A(n_530), .Y(n_1227) );
INVx1_ASAP7_75t_L g538 ( .A(n_531), .Y(n_538) );
BUFx3_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
BUFx2_ASAP7_75t_L g898 ( .A(n_533), .Y(n_898) );
INVx1_ASAP7_75t_L g1115 ( .A(n_533), .Y(n_1115) );
INVx2_ASAP7_75t_L g2018 ( .A(n_533), .Y(n_2018) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx2_ASAP7_75t_SL g1990 ( .A(n_536), .Y(n_1990) );
BUFx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
BUFx4f_ASAP7_75t_L g703 ( .A(n_537), .Y(n_703) );
INVx2_ASAP7_75t_L g985 ( .A(n_537), .Y(n_985) );
INVx1_ASAP7_75t_L g1021 ( .A(n_537), .Y(n_1021) );
INVx1_ASAP7_75t_L g1028 ( .A(n_537), .Y(n_1028) );
INVx1_ASAP7_75t_L g1155 ( .A(n_537), .Y(n_1155) );
AND2x2_ASAP7_75t_L g537 ( .A(n_538), .B(n_539), .Y(n_537) );
OR2x2_ASAP7_75t_L g542 ( .A(n_538), .B(n_539), .Y(n_542) );
OAI22xp5_ASAP7_75t_L g1015 ( .A1(n_540), .A2(n_997), .B1(n_1016), .B2(n_1017), .Y(n_1015) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx2_ASAP7_75t_L g696 ( .A(n_542), .Y(n_696) );
INVx1_ASAP7_75t_L g1064 ( .A(n_542), .Y(n_1064) );
BUFx2_ASAP7_75t_L g1151 ( .A(n_542), .Y(n_1151) );
OR2x2_ASAP7_75t_L g1974 ( .A(n_542), .B(n_1975), .Y(n_1974) );
INVx1_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
BUFx2_ASAP7_75t_L g824 ( .A(n_544), .Y(n_824) );
INVx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx2_ASAP7_75t_SL g616 ( .A(n_545), .Y(n_616) );
CKINVDCx5p33_ASAP7_75t_R g1024 ( .A(n_545), .Y(n_1024) );
HB1xp67_ASAP7_75t_L g1118 ( .A(n_545), .Y(n_1118) );
INVx1_ASAP7_75t_L g1468 ( .A(n_545), .Y(n_1468) );
OAI221xp5_ASAP7_75t_L g1634 ( .A1(n_545), .A2(n_1028), .B1(n_1209), .B2(n_1635), .C(n_1636), .Y(n_1634) );
OAI221xp5_ASAP7_75t_L g1953 ( .A1(n_545), .A2(n_1028), .B1(n_1209), .B2(n_1926), .C(n_1928), .Y(n_1953) );
INVx1_ASAP7_75t_L g2002 ( .A(n_546), .Y(n_2002) );
AOI221xp5_ASAP7_75t_L g547 ( .A1(n_548), .A2(n_557), .B1(n_563), .B2(n_565), .C(n_566), .Y(n_547) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx2_ASAP7_75t_L g982 ( .A(n_550), .Y(n_982) );
INVx2_ASAP7_75t_SL g1483 ( .A(n_550), .Y(n_1483) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx1_ASAP7_75t_L g1466 ( .A(n_552), .Y(n_1466) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
AND2x4_ASAP7_75t_L g607 ( .A(n_553), .B(n_608), .Y(n_607) );
BUFx6f_ASAP7_75t_L g823 ( .A(n_553), .Y(n_823) );
AOI22xp5_ASAP7_75t_L g1065 ( .A1(n_553), .A2(n_611), .B1(n_1059), .B2(n_1066), .Y(n_1065) );
INVx2_ASAP7_75t_SL g1070 ( .A(n_553), .Y(n_1070) );
BUFx3_ASAP7_75t_L g1405 ( .A(n_553), .Y(n_1405) );
BUFx4f_ASAP7_75t_L g1456 ( .A(n_553), .Y(n_1456) );
BUFx6f_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
BUFx6f_ASAP7_75t_L g569 ( .A(n_554), .Y(n_569) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
BUFx3_ASAP7_75t_L g601 ( .A(n_556), .Y(n_601) );
INVx2_ASAP7_75t_SL g705 ( .A(n_556), .Y(n_705) );
INVx2_ASAP7_75t_L g896 ( .A(n_556), .Y(n_896) );
INVx1_ASAP7_75t_L g1481 ( .A(n_556), .Y(n_1481) );
HB1xp67_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
BUFx6f_ASAP7_75t_L g604 ( .A(n_560), .Y(n_604) );
INVx2_ASAP7_75t_L g820 ( .A(n_560), .Y(n_820) );
INVx2_ASAP7_75t_SL g871 ( .A(n_560), .Y(n_871) );
INVx2_ASAP7_75t_L g882 ( .A(n_560), .Y(n_882) );
INVx1_ASAP7_75t_L g1467 ( .A(n_560), .Y(n_1467) );
HB1xp67_ASAP7_75t_L g2026 ( .A(n_560), .Y(n_2026) );
BUFx3_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g698 ( .A(n_562), .Y(n_698) );
BUFx6f_ASAP7_75t_L g1233 ( .A(n_562), .Y(n_1233) );
INVx1_ASAP7_75t_L g2020 ( .A(n_562), .Y(n_2020) );
INVx1_ASAP7_75t_L g799 ( .A(n_563), .Y(n_799) );
AOI221xp5_ASAP7_75t_L g872 ( .A1(n_563), .A2(n_566), .B1(n_873), .B2(n_874), .C(n_880), .Y(n_872) );
AOI221xp5_ASAP7_75t_L g1119 ( .A1(n_563), .A2(n_566), .B1(n_1120), .B2(n_1121), .C(n_1126), .Y(n_1119) );
AOI221xp5_ASAP7_75t_L g1282 ( .A1(n_563), .A2(n_566), .B1(n_1283), .B2(n_1286), .C(n_1287), .Y(n_1282) );
AOI221xp5_ASAP7_75t_L g1352 ( .A1(n_563), .A2(n_566), .B1(n_1340), .B2(n_1353), .C(n_1356), .Y(n_1352) );
BUFx6f_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx2_ASAP7_75t_SL g594 ( .A(n_564), .Y(n_594) );
HB1xp67_ASAP7_75t_L g1558 ( .A(n_564), .Y(n_1558) );
AOI221xp5_ASAP7_75t_L g1637 ( .A1(n_564), .A2(n_607), .B1(n_1638), .B2(n_1639), .C(n_1641), .Y(n_1637) );
HB1xp67_ASAP7_75t_L g1955 ( .A(n_564), .Y(n_1955) );
INVx1_ASAP7_75t_L g807 ( .A(n_566), .Y(n_807) );
AOI221xp5_ASAP7_75t_L g1557 ( .A1(n_566), .A2(n_1558), .B1(n_1559), .B2(n_1560), .C(n_1566), .Y(n_1557) );
AND2x4_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .Y(n_566) );
INVx1_ASAP7_75t_L g902 ( .A(n_568), .Y(n_902) );
INVx1_ASAP7_75t_L g1285 ( .A(n_568), .Y(n_1285) );
BUFx6f_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx2_ASAP7_75t_L g599 ( .A(n_569), .Y(n_599) );
INVx1_ASAP7_75t_L g879 ( .A(n_569), .Y(n_879) );
BUFx6f_ASAP7_75t_L g1077 ( .A(n_569), .Y(n_1077) );
AND2x4_ASAP7_75t_L g1992 ( .A(n_569), .B(n_1993), .Y(n_1992) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_571), .A2(n_572), .B1(n_574), .B2(n_575), .Y(n_570) );
AOI22xp5_ASAP7_75t_L g589 ( .A1(n_572), .A2(n_575), .B1(n_590), .B2(n_591), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g883 ( .A1(n_572), .A2(n_575), .B1(n_884), .B2(n_885), .Y(n_883) );
AOI22xp33_ASAP7_75t_L g1128 ( .A1(n_572), .A2(n_575), .B1(n_1129), .B2(n_1130), .Y(n_1128) );
AOI22xp33_ASAP7_75t_L g1288 ( .A1(n_572), .A2(n_575), .B1(n_1289), .B2(n_1290), .Y(n_1288) );
AOI22xp33_ASAP7_75t_L g1359 ( .A1(n_572), .A2(n_575), .B1(n_1342), .B2(n_1343), .Y(n_1359) );
AOI22xp33_ASAP7_75t_L g1570 ( .A1(n_572), .A2(n_575), .B1(n_1571), .B2(n_1572), .Y(n_1570) );
AOI22xp33_ASAP7_75t_L g1642 ( .A1(n_572), .A2(n_575), .B1(n_1643), .B2(n_1644), .Y(n_1642) );
AOI22xp33_ASAP7_75t_L g1958 ( .A1(n_572), .A2(n_575), .B1(n_1944), .B2(n_1946), .Y(n_1958) );
INVx6_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx4_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g1018 ( .A(n_577), .Y(n_1018) );
INVx2_ASAP7_75t_L g1358 ( .A(n_577), .Y(n_1358) );
AOI31xp33_ASAP7_75t_L g860 ( .A1(n_578), .A2(n_861), .A3(n_872), .B(n_883), .Y(n_860) );
INVx2_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
AOI22xp5_ASAP7_75t_L g587 ( .A1(n_579), .A2(n_588), .B1(n_626), .B2(n_627), .Y(n_587) );
CKINVDCx8_ASAP7_75t_R g579 ( .A(n_580), .Y(n_579) );
OAI31xp33_ASAP7_75t_L g1364 ( .A1(n_580), .A2(n_1365), .A3(n_1366), .B(n_1376), .Y(n_1364) );
XNOR2x1_ASAP7_75t_L g582 ( .A(n_583), .B(n_888), .Y(n_582) );
XNOR2xp5_ASAP7_75t_L g583 ( .A(n_584), .B(n_750), .Y(n_583) );
XOR2x2_ASAP7_75t_L g584 ( .A(n_585), .B(n_689), .Y(n_584) );
INVx1_ASAP7_75t_L g687 ( .A(n_586), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_587), .B(n_628), .Y(n_586) );
NAND3xp33_ASAP7_75t_L g588 ( .A(n_589), .B(n_592), .C(n_609), .Y(n_588) );
OAI22xp33_ASAP7_75t_L g681 ( .A1(n_590), .A2(n_595), .B1(n_682), .B2(n_683), .Y(n_681) );
OAI22xp5_ASAP7_75t_L g674 ( .A1(n_591), .A2(n_612), .B1(n_675), .B2(n_678), .Y(n_674) );
AOI221xp5_ASAP7_75t_L g592 ( .A1(n_593), .A2(n_595), .B1(n_596), .B2(n_602), .C(n_607), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx2_ASAP7_75t_L g876 ( .A(n_597), .Y(n_876) );
BUFx3_ASAP7_75t_L g1459 ( .A(n_597), .Y(n_1459) );
INVx1_ASAP7_75t_L g1563 ( .A(n_598), .Y(n_1563) );
INVx3_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx2_ASAP7_75t_L g1486 ( .A(n_599), .Y(n_1486) );
INVx3_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVxp67_ASAP7_75t_L g1071 ( .A(n_601), .Y(n_1071) );
INVx2_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx4_ASAP7_75t_L g1274 ( .A(n_604), .Y(n_1274) );
HB1xp67_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g620 ( .A(n_606), .Y(n_620) );
BUFx6f_ASAP7_75t_L g804 ( .A(n_606), .Y(n_804) );
INVx2_ASAP7_75t_L g906 ( .A(n_606), .Y(n_906) );
BUFx6f_ASAP7_75t_L g1079 ( .A(n_606), .Y(n_1079) );
INVx1_ASAP7_75t_L g1454 ( .A(n_606), .Y(n_1454) );
AND2x6_ASAP7_75t_L g1986 ( .A(n_606), .B(n_1987), .Y(n_1986) );
INVx1_ASAP7_75t_L g706 ( .A(n_607), .Y(n_706) );
AOI21xp5_ASAP7_75t_L g1067 ( .A1(n_607), .A2(n_1068), .B(n_1072), .Y(n_1067) );
AOI221xp5_ASAP7_75t_L g1954 ( .A1(n_607), .A2(n_1947), .B1(n_1955), .B2(n_1956), .C(n_1957), .Y(n_1954) );
BUFx3_ASAP7_75t_L g1032 ( .A(n_608), .Y(n_1032) );
AOI221xp5_ASAP7_75t_L g609 ( .A1(n_610), .A2(n_612), .B1(n_613), .B2(n_617), .C(n_621), .Y(n_609) );
INVx1_ASAP7_75t_L g708 ( .A(n_610), .Y(n_708) );
INVx1_ASAP7_75t_L g1211 ( .A(n_611), .Y(n_1211) );
BUFx2_ASAP7_75t_L g1225 ( .A(n_611), .Y(n_1225) );
BUFx2_ASAP7_75t_L g900 ( .A(n_614), .Y(n_900) );
AND2x2_ASAP7_75t_L g975 ( .A(n_614), .B(n_976), .Y(n_975) );
A2O1A1Ixp33_ASAP7_75t_L g1025 ( .A1(n_614), .A2(n_1026), .B(n_1027), .C(n_1032), .Y(n_1025) );
INVx2_ASAP7_75t_SL g614 ( .A(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g1127 ( .A(n_615), .Y(n_1127) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g1074 ( .A(n_620), .Y(n_1074) );
INVx1_ASAP7_75t_SL g622 ( .A(n_623), .Y(n_622) );
AOI22xp5_ASAP7_75t_L g709 ( .A1(n_623), .A2(n_625), .B1(n_710), .B2(n_711), .Y(n_709) );
INVx2_ASAP7_75t_L g864 ( .A(n_623), .Y(n_864) );
INVx4_ASAP7_75t_L g1448 ( .A(n_623), .Y(n_1448) );
INVx2_ASAP7_75t_SL g624 ( .A(n_625), .Y(n_624) );
AOI222xp33_ASAP7_75t_SL g1445 ( .A1(n_625), .A2(n_1080), .B1(n_1446), .B2(n_1447), .C1(n_1449), .C2(n_1450), .Y(n_1445) );
INVx2_ASAP7_75t_L g1632 ( .A(n_625), .Y(n_1632) );
NOR3xp33_ASAP7_75t_L g628 ( .A(n_629), .B(n_640), .C(n_652), .Y(n_628) );
NAND2xp5_ASAP7_75t_SL g629 ( .A(n_630), .B(n_636), .Y(n_629) );
AOI22xp33_ASAP7_75t_L g630 ( .A1(n_631), .A2(n_632), .B1(n_634), .B2(n_635), .Y(n_630) );
INVx2_ASAP7_75t_L g746 ( .A(n_632), .Y(n_746) );
INVx2_ASAP7_75t_L g730 ( .A(n_633), .Y(n_730) );
INVx1_ASAP7_75t_L g776 ( .A(n_633), .Y(n_776) );
INVx2_ASAP7_75t_L g1056 ( .A(n_633), .Y(n_1056) );
INVx1_ASAP7_75t_L g747 ( .A(n_635), .Y(n_747) );
INVxp67_ASAP7_75t_L g1442 ( .A(n_635), .Y(n_1442) );
INVx1_ASAP7_75t_L g1006 ( .A(n_639), .Y(n_1006) );
INVx1_ASAP7_75t_L g1425 ( .A(n_639), .Y(n_1425) );
INVx2_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx2_ASAP7_75t_SL g1324 ( .A(n_642), .Y(n_1324) );
INVx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
AOI22xp33_ASAP7_75t_L g966 ( .A1(n_644), .A2(n_648), .B1(n_914), .B2(n_919), .Y(n_966) );
NAND2x1p5_ASAP7_75t_L g1510 ( .A(n_644), .B(n_1511), .Y(n_1510) );
INVx2_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
BUFx4f_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
BUFx4f_ASAP7_75t_L g766 ( .A(n_647), .Y(n_766) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
OR2x6_ASAP7_75t_L g1203 ( .A(n_649), .B(n_961), .Y(n_1203) );
BUFx3_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
BUFx2_ASAP7_75t_L g767 ( .A(n_651), .Y(n_767) );
BUFx2_ASAP7_75t_L g1653 ( .A(n_651), .Y(n_1653) );
OAI33xp33_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_656), .A3(n_666), .B1(n_674), .B2(n_681), .B3(n_686), .Y(n_652) );
OAI33xp33_ASAP7_75t_L g768 ( .A1(n_653), .A2(n_769), .A3(n_778), .B1(n_783), .B2(n_789), .B3(n_795), .Y(n_768) );
OAI33xp33_ASAP7_75t_L g1325 ( .A1(n_653), .A2(n_795), .A3(n_1326), .B1(n_1331), .B2(n_1337), .B3(n_1341), .Y(n_1325) );
OAI33xp33_ASAP7_75t_L g1654 ( .A1(n_653), .A2(n_795), .A3(n_1655), .B1(n_1659), .B2(n_1664), .B3(n_1666), .Y(n_1654) );
OAI33xp33_ASAP7_75t_L g1931 ( .A1(n_653), .A2(n_795), .A3(n_1932), .B1(n_1936), .B2(n_1939), .B3(n_1945), .Y(n_1931) );
INVx1_ASAP7_75t_L g2043 ( .A(n_655), .Y(n_2043) );
OAI22xp33_ASAP7_75t_L g656 ( .A1(n_657), .A2(n_659), .B1(n_660), .B2(n_665), .Y(n_656) );
OAI221xp5_ASAP7_75t_L g1251 ( .A1(n_657), .A2(n_1220), .B1(n_1223), .B2(n_1252), .C(n_1254), .Y(n_1251) );
INVx2_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
OR2x2_ASAP7_75t_L g1189 ( .A(n_662), .B(n_961), .Y(n_1189) );
OR2x6_ASAP7_75t_L g1375 ( .A(n_662), .B(n_961), .Y(n_1375) );
OAI22xp33_ASAP7_75t_L g1431 ( .A1(n_662), .A2(n_1183), .B1(n_1432), .B2(n_1433), .Y(n_1431) );
INVx2_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx3_ASAP7_75t_L g793 ( .A(n_663), .Y(n_793) );
INVx2_ASAP7_75t_L g936 ( .A(n_663), .Y(n_936) );
BUFx2_ASAP7_75t_L g1253 ( .A(n_663), .Y(n_1253) );
OAI22xp5_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_671), .B1(n_672), .B2(n_673), .Y(n_666) );
OAI22xp5_ASAP7_75t_L g931 ( .A1(n_667), .A2(n_932), .B1(n_933), .B2(n_934), .Y(n_931) );
INVx2_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx2_ASAP7_75t_SL g945 ( .A(n_668), .Y(n_945) );
INVx2_ASAP7_75t_L g1429 ( .A(n_668), .Y(n_1429) );
BUFx3_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g1050 ( .A(n_669), .Y(n_1050) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g677 ( .A(n_670), .Y(n_677) );
BUFx2_ASAP7_75t_L g772 ( .A(n_670), .Y(n_772) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
HB1xp67_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g994 ( .A(n_677), .Y(n_994) );
INVx2_ASAP7_75t_L g1600 ( .A(n_677), .Y(n_1600) );
INVx1_ASAP7_75t_L g1662 ( .A(n_677), .Y(n_1662) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx2_ASAP7_75t_L g734 ( .A(n_680), .Y(n_734) );
OAI22xp33_ASAP7_75t_L g778 ( .A1(n_682), .A2(n_779), .B1(n_780), .B2(n_782), .Y(n_778) );
OAI22xp33_ASAP7_75t_L g789 ( .A1(n_682), .A2(n_790), .B1(n_791), .B2(n_794), .Y(n_789) );
BUFx2_ASAP7_75t_L g1327 ( .A(n_682), .Y(n_1327) );
OAI22xp33_ASAP7_75t_L g1666 ( .A1(n_682), .A2(n_936), .B1(n_1638), .B2(n_1643), .Y(n_1666) );
BUFx3_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
BUFx3_ASAP7_75t_L g781 ( .A(n_684), .Y(n_781) );
OAI221xp5_ASAP7_75t_L g950 ( .A1(n_684), .A2(n_951), .B1(n_952), .B2(n_954), .C(n_955), .Y(n_950) );
INVx2_ASAP7_75t_L g1441 ( .A(n_684), .Y(n_1441) );
BUFx6f_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g749 ( .A(n_690), .Y(n_749) );
NAND4xp75_ASAP7_75t_L g690 ( .A(n_691), .B(n_692), .C(n_721), .D(n_742), .Y(n_690) );
OAI31xp33_ASAP7_75t_L g692 ( .A1(n_693), .A2(n_707), .A3(n_717), .B(n_718), .Y(n_692) );
OAI22xp5_ASAP7_75t_L g694 ( .A1(n_695), .A2(n_697), .B1(n_698), .B2(n_699), .Y(n_694) );
OAI221xp5_ASAP7_75t_L g1228 ( .A1(n_695), .A2(n_714), .B1(n_1229), .B2(n_1230), .C(n_1231), .Y(n_1228) );
INVx2_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
HB1xp67_ASAP7_75t_L g802 ( .A(n_696), .Y(n_802) );
INVx2_ASAP7_75t_L g1117 ( .A(n_696), .Y(n_1117) );
INVx2_ASAP7_75t_L g1163 ( .A(n_696), .Y(n_1163) );
INVx1_ASAP7_75t_L g1209 ( .A(n_696), .Y(n_1209) );
INVx1_ASAP7_75t_L g1407 ( .A(n_698), .Y(n_1407) );
OAI21xp33_ASAP7_75t_L g700 ( .A1(n_701), .A2(n_702), .B(n_704), .Y(n_700) );
INVx2_ASAP7_75t_SL g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g714 ( .A(n_703), .Y(n_714) );
INVx2_ASAP7_75t_L g868 ( .A(n_703), .Y(n_868) );
INVx1_ASAP7_75t_L g1222 ( .A(n_703), .Y(n_1222) );
BUFx2_ASAP7_75t_L g806 ( .A(n_705), .Y(n_806) );
INVx1_ASAP7_75t_L g1125 ( .A(n_705), .Y(n_1125) );
OAI211xp5_ASAP7_75t_L g712 ( .A1(n_713), .A2(n_714), .B(n_715), .C(n_716), .Y(n_712) );
OAI31xp33_ASAP7_75t_L g797 ( .A1(n_718), .A2(n_798), .A3(n_808), .B(n_825), .Y(n_797) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
AOI31xp33_ASAP7_75t_SL g1060 ( .A1(n_719), .A2(n_1061), .A3(n_1067), .B(n_1075), .Y(n_1060) );
OAI31xp33_ASAP7_75t_SL g1176 ( .A1(n_719), .A2(n_1177), .A3(n_1180), .B(n_1190), .Y(n_1176) );
OAI31xp33_ASAP7_75t_L g1236 ( .A1(n_719), .A2(n_1237), .A3(n_1250), .B(n_1258), .Y(n_1236) );
AOI31xp33_ASAP7_75t_L g1271 ( .A1(n_719), .A2(n_1272), .A3(n_1282), .B(n_1288), .Y(n_1271) );
INVx2_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
NOR2xp67_ASAP7_75t_L g1145 ( .A(n_720), .B(n_959), .Y(n_1145) );
AOI22xp5_ASAP7_75t_L g1627 ( .A1(n_720), .A2(n_1545), .B1(n_1628), .B2(n_1645), .Y(n_1627) );
AND2x2_ASAP7_75t_SL g721 ( .A(n_722), .B(n_741), .Y(n_721) );
AOI33xp33_ASAP7_75t_L g722 ( .A1(n_723), .A2(n_724), .A3(n_726), .B1(n_731), .B2(n_735), .B3(n_739), .Y(n_722) );
AOI22xp5_ASAP7_75t_L g1040 ( .A1(n_723), .A2(n_1041), .B1(n_1046), .B2(n_1047), .Y(n_1040) );
BUFx2_ASAP7_75t_L g2010 ( .A(n_723), .Y(n_2010) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx2_ASAP7_75t_L g1943 ( .A(n_730), .Y(n_1943) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
OAI22xp5_ASAP7_75t_L g1501 ( .A1(n_733), .A2(n_1050), .B1(n_1502), .B2(n_1503), .Y(n_1501) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
AND2x4_ASAP7_75t_L g925 ( .A(n_734), .B(n_926), .Y(n_925) );
INVx2_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx2_ASAP7_75t_SL g1304 ( .A(n_737), .Y(n_1304) );
INVx3_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
BUFx6f_ASAP7_75t_L g845 ( .A(n_738), .Y(n_845) );
BUFx2_ASAP7_75t_L g1507 ( .A(n_738), .Y(n_1507) );
NAND3xp33_ASAP7_75t_L g1000 ( .A(n_739), .B(n_1001), .C(n_1002), .Y(n_1000) );
INVx2_ASAP7_75t_SL g956 ( .A(n_740), .Y(n_956) );
INVx1_ASAP7_75t_L g1197 ( .A(n_740), .Y(n_1197) );
OAI22xp5_ASAP7_75t_L g750 ( .A1(n_751), .A2(n_828), .B1(n_829), .B2(n_887), .Y(n_750) );
INVx1_ASAP7_75t_L g887 ( .A(n_751), .Y(n_887) );
INVx1_ASAP7_75t_L g826 ( .A(n_752), .Y(n_826) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
AOI21xp5_ASAP7_75t_L g858 ( .A1(n_754), .A2(n_859), .B(n_860), .Y(n_858) );
AOI21xp5_ASAP7_75t_L g1107 ( .A1(n_754), .A2(n_1108), .B(n_1109), .Y(n_1107) );
AOI21xp5_ASAP7_75t_L g1269 ( .A1(n_754), .A2(n_1270), .B(n_1271), .Y(n_1269) );
AOI21xp33_ASAP7_75t_SL g1344 ( .A1(n_754), .A2(n_1345), .B(n_1346), .Y(n_1344) );
NOR3xp33_ASAP7_75t_L g755 ( .A(n_756), .B(n_765), .C(n_768), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_757), .B(n_761), .Y(n_756) );
OAI221xp5_ASAP7_75t_L g814 ( .A1(n_758), .A2(n_763), .B1(n_803), .B2(n_815), .C(n_817), .Y(n_814) );
INVx1_ASAP7_75t_L g1472 ( .A(n_759), .Y(n_1472) );
OAI22xp5_ASAP7_75t_L g769 ( .A1(n_770), .A2(n_773), .B1(n_774), .B2(n_777), .Y(n_769) );
OAI22xp5_ASAP7_75t_L g783 ( .A1(n_770), .A2(n_784), .B1(n_785), .B2(n_788), .Y(n_783) );
OAI22xp5_ASAP7_75t_L g1434 ( .A1(n_770), .A2(n_776), .B1(n_1435), .B2(n_1436), .Y(n_1434) );
OAI22xp5_ASAP7_75t_L g1611 ( .A1(n_770), .A2(n_774), .B1(n_1612), .B2(n_1613), .Y(n_1611) );
INVx2_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
INVx2_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
OR2x2_ASAP7_75t_L g2048 ( .A(n_772), .B(n_2049), .Y(n_2048) );
OAI22xp5_ASAP7_75t_L g1185 ( .A1(n_774), .A2(n_1186), .B1(n_1187), .B2(n_1188), .Y(n_1185) );
INVx2_ASAP7_75t_SL g774 ( .A(n_775), .Y(n_774) );
INVx1_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
OAI221xp5_ASAP7_75t_L g800 ( .A1(n_777), .A2(n_779), .B1(n_801), .B2(n_803), .C(n_805), .Y(n_800) );
BUFx3_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
OAI22xp33_ASAP7_75t_L g1655 ( .A1(n_781), .A2(n_1656), .B1(n_1657), .B2(n_1658), .Y(n_1655) );
INVx1_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
INVx3_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
INVx2_ASAP7_75t_L g948 ( .A(n_787), .Y(n_948) );
INVx2_ASAP7_75t_L g1335 ( .A(n_787), .Y(n_1335) );
INVx1_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
INVx1_ASAP7_75t_L g1329 ( .A(n_792), .Y(n_1329) );
INVx1_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
AOI21xp33_ASAP7_75t_L g965 ( .A1(n_793), .A2(n_961), .B(n_966), .Y(n_965) );
BUFx2_ASAP7_75t_L g1182 ( .A(n_793), .Y(n_1182) );
OAI21xp5_ASAP7_75t_SL g1498 ( .A1(n_793), .A2(n_1499), .B(n_1500), .Y(n_1498) );
INVx1_ASAP7_75t_L g1543 ( .A(n_795), .Y(n_1543) );
CKINVDCx8_ASAP7_75t_R g795 ( .A(n_796), .Y(n_795) );
NAND3xp33_ASAP7_75t_L g2011 ( .A(n_796), .B(n_2012), .C(n_2013), .Y(n_2011) );
INVx1_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
INVx2_ASAP7_75t_SL g803 ( .A(n_804), .Y(n_803) );
INVx1_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
INVx2_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
INVx1_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
BUFx6f_ASAP7_75t_L g1073 ( .A(n_820), .Y(n_1073) );
INVx1_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
INVx1_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
INVx1_ASAP7_75t_L g1123 ( .A(n_823), .Y(n_1123) );
NAND2xp5_ASAP7_75t_L g1411 ( .A(n_823), .B(n_921), .Y(n_1411) );
INVx2_ASAP7_75t_SL g828 ( .A(n_829), .Y(n_828) );
XNOR2x1_ASAP7_75t_L g829 ( .A(n_830), .B(n_886), .Y(n_829) );
AND2x2_ASAP7_75t_L g830 ( .A(n_831), .B(n_858), .Y(n_830) );
AND4x1_ASAP7_75t_L g831 ( .A(n_832), .B(n_835), .C(n_839), .D(n_842), .Y(n_831) );
OAI211xp5_ASAP7_75t_L g867 ( .A1(n_838), .A2(n_868), .B(n_869), .C(n_870), .Y(n_867) );
HB1xp67_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
INVx1_ASAP7_75t_L g855 ( .A(n_845), .Y(n_855) );
INVx1_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
INVx1_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
INVx1_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
INVx2_ASAP7_75t_L g856 ( .A(n_857), .Y(n_856) );
INVx2_ASAP7_75t_SL g1305 ( .A(n_857), .Y(n_1305) );
INVx3_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
INVx1_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
INVx2_ASAP7_75t_SL g1350 ( .A(n_876), .Y(n_1350) );
HB1xp67_ASAP7_75t_L g877 ( .A(n_878), .Y(n_877) );
AND2x2_ASAP7_75t_L g920 ( .A(n_878), .B(n_921), .Y(n_920) );
INVx1_ASAP7_75t_L g878 ( .A(n_879), .Y(n_878) );
BUFx3_ASAP7_75t_L g881 ( .A(n_882), .Y(n_881) );
HB1xp67_ASAP7_75t_L g1402 ( .A(n_882), .Y(n_1402) );
AO22x2_ASAP7_75t_L g888 ( .A1(n_889), .A2(n_1086), .B1(n_1133), .B2(n_1134), .Y(n_888) );
INVx1_ASAP7_75t_L g1133 ( .A(n_889), .Y(n_1133) );
XNOR2xp5_ASAP7_75t_L g889 ( .A(n_890), .B(n_986), .Y(n_889) );
NAND4xp75_ASAP7_75t_L g891 ( .A(n_892), .B(n_922), .C(n_974), .D(n_980), .Y(n_891) );
AND2x2_ASAP7_75t_SL g892 ( .A(n_893), .B(n_910), .Y(n_892) );
AOI33xp33_ASAP7_75t_L g893 ( .A1(n_894), .A2(n_897), .A3(n_899), .B1(n_903), .B2(n_904), .B3(n_907), .Y(n_893) );
CKINVDCx5p33_ASAP7_75t_R g894 ( .A(n_895), .Y(n_894) );
INVx2_ASAP7_75t_L g1149 ( .A(n_895), .Y(n_1149) );
OAI22xp5_ASAP7_75t_L g1217 ( .A1(n_895), .A2(n_908), .B1(n_1218), .B2(n_1228), .Y(n_1217) );
CKINVDCx5p33_ASAP7_75t_R g1399 ( .A(n_895), .Y(n_1399) );
INVx1_ASAP7_75t_L g1565 ( .A(n_896), .Y(n_1565) );
INVx1_ASAP7_75t_L g901 ( .A(n_902), .Y(n_901) );
INVx1_ASAP7_75t_L g905 ( .A(n_906), .Y(n_905) );
INVx1_ASAP7_75t_L g907 ( .A(n_908), .Y(n_907) );
OAI22xp33_ASAP7_75t_L g1147 ( .A1(n_908), .A2(n_1148), .B1(n_1150), .B2(n_1162), .Y(n_1147) );
OAI22xp5_ASAP7_75t_L g1585 ( .A1(n_908), .A2(n_1148), .B1(n_1586), .B2(n_1591), .Y(n_1585) );
INVx4_ASAP7_75t_L g908 ( .A(n_909), .Y(n_908) );
BUFx4f_ASAP7_75t_L g1408 ( .A(n_909), .Y(n_1408) );
AOI221xp5_ASAP7_75t_L g910 ( .A1(n_911), .A2(n_914), .B1(n_915), .B2(n_919), .C(n_920), .Y(n_910) );
AOI22xp5_ASAP7_75t_L g1397 ( .A1(n_911), .A2(n_1174), .B1(n_1387), .B2(n_1389), .Y(n_1397) );
AOI221xp5_ASAP7_75t_L g1489 ( .A1(n_911), .A2(n_920), .B1(n_1490), .B2(n_1491), .C(n_1492), .Y(n_1489) );
INVx2_ASAP7_75t_L g911 ( .A(n_912), .Y(n_911) );
INVx2_ASAP7_75t_SL g918 ( .A(n_913), .Y(n_918) );
INVx1_ASAP7_75t_L g921 ( .A(n_913), .Y(n_921) );
INVx1_ASAP7_75t_L g915 ( .A(n_916), .Y(n_915) );
INVx2_ASAP7_75t_L g1174 ( .A(n_916), .Y(n_1174) );
HB1xp67_ASAP7_75t_L g1235 ( .A(n_916), .Y(n_1235) );
INVx2_ASAP7_75t_L g1490 ( .A(n_916), .Y(n_1490) );
NAND2x1p5_ASAP7_75t_L g916 ( .A(n_917), .B(n_918), .Y(n_916) );
BUFx2_ASAP7_75t_L g1171 ( .A(n_920), .Y(n_1171) );
OAI31xp33_ASAP7_75t_L g922 ( .A1(n_923), .A2(n_930), .A3(n_967), .B(n_972), .Y(n_922) );
INVx3_ASAP7_75t_L g924 ( .A(n_925), .Y(n_924) );
INVx3_ASAP7_75t_L g1179 ( .A(n_925), .Y(n_1179) );
AOI221x1_ASAP7_75t_L g1494 ( .A1(n_925), .A2(n_971), .B1(n_1495), .B2(n_1496), .C(n_1497), .Y(n_1494) );
INVx1_ASAP7_75t_L g926 ( .A(n_927), .Y(n_926) );
INVx8_ASAP7_75t_L g928 ( .A(n_929), .Y(n_928) );
AOI221xp5_ASAP7_75t_SL g1504 ( .A1(n_929), .A2(n_1505), .B1(n_1506), .B2(n_1508), .C(n_1509), .Y(n_1504) );
OAI221xp5_ASAP7_75t_L g930 ( .A1(n_931), .A2(n_935), .B1(n_944), .B2(n_950), .C(n_957), .Y(n_930) );
OAI221xp5_ASAP7_75t_L g1191 ( .A1(n_934), .A2(n_1192), .B1(n_1194), .B2(n_1195), .C(n_1196), .Y(n_1191) );
OAI221xp5_ASAP7_75t_L g935 ( .A1(n_936), .A2(n_937), .B1(n_938), .B2(n_941), .C(n_942), .Y(n_935) );
INVx1_ASAP7_75t_L g938 ( .A(n_939), .Y(n_938) );
INVx1_ASAP7_75t_L g1657 ( .A(n_939), .Y(n_1657) );
INVx2_ASAP7_75t_SL g939 ( .A(n_940), .Y(n_939) );
OAI221xp5_ASAP7_75t_L g1181 ( .A1(n_942), .A2(n_1152), .B1(n_1156), .B2(n_1182), .C(n_1183), .Y(n_1181) );
OAI221xp5_ASAP7_75t_L g1609 ( .A1(n_942), .A2(n_1183), .B1(n_1587), .B2(n_1588), .C(n_1610), .Y(n_1609) );
INVx2_ASAP7_75t_L g942 ( .A(n_943), .Y(n_942) );
OAI22xp5_ASAP7_75t_L g944 ( .A1(n_945), .A2(n_946), .B1(n_947), .B2(n_949), .Y(n_944) );
BUFx2_ASAP7_75t_L g1186 ( .A(n_945), .Y(n_1186) );
AOI22xp5_ASAP7_75t_L g980 ( .A1(n_946), .A2(n_951), .B1(n_981), .B2(n_983), .Y(n_980) );
OAI22xp5_ASAP7_75t_L g1659 ( .A1(n_947), .A2(n_1660), .B1(n_1661), .B2(n_1663), .Y(n_1659) );
OAI22xp5_ASAP7_75t_L g1936 ( .A1(n_947), .A2(n_1661), .B1(n_1937), .B2(n_1938), .Y(n_1936) );
INVx1_ASAP7_75t_L g947 ( .A(n_948), .Y(n_947) );
OAI22xp5_ASAP7_75t_SL g1437 ( .A1(n_952), .A2(n_1438), .B1(n_1439), .B2(n_1440), .Y(n_1437) );
INVx2_ASAP7_75t_L g952 ( .A(n_953), .Y(n_952) );
INVx1_ASAP7_75t_L g1379 ( .A(n_953), .Y(n_1379) );
OAI221xp5_ASAP7_75t_L g1377 ( .A1(n_955), .A2(n_1252), .B1(n_1378), .B2(n_1379), .C(n_1380), .Y(n_1377) );
INVx1_ASAP7_75t_L g955 ( .A(n_956), .Y(n_955) );
AOI21xp5_ASAP7_75t_L g957 ( .A1(n_958), .A2(n_964), .B(n_965), .Y(n_957) );
INVx1_ASAP7_75t_L g958 ( .A(n_959), .Y(n_958) );
NAND2xp5_ASAP7_75t_L g959 ( .A(n_960), .B(n_963), .Y(n_959) );
INVx1_ASAP7_75t_L g960 ( .A(n_961), .Y(n_960) );
INVx1_ASAP7_75t_L g1511 ( .A(n_961), .Y(n_1511) );
INVx2_ASAP7_75t_L g961 ( .A(n_962), .Y(n_961) );
BUFx2_ASAP7_75t_L g1244 ( .A(n_963), .Y(n_1244) );
CKINVDCx6p67_ASAP7_75t_R g968 ( .A(n_969), .Y(n_968) );
INVx3_ASAP7_75t_L g970 ( .A(n_971), .Y(n_970) );
INVx3_ASAP7_75t_L g1178 ( .A(n_971), .Y(n_1178) );
INVx2_ASAP7_75t_L g1033 ( .A(n_972), .Y(n_1033) );
AOI31xp33_ASAP7_75t_L g1547 ( .A1(n_972), .A2(n_1548), .A3(n_1557), .B(n_1570), .Y(n_1547) );
BUFx8_ASAP7_75t_SL g1617 ( .A(n_972), .Y(n_1617) );
INVx2_ASAP7_75t_L g972 ( .A(n_973), .Y(n_972) );
BUFx2_ASAP7_75t_L g1132 ( .A(n_973), .Y(n_1132) );
AND2x4_ASAP7_75t_L g2001 ( .A(n_973), .B(n_2002), .Y(n_2001) );
AOI22xp33_ASAP7_75t_L g1395 ( .A1(n_975), .A2(n_981), .B1(n_1380), .B2(n_1384), .Y(n_1395) );
AND2x2_ASAP7_75t_L g981 ( .A(n_976), .B(n_982), .Y(n_981) );
INVx1_ASAP7_75t_L g976 ( .A(n_977), .Y(n_976) );
OR2x6_ASAP7_75t_L g984 ( .A(n_977), .B(n_985), .Y(n_984) );
OR2x2_ASAP7_75t_L g1208 ( .A(n_977), .B(n_1209), .Y(n_1208) );
OR2x2_ASAP7_75t_L g1210 ( .A(n_977), .B(n_1211), .Y(n_1210) );
AOI22xp33_ASAP7_75t_L g1394 ( .A1(n_978), .A2(n_983), .B1(n_1378), .B2(n_1385), .Y(n_1394) );
CKINVDCx6p67_ASAP7_75t_R g978 ( .A(n_979), .Y(n_978) );
CKINVDCx6p67_ASAP7_75t_R g983 ( .A(n_984), .Y(n_983) );
OAI21xp33_ASAP7_75t_L g1012 ( .A1(n_985), .A2(n_1013), .B(n_1014), .Y(n_1012) );
OAI221xp5_ASAP7_75t_L g1116 ( .A1(n_985), .A2(n_1098), .B1(n_1100), .B2(n_1117), .C(n_1118), .Y(n_1116) );
INVx1_ASAP7_75t_L g1166 ( .A(n_985), .Y(n_1166) );
XNOR2xp5_ASAP7_75t_L g986 ( .A(n_987), .B(n_1034), .Y(n_986) );
NAND3xp33_ASAP7_75t_L g988 ( .A(n_989), .B(n_1004), .C(n_1008), .Y(n_988) );
NOR2xp33_ASAP7_75t_L g989 ( .A(n_990), .B(n_1003), .Y(n_989) );
INVx1_ASAP7_75t_L g991 ( .A(n_992), .Y(n_991) );
OAI221xp5_ASAP7_75t_L g993 ( .A1(n_994), .A2(n_995), .B1(n_996), .B2(n_997), .C(n_998), .Y(n_993) );
INVx1_ASAP7_75t_L g1383 ( .A(n_994), .Y(n_1383) );
BUFx2_ASAP7_75t_L g1245 ( .A(n_999), .Y(n_1245) );
INVx2_ASAP7_75t_SL g2009 ( .A(n_999), .Y(n_2009) );
AOI222xp33_ASAP7_75t_L g2031 ( .A1(n_999), .A2(n_1998), .B1(n_2000), .B2(n_2032), .C1(n_2033), .C2(n_2034), .Y(n_2031) );
NOR2xp33_ASAP7_75t_SL g1004 ( .A(n_1005), .B(n_1007), .Y(n_1004) );
OAI31xp33_ASAP7_75t_SL g1008 ( .A1(n_1009), .A2(n_1010), .A3(n_1011), .B(n_1033), .Y(n_1008) );
OAI211xp5_ASAP7_75t_SL g1011 ( .A1(n_1012), .A2(n_1015), .B(n_1019), .C(n_1025), .Y(n_1011) );
INVx1_ASAP7_75t_L g1017 ( .A(n_1018), .Y(n_1017) );
OAI211xp5_ASAP7_75t_L g1019 ( .A1(n_1020), .A2(n_1021), .B(n_1022), .C(n_1023), .Y(n_1019) );
OAI221xp5_ASAP7_75t_L g1351 ( .A1(n_1021), .A2(n_1117), .B1(n_1118), .B2(n_1319), .C(n_1321), .Y(n_1351) );
NAND2xp33_ASAP7_75t_L g1027 ( .A(n_1028), .B(n_1029), .Y(n_1027) );
INVx1_ASAP7_75t_L g1555 ( .A(n_1028), .Y(n_1555) );
AOI22xp5_ASAP7_75t_L g1948 ( .A1(n_1033), .A2(n_1545), .B1(n_1949), .B2(n_1959), .Y(n_1948) );
NAND2xp5_ASAP7_75t_SL g1034 ( .A(n_1035), .B(n_1082), .Y(n_1034) );
INVx1_ASAP7_75t_L g1084 ( .A(n_1036), .Y(n_1084) );
NAND3xp33_ASAP7_75t_SL g1036 ( .A(n_1037), .B(n_1040), .C(n_1048), .Y(n_1036) );
AOI22xp5_ASAP7_75t_L g1075 ( .A1(n_1046), .A2(n_1076), .B1(n_1078), .B2(n_1080), .Y(n_1075) );
INVx2_ASAP7_75t_L g1193 ( .A(n_1050), .Y(n_1193) );
INVx1_ASAP7_75t_L g1241 ( .A(n_1055), .Y(n_1241) );
INVx2_ASAP7_75t_L g1055 ( .A(n_1056), .Y(n_1055) );
INVx1_ASAP7_75t_L g1083 ( .A(n_1060), .Y(n_1083) );
BUFx2_ASAP7_75t_L g1219 ( .A(n_1063), .Y(n_1219) );
OAI221xp5_ASAP7_75t_SL g1453 ( .A1(n_1063), .A2(n_1430), .B1(n_1433), .B2(n_1454), .C(n_1455), .Y(n_1453) );
INVx2_ASAP7_75t_L g1063 ( .A(n_1064), .Y(n_1063) );
INVx1_ASAP7_75t_L g1069 ( .A(n_1070), .Y(n_1069) );
INVx2_ASAP7_75t_L g1403 ( .A(n_1070), .Y(n_1403) );
INVx1_ASAP7_75t_L g1640 ( .A(n_1070), .Y(n_1640) );
HB1xp67_ASAP7_75t_L g1355 ( .A(n_1077), .Y(n_1355) );
INVx1_ASAP7_75t_L g1161 ( .A(n_1079), .Y(n_1161) );
INVx2_ASAP7_75t_L g1080 ( .A(n_1081), .Y(n_1080) );
NAND3xp33_ASAP7_75t_L g1082 ( .A(n_1083), .B(n_1084), .C(n_1085), .Y(n_1082) );
INVx2_ASAP7_75t_L g1134 ( .A(n_1086), .Y(n_1134) );
NAND2xp5_ASAP7_75t_L g1087 ( .A(n_1088), .B(n_1107), .Y(n_1087) );
AND4x1_ASAP7_75t_L g1088 ( .A(n_1089), .B(n_1095), .C(n_1099), .D(n_1102), .Y(n_1088) );
INVx1_ASAP7_75t_L g1092 ( .A(n_1093), .Y(n_1092) );
AOI31xp33_ASAP7_75t_L g1109 ( .A1(n_1110), .A2(n_1119), .A3(n_1128), .B(n_1131), .Y(n_1109) );
INVx1_ASAP7_75t_L g1114 ( .A(n_1115), .Y(n_1114) );
INVx1_ASAP7_75t_L g1122 ( .A(n_1123), .Y(n_1122) );
INVx1_ASAP7_75t_L g1124 ( .A(n_1125), .Y(n_1124) );
AOI31xp33_ASAP7_75t_L g1346 ( .A1(n_1131), .A2(n_1347), .A3(n_1352), .B(n_1359), .Y(n_1346) );
INVx1_ASAP7_75t_L g1469 ( .A(n_1131), .Y(n_1469) );
INVx2_ASAP7_75t_L g1131 ( .A(n_1132), .Y(n_1131) );
AOI21x1_ASAP7_75t_L g1493 ( .A1(n_1132), .A2(n_1494), .B(n_1504), .Y(n_1493) );
INVx1_ASAP7_75t_L g1415 ( .A(n_1135), .Y(n_1415) );
OAI22xp5_ASAP7_75t_L g1135 ( .A1(n_1136), .A2(n_1137), .B1(n_1311), .B2(n_1414), .Y(n_1135) );
INVx1_ASAP7_75t_L g1136 ( .A(n_1137), .Y(n_1136) );
XNOR2xp5_ASAP7_75t_L g1137 ( .A(n_1138), .B(n_1212), .Y(n_1137) );
INVx1_ASAP7_75t_L g1138 ( .A(n_1139), .Y(n_1138) );
XNOR2xp5_ASAP7_75t_L g1139 ( .A(n_1140), .B(n_1141), .Y(n_1139) );
AND4x1_ASAP7_75t_L g1141 ( .A(n_1142), .B(n_1146), .C(n_1176), .D(n_1205), .Y(n_1141) );
NAND2xp5_ASAP7_75t_L g1142 ( .A(n_1143), .B(n_1144), .Y(n_1142) );
NAND2xp5_ASAP7_75t_L g1259 ( .A(n_1144), .B(n_1260), .Y(n_1259) );
NAND2xp5_ASAP7_75t_L g1390 ( .A(n_1144), .B(n_1391), .Y(n_1390) );
NAND2xp5_ASAP7_75t_L g1582 ( .A(n_1144), .B(n_1583), .Y(n_1582) );
NOR3xp33_ASAP7_75t_L g1146 ( .A(n_1147), .B(n_1171), .C(n_1172), .Y(n_1146) );
INVx1_ASAP7_75t_L g1148 ( .A(n_1149), .Y(n_1148) );
OAI221xp5_ASAP7_75t_L g1150 ( .A1(n_1151), .A2(n_1152), .B1(n_1153), .B2(n_1156), .C(n_1157), .Y(n_1150) );
OAI221xp5_ASAP7_75t_L g1553 ( .A1(n_1151), .A2(n_1526), .B1(n_1529), .B2(n_1554), .C(n_1556), .Y(n_1553) );
OAI221xp5_ASAP7_75t_L g1591 ( .A1(n_1151), .A2(n_1165), .B1(n_1592), .B2(n_1593), .C(n_1594), .Y(n_1591) );
OAI221xp5_ASAP7_75t_L g1586 ( .A1(n_1153), .A2(n_1163), .B1(n_1587), .B2(n_1588), .C(n_1589), .Y(n_1586) );
INVx2_ASAP7_75t_L g1153 ( .A(n_1154), .Y(n_1153) );
INVx1_ASAP7_75t_L g1154 ( .A(n_1155), .Y(n_1154) );
INVx1_ASAP7_75t_L g1158 ( .A(n_1159), .Y(n_1158) );
INVx1_ASAP7_75t_L g1276 ( .A(n_1159), .Y(n_1276) );
INVx1_ASAP7_75t_L g1354 ( .A(n_1159), .Y(n_1354) );
INVx1_ASAP7_75t_L g1160 ( .A(n_1161), .Y(n_1160) );
OAI221xp5_ASAP7_75t_L g1162 ( .A1(n_1163), .A2(n_1164), .B1(n_1165), .B2(n_1167), .C(n_1168), .Y(n_1162) );
INVx2_ASAP7_75t_L g1165 ( .A(n_1166), .Y(n_1165) );
BUFx3_ASAP7_75t_L g1169 ( .A(n_1170), .Y(n_1169) );
NOR3xp33_ASAP7_75t_L g1216 ( .A(n_1171), .B(n_1217), .C(n_1234), .Y(n_1216) );
NOR3xp33_ASAP7_75t_SL g1584 ( .A(n_1171), .B(n_1585), .C(n_1595), .Y(n_1584) );
INVx1_ASAP7_75t_L g1173 ( .A(n_1174), .Y(n_1173) );
OAI22xp5_ASAP7_75t_L g1337 ( .A1(n_1182), .A2(n_1338), .B1(n_1339), .B2(n_1340), .Y(n_1337) );
OAI221xp5_ASAP7_75t_L g1371 ( .A1(n_1183), .A2(n_1254), .B1(n_1372), .B2(n_1373), .C(n_1374), .Y(n_1371) );
INVx3_ASAP7_75t_L g1183 ( .A(n_1184), .Y(n_1183) );
OAI22xp5_ASAP7_75t_L g1331 ( .A1(n_1192), .A2(n_1332), .B1(n_1333), .B2(n_1336), .Y(n_1331) );
OAI22xp5_ASAP7_75t_L g1367 ( .A1(n_1192), .A2(n_1368), .B1(n_1369), .B2(n_1370), .Y(n_1367) );
INVx2_ASAP7_75t_L g1192 ( .A(n_1193), .Y(n_1192) );
INVx1_ASAP7_75t_L g1239 ( .A(n_1193), .Y(n_1239) );
INVx2_ASAP7_75t_L g1338 ( .A(n_1193), .Y(n_1338) );
INVx2_ASAP7_75t_L g1665 ( .A(n_1193), .Y(n_1665) );
INVx1_ASAP7_75t_L g1940 ( .A(n_1193), .Y(n_1940) );
AOI22xp33_ASAP7_75t_L g1198 ( .A1(n_1199), .A2(n_1201), .B1(n_1202), .B2(n_1204), .Y(n_1198) );
AOI22xp33_ASAP7_75t_L g1605 ( .A1(n_1199), .A2(n_1202), .B1(n_1606), .B2(n_1607), .Y(n_1605) );
HB1xp67_ASAP7_75t_L g1199 ( .A(n_1200), .Y(n_1199) );
AOI22xp33_ASAP7_75t_L g1247 ( .A1(n_1200), .A2(n_1202), .B1(n_1248), .B2(n_1249), .Y(n_1247) );
AOI22xp33_ASAP7_75t_L g1386 ( .A1(n_1202), .A2(n_1387), .B1(n_1388), .B2(n_1389), .Y(n_1386) );
CKINVDCx11_ASAP7_75t_R g1202 ( .A(n_1203), .Y(n_1202) );
NOR2xp33_ASAP7_75t_L g1205 ( .A(n_1206), .B(n_1207), .Y(n_1205) );
AO22x1_ASAP7_75t_L g1212 ( .A1(n_1213), .A2(n_1214), .B1(n_1265), .B2(n_1310), .Y(n_1212) );
INVx1_ASAP7_75t_L g1213 ( .A(n_1214), .Y(n_1213) );
AND4x1_ASAP7_75t_L g1215 ( .A(n_1216), .B(n_1236), .C(n_1259), .D(n_1261), .Y(n_1215) );
OAI221xp5_ASAP7_75t_L g1218 ( .A1(n_1219), .A2(n_1220), .B1(n_1221), .B2(n_1223), .C(n_1224), .Y(n_1218) );
BUFx2_ASAP7_75t_L g1221 ( .A(n_1222), .Y(n_1221) );
INVx1_ASAP7_75t_L g1226 ( .A(n_1227), .Y(n_1226) );
INVx1_ASAP7_75t_L g1569 ( .A(n_1227), .Y(n_1569) );
INVx1_ASAP7_75t_L g2028 ( .A(n_1227), .Y(n_2028) );
OAI221xp5_ASAP7_75t_L g1238 ( .A1(n_1239), .A2(n_1240), .B1(n_1241), .B2(n_1242), .C(n_1243), .Y(n_1238) );
INVx2_ASAP7_75t_L g1252 ( .A(n_1253), .Y(n_1252) );
INVx1_ASAP7_75t_L g1372 ( .A(n_1253), .Y(n_1372) );
INVx1_ASAP7_75t_L g1935 ( .A(n_1253), .Y(n_1935) );
NOR2xp33_ASAP7_75t_L g1261 ( .A(n_1262), .B(n_1264), .Y(n_1261) );
INVx1_ASAP7_75t_L g1310 ( .A(n_1265), .Y(n_1310) );
INVx1_ASAP7_75t_L g1265 ( .A(n_1266), .Y(n_1265) );
XNOR2x1_ASAP7_75t_SL g1266 ( .A(n_1267), .B(n_1268), .Y(n_1266) );
AND2x2_ASAP7_75t_L g1268 ( .A(n_1269), .B(n_1291), .Y(n_1268) );
INVx2_ASAP7_75t_SL g1280 ( .A(n_1281), .Y(n_1280) );
INVx1_ASAP7_75t_L g1284 ( .A(n_1285), .Y(n_1284) );
AND4x1_ASAP7_75t_L g1291 ( .A(n_1292), .B(n_1295), .C(n_1298), .D(n_1302), .Y(n_1291) );
AOI22xp33_ASAP7_75t_L g1524 ( .A1(n_1301), .A2(n_1525), .B1(n_1526), .B2(n_1527), .Y(n_1524) );
INVx1_ASAP7_75t_L g1414 ( .A(n_1311), .Y(n_1414) );
AOI22xp5_ASAP7_75t_L g1311 ( .A1(n_1312), .A2(n_1313), .B1(n_1361), .B2(n_1413), .Y(n_1311) );
INVx2_ASAP7_75t_L g1312 ( .A(n_1313), .Y(n_1312) );
XNOR2x1_ASAP7_75t_L g1313 ( .A(n_1314), .B(n_1360), .Y(n_1313) );
AND2x2_ASAP7_75t_L g1314 ( .A(n_1315), .B(n_1344), .Y(n_1314) );
NOR3xp33_ASAP7_75t_L g1315 ( .A(n_1316), .B(n_1323), .C(n_1325), .Y(n_1315) );
NAND2xp5_ASAP7_75t_L g1316 ( .A(n_1317), .B(n_1320), .Y(n_1316) );
OAI22xp33_ASAP7_75t_L g1326 ( .A1(n_1327), .A2(n_1328), .B1(n_1329), .B2(n_1330), .Y(n_1326) );
INVx1_ASAP7_75t_L g1333 ( .A(n_1334), .Y(n_1333) );
HB1xp67_ASAP7_75t_L g1334 ( .A(n_1335), .Y(n_1334) );
HB1xp67_ASAP7_75t_L g1590 ( .A(n_1357), .Y(n_1590) );
BUFx2_ASAP7_75t_L g1357 ( .A(n_1358), .Y(n_1357) );
INVx2_ASAP7_75t_L g1463 ( .A(n_1358), .Y(n_1463) );
INVx1_ASAP7_75t_L g1413 ( .A(n_1361), .Y(n_1413) );
INVx1_ASAP7_75t_L g1362 ( .A(n_1363), .Y(n_1362) );
NAND3xp33_ASAP7_75t_SL g1363 ( .A(n_1364), .B(n_1390), .C(n_1392), .Y(n_1363) );
OAI21xp5_ASAP7_75t_L g1497 ( .A1(n_1375), .A2(n_1498), .B(n_1501), .Y(n_1497) );
INVx1_ASAP7_75t_L g1382 ( .A(n_1383), .Y(n_1382) );
NOR2xp33_ASAP7_75t_L g1392 ( .A(n_1393), .B(n_1396), .Y(n_1392) );
NAND2xp5_ASAP7_75t_L g1393 ( .A(n_1394), .B(n_1395), .Y(n_1393) );
NAND3xp33_ASAP7_75t_SL g1396 ( .A(n_1397), .B(n_1398), .C(n_1409), .Y(n_1396) );
AOI33xp33_ASAP7_75t_L g1398 ( .A1(n_1399), .A2(n_1400), .A3(n_1401), .B1(n_1404), .B2(n_1406), .B3(n_1408), .Y(n_1398) );
NAND3xp33_ASAP7_75t_L g2023 ( .A(n_1408), .B(n_2024), .C(n_2027), .Y(n_2023) );
INVx1_ASAP7_75t_L g1409 ( .A(n_1410), .Y(n_1409) );
INVx1_ASAP7_75t_L g1410 ( .A(n_1411), .Y(n_1410) );
XNOR2xp5_ASAP7_75t_L g1416 ( .A(n_1417), .B(n_1575), .Y(n_1416) );
HB1xp67_ASAP7_75t_L g1417 ( .A(n_1418), .Y(n_1417) );
OAI22xp5_ASAP7_75t_L g1418 ( .A1(n_1419), .A2(n_1420), .B1(n_1518), .B2(n_1574), .Y(n_1418) );
INVx1_ASAP7_75t_L g1419 ( .A(n_1420), .Y(n_1419) );
AO22x2_ASAP7_75t_L g1420 ( .A1(n_1421), .A2(n_1474), .B1(n_1475), .B2(n_1517), .Y(n_1420) );
INVx1_ASAP7_75t_L g1517 ( .A(n_1421), .Y(n_1517) );
AND2x2_ASAP7_75t_L g1422 ( .A(n_1423), .B(n_1443), .Y(n_1422) );
NOR2xp33_ASAP7_75t_L g1423 ( .A(n_1424), .B(n_1426), .Y(n_1423) );
OAI22xp33_ASAP7_75t_L g1945 ( .A1(n_1440), .A2(n_1657), .B1(n_1946), .B2(n_1947), .Y(n_1945) );
INVx2_ASAP7_75t_L g1440 ( .A(n_1441), .Y(n_1440) );
INVx1_ASAP7_75t_L g1610 ( .A(n_1441), .Y(n_1610) );
AOI21xp5_ASAP7_75t_SL g1443 ( .A1(n_1444), .A2(n_1469), .B(n_1470), .Y(n_1443) );
NAND4xp25_ASAP7_75t_SL g1444 ( .A(n_1445), .B(n_1451), .C(n_1453), .D(n_1457), .Y(n_1444) );
INVx1_ASAP7_75t_L g1447 ( .A(n_1448), .Y(n_1447) );
OAI221xp5_ASAP7_75t_L g1457 ( .A1(n_1458), .A2(n_1460), .B1(n_1461), .B2(n_1464), .C(n_1465), .Y(n_1457) );
INVx1_ASAP7_75t_L g1458 ( .A(n_1459), .Y(n_1458) );
INVx1_ASAP7_75t_L g1461 ( .A(n_1462), .Y(n_1461) );
INVx1_ASAP7_75t_L g1462 ( .A(n_1463), .Y(n_1462) );
INVx1_ASAP7_75t_L g1556 ( .A(n_1468), .Y(n_1556) );
INVx1_ASAP7_75t_L g1474 ( .A(n_1475), .Y(n_1474) );
NOR4xp75_ASAP7_75t_L g1476 ( .A(n_1477), .B(n_1493), .C(n_1515), .D(n_1516), .Y(n_1476) );
NAND2xp5_ASAP7_75t_L g1477 ( .A(n_1478), .B(n_1489), .Y(n_1477) );
AOI33xp33_ASAP7_75t_L g1478 ( .A1(n_1479), .A2(n_1482), .A3(n_1484), .B1(n_1485), .B2(n_1487), .B3(n_1488), .Y(n_1478) );
INVx3_ASAP7_75t_L g1479 ( .A(n_1480), .Y(n_1479) );
INVx2_ASAP7_75t_L g1596 ( .A(n_1490), .Y(n_1596) );
NAND2xp5_ASAP7_75t_L g1512 ( .A(n_1513), .B(n_1514), .Y(n_1512) );
BUFx3_ASAP7_75t_L g1535 ( .A(n_1514), .Y(n_1535) );
INVx2_ASAP7_75t_L g1574 ( .A(n_1518), .Y(n_1574) );
XOR2x2_ASAP7_75t_L g1518 ( .A(n_1519), .B(n_1573), .Y(n_1518) );
NAND2xp5_ASAP7_75t_L g1519 ( .A(n_1520), .B(n_1544), .Y(n_1519) );
AND4x1_ASAP7_75t_L g1520 ( .A(n_1521), .B(n_1524), .C(n_1528), .D(n_1533), .Y(n_1520) );
AOI22xp33_ASAP7_75t_L g1528 ( .A1(n_1529), .A2(n_1530), .B1(n_1531), .B2(n_1532), .Y(n_1528) );
INVx1_ASAP7_75t_L g1536 ( .A(n_1537), .Y(n_1536) );
CKINVDCx5p33_ASAP7_75t_R g1537 ( .A(n_1538), .Y(n_1537) );
AOI21xp5_ASAP7_75t_L g1544 ( .A1(n_1545), .A2(n_1546), .B(n_1547), .Y(n_1544) );
INVx1_ASAP7_75t_L g1554 ( .A(n_1555), .Y(n_1554) );
INVx1_ASAP7_75t_L g1562 ( .A(n_1563), .Y(n_1562) );
INVx1_ASAP7_75t_L g1564 ( .A(n_1565), .Y(n_1564) );
HB1xp67_ASAP7_75t_L g1567 ( .A(n_1568), .Y(n_1567) );
OAI22xp5_ASAP7_75t_L g1718 ( .A1(n_1573), .A2(n_1719), .B1(n_1720), .B2(n_1722), .Y(n_1718) );
XNOR2xp5_ASAP7_75t_L g1575 ( .A(n_1576), .B(n_1621), .Y(n_1575) );
INVx1_ASAP7_75t_L g1576 ( .A(n_1577), .Y(n_1576) );
INVx1_ASAP7_75t_L g1577 ( .A(n_1578), .Y(n_1577) );
INVx1_ASAP7_75t_L g1578 ( .A(n_1579), .Y(n_1578) );
XNOR2xp5_ASAP7_75t_L g1579 ( .A(n_1580), .B(n_1581), .Y(n_1579) );
AND4x1_ASAP7_75t_L g1581 ( .A(n_1582), .B(n_1584), .C(n_1597), .D(n_1618), .Y(n_1581) );
OAI31xp33_ASAP7_75t_L g1597 ( .A1(n_1598), .A2(n_1608), .A3(n_1614), .B(n_1615), .Y(n_1597) );
INVx1_ASAP7_75t_SL g1615 ( .A(n_1616), .Y(n_1615) );
INVx5_ASAP7_75t_L g1616 ( .A(n_1617), .Y(n_1616) );
NOR2xp33_ASAP7_75t_L g1618 ( .A(n_1619), .B(n_1620), .Y(n_1618) );
INVx1_ASAP7_75t_L g1621 ( .A(n_1622), .Y(n_1621) );
INVx1_ASAP7_75t_L g1622 ( .A(n_1623), .Y(n_1622) );
HB1xp67_ASAP7_75t_L g1623 ( .A(n_1624), .Y(n_1623) );
INVx1_ASAP7_75t_L g1624 ( .A(n_1625), .Y(n_1624) );
AND2x2_ASAP7_75t_L g1626 ( .A(n_1627), .B(n_1646), .Y(n_1626) );
NAND3xp33_ASAP7_75t_L g1628 ( .A(n_1629), .B(n_1637), .C(n_1642), .Y(n_1628) );
NOR3xp33_ASAP7_75t_SL g1646 ( .A(n_1647), .B(n_1652), .C(n_1654), .Y(n_1646) );
NAND2xp5_ASAP7_75t_L g1647 ( .A(n_1648), .B(n_1650), .Y(n_1647) );
OAI22xp33_ASAP7_75t_L g1932 ( .A1(n_1657), .A2(n_1933), .B1(n_1934), .B2(n_1935), .Y(n_1932) );
BUFx2_ASAP7_75t_L g1661 ( .A(n_1662), .Y(n_1661) );
OAI221xp5_ASAP7_75t_L g1668 ( .A1(n_1669), .A2(n_1918), .B1(n_1920), .B2(n_1960), .C(n_1964), .Y(n_1668) );
O2A1O1Ixp33_ASAP7_75t_L g1669 ( .A1(n_1670), .A2(n_1800), .B(n_1836), .C(n_1886), .Y(n_1669) );
NAND5xp2_ASAP7_75t_L g1670 ( .A(n_1671), .B(n_1757), .C(n_1785), .D(n_1794), .E(n_1798), .Y(n_1670) );
AOI221xp5_ASAP7_75t_L g1671 ( .A1(n_1672), .A2(n_1708), .B1(n_1732), .B2(n_1739), .C(n_1746), .Y(n_1671) );
INVxp67_ASAP7_75t_SL g1672 ( .A(n_1673), .Y(n_1672) );
NOR2xp33_ASAP7_75t_L g1673 ( .A(n_1674), .B(n_1698), .Y(n_1673) );
AOI221xp5_ASAP7_75t_L g1887 ( .A1(n_1674), .A2(n_1715), .B1(n_1821), .B2(n_1888), .C(n_1889), .Y(n_1887) );
AND2x2_ASAP7_75t_L g1674 ( .A(n_1675), .B(n_1694), .Y(n_1674) );
INVx2_ASAP7_75t_L g1701 ( .A(n_1675), .Y(n_1701) );
AND2x2_ASAP7_75t_L g1737 ( .A(n_1675), .B(n_1738), .Y(n_1737) );
AND2x2_ASAP7_75t_L g1752 ( .A(n_1675), .B(n_1702), .Y(n_1752) );
OR2x2_ASAP7_75t_L g1788 ( .A(n_1675), .B(n_1702), .Y(n_1788) );
NOR2xp33_ASAP7_75t_L g1842 ( .A(n_1675), .B(n_1694), .Y(n_1842) );
AND2x2_ASAP7_75t_L g1675 ( .A(n_1676), .B(n_1688), .Y(n_1675) );
AND2x4_ASAP7_75t_L g1677 ( .A(n_1678), .B(n_1683), .Y(n_1677) );
INVx1_ASAP7_75t_L g1678 ( .A(n_1679), .Y(n_1678) );
OR2x2_ASAP7_75t_L g1705 ( .A(n_1679), .B(n_1684), .Y(n_1705) );
NAND2xp5_ASAP7_75t_L g1679 ( .A(n_1680), .B(n_1682), .Y(n_1679) );
INVx1_ASAP7_75t_L g1680 ( .A(n_1681), .Y(n_1680) );
INVx1_ASAP7_75t_L g1692 ( .A(n_1682), .Y(n_1692) );
AND2x4_ASAP7_75t_L g1685 ( .A(n_1683), .B(n_1686), .Y(n_1685) );
INVx1_ASAP7_75t_L g1683 ( .A(n_1684), .Y(n_1683) );
OR2x2_ASAP7_75t_L g1707 ( .A(n_1684), .B(n_1687), .Y(n_1707) );
BUFx2_ASAP7_75t_L g1743 ( .A(n_1685), .Y(n_1743) );
HB1xp67_ASAP7_75t_L g2058 ( .A(n_1686), .Y(n_2058) );
INVx1_ASAP7_75t_L g1686 ( .A(n_1687), .Y(n_1686) );
AND2x2_ASAP7_75t_L g1689 ( .A(n_1690), .B(n_1691), .Y(n_1689) );
AND2x4_ASAP7_75t_L g1693 ( .A(n_1690), .B(n_1692), .Y(n_1693) );
AND2x4_ASAP7_75t_L g1714 ( .A(n_1690), .B(n_1691), .Y(n_1714) );
INVx1_ASAP7_75t_L g1691 ( .A(n_1692), .Y(n_1691) );
INVx2_ASAP7_75t_L g1726 ( .A(n_1693), .Y(n_1726) );
OR2x2_ASAP7_75t_L g1751 ( .A(n_1694), .B(n_1711), .Y(n_1751) );
OR2x2_ASAP7_75t_L g1761 ( .A(n_1694), .B(n_1762), .Y(n_1761) );
NAND2xp5_ASAP7_75t_L g1763 ( .A(n_1694), .B(n_1701), .Y(n_1763) );
AND2x2_ASAP7_75t_L g1776 ( .A(n_1694), .B(n_1737), .Y(n_1776) );
AND2x2_ASAP7_75t_L g1848 ( .A(n_1694), .B(n_1849), .Y(n_1848) );
OAI322xp33_ASAP7_75t_L g1858 ( .A1(n_1694), .A2(n_1844), .A3(n_1859), .B1(n_1860), .B2(n_1861), .C1(n_1862), .C2(n_1864), .Y(n_1858) );
AND2x2_ASAP7_75t_L g1863 ( .A(n_1694), .B(n_1738), .Y(n_1863) );
BUFx3_ASAP7_75t_L g1694 ( .A(n_1695), .Y(n_1694) );
INVxp67_ASAP7_75t_L g1699 ( .A(n_1695), .Y(n_1699) );
BUFx2_ASAP7_75t_L g1768 ( .A(n_1695), .Y(n_1768) );
OR2x2_ASAP7_75t_L g1805 ( .A(n_1695), .B(n_1702), .Y(n_1805) );
AND2x2_ASAP7_75t_L g1814 ( .A(n_1695), .B(n_1815), .Y(n_1814) );
AND2x2_ASAP7_75t_L g1695 ( .A(n_1696), .B(n_1697), .Y(n_1695) );
AND2x2_ASAP7_75t_L g1797 ( .A(n_1698), .B(n_1773), .Y(n_1797) );
NAND2xp5_ASAP7_75t_L g1822 ( .A(n_1698), .B(n_1711), .Y(n_1822) );
AND2x2_ASAP7_75t_L g1698 ( .A(n_1699), .B(n_1700), .Y(n_1698) );
NAND2xp5_ASAP7_75t_L g1736 ( .A(n_1699), .B(n_1737), .Y(n_1736) );
AND2x2_ASAP7_75t_L g1786 ( .A(n_1699), .B(n_1787), .Y(n_1786) );
AND2x2_ASAP7_75t_L g1900 ( .A(n_1699), .B(n_1820), .Y(n_1900) );
AND2x2_ASAP7_75t_L g1914 ( .A(n_1699), .B(n_1815), .Y(n_1914) );
AND2x2_ASAP7_75t_L g1754 ( .A(n_1700), .B(n_1710), .Y(n_1754) );
INVx1_ASAP7_75t_L g1829 ( .A(n_1700), .Y(n_1829) );
AND2x2_ASAP7_75t_L g1853 ( .A(n_1700), .B(n_1768), .Y(n_1853) );
AND2x2_ASAP7_75t_L g1700 ( .A(n_1701), .B(n_1702), .Y(n_1700) );
INVx2_ASAP7_75t_SL g1738 ( .A(n_1702), .Y(n_1738) );
OAI22xp5_ASAP7_75t_L g1703 ( .A1(n_1704), .A2(n_1705), .B1(n_1706), .B2(n_1707), .Y(n_1703) );
BUFx6f_ASAP7_75t_L g1719 ( .A(n_1705), .Y(n_1719) );
INVx1_ASAP7_75t_L g1721 ( .A(n_1707), .Y(n_1721) );
INVx1_ASAP7_75t_L g1708 ( .A(n_1709), .Y(n_1708) );
NAND2xp5_ASAP7_75t_L g1709 ( .A(n_1710), .B(n_1715), .Y(n_1709) );
NOR2xp33_ASAP7_75t_L g1787 ( .A(n_1710), .B(n_1788), .Y(n_1787) );
AND2x2_ASAP7_75t_L g1828 ( .A(n_1710), .B(n_1815), .Y(n_1828) );
AND2x2_ASAP7_75t_L g1849 ( .A(n_1710), .B(n_1752), .Y(n_1849) );
NOR2xp33_ASAP7_75t_L g1902 ( .A(n_1710), .B(n_1775), .Y(n_1902) );
INVx2_ASAP7_75t_L g1710 ( .A(n_1711), .Y(n_1710) );
BUFx2_ASAP7_75t_L g1735 ( .A(n_1711), .Y(n_1735) );
AND2x2_ASAP7_75t_L g1767 ( .A(n_1711), .B(n_1768), .Y(n_1767) );
INVx2_ASAP7_75t_L g1774 ( .A(n_1711), .Y(n_1774) );
AND2x2_ASAP7_75t_L g1820 ( .A(n_1711), .B(n_1752), .Y(n_1820) );
NAND2xp5_ASAP7_75t_L g1859 ( .A(n_1711), .B(n_1793), .Y(n_1859) );
NAND2xp5_ASAP7_75t_L g1872 ( .A(n_1711), .B(n_1716), .Y(n_1872) );
AND2x2_ASAP7_75t_L g1881 ( .A(n_1711), .B(n_1796), .Y(n_1881) );
AND2x2_ASAP7_75t_L g1711 ( .A(n_1712), .B(n_1713), .Y(n_1711) );
INVx1_ASAP7_75t_L g1724 ( .A(n_1714), .Y(n_1724) );
BUFx3_ASAP7_75t_L g1779 ( .A(n_1714), .Y(n_1779) );
AND2x2_ASAP7_75t_L g1789 ( .A(n_1715), .B(n_1790), .Y(n_1789) );
INVx1_ASAP7_75t_L g1876 ( .A(n_1715), .Y(n_1876) );
AND2x4_ASAP7_75t_L g1715 ( .A(n_1716), .B(n_1728), .Y(n_1715) );
AND2x2_ASAP7_75t_L g1748 ( .A(n_1716), .B(n_1729), .Y(n_1748) );
HB1xp67_ASAP7_75t_L g1765 ( .A(n_1716), .Y(n_1765) );
AND2x2_ASAP7_75t_L g1773 ( .A(n_1716), .B(n_1774), .Y(n_1773) );
INVx2_ASAP7_75t_SL g1811 ( .A(n_1716), .Y(n_1811) );
INVx1_ASAP7_75t_L g1831 ( .A(n_1716), .Y(n_1831) );
NAND2xp5_ASAP7_75t_L g1857 ( .A(n_1716), .B(n_1790), .Y(n_1857) );
NOR2xp33_ASAP7_75t_L g1868 ( .A(n_1716), .B(n_1774), .Y(n_1868) );
CKINVDCx5p33_ASAP7_75t_R g1716 ( .A(n_1717), .Y(n_1716) );
AND2x2_ASAP7_75t_L g1793 ( .A(n_1717), .B(n_1728), .Y(n_1793) );
AND2x2_ASAP7_75t_L g1878 ( .A(n_1717), .B(n_1729), .Y(n_1878) );
OR2x2_ASAP7_75t_L g1717 ( .A(n_1718), .B(n_1723), .Y(n_1717) );
BUFx3_ASAP7_75t_L g1782 ( .A(n_1719), .Y(n_1782) );
HB1xp67_ASAP7_75t_L g1784 ( .A(n_1720), .Y(n_1784) );
INVx1_ASAP7_75t_L g1720 ( .A(n_1721), .Y(n_1720) );
OAI22xp5_ASAP7_75t_L g1723 ( .A1(n_1724), .A2(n_1725), .B1(n_1726), .B2(n_1727), .Y(n_1723) );
INVx2_ASAP7_75t_L g1745 ( .A(n_1726), .Y(n_1745) );
AND2x2_ASAP7_75t_L g1756 ( .A(n_1728), .B(n_1741), .Y(n_1756) );
OR2x2_ASAP7_75t_L g1770 ( .A(n_1728), .B(n_1771), .Y(n_1770) );
AOI22xp5_ASAP7_75t_L g1802 ( .A1(n_1728), .A2(n_1803), .B1(n_1804), .B2(n_1806), .Y(n_1802) );
INVx1_ASAP7_75t_L g1817 ( .A(n_1728), .Y(n_1817) );
NAND3xp33_ASAP7_75t_L g1867 ( .A(n_1728), .B(n_1815), .C(n_1868), .Y(n_1867) );
NOR2xp33_ASAP7_75t_L g1871 ( .A(n_1728), .B(n_1872), .Y(n_1871) );
INVx3_ASAP7_75t_L g1728 ( .A(n_1729), .Y(n_1728) );
AND2x2_ASAP7_75t_L g1739 ( .A(n_1729), .B(n_1740), .Y(n_1739) );
OR2x2_ASAP7_75t_L g1812 ( .A(n_1729), .B(n_1741), .Y(n_1812) );
AND2x2_ASAP7_75t_L g1729 ( .A(n_1730), .B(n_1731), .Y(n_1729) );
AOI211xp5_ASAP7_75t_L g1891 ( .A1(n_1732), .A2(n_1748), .B(n_1892), .C(n_1903), .Y(n_1891) );
INVx1_ASAP7_75t_L g1732 ( .A(n_1733), .Y(n_1732) );
OR2x2_ASAP7_75t_L g1733 ( .A(n_1734), .B(n_1736), .Y(n_1733) );
NAND2xp5_ASAP7_75t_L g1759 ( .A(n_1734), .B(n_1739), .Y(n_1759) );
NAND2xp5_ASAP7_75t_L g1841 ( .A(n_1734), .B(n_1842), .Y(n_1841) );
NAND2xp5_ASAP7_75t_L g1852 ( .A(n_1734), .B(n_1853), .Y(n_1852) );
OAI21xp33_ASAP7_75t_L g1915 ( .A1(n_1734), .A2(n_1829), .B(n_1916), .Y(n_1915) );
INVx2_ASAP7_75t_L g1734 ( .A(n_1735), .Y(n_1734) );
NAND2xp5_ASAP7_75t_L g1884 ( .A(n_1735), .B(n_1737), .Y(n_1884) );
NAND2xp5_ASAP7_75t_L g1896 ( .A(n_1735), .B(n_1817), .Y(n_1896) );
INVx1_ASAP7_75t_L g1875 ( .A(n_1737), .Y(n_1875) );
NOR2x1_ASAP7_75t_L g1911 ( .A(n_1738), .B(n_1768), .Y(n_1911) );
NAND2xp5_ASAP7_75t_L g1830 ( .A(n_1739), .B(n_1831), .Y(n_1830) );
AOI22xp5_ASAP7_75t_L g1847 ( .A1(n_1739), .A2(n_1797), .B1(n_1817), .B2(n_1848), .Y(n_1847) );
AOI322xp5_ASAP7_75t_L g1912 ( .A1(n_1739), .A2(n_1804), .A3(n_1839), .B1(n_1913), .B2(n_1914), .C1(n_1915), .C2(n_1917), .Y(n_1912) );
INVx1_ASAP7_75t_L g1790 ( .A(n_1740), .Y(n_1790) );
INVx1_ASAP7_75t_L g1801 ( .A(n_1740), .Y(n_1801) );
INVx1_ASAP7_75t_L g1740 ( .A(n_1741), .Y(n_1740) );
INVx1_ASAP7_75t_L g1771 ( .A(n_1741), .Y(n_1771) );
INVx1_ASAP7_75t_L g1796 ( .A(n_1741), .Y(n_1796) );
AND2x2_ASAP7_75t_L g1741 ( .A(n_1742), .B(n_1744), .Y(n_1741) );
OAI22xp5_ASAP7_75t_L g1746 ( .A1(n_1747), .A2(n_1749), .B1(n_1753), .B2(n_1755), .Y(n_1746) );
INVx1_ASAP7_75t_L g1747 ( .A(n_1748), .Y(n_1747) );
NAND2xp5_ASAP7_75t_L g1749 ( .A(n_1750), .B(n_1752), .Y(n_1749) );
OAI211xp5_ASAP7_75t_SL g1906 ( .A1(n_1750), .A2(n_1849), .B(n_1907), .C(n_1910), .Y(n_1906) );
INVx1_ASAP7_75t_L g1750 ( .A(n_1751), .Y(n_1750) );
OR2x2_ASAP7_75t_L g1855 ( .A(n_1751), .B(n_1788), .Y(n_1855) );
OR2x2_ASAP7_75t_L g1874 ( .A(n_1751), .B(n_1875), .Y(n_1874) );
INVx1_ASAP7_75t_L g1762 ( .A(n_1752), .Y(n_1762) );
NAND2xp5_ASAP7_75t_L g1766 ( .A(n_1752), .B(n_1767), .Y(n_1766) );
AND2x2_ASAP7_75t_L g1806 ( .A(n_1752), .B(n_1768), .Y(n_1806) );
INVx1_ASAP7_75t_L g1753 ( .A(n_1754), .Y(n_1753) );
OAI21xp33_ASAP7_75t_L g1901 ( .A1(n_1754), .A2(n_1789), .B(n_1902), .Y(n_1901) );
NAND2xp5_ASAP7_75t_L g1813 ( .A(n_1755), .B(n_1814), .Y(n_1813) );
INVx1_ASAP7_75t_L g1755 ( .A(n_1756), .Y(n_1755) );
AOI221xp5_ASAP7_75t_L g1837 ( .A1(n_1756), .A2(n_1838), .B1(n_1839), .B2(n_1840), .C(n_1843), .Y(n_1837) );
NAND2xp5_ASAP7_75t_L g1861 ( .A(n_1756), .B(n_1831), .Y(n_1861) );
AOI211xp5_ASAP7_75t_SL g1757 ( .A1(n_1758), .A2(n_1760), .B(n_1764), .C(n_1769), .Y(n_1757) );
INVxp67_ASAP7_75t_SL g1758 ( .A(n_1759), .Y(n_1758) );
NAND2xp5_ASAP7_75t_L g1760 ( .A(n_1761), .B(n_1763), .Y(n_1760) );
INVx1_ASAP7_75t_L g1838 ( .A(n_1761), .Y(n_1838) );
NOR2xp33_ASAP7_75t_L g1791 ( .A(n_1763), .B(n_1792), .Y(n_1791) );
INVx1_ASAP7_75t_L g1894 ( .A(n_1763), .Y(n_1894) );
NOR2xp33_ASAP7_75t_L g1764 ( .A(n_1765), .B(n_1766), .Y(n_1764) );
A2O1A1Ixp33_ASAP7_75t_L g1904 ( .A1(n_1765), .A2(n_1820), .B(n_1854), .C(n_1905), .Y(n_1904) );
NAND2xp5_ASAP7_75t_L g1818 ( .A(n_1766), .B(n_1819), .Y(n_1818) );
AND2x2_ASAP7_75t_L g1898 ( .A(n_1767), .B(n_1815), .Y(n_1898) );
AOI321xp33_ASAP7_75t_L g1879 ( .A1(n_1768), .A2(n_1880), .A3(n_1881), .B1(n_1882), .B2(n_1883), .C(n_1885), .Y(n_1879) );
A2O1A1Ixp33_ASAP7_75t_L g1769 ( .A1(n_1770), .A2(n_1772), .B(n_1775), .C(n_1777), .Y(n_1769) );
INVx1_ASAP7_75t_L g1905 ( .A(n_1770), .Y(n_1905) );
INVx1_ASAP7_75t_L g1772 ( .A(n_1773), .Y(n_1772) );
NAND2xp5_ASAP7_75t_L g1792 ( .A(n_1774), .B(n_1793), .Y(n_1792) );
INVx1_ASAP7_75t_L g1775 ( .A(n_1776), .Y(n_1775) );
INVx3_ASAP7_75t_L g1777 ( .A(n_1778), .Y(n_1777) );
INVx3_ASAP7_75t_L g1885 ( .A(n_1778), .Y(n_1885) );
OAI22xp33_ASAP7_75t_L g1780 ( .A1(n_1781), .A2(n_1782), .B1(n_1783), .B2(n_1784), .Y(n_1780) );
BUFx2_ASAP7_75t_SL g1919 ( .A(n_1784), .Y(n_1919) );
AOI21xp5_ASAP7_75t_L g1785 ( .A1(n_1786), .A2(n_1789), .B(n_1791), .Y(n_1785) );
INVx1_ASAP7_75t_L g1864 ( .A(n_1787), .Y(n_1864) );
NOR2xp33_ASAP7_75t_L g1799 ( .A(n_1788), .B(n_1792), .Y(n_1799) );
INVx1_ASAP7_75t_L g1815 ( .A(n_1788), .Y(n_1815) );
AND2x2_ASAP7_75t_L g1845 ( .A(n_1790), .B(n_1831), .Y(n_1845) );
INVx2_ASAP7_75t_L g1860 ( .A(n_1790), .Y(n_1860) );
INVx1_ASAP7_75t_L g1803 ( .A(n_1792), .Y(n_1803) );
AND2x2_ASAP7_75t_L g1839 ( .A(n_1793), .B(n_1796), .Y(n_1839) );
NAND2xp5_ASAP7_75t_L g1794 ( .A(n_1795), .B(n_1797), .Y(n_1794) );
INVx1_ASAP7_75t_L g1795 ( .A(n_1796), .Y(n_1795) );
NAND2xp5_ASAP7_75t_L g1825 ( .A(n_1796), .B(n_1826), .Y(n_1825) );
INVxp67_ASAP7_75t_L g1798 ( .A(n_1799), .Y(n_1798) );
OAI211xp5_ASAP7_75t_L g1800 ( .A1(n_1801), .A2(n_1802), .B(n_1807), .C(n_1832), .Y(n_1800) );
INVx1_ASAP7_75t_L g1823 ( .A(n_1801), .Y(n_1823) );
OAI211xp5_ASAP7_75t_SL g1886 ( .A1(n_1801), .A2(n_1887), .B(n_1891), .C(n_1912), .Y(n_1886) );
INVx1_ASAP7_75t_L g1909 ( .A(n_1801), .Y(n_1909) );
NAND2xp5_ASAP7_75t_L g1870 ( .A(n_1804), .B(n_1871), .Y(n_1870) );
INVx1_ASAP7_75t_L g1804 ( .A(n_1805), .Y(n_1804) );
INVx1_ASAP7_75t_L g1890 ( .A(n_1806), .Y(n_1890) );
AOI221xp5_ASAP7_75t_L g1807 ( .A1(n_1808), .A2(n_1820), .B1(n_1821), .B2(n_1823), .C(n_1824), .Y(n_1807) );
NAND3xp33_ASAP7_75t_L g1808 ( .A(n_1809), .B(n_1813), .C(n_1816), .Y(n_1808) );
INVx1_ASAP7_75t_L g1809 ( .A(n_1810), .Y(n_1809) );
NOR2xp33_ASAP7_75t_L g1810 ( .A(n_1811), .B(n_1812), .Y(n_1810) );
INVx2_ASAP7_75t_L g1819 ( .A(n_1811), .Y(n_1819) );
INVx1_ASAP7_75t_L g1826 ( .A(n_1811), .Y(n_1826) );
AND2x2_ASAP7_75t_L g1897 ( .A(n_1811), .B(n_1898), .Y(n_1897) );
INVxp67_ASAP7_75t_L g1834 ( .A(n_1813), .Y(n_1834) );
INVx1_ASAP7_75t_L g1846 ( .A(n_1814), .Y(n_1846) );
INVxp67_ASAP7_75t_L g1833 ( .A(n_1816), .Y(n_1833) );
NAND2xp5_ASAP7_75t_L g1816 ( .A(n_1817), .B(n_1818), .Y(n_1816) );
INVx1_ASAP7_75t_L g1821 ( .A(n_1822), .Y(n_1821) );
OAI22xp5_ASAP7_75t_L g1824 ( .A1(n_1825), .A2(n_1827), .B1(n_1829), .B2(n_1830), .Y(n_1824) );
INVx1_ASAP7_75t_L g1882 ( .A(n_1825), .Y(n_1882) );
INVx1_ASAP7_75t_L g1827 ( .A(n_1828), .Y(n_1827) );
NAND2xp5_ASAP7_75t_L g1880 ( .A(n_1829), .B(n_1875), .Y(n_1880) );
INVx1_ASAP7_75t_L g1917 ( .A(n_1830), .Y(n_1917) );
INVx1_ASAP7_75t_L g1835 ( .A(n_1831), .Y(n_1835) );
OAI21xp5_ASAP7_75t_L g1832 ( .A1(n_1833), .A2(n_1834), .B(n_1835), .Y(n_1832) );
NAND5xp2_ASAP7_75t_L g1836 ( .A(n_1837), .B(n_1847), .C(n_1850), .D(n_1865), .E(n_1879), .Y(n_1836) );
INVx1_ASAP7_75t_L g1840 ( .A(n_1841), .Y(n_1840) );
NOR2xp33_ASAP7_75t_L g1843 ( .A(n_1844), .B(n_1846), .Y(n_1843) );
INVx1_ASAP7_75t_L g1844 ( .A(n_1845), .Y(n_1844) );
O2A1O1Ixp33_ASAP7_75t_L g1850 ( .A1(n_1851), .A2(n_1854), .B(n_1856), .C(n_1858), .Y(n_1850) );
INVx1_ASAP7_75t_L g1851 ( .A(n_1852), .Y(n_1851) );
INVx1_ASAP7_75t_L g1916 ( .A(n_1853), .Y(n_1916) );
INVx1_ASAP7_75t_L g1854 ( .A(n_1855), .Y(n_1854) );
OAI22xp33_ASAP7_75t_L g1873 ( .A1(n_1855), .A2(n_1874), .B1(n_1876), .B2(n_1877), .Y(n_1873) );
INVx1_ASAP7_75t_L g1856 ( .A(n_1857), .Y(n_1856) );
INVx1_ASAP7_75t_L g1888 ( .A(n_1859), .Y(n_1888) );
OAI221xp5_ASAP7_75t_L g1892 ( .A1(n_1860), .A2(n_1861), .B1(n_1893), .B2(n_1899), .C(n_1901), .Y(n_1892) );
INVx1_ASAP7_75t_L g1862 ( .A(n_1863), .Y(n_1862) );
NOR3xp33_ASAP7_75t_SL g1865 ( .A(n_1866), .B(n_1869), .C(n_1873), .Y(n_1865) );
INVxp67_ASAP7_75t_L g1866 ( .A(n_1867), .Y(n_1866) );
INVxp67_ASAP7_75t_SL g1869 ( .A(n_1870), .Y(n_1869) );
INVx1_ASAP7_75t_L g1913 ( .A(n_1872), .Y(n_1913) );
NOR2xp33_ASAP7_75t_L g1889 ( .A(n_1876), .B(n_1890), .Y(n_1889) );
OR2x2_ASAP7_75t_L g1908 ( .A(n_1877), .B(n_1909), .Y(n_1908) );
CKINVDCx5p33_ASAP7_75t_R g1877 ( .A(n_1878), .Y(n_1877) );
INVx1_ASAP7_75t_L g1883 ( .A(n_1884), .Y(n_1883) );
AOI21xp33_ASAP7_75t_L g1893 ( .A1(n_1894), .A2(n_1895), .B(n_1897), .Y(n_1893) );
INVx1_ASAP7_75t_L g1895 ( .A(n_1896), .Y(n_1895) );
INVx1_ASAP7_75t_L g1899 ( .A(n_1900), .Y(n_1899) );
NAND2xp5_ASAP7_75t_SL g1903 ( .A(n_1904), .B(n_1906), .Y(n_1903) );
INVx1_ASAP7_75t_L g1907 ( .A(n_1908), .Y(n_1907) );
INVx1_ASAP7_75t_L g1910 ( .A(n_1911), .Y(n_1910) );
HB1xp67_ASAP7_75t_L g1918 ( .A(n_1919), .Y(n_1918) );
AND2x2_ASAP7_75t_L g1921 ( .A(n_1922), .B(n_1948), .Y(n_1921) );
NOR3xp33_ASAP7_75t_L g1922 ( .A(n_1923), .B(n_1930), .C(n_1931), .Y(n_1922) );
NAND2xp5_ASAP7_75t_L g1923 ( .A(n_1924), .B(n_1927), .Y(n_1923) );
OAI22xp5_ASAP7_75t_L g1939 ( .A1(n_1940), .A2(n_1941), .B1(n_1942), .B2(n_1944), .Y(n_1939) );
INVx1_ASAP7_75t_L g1942 ( .A(n_1943), .Y(n_1942) );
NAND3xp33_ASAP7_75t_L g1949 ( .A(n_1950), .B(n_1954), .C(n_1958), .Y(n_1949) );
CKINVDCx5p33_ASAP7_75t_R g1960 ( .A(n_1961), .Y(n_1960) );
BUFx2_ASAP7_75t_L g1961 ( .A(n_1962), .Y(n_1961) );
OAI21xp5_ASAP7_75t_L g2057 ( .A1(n_1963), .A2(n_2058), .B(n_2059), .Y(n_2057) );
BUFx3_ASAP7_75t_L g1965 ( .A(n_1966), .Y(n_1965) );
BUFx2_ASAP7_75t_L g1966 ( .A(n_1967), .Y(n_1966) );
INVx1_ASAP7_75t_L g1968 ( .A(n_1969), .Y(n_1968) );
INVx1_ASAP7_75t_L g1969 ( .A(n_1970), .Y(n_1969) );
NAND3x1_ASAP7_75t_L g1971 ( .A(n_1972), .B(n_2003), .C(n_2029), .Y(n_1971) );
OAI31xp33_ASAP7_75t_L g1972 ( .A1(n_1973), .A2(n_1980), .A3(n_1989), .B(n_2001), .Y(n_1972) );
INVx1_ASAP7_75t_L g1975 ( .A(n_1976), .Y(n_1975) );
INVx1_ASAP7_75t_L g1993 ( .A(n_1976), .Y(n_1993) );
INVx1_ASAP7_75t_L g1976 ( .A(n_1977), .Y(n_1976) );
CKINVDCx6p67_ASAP7_75t_R g1978 ( .A(n_1979), .Y(n_1978) );
INVx4_ASAP7_75t_L g1981 ( .A(n_1982), .Y(n_1981) );
AND2x4_ASAP7_75t_L g1995 ( .A(n_1983), .B(n_1996), .Y(n_1995) );
INVx1_ASAP7_75t_L g1983 ( .A(n_1984), .Y(n_1983) );
INVx4_ASAP7_75t_L g1985 ( .A(n_1986), .Y(n_1985) );
INVx1_ASAP7_75t_SL g1987 ( .A(n_1988), .Y(n_1987) );
CKINVDCx8_ASAP7_75t_R g1991 ( .A(n_1992), .Y(n_1991) );
AOI22xp33_ASAP7_75t_SL g1994 ( .A1(n_1995), .A2(n_1998), .B1(n_1999), .B2(n_2000), .Y(n_1994) );
INVx1_ASAP7_75t_L g1996 ( .A(n_1997), .Y(n_1996) );
AND4x1_ASAP7_75t_L g2003 ( .A(n_2004), .B(n_2011), .C(n_2014), .D(n_2023), .Y(n_2003) );
NAND3xp33_ASAP7_75t_L g2004 ( .A(n_2005), .B(n_2007), .C(n_2010), .Y(n_2004) );
INVx2_ASAP7_75t_L g2008 ( .A(n_2009), .Y(n_2008) );
NAND3xp33_ASAP7_75t_L g2014 ( .A(n_2015), .B(n_2016), .C(n_2021), .Y(n_2014) );
INVx1_ASAP7_75t_L g2017 ( .A(n_2018), .Y(n_2017) );
INVx1_ASAP7_75t_L g2019 ( .A(n_2020), .Y(n_2019) );
INVx1_ASAP7_75t_SL g2021 ( .A(n_2022), .Y(n_2021) );
INVx1_ASAP7_75t_L g2025 ( .A(n_2026), .Y(n_2025) );
OAI21xp5_ASAP7_75t_L g2029 ( .A1(n_2030), .A2(n_2047), .B(n_2054), .Y(n_2029) );
NAND3xp33_ASAP7_75t_L g2030 ( .A(n_2031), .B(n_2037), .C(n_2044), .Y(n_2030) );
INVxp67_ASAP7_75t_L g2035 ( .A(n_2036), .Y(n_2035) );
INVx1_ASAP7_75t_L g2046 ( .A(n_2036), .Y(n_2046) );
AOI22xp33_ASAP7_75t_L g2037 ( .A1(n_2038), .A2(n_2039), .B1(n_2040), .B2(n_2041), .Y(n_2037) );
INVx4_ASAP7_75t_L g2041 ( .A(n_2042), .Y(n_2041) );
INVx1_ASAP7_75t_L g2049 ( .A(n_2043), .Y(n_2049) );
AND2x4_ASAP7_75t_L g2051 ( .A(n_2043), .B(n_2052), .Y(n_2051) );
CKINVDCx11_ASAP7_75t_R g2044 ( .A(n_2045), .Y(n_2044) );
INVx5_ASAP7_75t_SL g2050 ( .A(n_2051), .Y(n_2050) );
INVx1_ASAP7_75t_L g2052 ( .A(n_2053), .Y(n_2052) );
CKINVDCx16_ASAP7_75t_R g2054 ( .A(n_2055), .Y(n_2054) );
BUFx2_ASAP7_75t_L g2056 ( .A(n_2057), .Y(n_2056) );
endmodule