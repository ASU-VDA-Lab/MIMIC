module real_aes_6928_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_555;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_552;
wire n_402;
wire n_617;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_193;
wire n_293;
wire n_162;
wire n_749;
wire n_385;
wire n_275;
wire n_214;
wire n_358;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_729;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g554 ( .A1(n_0), .A2(n_161), .B(n_555), .C(n_558), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_1), .B(n_499), .Y(n_559) );
NAND3xp33_ASAP7_75t_SL g107 ( .A(n_2), .B(n_108), .C(n_109), .Y(n_107) );
INVx1_ASAP7_75t_L g123 ( .A(n_2), .Y(n_123) );
INVx1_ASAP7_75t_L g195 ( .A(n_3), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g533 ( .A(n_4), .B(n_153), .Y(n_533) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_5), .A2(n_468), .B(n_493), .Y(n_492) );
AO21x2_ASAP7_75t_L g483 ( .A1(n_6), .A2(n_138), .B(n_484), .Y(n_483) );
AOI22xp33_ASAP7_75t_L g224 ( .A1(n_7), .A2(n_35), .B1(n_147), .B2(n_225), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_8), .B(n_138), .Y(n_164) );
AND2x6_ASAP7_75t_L g162 ( .A(n_9), .B(n_163), .Y(n_162) );
A2O1A1Ixp33_ASAP7_75t_L g457 ( .A1(n_10), .A2(n_162), .B(n_458), .C(n_460), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_11), .B(n_106), .Y(n_105) );
NOR2xp33_ASAP7_75t_L g124 ( .A(n_11), .B(n_36), .Y(n_124) );
INVx1_ASAP7_75t_L g143 ( .A(n_12), .Y(n_143) );
INVx1_ASAP7_75t_L g188 ( .A(n_13), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_14), .B(n_151), .Y(n_231) );
NAND2xp5_ASAP7_75t_SL g489 ( .A(n_15), .B(n_153), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_16), .B(n_139), .Y(n_200) );
AO32x2_ASAP7_75t_L g222 ( .A1(n_17), .A2(n_138), .A3(n_168), .B1(n_179), .B2(n_223), .Y(n_222) );
NAND2xp5_ASAP7_75t_SL g235 ( .A(n_18), .B(n_147), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_19), .B(n_139), .Y(n_197) );
AOI22xp33_ASAP7_75t_L g226 ( .A1(n_20), .A2(n_53), .B1(n_147), .B2(n_225), .Y(n_226) );
AOI22xp33_ASAP7_75t_SL g247 ( .A1(n_21), .A2(n_80), .B1(n_147), .B2(n_151), .Y(n_247) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_22), .B(n_147), .Y(n_217) );
A2O1A1Ixp33_ASAP7_75t_L g518 ( .A1(n_23), .A2(n_179), .B(n_458), .C(n_519), .Y(n_518) );
A2O1A1Ixp33_ASAP7_75t_L g486 ( .A1(n_24), .A2(n_179), .B(n_458), .C(n_487), .Y(n_486) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_25), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_26), .B(n_181), .Y(n_180) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_27), .Y(n_125) );
AOI21xp5_ASAP7_75t_L g551 ( .A1(n_28), .A2(n_468), .B(n_552), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_29), .B(n_181), .Y(n_219) );
INVx2_ASAP7_75t_L g149 ( .A(n_30), .Y(n_149) );
A2O1A1Ixp33_ASAP7_75t_L g506 ( .A1(n_31), .A2(n_470), .B(n_478), .C(n_507), .Y(n_506) );
NAND2xp5_ASAP7_75t_SL g171 ( .A(n_32), .B(n_147), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_33), .B(n_181), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_34), .B(n_233), .Y(n_488) );
INVx1_ASAP7_75t_L g106 ( .A(n_36), .Y(n_106) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_37), .B(n_517), .Y(n_516) );
CKINVDCx20_ASAP7_75t_R g464 ( .A(n_38), .Y(n_464) );
AOI222xp33_ASAP7_75t_SL g126 ( .A1(n_39), .A2(n_78), .B1(n_127), .B2(n_732), .C1(n_733), .C2(n_737), .Y(n_126) );
CKINVDCx16_ASAP7_75t_R g732 ( .A(n_39), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_40), .B(n_153), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_41), .B(n_468), .Y(n_485) );
OAI22xp5_ASAP7_75t_SL g747 ( .A1(n_42), .A2(n_77), .B1(n_441), .B2(n_748), .Y(n_747) );
CKINVDCx20_ASAP7_75t_R g748 ( .A(n_42), .Y(n_748) );
A2O1A1Ixp33_ASAP7_75t_L g469 ( .A1(n_43), .A2(n_470), .B(n_472), .C(n_478), .Y(n_469) );
AOI22xp33_ASAP7_75t_L g100 ( .A1(n_44), .A2(n_101), .B1(n_112), .B2(n_751), .Y(n_100) );
NAND2xp5_ASAP7_75t_SL g146 ( .A(n_45), .B(n_147), .Y(n_146) );
INVx1_ASAP7_75t_L g556 ( .A(n_46), .Y(n_556) );
AOI22xp33_ASAP7_75t_L g245 ( .A1(n_47), .A2(n_89), .B1(n_225), .B2(n_246), .Y(n_245) );
INVx1_ASAP7_75t_L g473 ( .A(n_48), .Y(n_473) );
NAND2xp5_ASAP7_75t_SL g157 ( .A(n_49), .B(n_147), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_50), .B(n_147), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_51), .B(n_468), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_52), .B(n_159), .Y(n_158) );
AOI22xp33_ASAP7_75t_SL g204 ( .A1(n_54), .A2(n_58), .B1(n_147), .B2(n_151), .Y(n_204) );
CKINVDCx20_ASAP7_75t_R g524 ( .A(n_55), .Y(n_524) );
NAND2xp5_ASAP7_75t_SL g176 ( .A(n_56), .B(n_147), .Y(n_176) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_57), .B(n_147), .Y(n_230) );
INVx1_ASAP7_75t_L g163 ( .A(n_59), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_60), .B(n_468), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_61), .B(n_499), .Y(n_498) );
A2O1A1Ixp33_ASAP7_75t_L g495 ( .A1(n_62), .A2(n_159), .B(n_191), .C(n_496), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_63), .B(n_147), .Y(n_196) );
INVx1_ASAP7_75t_L g142 ( .A(n_64), .Y(n_142) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_65), .Y(n_117) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_66), .B(n_153), .Y(n_509) );
AO32x2_ASAP7_75t_L g243 ( .A1(n_67), .A2(n_138), .A3(n_179), .B1(n_244), .B2(n_248), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_68), .B(n_154), .Y(n_461) );
INVx1_ASAP7_75t_L g174 ( .A(n_69), .Y(n_174) );
INVx1_ASAP7_75t_L g214 ( .A(n_70), .Y(n_214) );
CKINVDCx16_ASAP7_75t_R g553 ( .A(n_71), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_72), .B(n_475), .Y(n_520) );
A2O1A1Ixp33_ASAP7_75t_L g530 ( .A1(n_73), .A2(n_458), .B(n_478), .C(n_531), .Y(n_530) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_74), .B(n_151), .Y(n_215) );
CKINVDCx16_ASAP7_75t_R g494 ( .A(n_75), .Y(n_494) );
INVx1_ASAP7_75t_L g111 ( .A(n_76), .Y(n_111) );
OAI22xp5_ASAP7_75t_SL g129 ( .A1(n_77), .A2(n_130), .B1(n_440), .B2(n_441), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g441 ( .A(n_77), .Y(n_441) );
NAND2xp5_ASAP7_75t_SL g521 ( .A(n_79), .B(n_474), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_81), .B(n_225), .Y(n_236) );
CKINVDCx20_ASAP7_75t_R g511 ( .A(n_82), .Y(n_511) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_83), .B(n_151), .Y(n_218) );
INVx2_ASAP7_75t_L g140 ( .A(n_84), .Y(n_140) );
CKINVDCx20_ASAP7_75t_R g537 ( .A(n_85), .Y(n_537) );
NAND2xp5_ASAP7_75t_SL g462 ( .A(n_86), .B(n_178), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_87), .B(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g108 ( .A(n_88), .Y(n_108) );
OR2x2_ASAP7_75t_L g120 ( .A(n_88), .B(n_121), .Y(n_120) );
OR2x2_ASAP7_75t_L g444 ( .A(n_88), .B(n_122), .Y(n_444) );
AOI22xp33_ASAP7_75t_L g203 ( .A1(n_90), .A2(n_99), .B1(n_151), .B2(n_152), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_91), .B(n_468), .Y(n_505) );
INVx1_ASAP7_75t_L g508 ( .A(n_92), .Y(n_508) );
INVxp67_ASAP7_75t_L g497 ( .A(n_93), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_94), .B(n_151), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_95), .B(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g454 ( .A(n_96), .Y(n_454) );
INVx1_ASAP7_75t_L g532 ( .A(n_97), .Y(n_532) );
AND2x2_ASAP7_75t_L g480 ( .A(n_98), .B(n_181), .Y(n_480) );
INVx1_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
CKINVDCx12_ASAP7_75t_R g103 ( .A(n_104), .Y(n_103) );
INVx1_ASAP7_75t_SL g752 ( .A(n_104), .Y(n_752) );
OR2x2_ASAP7_75t_L g104 ( .A(n_105), .B(n_107), .Y(n_104) );
OR2x2_ASAP7_75t_L g731 ( .A(n_108), .B(n_122), .Y(n_731) );
NOR2x2_ASAP7_75t_L g739 ( .A(n_108), .B(n_121), .Y(n_739) );
INVx1_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
AOI22x1_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_126), .B1(n_740), .B2(n_741), .Y(n_112) );
NOR2xp33_ASAP7_75t_L g113 ( .A(n_114), .B(n_118), .Y(n_113) );
INVx1_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
BUFx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_SL g740 ( .A(n_116), .Y(n_740) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
AOI21xp5_ASAP7_75t_L g741 ( .A1(n_118), .A2(n_742), .B(n_749), .Y(n_741) );
NOR2xp33_ASAP7_75t_SL g118 ( .A(n_119), .B(n_125), .Y(n_118) );
HB1xp67_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx1_ASAP7_75t_SL g750 ( .A(n_120), .Y(n_750) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
AND2x2_ASAP7_75t_L g122 ( .A(n_123), .B(n_124), .Y(n_122) );
OAI22xp5_ASAP7_75t_SL g127 ( .A1(n_128), .A2(n_442), .B1(n_445), .B2(n_729), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
OAI22xp5_ASAP7_75t_SL g733 ( .A1(n_129), .A2(n_734), .B1(n_735), .B2(n_736), .Y(n_733) );
INVx2_ASAP7_75t_L g440 ( .A(n_130), .Y(n_440) );
OAI22xp5_ASAP7_75t_L g745 ( .A1(n_130), .A2(n_440), .B1(n_746), .B2(n_747), .Y(n_745) );
NAND2x1p5_ASAP7_75t_L g130 ( .A(n_131), .B(n_364), .Y(n_130) );
AND2x2_ASAP7_75t_SL g131 ( .A(n_132), .B(n_322), .Y(n_131) );
NOR4xp25_ASAP7_75t_L g132 ( .A(n_133), .B(n_262), .C(n_298), .D(n_312), .Y(n_132) );
OAI221xp5_ASAP7_75t_SL g133 ( .A1(n_134), .A2(n_206), .B1(n_238), .B2(n_249), .C(n_253), .Y(n_133) );
NAND2xp5_ASAP7_75t_SL g396 ( .A(n_134), .B(n_397), .Y(n_396) );
OR2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_182), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
AND2x2_ASAP7_75t_L g136 ( .A(n_137), .B(n_165), .Y(n_136) );
AND2x2_ASAP7_75t_L g259 ( .A(n_137), .B(n_166), .Y(n_259) );
INVx3_ASAP7_75t_L g267 ( .A(n_137), .Y(n_267) );
AND2x2_ASAP7_75t_L g321 ( .A(n_137), .B(n_185), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_137), .B(n_184), .Y(n_357) );
AND2x2_ASAP7_75t_L g415 ( .A(n_137), .B(n_277), .Y(n_415) );
OA21x2_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_144), .B(n_164), .Y(n_137) );
INVx4_ASAP7_75t_L g205 ( .A(n_138), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_138), .A2(n_485), .B(n_486), .Y(n_484) );
HB1xp67_ASAP7_75t_L g491 ( .A(n_138), .Y(n_491) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx1_ASAP7_75t_L g168 ( .A(n_139), .Y(n_168) );
AND2x2_ASAP7_75t_L g139 ( .A(n_140), .B(n_141), .Y(n_139) );
AND2x2_ASAP7_75t_SL g181 ( .A(n_140), .B(n_141), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_142), .B(n_143), .Y(n_141) );
OAI21xp5_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_156), .B(n_162), .Y(n_144) );
AOI21xp5_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_150), .B(n_153), .Y(n_145) );
INVx3_ASAP7_75t_L g213 ( .A(n_147), .Y(n_213) );
HB1xp67_ASAP7_75t_L g534 ( .A(n_147), .Y(n_534) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx1_ASAP7_75t_L g225 ( .A(n_148), .Y(n_225) );
BUFx3_ASAP7_75t_L g246 ( .A(n_148), .Y(n_246) );
AND2x6_ASAP7_75t_L g458 ( .A(n_148), .B(n_459), .Y(n_458) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g152 ( .A(n_149), .Y(n_152) );
INVx1_ASAP7_75t_L g160 ( .A(n_149), .Y(n_160) );
INVx2_ASAP7_75t_L g189 ( .A(n_151), .Y(n_189) );
INVx3_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g161 ( .A(n_153), .Y(n_161) );
AOI21xp5_ASAP7_75t_L g170 ( .A1(n_153), .A2(n_171), .B(n_172), .Y(n_170) );
O2A1O1Ixp5_ASAP7_75t_SL g212 ( .A1(n_153), .A2(n_213), .B(n_214), .C(n_215), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_153), .B(n_497), .Y(n_496) );
INVx5_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
OAI22xp5_ASAP7_75t_SL g244 ( .A1(n_154), .A2(n_178), .B1(n_245), .B2(n_247), .Y(n_244) );
INVx3_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
BUFx6f_ASAP7_75t_L g178 ( .A(n_155), .Y(n_178) );
BUFx6f_ASAP7_75t_L g193 ( .A(n_155), .Y(n_193) );
INVx1_ASAP7_75t_L g233 ( .A(n_155), .Y(n_233) );
AND2x2_ASAP7_75t_L g456 ( .A(n_155), .B(n_160), .Y(n_456) );
INVx1_ASAP7_75t_L g459 ( .A(n_155), .Y(n_459) );
AOI21xp5_ASAP7_75t_L g156 ( .A1(n_157), .A2(n_158), .B(n_161), .Y(n_156) );
INVx2_ASAP7_75t_L g175 ( .A(n_159), .Y(n_175) );
INVx1_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
O2A1O1Ixp33_ASAP7_75t_L g194 ( .A1(n_161), .A2(n_175), .B(n_195), .C(n_196), .Y(n_194) );
OAI22xp5_ASAP7_75t_L g202 ( .A1(n_161), .A2(n_178), .B1(n_203), .B2(n_204), .Y(n_202) );
OAI22xp5_ASAP7_75t_L g223 ( .A1(n_161), .A2(n_178), .B1(n_224), .B2(n_226), .Y(n_223) );
BUFx3_ASAP7_75t_L g179 ( .A(n_162), .Y(n_179) );
OAI21xp5_ASAP7_75t_L g186 ( .A1(n_162), .A2(n_187), .B(n_194), .Y(n_186) );
OAI21xp5_ASAP7_75t_L g211 ( .A1(n_162), .A2(n_212), .B(n_216), .Y(n_211) );
OAI21xp5_ASAP7_75t_L g228 ( .A1(n_162), .A2(n_229), .B(n_234), .Y(n_228) );
NAND2x1p5_ASAP7_75t_L g455 ( .A(n_162), .B(n_456), .Y(n_455) );
AND2x4_ASAP7_75t_L g468 ( .A(n_162), .B(n_456), .Y(n_468) );
INVx4_ASAP7_75t_SL g479 ( .A(n_162), .Y(n_479) );
AND2x2_ASAP7_75t_L g250 ( .A(n_165), .B(n_251), .Y(n_250) );
AND2x2_ASAP7_75t_L g264 ( .A(n_165), .B(n_185), .Y(n_264) );
INVx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_166), .B(n_185), .Y(n_279) );
AND2x2_ASAP7_75t_L g291 ( .A(n_166), .B(n_267), .Y(n_291) );
OR2x2_ASAP7_75t_L g293 ( .A(n_166), .B(n_251), .Y(n_293) );
AND2x2_ASAP7_75t_L g328 ( .A(n_166), .B(n_251), .Y(n_328) );
HB1xp67_ASAP7_75t_L g373 ( .A(n_166), .Y(n_373) );
INVx1_ASAP7_75t_L g381 ( .A(n_166), .Y(n_381) );
OA21x2_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_169), .B(n_180), .Y(n_166) );
OA21x2_ASAP7_75t_L g185 ( .A1(n_167), .A2(n_186), .B(n_197), .Y(n_185) );
INVx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
NOR2xp33_ASAP7_75t_L g463 ( .A(n_168), .B(n_464), .Y(n_463) );
OAI21xp5_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_173), .B(n_179), .Y(n_169) );
O2A1O1Ixp5_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_175), .B(n_176), .C(n_177), .Y(n_173) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_175), .A2(n_520), .B(n_521), .Y(n_519) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_177), .A2(n_235), .B(n_236), .Y(n_234) );
INVx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVx4_ASAP7_75t_L g557 ( .A(n_178), .Y(n_557) );
NAND3xp33_ASAP7_75t_L g201 ( .A(n_179), .B(n_202), .C(n_205), .Y(n_201) );
OA21x2_ASAP7_75t_L g210 ( .A1(n_181), .A2(n_211), .B(n_219), .Y(n_210) );
OA21x2_ASAP7_75t_L g227 ( .A1(n_181), .A2(n_228), .B(n_237), .Y(n_227) );
INVx2_ASAP7_75t_L g248 ( .A(n_181), .Y(n_248) );
AOI21xp5_ASAP7_75t_L g466 ( .A1(n_181), .A2(n_467), .B(n_469), .Y(n_466) );
AOI21xp5_ASAP7_75t_L g504 ( .A1(n_181), .A2(n_505), .B(n_506), .Y(n_504) );
INVx1_ASAP7_75t_L g525 ( .A(n_181), .Y(n_525) );
OAI221xp5_ASAP7_75t_L g298 ( .A1(n_182), .A2(n_299), .B1(n_303), .B2(n_307), .C(n_308), .Y(n_298) );
INVx1_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
AND2x2_ASAP7_75t_L g258 ( .A(n_183), .B(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g183 ( .A(n_184), .B(n_198), .Y(n_183) );
INVx2_ASAP7_75t_L g257 ( .A(n_184), .Y(n_257) );
AND2x2_ASAP7_75t_L g310 ( .A(n_184), .B(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g329 ( .A(n_184), .B(n_267), .Y(n_329) );
INVx2_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
AND2x2_ASAP7_75t_L g392 ( .A(n_185), .B(n_267), .Y(n_392) );
O2A1O1Ixp33_ASAP7_75t_L g187 ( .A1(n_188), .A2(n_189), .B(n_190), .C(n_191), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g460 ( .A1(n_189), .A2(n_461), .B(n_462), .Y(n_460) );
AOI21xp5_ASAP7_75t_L g487 ( .A1(n_189), .A2(n_488), .B(n_489), .Y(n_487) );
O2A1O1Ixp33_ASAP7_75t_L g531 ( .A1(n_191), .A2(n_532), .B(n_533), .C(n_534), .Y(n_531) );
INVx1_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_192), .A2(n_217), .B(n_218), .Y(n_216) );
INVx4_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
INVx2_ASAP7_75t_L g475 ( .A(n_193), .Y(n_475) );
AND2x2_ASAP7_75t_L g314 ( .A(n_198), .B(n_259), .Y(n_314) );
OAI322xp33_ASAP7_75t_L g382 ( .A1(n_198), .A2(n_338), .A3(n_383), .B1(n_385), .B2(n_388), .C1(n_390), .C2(n_394), .Y(n_382) );
INVx3_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
NOR2x1_ASAP7_75t_L g265 ( .A(n_199), .B(n_266), .Y(n_265) );
INVx2_ASAP7_75t_L g278 ( .A(n_199), .Y(n_278) );
AND2x2_ASAP7_75t_L g387 ( .A(n_199), .B(n_267), .Y(n_387) );
AND2x2_ASAP7_75t_L g419 ( .A(n_199), .B(n_291), .Y(n_419) );
OR2x2_ASAP7_75t_L g422 ( .A(n_199), .B(n_423), .Y(n_422) );
AND2x4_ASAP7_75t_L g199 ( .A(n_200), .B(n_201), .Y(n_199) );
INVx1_ASAP7_75t_L g252 ( .A(n_200), .Y(n_252) );
AO21x1_ASAP7_75t_L g251 ( .A1(n_202), .A2(n_205), .B(n_252), .Y(n_251) );
AO21x2_ASAP7_75t_L g452 ( .A1(n_205), .A2(n_453), .B(n_463), .Y(n_452) );
INVx3_ASAP7_75t_L g499 ( .A(n_205), .Y(n_499) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_205), .B(n_511), .Y(n_510) );
AO21x2_ASAP7_75t_L g528 ( .A1(n_205), .A2(n_529), .B(n_536), .Y(n_528) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_205), .B(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
AND2x2_ASAP7_75t_L g207 ( .A(n_208), .B(n_220), .Y(n_207) );
INVx1_ASAP7_75t_L g435 ( .A(n_208), .Y(n_435) );
INVx1_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
OR2x2_ASAP7_75t_L g240 ( .A(n_209), .B(n_227), .Y(n_240) );
INVx2_ASAP7_75t_L g275 ( .A(n_209), .Y(n_275) );
INVx2_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
INVx2_ASAP7_75t_L g297 ( .A(n_210), .Y(n_297) );
HB1xp67_ASAP7_75t_L g305 ( .A(n_210), .Y(n_305) );
OR2x2_ASAP7_75t_L g429 ( .A(n_210), .B(n_430), .Y(n_429) );
AND2x2_ASAP7_75t_L g254 ( .A(n_220), .B(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g294 ( .A(n_220), .B(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g346 ( .A(n_220), .B(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g220 ( .A(n_221), .B(n_227), .Y(n_220) );
AND2x2_ASAP7_75t_L g241 ( .A(n_221), .B(n_242), .Y(n_241) );
NOR2xp67_ASAP7_75t_L g301 ( .A(n_221), .B(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g355 ( .A(n_221), .B(n_243), .Y(n_355) );
OR2x2_ASAP7_75t_L g363 ( .A(n_221), .B(n_297), .Y(n_363) );
INVx2_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
BUFx2_ASAP7_75t_L g272 ( .A(n_222), .Y(n_272) );
AND2x2_ASAP7_75t_L g282 ( .A(n_222), .B(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g306 ( .A(n_222), .B(n_227), .Y(n_306) );
AND2x2_ASAP7_75t_L g370 ( .A(n_222), .B(n_243), .Y(n_370) );
NOR2xp33_ASAP7_75t_L g260 ( .A(n_227), .B(n_261), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_227), .B(n_275), .Y(n_274) );
INVx2_ASAP7_75t_L g283 ( .A(n_227), .Y(n_283) );
INVx1_ASAP7_75t_L g288 ( .A(n_227), .Y(n_288) );
AND2x2_ASAP7_75t_L g300 ( .A(n_227), .B(n_301), .Y(n_300) );
HB1xp67_ASAP7_75t_L g378 ( .A(n_227), .Y(n_378) );
INVx1_ASAP7_75t_L g430 ( .A(n_227), .Y(n_430) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_230), .A2(n_231), .B(n_232), .Y(n_229) );
INVx1_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_239), .B(n_241), .Y(n_238) );
AND2x2_ASAP7_75t_L g407 ( .A(n_239), .B(n_316), .Y(n_407) );
INVx2_ASAP7_75t_SL g239 ( .A(n_240), .Y(n_239) );
AND2x2_ASAP7_75t_L g334 ( .A(n_241), .B(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g433 ( .A(n_241), .B(n_368), .Y(n_433) );
INVx1_ASAP7_75t_L g255 ( .A(n_242), .Y(n_255) );
AND2x2_ASAP7_75t_L g281 ( .A(n_242), .B(n_275), .Y(n_281) );
BUFx2_ASAP7_75t_L g340 ( .A(n_242), .Y(n_340) );
INVx1_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
BUFx6f_ASAP7_75t_L g261 ( .A(n_243), .Y(n_261) );
INVx1_ASAP7_75t_L g271 ( .A(n_243), .Y(n_271) );
HB1xp67_ASAP7_75t_L g477 ( .A(n_246), .Y(n_477) );
INVx2_ASAP7_75t_L g558 ( .A(n_246), .Y(n_558) );
INVx1_ASAP7_75t_L g522 ( .A(n_248), .Y(n_522) );
NOR2xp67_ASAP7_75t_L g409 ( .A(n_249), .B(n_256), .Y(n_409) );
INVx2_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
AOI32xp33_ASAP7_75t_L g253 ( .A1(n_250), .A2(n_254), .A3(n_256), .B1(n_258), .B2(n_260), .Y(n_253) );
AND2x2_ASAP7_75t_L g393 ( .A(n_250), .B(n_266), .Y(n_393) );
AND2x2_ASAP7_75t_L g431 ( .A(n_250), .B(n_329), .Y(n_431) );
INVx1_ASAP7_75t_L g311 ( .A(n_251), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_255), .B(n_317), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_256), .B(n_291), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_256), .B(n_259), .Y(n_307) );
NAND2xp5_ASAP7_75t_SL g410 ( .A(n_256), .B(n_328), .Y(n_410) );
OR2x2_ASAP7_75t_L g424 ( .A(n_256), .B(n_293), .Y(n_424) );
INVx3_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
AND2x2_ASAP7_75t_L g351 ( .A(n_257), .B(n_259), .Y(n_351) );
OR2x2_ASAP7_75t_L g360 ( .A(n_257), .B(n_347), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_259), .B(n_310), .Y(n_332) );
INVx2_ASAP7_75t_L g347 ( .A(n_261), .Y(n_347) );
OR2x2_ASAP7_75t_L g362 ( .A(n_261), .B(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_L g377 ( .A(n_261), .B(n_378), .Y(n_377) );
A2O1A1Ixp33_ASAP7_75t_L g434 ( .A1(n_261), .A2(n_354), .B(n_435), .C(n_436), .Y(n_434) );
OAI321xp33_ASAP7_75t_L g262 ( .A1(n_263), .A2(n_268), .A3(n_273), .B1(n_276), .B2(n_280), .C(n_284), .Y(n_262) );
INVx1_ASAP7_75t_L g375 ( .A(n_263), .Y(n_375) );
NAND2x1p5_ASAP7_75t_L g263 ( .A(n_264), .B(n_265), .Y(n_263) );
AND2x2_ASAP7_75t_L g386 ( .A(n_264), .B(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g338 ( .A(n_266), .Y(n_338) );
INVx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_267), .B(n_381), .Y(n_398) );
OAI221xp5_ASAP7_75t_L g405 ( .A1(n_268), .A2(n_406), .B1(n_408), .B2(n_410), .C(n_411), .Y(n_405) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_272), .Y(n_269) );
AND2x2_ASAP7_75t_L g343 ( .A(n_270), .B(n_317), .Y(n_343) );
HB1xp67_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_271), .B(n_297), .Y(n_296) );
INVx2_ASAP7_75t_L g316 ( .A(n_272), .Y(n_316) );
A2O1A1Ixp33_ASAP7_75t_L g358 ( .A1(n_273), .A2(n_314), .B(n_359), .C(n_361), .Y(n_358) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g325 ( .A(n_275), .B(n_282), .Y(n_325) );
BUFx2_ASAP7_75t_L g335 ( .A(n_275), .Y(n_335) );
INVx1_ASAP7_75t_L g350 ( .A(n_275), .Y(n_350) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
NOR2xp33_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
OR2x2_ASAP7_75t_L g356 ( .A(n_278), .B(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g439 ( .A(n_278), .Y(n_439) );
INVx1_ASAP7_75t_L g432 ( .A(n_279), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_281), .B(n_282), .Y(n_280) );
AND2x2_ASAP7_75t_L g285 ( .A(n_281), .B(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g389 ( .A(n_281), .B(n_306), .Y(n_389) );
INVx1_ASAP7_75t_L g318 ( .A(n_282), .Y(n_318) );
AOI22xp5_ASAP7_75t_L g284 ( .A1(n_285), .A2(n_289), .B1(n_292), .B2(n_294), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_286), .B(n_402), .Y(n_401) );
INVxp67_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
AND2x4_ASAP7_75t_L g354 ( .A(n_287), .B(n_355), .Y(n_354) );
BUFx3_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_SL g317 ( .A(n_288), .B(n_297), .Y(n_317) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g309 ( .A(n_291), .B(n_310), .Y(n_309) );
INVx1_ASAP7_75t_SL g292 ( .A(n_293), .Y(n_292) );
OR2x2_ASAP7_75t_L g319 ( .A(n_293), .B(n_320), .Y(n_319) );
INVx1_ASAP7_75t_SL g295 ( .A(n_296), .Y(n_295) );
OAI221xp5_ASAP7_75t_L g413 ( .A1(n_296), .A2(n_414), .B1(n_416), .B2(n_417), .C(n_418), .Y(n_413) );
INVx1_ASAP7_75t_L g302 ( .A(n_297), .Y(n_302) );
HB1xp67_ASAP7_75t_L g368 ( .A(n_297), .Y(n_368) );
INVx1_ASAP7_75t_SL g299 ( .A(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_300), .B(n_419), .Y(n_418) );
OAI21xp5_ASAP7_75t_L g308 ( .A1(n_301), .A2(n_306), .B(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_304), .B(n_314), .Y(n_411) );
AND2x2_ASAP7_75t_L g304 ( .A(n_305), .B(n_306), .Y(n_304) );
INVx1_ASAP7_75t_L g380 ( .A(n_305), .Y(n_380) );
AND2x2_ASAP7_75t_L g339 ( .A(n_306), .B(n_340), .Y(n_339) );
INVx2_ASAP7_75t_L g428 ( .A(n_306), .Y(n_428) );
INVx1_ASAP7_75t_L g344 ( .A(n_309), .Y(n_344) );
INVx1_ASAP7_75t_L g399 ( .A(n_310), .Y(n_399) );
OAI22xp5_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_315), .B1(n_318), .B2(n_319), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_316), .B(n_350), .Y(n_349) );
INVx2_ASAP7_75t_L g384 ( .A(n_317), .Y(n_384) );
NAND2xp5_ASAP7_75t_SL g421 ( .A(n_317), .B(n_355), .Y(n_421) );
OR2x2_ASAP7_75t_L g394 ( .A(n_318), .B(n_347), .Y(n_394) );
INVx1_ASAP7_75t_L g333 ( .A(n_319), .Y(n_333) );
INVx1_ASAP7_75t_SL g320 ( .A(n_321), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_321), .B(n_372), .Y(n_371) );
NOR3xp33_ASAP7_75t_L g322 ( .A(n_323), .B(n_341), .C(n_352), .Y(n_322) );
OAI211xp5_ASAP7_75t_L g323 ( .A1(n_324), .A2(n_326), .B(n_330), .C(n_336), .Y(n_323) );
INVxp67_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
AOI221xp5_ASAP7_75t_L g395 ( .A1(n_325), .A2(n_396), .B1(n_400), .B2(n_403), .C(n_405), .Y(n_395) );
INVx1_ASAP7_75t_SL g326 ( .A(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g327 ( .A(n_328), .B(n_329), .Y(n_327) );
AND2x2_ASAP7_75t_L g337 ( .A(n_328), .B(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g391 ( .A(n_328), .B(n_392), .Y(n_391) );
OAI211xp5_ASAP7_75t_L g376 ( .A1(n_329), .A2(n_377), .B(n_379), .C(n_381), .Y(n_376) );
INVx2_ASAP7_75t_L g423 ( .A(n_329), .Y(n_423) );
OAI21xp5_ASAP7_75t_SL g330 ( .A1(n_331), .A2(n_333), .B(n_334), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g402 ( .A(n_335), .B(n_355), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_337), .B(n_339), .Y(n_336) );
OAI21xp5_ASAP7_75t_SL g341 ( .A1(n_342), .A2(n_344), .B(n_345), .Y(n_341) );
INVxp67_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
OAI21xp5_ASAP7_75t_SL g345 ( .A1(n_346), .A2(n_348), .B(n_351), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_346), .B(n_375), .Y(n_374) );
INVxp67_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_351), .B(n_438), .Y(n_437) );
OAI21xp33_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_356), .B(n_358), .Y(n_352) );
INVx1_ASAP7_75t_SL g353 ( .A(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g379 ( .A(n_355), .B(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
AND4x1_ASAP7_75t_L g364 ( .A(n_365), .B(n_395), .C(n_412), .D(n_434), .Y(n_364) );
NOR2xp33_ASAP7_75t_L g365 ( .A(n_366), .B(n_382), .Y(n_365) );
OAI211xp5_ASAP7_75t_SL g366 ( .A1(n_367), .A2(n_371), .B(n_374), .C(n_376), .Y(n_366) );
OR2x2_ASAP7_75t_L g367 ( .A(n_368), .B(n_369), .Y(n_367) );
INVx1_ASAP7_75t_SL g369 ( .A(n_370), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_370), .B(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
NOR2xp33_ASAP7_75t_L g403 ( .A(n_381), .B(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
NOR2xp33_ASAP7_75t_L g390 ( .A(n_391), .B(n_393), .Y(n_390) );
INVx1_ASAP7_75t_L g416 ( .A(n_391), .Y(n_416) );
INVx2_ASAP7_75t_SL g404 ( .A(n_392), .Y(n_404) );
OR2x2_ASAP7_75t_L g397 ( .A(n_398), .B(n_399), .Y(n_397) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g417 ( .A(n_402), .Y(n_417) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
NOR2xp33_ASAP7_75t_SL g412 ( .A(n_413), .B(n_420), .Y(n_412) );
INVx1_ASAP7_75t_SL g414 ( .A(n_415), .Y(n_414) );
OAI221xp5_ASAP7_75t_SL g420 ( .A1(n_421), .A2(n_422), .B1(n_424), .B2(n_425), .C(n_426), .Y(n_420) );
AOI22xp5_ASAP7_75t_L g426 ( .A1(n_427), .A2(n_431), .B1(n_432), .B2(n_433), .Y(n_426) );
NAND2xp5_ASAP7_75t_SL g427 ( .A(n_428), .B(n_429), .Y(n_427) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx2_ASAP7_75t_L g734 ( .A(n_443), .Y(n_734) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g735 ( .A(n_445), .Y(n_735) );
OR3x1_ASAP7_75t_L g445 ( .A(n_446), .B(n_627), .C(n_692), .Y(n_445) );
NAND4xp25_ASAP7_75t_SL g446 ( .A(n_447), .B(n_568), .C(n_594), .D(n_617), .Y(n_446) );
AOI221xp5_ASAP7_75t_L g447 ( .A1(n_448), .A2(n_500), .B1(n_538), .B2(n_545), .C(n_560), .Y(n_447) );
CKINVDCx14_ASAP7_75t_R g448 ( .A(n_449), .Y(n_448) );
OAI22xp5_ASAP7_75t_L g715 ( .A1(n_449), .A2(n_561), .B1(n_585), .B2(n_716), .Y(n_715) );
OR2x2_ASAP7_75t_L g449 ( .A(n_450), .B(n_481), .Y(n_449) );
INVx1_ASAP7_75t_SL g621 ( .A(n_450), .Y(n_621) );
OR2x2_ASAP7_75t_L g450 ( .A(n_451), .B(n_465), .Y(n_450) );
OR2x2_ASAP7_75t_L g543 ( .A(n_451), .B(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_L g563 ( .A(n_451), .B(n_482), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_451), .B(n_490), .Y(n_576) );
AND2x2_ASAP7_75t_L g593 ( .A(n_451), .B(n_465), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_451), .B(n_541), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_451), .B(n_592), .Y(n_704) );
NOR2xp33_ASAP7_75t_L g714 ( .A(n_451), .B(n_481), .Y(n_714) );
AOI211xp5_ASAP7_75t_SL g725 ( .A1(n_451), .A2(n_631), .B(n_726), .C(n_727), .Y(n_725) );
INVx5_ASAP7_75t_SL g451 ( .A(n_452), .Y(n_451) );
NAND2xp5_ASAP7_75t_SL g597 ( .A(n_452), .B(n_482), .Y(n_597) );
AND2x2_ASAP7_75t_L g600 ( .A(n_452), .B(n_483), .Y(n_600) );
OR2x2_ASAP7_75t_L g645 ( .A(n_452), .B(n_482), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_452), .B(n_490), .Y(n_654) );
OAI21xp5_ASAP7_75t_L g453 ( .A1(n_454), .A2(n_455), .B(n_457), .Y(n_453) );
INVx5_ASAP7_75t_L g471 ( .A(n_458), .Y(n_471) );
INVx5_ASAP7_75t_SL g544 ( .A(n_465), .Y(n_544) );
AND2x2_ASAP7_75t_L g562 ( .A(n_465), .B(n_563), .Y(n_562) );
NOR2xp33_ASAP7_75t_L g644 ( .A(n_465), .B(n_645), .Y(n_644) );
AND2x2_ASAP7_75t_L g648 ( .A(n_465), .B(n_649), .Y(n_648) );
AND2x2_ASAP7_75t_L g680 ( .A(n_465), .B(n_490), .Y(n_680) );
OR2x2_ASAP7_75t_L g686 ( .A(n_465), .B(n_576), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_465), .B(n_636), .Y(n_695) );
OR2x6_ASAP7_75t_L g465 ( .A(n_466), .B(n_480), .Y(n_465) );
BUFx2_ASAP7_75t_L g517 ( .A(n_468), .Y(n_517) );
INVx2_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
O2A1O1Ixp33_ASAP7_75t_L g493 ( .A1(n_471), .A2(n_479), .B(n_494), .C(n_495), .Y(n_493) );
O2A1O1Ixp33_ASAP7_75t_SL g552 ( .A1(n_471), .A2(n_479), .B(n_553), .C(n_554), .Y(n_552) );
O2A1O1Ixp33_ASAP7_75t_L g472 ( .A1(n_473), .A2(n_474), .B(n_476), .C(n_477), .Y(n_472) );
O2A1O1Ixp33_ASAP7_75t_L g507 ( .A1(n_474), .A2(n_477), .B(n_508), .C(n_509), .Y(n_507) );
INVx2_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_482), .B(n_490), .Y(n_481) );
AND2x2_ASAP7_75t_L g577 ( .A(n_482), .B(n_544), .Y(n_577) );
INVx1_ASAP7_75t_SL g590 ( .A(n_482), .Y(n_590) );
OR2x2_ASAP7_75t_L g625 ( .A(n_482), .B(n_626), .Y(n_625) );
OR2x2_ASAP7_75t_L g631 ( .A(n_482), .B(n_490), .Y(n_631) );
AND2x2_ASAP7_75t_L g689 ( .A(n_482), .B(n_541), .Y(n_689) );
INVx2_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_483), .B(n_544), .Y(n_616) );
INVx3_ASAP7_75t_L g541 ( .A(n_490), .Y(n_541) );
OR2x2_ASAP7_75t_L g582 ( .A(n_490), .B(n_544), .Y(n_582) );
AND2x2_ASAP7_75t_L g592 ( .A(n_490), .B(n_590), .Y(n_592) );
HB1xp67_ASAP7_75t_L g640 ( .A(n_490), .Y(n_640) );
AND2x2_ASAP7_75t_L g649 ( .A(n_490), .B(n_563), .Y(n_649) );
OA21x2_ASAP7_75t_L g490 ( .A1(n_491), .A2(n_492), .B(n_498), .Y(n_490) );
OA21x2_ASAP7_75t_L g550 ( .A1(n_499), .A2(n_551), .B(n_559), .Y(n_550) );
AOI221xp5_ASAP7_75t_L g665 ( .A1(n_500), .A2(n_666), .B1(n_668), .B2(n_670), .C(n_673), .Y(n_665) );
INVx2_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
OR2x2_ASAP7_75t_L g501 ( .A(n_502), .B(n_512), .Y(n_501) );
AND2x2_ASAP7_75t_L g639 ( .A(n_502), .B(n_620), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_502), .B(n_698), .Y(n_702) );
OR2x2_ASAP7_75t_L g723 ( .A(n_502), .B(n_724), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_502), .B(n_728), .Y(n_727) );
BUFx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx5_ASAP7_75t_L g570 ( .A(n_503), .Y(n_570) );
AND2x2_ASAP7_75t_L g647 ( .A(n_503), .B(n_514), .Y(n_647) );
AND2x2_ASAP7_75t_L g708 ( .A(n_503), .B(n_587), .Y(n_708) );
AND2x2_ASAP7_75t_L g721 ( .A(n_503), .B(n_541), .Y(n_721) );
OR2x6_ASAP7_75t_L g503 ( .A(n_504), .B(n_510), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_513), .B(n_526), .Y(n_512) );
AND2x4_ASAP7_75t_L g548 ( .A(n_513), .B(n_549), .Y(n_548) );
AND2x2_ASAP7_75t_L g566 ( .A(n_513), .B(n_567), .Y(n_566) );
INVx2_ASAP7_75t_L g573 ( .A(n_513), .Y(n_573) );
AND2x2_ASAP7_75t_L g642 ( .A(n_513), .B(n_620), .Y(n_642) );
AND2x2_ASAP7_75t_L g652 ( .A(n_513), .B(n_570), .Y(n_652) );
HB1xp67_ASAP7_75t_L g660 ( .A(n_513), .Y(n_660) );
AND2x2_ASAP7_75t_L g672 ( .A(n_513), .B(n_550), .Y(n_672) );
NOR2xp33_ASAP7_75t_L g676 ( .A(n_513), .B(n_604), .Y(n_676) );
AND2x2_ASAP7_75t_L g713 ( .A(n_513), .B(n_708), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_513), .B(n_587), .Y(n_724) );
OR2x2_ASAP7_75t_L g726 ( .A(n_513), .B(n_662), .Y(n_726) );
INVx5_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
AND2x2_ASAP7_75t_L g612 ( .A(n_514), .B(n_613), .Y(n_612) );
AND2x2_ASAP7_75t_L g622 ( .A(n_514), .B(n_567), .Y(n_622) );
AND2x2_ASAP7_75t_L g634 ( .A(n_514), .B(n_550), .Y(n_634) );
HB1xp67_ASAP7_75t_L g664 ( .A(n_514), .Y(n_664) );
AND2x4_ASAP7_75t_L g698 ( .A(n_514), .B(n_549), .Y(n_698) );
OR2x6_ASAP7_75t_L g514 ( .A(n_515), .B(n_523), .Y(n_514) );
AOI21xp5_ASAP7_75t_SL g515 ( .A1(n_516), .A2(n_518), .B(n_522), .Y(n_515) );
NOR2xp33_ASAP7_75t_L g523 ( .A(n_524), .B(n_525), .Y(n_523) );
BUFx2_ASAP7_75t_L g547 ( .A(n_526), .Y(n_547) );
HB1xp67_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx2_ASAP7_75t_L g587 ( .A(n_527), .Y(n_587) );
AND2x2_ASAP7_75t_L g620 ( .A(n_527), .B(n_550), .Y(n_620) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
AND2x2_ASAP7_75t_L g567 ( .A(n_528), .B(n_550), .Y(n_567) );
BUFx2_ASAP7_75t_L g613 ( .A(n_528), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_530), .B(n_535), .Y(n_529) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_540), .B(n_542), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_540), .B(n_621), .Y(n_700) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_541), .B(n_563), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_541), .B(n_544), .Y(n_602) );
AND2x2_ASAP7_75t_L g657 ( .A(n_541), .B(n_593), .Y(n_657) );
AOI221xp5_ASAP7_75t_SL g594 ( .A1(n_542), .A2(n_595), .B1(n_603), .B2(n_605), .C(n_609), .Y(n_594) );
INVx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
OR2x2_ASAP7_75t_L g589 ( .A(n_543), .B(n_590), .Y(n_589) );
OR2x2_ASAP7_75t_L g630 ( .A(n_543), .B(n_631), .Y(n_630) );
OAI321xp33_ASAP7_75t_L g637 ( .A1(n_543), .A2(n_596), .A3(n_638), .B1(n_640), .B2(n_641), .C(n_643), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_544), .B(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_547), .B(n_548), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_547), .B(n_698), .Y(n_716) );
AND2x2_ASAP7_75t_L g603 ( .A(n_548), .B(n_604), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_548), .B(n_607), .Y(n_606) );
HB1xp67_ASAP7_75t_L g579 ( .A(n_549), .Y(n_579) );
AND2x2_ASAP7_75t_L g586 ( .A(n_549), .B(n_587), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_549), .B(n_661), .Y(n_691) );
INVx1_ASAP7_75t_L g728 ( .A(n_549), .Y(n_728) );
INVx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
NOR2xp33_ASAP7_75t_L g555 ( .A(n_556), .B(n_557), .Y(n_555) );
AOI21xp5_ASAP7_75t_L g560 ( .A1(n_561), .A2(n_564), .B(n_565), .Y(n_560) );
INVx1_ASAP7_75t_SL g561 ( .A(n_562), .Y(n_561) );
A2O1A1Ixp33_ASAP7_75t_L g720 ( .A1(n_562), .A2(n_672), .B(n_721), .C(n_722), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_563), .B(n_581), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_563), .B(n_601), .Y(n_667) );
INVx1_ASAP7_75t_SL g565 ( .A(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g610 ( .A(n_567), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_567), .B(n_570), .Y(n_624) );
NOR2xp33_ASAP7_75t_L g633 ( .A(n_567), .B(n_634), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_567), .B(n_652), .Y(n_651) );
AOI22xp33_ASAP7_75t_L g568 ( .A1(n_569), .A2(n_571), .B1(n_583), .B2(n_588), .Y(n_568) );
HB1xp67_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
OR2x2_ASAP7_75t_L g584 ( .A(n_570), .B(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_L g607 ( .A(n_570), .B(n_608), .Y(n_607) );
AND2x2_ASAP7_75t_L g619 ( .A(n_570), .B(n_620), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_570), .B(n_613), .Y(n_655) );
OR2x2_ASAP7_75t_L g662 ( .A(n_570), .B(n_587), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_570), .B(n_672), .Y(n_671) );
AND2x2_ASAP7_75t_L g712 ( .A(n_570), .B(n_698), .Y(n_712) );
OAI22xp33_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_574), .B1(n_578), .B2(n_580), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g618 ( .A(n_573), .B(n_619), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_575), .B(n_577), .Y(n_574) );
INVx1_ASAP7_75t_SL g575 ( .A(n_576), .Y(n_575) );
OAI22xp33_ASAP7_75t_L g658 ( .A1(n_576), .A2(n_591), .B1(n_659), .B2(n_663), .Y(n_658) );
INVx1_ASAP7_75t_L g706 ( .A(n_577), .Y(n_706) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
AOI221xp5_ASAP7_75t_L g617 ( .A1(n_581), .A2(n_618), .B1(n_621), .B2(n_622), .C(n_623), .Y(n_617) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
OR2x2_ASAP7_75t_L g596 ( .A(n_582), .B(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_586), .B(n_652), .Y(n_684) );
HB1xp67_ASAP7_75t_L g604 ( .A(n_587), .Y(n_604) );
INVx1_ASAP7_75t_L g608 ( .A(n_587), .Y(n_608) );
NAND2xp33_ASAP7_75t_L g588 ( .A(n_589), .B(n_591), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .Y(n_591) );
INVx1_ASAP7_75t_L g626 ( .A(n_593), .Y(n_626) );
AND2x2_ASAP7_75t_L g635 ( .A(n_593), .B(n_636), .Y(n_635) );
NAND2xp33_ASAP7_75t_L g595 ( .A(n_596), .B(n_598), .Y(n_595) );
INVx2_ASAP7_75t_SL g598 ( .A(n_599), .Y(n_598) );
AND2x4_ASAP7_75t_L g599 ( .A(n_600), .B(n_601), .Y(n_599) );
AND2x2_ASAP7_75t_L g679 ( .A(n_600), .B(n_680), .Y(n_679) );
INVx2_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
AOI221xp5_ASAP7_75t_L g628 ( .A1(n_603), .A2(n_629), .B1(n_632), .B2(n_635), .C(n_637), .Y(n_628) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_607), .B(n_664), .Y(n_663) );
AOI21xp33_ASAP7_75t_SL g609 ( .A1(n_610), .A2(n_611), .B(n_614), .Y(n_609) );
INVx2_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
CKINVDCx16_ASAP7_75t_R g711 ( .A(n_614), .Y(n_711) );
OR2x2_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
OR2x2_ASAP7_75t_L g653 ( .A(n_616), .B(n_654), .Y(n_653) );
INVx1_ASAP7_75t_SL g674 ( .A(n_619), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_619), .B(n_679), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_622), .B(n_644), .Y(n_643) );
NOR2xp33_ASAP7_75t_L g623 ( .A(n_624), .B(n_625), .Y(n_623) );
NAND4xp25_ASAP7_75t_L g627 ( .A(n_628), .B(n_646), .C(n_665), .D(n_678), .Y(n_627) );
INVx1_ASAP7_75t_SL g629 ( .A(n_630), .Y(n_629) );
INVx1_ASAP7_75t_SL g636 ( .A(n_631), .Y(n_636) );
INVxp67_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
OR2x2_ASAP7_75t_L g669 ( .A(n_640), .B(n_645), .Y(n_669) );
INVxp67_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
AOI211xp5_ASAP7_75t_L g646 ( .A1(n_647), .A2(n_648), .B(n_650), .C(n_658), .Y(n_646) );
AOI211xp5_ASAP7_75t_L g717 ( .A1(n_648), .A2(n_690), .B(n_718), .C(n_725), .Y(n_717) );
INVx1_ASAP7_75t_SL g677 ( .A(n_649), .Y(n_677) );
OAI22xp5_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_653), .B1(n_655), .B2(n_656), .Y(n_650) );
INVx1_ASAP7_75t_L g681 ( .A(n_655), .Y(n_681) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_660), .B(n_661), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_661), .B(n_698), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_661), .B(n_672), .Y(n_705) );
INVx2_ASAP7_75t_SL g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_SL g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g682 ( .A(n_672), .Y(n_682) );
AOI21xp33_ASAP7_75t_L g673 ( .A1(n_674), .A2(n_675), .B(n_677), .Y(n_673) );
INVxp33_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
AOI322xp5_ASAP7_75t_L g678 ( .A1(n_679), .A2(n_681), .A3(n_682), .B1(n_683), .B2(n_685), .C1(n_687), .C2(n_690), .Y(n_678) );
INVxp67_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
NAND3xp33_ASAP7_75t_SL g692 ( .A(n_693), .B(n_710), .C(n_717), .Y(n_692) );
AOI221xp5_ASAP7_75t_L g693 ( .A1(n_694), .A2(n_696), .B1(n_699), .B2(n_701), .C(n_703), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_SL g709 ( .A(n_698), .Y(n_709) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVxp67_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
OAI22xp33_ASAP7_75t_L g703 ( .A1(n_704), .A2(n_705), .B1(n_706), .B2(n_707), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_708), .B(n_709), .Y(n_707) );
AOI221xp5_ASAP7_75t_L g710 ( .A1(n_711), .A2(n_712), .B1(n_713), .B2(n_714), .C(n_715), .Y(n_710) );
NAND2xp33_ASAP7_75t_L g718 ( .A(n_719), .B(n_720), .Y(n_718) );
INVxp67_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx2_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx2_ASAP7_75t_L g736 ( .A(n_730), .Y(n_736) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_SL g737 ( .A(n_738), .Y(n_737) );
INVx3_ASAP7_75t_SL g738 ( .A(n_739), .Y(n_738) );
INVxp67_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
HB1xp67_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_SL g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
endmodule