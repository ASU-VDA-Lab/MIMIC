module real_jpeg_16660_n_13 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_13);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_13;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI21xp5_ASAP7_75t_L g13 ( 
.A1(n_0),
.A2(n_14),
.B(n_345),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_0),
.B(n_346),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_1),
.Y(n_56)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_1),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_1),
.Y(n_69)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_1),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_2),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_2),
.Y(n_123)
);

BUFx5_ASAP7_75t_L g130 ( 
.A(n_2),
.Y(n_130)
);

BUFx5_ASAP7_75t_L g268 ( 
.A(n_2),
.Y(n_268)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_3),
.Y(n_90)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_3),
.Y(n_103)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_4),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_4),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_4),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_4),
.Y(n_132)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_4),
.Y(n_198)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_4),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_5),
.A2(n_105),
.B1(n_108),
.B2(n_109),
.Y(n_104)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_5),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_5),
.A2(n_108),
.B1(n_196),
.B2(n_199),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_6),
.Y(n_163)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_7),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_8),
.A2(n_141),
.B1(n_145),
.B2(n_146),
.Y(n_140)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_8),
.Y(n_145)
);

OAI22xp33_ASAP7_75t_SL g337 ( 
.A1(n_8),
.A2(n_145),
.B1(n_338),
.B2(n_339),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_10),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_10),
.Y(n_99)
);

BUFx4f_ASAP7_75t_L g107 ( 
.A(n_10),
.Y(n_107)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_10),
.Y(n_125)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_11),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_11),
.A2(n_26),
.B1(n_92),
.B2(n_95),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_11),
.A2(n_26),
.B1(n_113),
.B2(n_115),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_11),
.B(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_11),
.B(n_52),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_11),
.B(n_266),
.C(n_269),
.Y(n_265)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_12),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_323),
.Y(n_14)
);

AO21x1_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_207),
.B(n_321),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_185),
.Y(n_18)
);

OR2x2_ASAP7_75t_L g322 ( 
.A(n_19),
.B(n_185),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_134),
.C(n_149),
.Y(n_19)
);

HB1xp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_21),
.B(n_134),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_80),
.B2(n_133),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

OAI22x1_ASAP7_75t_L g203 ( 
.A1(n_23),
.A2(n_204),
.B1(n_205),
.B2(n_206),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_23),
.Y(n_204)
);

XNOR2x1_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_51),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_24),
.B(n_51),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_24),
.B(n_51),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_24),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_24),
.B(n_111),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_24),
.Y(n_333)
);

AND2x4_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_33),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B(n_30),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_26),
.B(n_31),
.Y(n_30)
);

OAI21xp33_ASAP7_75t_L g73 ( 
.A1(n_26),
.A2(n_74),
.B(n_76),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_26),
.B(n_77),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_26),
.B(n_119),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_26),
.B(n_284),
.Y(n_283)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_29),
.A2(n_45),
.B1(n_46),
.B2(n_49),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_30),
.Y(n_176)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_35),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_44),
.Y(n_34)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_35),
.Y(n_216)
);

OA22x2_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_38),
.Y(n_175)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_43),
.Y(n_157)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_47),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g214 ( 
.A(n_51),
.Y(n_214)
);

BUFx2_ASAP7_75t_L g223 ( 
.A(n_51),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_51),
.B(n_111),
.Y(n_255)
);

OA21x2_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_62),
.B(n_73),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_63),
.Y(n_62)
);

OA22x2_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_57),
.B1(n_59),
.B2(n_61),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_56),
.Y(n_61)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_57),
.Y(n_114)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_58),
.Y(n_117)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_67),
.B1(n_68),
.B2(n_70),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_72),
.Y(n_75)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

OAI32xp33_ASAP7_75t_L g231 ( 
.A1(n_76),
.A2(n_232),
.A3(n_234),
.B1(n_237),
.B2(n_243),
.Y(n_231)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_80),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_80),
.A2(n_181),
.B(n_182),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_111),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_81),
.A2(n_111),
.B1(n_147),
.B2(n_306),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_81),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_91),
.B1(n_100),
.B2(n_104),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_82),
.A2(n_104),
.B1(n_136),
.B2(n_139),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_87),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_86),
.Y(n_94)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_86),
.Y(n_110)
);

OA22x2_ASAP7_75t_L g119 ( 
.A1(n_86),
.A2(n_120),
.B1(n_122),
.B2(n_124),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_86),
.Y(n_269)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g178 ( 
.A(n_91),
.B(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_93),
.B(n_180),
.Y(n_179)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_98),
.Y(n_282)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_101),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_101),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_103),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_107),
.Y(n_144)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_109),
.Y(n_146)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_111),
.A2(n_135),
.B1(n_147),
.B2(n_148),
.Y(n_134)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_111),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_111),
.B(n_135),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_111),
.A2(n_147),
.B1(n_214),
.B2(n_223),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_111),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_111),
.A2(n_147),
.B1(n_229),
.B2(n_230),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_111),
.A2(n_147),
.B1(n_261),
.B2(n_262),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_111),
.A2(n_147),
.B1(n_264),
.B2(n_289),
.Y(n_288)
);

AND2x4_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_118),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_112),
.A2(n_193),
.B1(n_194),
.B2(n_195),
.Y(n_192)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_114),
.Y(n_338)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_126),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_119),
.B(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_119),
.Y(n_194)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_123),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_126),
.Y(n_193)
);

OAI22xp33_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_130),
.B1(n_131),
.B2(n_132),
.Y(n_127)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_128),
.Y(n_340)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_129),
.Y(n_236)
);

BUFx12f_ASAP7_75t_L g246 ( 
.A(n_129),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_135),
.Y(n_148)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_140),
.B(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

A2O1A1Ixp33_ASAP7_75t_L g252 ( 
.A1(n_147),
.A2(n_214),
.B(n_253),
.C(n_255),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_147),
.B(n_264),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_147),
.B(n_217),
.C(n_262),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_149),
.B(n_314),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_181),
.B(n_182),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_150),
.B(n_204),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_177),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_151),
.A2(n_177),
.B1(n_217),
.B2(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_151),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_158),
.B(n_168),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

HB1xp67_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_157),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_159),
.B(n_164),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx8_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_171),
.B(n_176),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_177),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_177),
.A2(n_178),
.B1(n_215),
.B2(n_227),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_177),
.B(n_231),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_177),
.B(n_275),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_177),
.B(n_277),
.Y(n_276)
);

AND2x2_ASAP7_75t_SL g287 ( 
.A(n_177),
.B(n_288),
.Y(n_287)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_179),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_181),
.A2(n_182),
.B(n_205),
.Y(n_327)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

AND3x1_ASAP7_75t_L g308 ( 
.A(n_184),
.B(n_255),
.C(n_309),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_186),
.B(n_188),
.C(n_203),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_203),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_191),
.B1(n_192),
.B2(n_202),
.Y(n_188)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_189),
.Y(n_202)
);

NOR2xp67_ASAP7_75t_R g331 ( 
.A(n_189),
.B(n_192),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_189),
.A2(n_202),
.B1(n_221),
.B2(n_333),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_193),
.A2(n_194),
.B1(n_195),
.B2(n_337),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_205),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_298),
.B(n_315),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

AO21x2_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_248),
.B(n_297),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_211),
.B(n_224),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_211),
.B(n_224),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_220),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_218),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_213),
.B(n_218),
.C(n_220),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.C(n_217),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_214),
.A2(n_223),
.B1(n_226),
.B2(n_228),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_214),
.A2(n_336),
.B(n_341),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_214),
.B(n_336),
.Y(n_341)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_215),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_217),
.B(n_231),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_217),
.B(n_260),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_222),
.A2(n_253),
.B1(n_254),
.B2(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_222),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_229),
.C(n_247),
.Y(n_224)
);

XOR2x2_ASAP7_75t_SL g250 ( 
.A(n_225),
.B(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_226),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g244 ( 
.A(n_239),
.Y(n_244)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_246),
.Y(n_271)
);

OAI21x1_ASAP7_75t_SL g248 ( 
.A1(n_249),
.A2(n_256),
.B(n_296),
.Y(n_248)
);

NOR2xp67_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_252),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_250),
.B(n_252),
.Y(n_296)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

AOI21x1_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_291),
.B(n_295),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_258),
.A2(n_272),
.B(n_290),
.Y(n_257)
);

NOR2x1_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_263),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_259),
.B(n_263),
.Y(n_290)
);

INVxp67_ASAP7_75t_SL g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_264),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_265),
.B(n_270),
.Y(n_264)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

NOR2x1_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_287),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_276),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_283),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

OR2x2_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_292),
.B(n_293),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_311),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_301),
.B(n_310),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_301),
.B(n_310),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_SL g301 ( 
.A(n_302),
.B(n_303),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_302),
.B(n_305),
.C(n_307),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_304),
.A2(n_305),
.B1(n_307),
.B2(n_308),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g316 ( 
.A(n_311),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_313),
.Y(n_311)
);

OR2x2_ASAP7_75t_L g320 ( 
.A(n_312),
.B(n_313),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_316),
.A2(n_317),
.B(n_319),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_342),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_326),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_325),
.B(n_326),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_329),
.A2(n_330),
.B1(n_334),
.B2(n_335),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_332),
.Y(n_330)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVxp33_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

HB1xp67_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);


endmodule