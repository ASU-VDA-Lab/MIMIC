module fake_jpeg_12768_n_141 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_141);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_141;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx4_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_39),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_24),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_41),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_42),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_9),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_0),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_0),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

CKINVDCx11_ASAP7_75t_R g59 ( 
.A(n_44),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_7),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_17),
.B(n_6),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_14),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_11),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_45),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_10),
.B(n_43),
.Y(n_65)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_1),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_68),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_61),
.B(n_20),
.C(n_40),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_70),
.Y(n_78)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_71),
.Y(n_75)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_77),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_63),
.Y(n_79)
);

INVx6_ASAP7_75t_SL g81 ( 
.A(n_70),
.Y(n_81)
);

INVx13_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_46),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_82),
.B(n_1),
.Y(n_101)
);

AND2x2_ASAP7_75t_SL g83 ( 
.A(n_68),
.B(n_51),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_49),
.C(n_48),
.Y(n_97)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_82),
.A2(n_55),
.B1(n_60),
.B2(n_57),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_86),
.A2(n_90),
.B1(n_96),
.B2(n_102),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_79),
.A2(n_57),
.B(n_51),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_87),
.A2(n_8),
.B(n_10),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_88),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_80),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_89),
.B(n_94),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_75),
.A2(n_55),
.B1(n_60),
.B2(n_47),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_81),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_92),
.B(n_8),
.Y(n_114)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_95),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_76),
.A2(n_65),
.B(n_64),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_62),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_84),
.A2(n_47),
.B1(n_53),
.B2(n_52),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_97),
.B(n_100),
.C(n_4),
.Y(n_105)
);

BUFx12_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_98),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_59),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_101),
.B(n_5),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_75),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_105),
.B(n_114),
.C(n_115),
.Y(n_122)
);

AND2x6_ASAP7_75t_L g106 ( 
.A(n_98),
.B(n_25),
.Y(n_106)
);

AND2x6_ASAP7_75t_L g119 ( 
.A(n_106),
.B(n_18),
.Y(n_119)
);

OAI21xp33_ASAP7_75t_L g107 ( 
.A1(n_99),
.A2(n_85),
.B(n_23),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_107),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_90),
.A2(n_85),
.B1(n_6),
.B2(n_7),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_108),
.A2(n_19),
.B1(n_22),
.B2(n_26),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_110),
.B(n_111),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_98),
.B(n_5),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_112),
.A2(n_88),
.B1(n_89),
.B2(n_93),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_91),
.B(n_12),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_13),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_116),
.B(n_118),
.C(n_32),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_SL g118 ( 
.A(n_89),
.B(n_15),
.C(n_16),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_119),
.A2(n_124),
.B(n_107),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_121),
.A2(n_126),
.B1(n_106),
.B2(n_38),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_123),
.A2(n_128),
.B1(n_113),
.B2(n_103),
.Y(n_131)
);

FAx1_ASAP7_75t_L g124 ( 
.A(n_112),
.B(n_28),
.CI(n_29),
.CON(n_124),
.SN(n_124)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_117),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_127),
.B(n_118),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_104),
.A2(n_34),
.B1(n_35),
.B2(n_37),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_129),
.A2(n_131),
.B1(n_133),
.B2(n_125),
.Y(n_134)
);

MAJx2_ASAP7_75t_L g130 ( 
.A(n_122),
.B(n_105),
.C(n_109),
.Y(n_130)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_130),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_132),
.Y(n_136)
);

OAI21x1_ASAP7_75t_L g137 ( 
.A1(n_134),
.A2(n_125),
.B(n_124),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_137),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_138),
.A2(n_135),
.B1(n_136),
.B2(n_131),
.Y(n_139)
);

AOI21xp33_ASAP7_75t_SL g140 ( 
.A1(n_139),
.A2(n_124),
.B(n_135),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_120),
.Y(n_141)
);


endmodule