module fake_jpeg_18305_n_110 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_110);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_110;

wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx3_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_8),
.B(n_5),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

BUFx2_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_8),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_19),
.B(n_20),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_13),
.B(n_0),
.Y(n_20)
);

INVx4_ASAP7_75t_SL g21 ( 
.A(n_12),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_21),
.B(n_22),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_24),
.B(n_25),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_21),
.A2(n_17),
.B1(n_18),
.B2(n_16),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_27),
.A2(n_11),
.B1(n_14),
.B2(n_15),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_20),
.A2(n_17),
.B1(n_10),
.B2(n_11),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_28),
.A2(n_30),
.B1(n_10),
.B2(n_18),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g30 ( 
.A1(n_21),
.A2(n_17),
.B1(n_12),
.B2(n_10),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_27),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_33),
.B(n_34),
.Y(n_47)
);

AND2x6_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_20),
.Y(n_34)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_36),
.A2(n_41),
.B1(n_15),
.B2(n_26),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_25),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_32),
.C(n_19),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_16),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_39),
.Y(n_45)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_14),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_40),
.B(n_42),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_28),
.B(n_25),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_33),
.A2(n_26),
.B1(n_31),
.B2(n_29),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_43),
.A2(n_49),
.B1(n_36),
.B2(n_26),
.Y(n_59)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_39),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_37),
.C(n_32),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_34),
.B(n_30),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_SL g57 ( 
.A1(n_50),
.A2(n_52),
.B(n_44),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_35),
.B(n_32),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_SL g53 ( 
.A1(n_47),
.A2(n_42),
.B(n_37),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_53),
.A2(n_63),
.B(n_12),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_54),
.A2(n_25),
.B1(n_24),
.B2(n_22),
.Y(n_71)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_52),
.Y(n_55)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_58),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_59),
.A2(n_61),
.B1(n_45),
.B2(n_48),
.Y(n_67)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_60),
.B(n_46),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_49),
.A2(n_39),
.B1(n_26),
.B2(n_23),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

NOR3xp33_ASAP7_75t_L g75 ( 
.A(n_62),
.B(n_61),
.C(n_59),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_50),
.A2(n_0),
.B(n_1),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_63),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_64),
.B(n_69),
.Y(n_85)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_67),
.A2(n_72),
.B1(n_75),
.B2(n_19),
.Y(n_78)
);

AOI322xp5_ASAP7_75t_SL g69 ( 
.A1(n_53),
.A2(n_44),
.A3(n_7),
.B1(n_6),
.B2(n_3),
.C1(n_4),
.C2(n_5),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_74),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_54),
.A2(n_24),
.B1(n_22),
.B2(n_19),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_73),
.A2(n_12),
.B(n_1),
.Y(n_79)
);

MAJx2_ASAP7_75t_L g74 ( 
.A(n_62),
.B(n_24),
.C(n_22),
.Y(n_74)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_78),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_79),
.A2(n_84),
.B(n_72),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

BUFx12_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_81),
.B(n_83),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_68),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_82),
.B(n_71),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_86),
.B(n_88),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_82),
.A2(n_67),
.B(n_74),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_90),
.Y(n_97)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_92),
.Y(n_94)
);

NOR2x1_ASAP7_75t_SL g93 ( 
.A(n_86),
.B(n_81),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_93),
.B(n_95),
.Y(n_99)
);

AOI21xp33_ASAP7_75t_L g95 ( 
.A1(n_87),
.A2(n_85),
.B(n_77),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_94),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_98),
.A2(n_102),
.B(n_76),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_97),
.B(n_80),
.Y(n_100)
);

INVxp33_ASAP7_75t_L g104 ( 
.A(n_100),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_96),
.A2(n_81),
.B1(n_79),
.B2(n_89),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_97),
.B(n_91),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_103),
.Y(n_107)
);

NOR2x1_ASAP7_75t_L g105 ( 
.A(n_99),
.B(n_7),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_101),
.C(n_1),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_106),
.B(n_104),
.C(n_1),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_108),
.B(n_109),
.Y(n_110)
);

AOI221xp5_ASAP7_75t_L g109 ( 
.A1(n_107),
.A2(n_0),
.B1(n_2),
.B2(n_99),
.C(n_98),
.Y(n_109)
);


endmodule