module real_jpeg_16475_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_556;
wire n_507;
wire n_57;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_470;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_548;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_546;
wire n_285;
wire n_531;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_549;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_0),
.A2(n_19),
.B(n_556),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_0),
.B(n_557),
.Y(n_556)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_1),
.Y(n_400)
);

OAI32xp33_ASAP7_75t_L g78 ( 
.A1(n_2),
.A2(n_79),
.A3(n_83),
.B1(n_88),
.B2(n_93),
.Y(n_78)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_2),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_2),
.A2(n_92),
.B1(n_268),
.B2(n_272),
.Y(n_267)
);

OAI32xp33_ASAP7_75t_L g290 ( 
.A1(n_2),
.A2(n_79),
.A3(n_83),
.B1(n_88),
.B2(n_93),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_2),
.B(n_143),
.Y(n_299)
);

OAI32xp33_ASAP7_75t_L g380 ( 
.A1(n_2),
.A2(n_381),
.A3(n_385),
.B1(n_389),
.B2(n_392),
.Y(n_380)
);

AOI22xp33_ASAP7_75t_SL g418 ( 
.A1(n_2),
.A2(n_79),
.B1(n_92),
.B2(n_419),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_2),
.B(n_29),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_2),
.B(n_507),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_2),
.B(n_265),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_3),
.A2(n_56),
.B1(n_62),
.B2(n_63),
.Y(n_55)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_3),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_3),
.A2(n_62),
.B1(n_136),
.B2(n_162),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g410 ( 
.A1(n_3),
.A2(n_62),
.B1(n_411),
.B2(n_414),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_3),
.A2(n_62),
.B1(n_470),
.B2(n_472),
.Y(n_469)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_4),
.Y(n_200)
);

BUFx5_ASAP7_75t_L g202 ( 
.A(n_4),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_4),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_4),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_5),
.A2(n_126),
.B1(n_130),
.B2(n_132),
.Y(n_125)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_5),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g245 ( 
.A1(n_5),
.A2(n_132),
.B1(n_190),
.B2(n_246),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_5),
.A2(n_132),
.B1(n_345),
.B2(n_348),
.Y(n_344)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_6),
.A2(n_113),
.B1(n_118),
.B2(n_121),
.Y(n_112)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_6),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_6),
.A2(n_121),
.B1(n_184),
.B2(n_189),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g321 ( 
.A1(n_6),
.A2(n_121),
.B1(n_322),
.B2(n_324),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_SL g539 ( 
.A1(n_6),
.A2(n_121),
.B1(n_540),
.B2(n_542),
.Y(n_539)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_7),
.Y(n_111)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_7),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g237 ( 
.A(n_7),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_8),
.A2(n_70),
.B1(n_73),
.B2(n_74),
.Y(n_69)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_8),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_8),
.A2(n_73),
.B1(n_130),
.B2(n_239),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_8),
.A2(n_73),
.B1(n_257),
.B2(n_259),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_8),
.A2(n_73),
.B1(n_271),
.B2(n_329),
.Y(n_328)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_9),
.A2(n_136),
.B1(n_138),
.B2(n_139),
.Y(n_135)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_9),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g293 ( 
.A1(n_9),
.A2(n_138),
.B1(n_294),
.B2(n_297),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g458 ( 
.A1(n_9),
.A2(n_138),
.B1(n_459),
.B2(n_464),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_9),
.A2(n_138),
.B1(n_498),
.B2(n_502),
.Y(n_497)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_10),
.Y(n_188)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_10),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_10),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_10),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g263 ( 
.A(n_10),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g447 ( 
.A(n_10),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_11),
.A2(n_114),
.B1(n_177),
.B2(n_178),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_11),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_11),
.A2(n_177),
.B1(n_217),
.B2(n_218),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_11),
.A2(n_177),
.B1(n_228),
.B2(n_230),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_11),
.A2(n_137),
.B1(n_177),
.B2(n_363),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_12),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_12),
.Y(n_145)
);

BUFx5_ASAP7_75t_L g148 ( 
.A(n_12),
.Y(n_148)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_13),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_14),
.Y(n_61)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_15),
.Y(n_107)
);

BUFx4f_ASAP7_75t_L g117 ( 
.A(n_15),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g131 ( 
.A(n_15),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_15),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g159 ( 
.A(n_16),
.Y(n_159)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_17),
.Y(n_87)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_17),
.Y(n_96)
);

BUFx8_ASAP7_75t_L g140 ( 
.A(n_17),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_17),
.Y(n_163)
);

BUFx5_ASAP7_75t_L g364 ( 
.A(n_17),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_528),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_369),
.Y(n_21)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_304),
.B(n_332),
.C(n_333),
.D(n_368),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_251),
.C(n_284),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_24),
.B(n_251),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_165),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_25),
.B(n_166),
.C(n_250),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_77),
.C(n_133),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_26),
.B(n_133),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_54),
.B(n_67),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_27),
.A2(n_29),
.B1(n_343),
.B2(n_344),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g547 ( 
.A1(n_27),
.A2(n_344),
.B(n_548),
.Y(n_547)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI21x1_ASAP7_75t_L g225 ( 
.A1(n_28),
.A2(n_69),
.B(n_226),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_28),
.A2(n_55),
.B1(n_68),
.B2(n_275),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_28),
.A2(n_68),
.B1(n_275),
.B2(n_293),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_28),
.A2(n_68),
.B1(n_320),
.B2(n_321),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_28),
.A2(n_68),
.B1(n_293),
.B2(n_418),
.Y(n_417)
);

OR2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_40),
.Y(n_28)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_29),
.B(n_227),
.Y(n_226)
);

AO22x2_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_34),
.B1(n_37),
.B2(n_38),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_35),
.Y(n_220)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_37),
.Y(n_217)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_44),
.B1(n_49),
.B2(n_52),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g347 ( 
.A(n_46),
.Y(n_347)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_48),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_48),
.Y(n_282)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_59),
.Y(n_323)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_60),
.Y(n_146)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_60),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_69),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_72),
.Y(n_279)
);

INVxp67_ASAP7_75t_SL g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_76),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_77),
.B(n_253),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_101),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_82),
.Y(n_231)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_86),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_87),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_92),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

AO22x2_ASAP7_75t_L g143 ( 
.A1(n_91),
.A2(n_144),
.B1(n_146),
.B2(n_147),
.Y(n_143)
);

INVx2_ASAP7_75t_SL g351 ( 
.A(n_91),
.Y(n_351)
);

HB1xp67_ASAP7_75t_L g395 ( 
.A(n_91),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_SL g389 ( 
.A(n_92),
.B(n_390),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_92),
.B(n_446),
.Y(n_445)
);

OAI21xp33_ASAP7_75t_SL g455 ( 
.A1(n_92),
.A2(n_445),
.B(n_456),
.Y(n_455)
);

AOI22xp33_ASAP7_75t_L g495 ( 
.A1(n_92),
.A2(n_103),
.B1(n_496),
.B2(n_497),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_97),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_100),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_101),
.B(n_290),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_112),
.B1(n_122),
.B2(n_125),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_102),
.A2(n_125),
.B(n_170),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g401 ( 
.A1(n_102),
.A2(n_170),
.B(n_402),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_102),
.A2(n_122),
.B1(n_483),
.B2(n_490),
.Y(n_482)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_103),
.B(n_176),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_103),
.A2(n_238),
.B(n_310),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g468 ( 
.A1(n_103),
.A2(n_469),
.B(n_476),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_103),
.A2(n_484),
.B1(n_497),
.B2(n_510),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_108),
.Y(n_103)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g471 ( 
.A(n_105),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_106),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_107),
.Y(n_120)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_108),
.Y(n_496)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx4_ASAP7_75t_L g507 ( 
.A(n_110),
.Y(n_507)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_112),
.A2(n_241),
.B(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_117),
.Y(n_487)
);

INVx3_ASAP7_75t_L g501 ( 
.A(n_117),
.Y(n_501)
);

BUFx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_119),
.Y(n_502)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_120),
.Y(n_452)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_120),
.Y(n_475)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_124),
.Y(n_175)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_129),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_131),
.Y(n_180)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_131),
.Y(n_201)
);

INVx4_ASAP7_75t_L g505 ( 
.A(n_131),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_141),
.B1(n_143),
.B2(n_156),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_135),
.A2(n_142),
.B1(n_223),
.B2(n_267),
.Y(n_266)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_139),
.Y(n_158)
);

BUFx12f_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_140),
.Y(n_153)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_140),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_141),
.B(n_362),
.Y(n_543)
);

INVx1_ASAP7_75t_SL g141 ( 
.A(n_142),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_142),
.A2(n_157),
.B1(n_223),
.B2(n_224),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_142),
.A2(n_224),
.B(n_327),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g359 ( 
.A1(n_142),
.A2(n_360),
.B(n_361),
.Y(n_359)
);

OR2x6_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_149),
.Y(n_142)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_143),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_143),
.B(n_328),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_143),
.B(n_362),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_145),
.Y(n_155)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_150),
.A2(n_151),
.B1(n_153),
.B2(n_154),
.Y(n_149)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_151),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_151),
.Y(n_541)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_158),
.A2(n_159),
.B1(n_160),
.B2(n_164),
.Y(n_157)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_159),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_159),
.A2(n_164),
.B1(n_276),
.B2(n_280),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_159),
.A2(n_164),
.B1(n_406),
.B2(n_408),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_159),
.A2(n_164),
.B1(n_485),
.B2(n_488),
.Y(n_484)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_163),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_167),
.B1(n_232),
.B2(n_250),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_221),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_168),
.B(n_222),
.C(n_225),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_181),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_169),
.B(n_181),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_176),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx4_ASAP7_75t_SL g301 ( 
.A(n_174),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_175),
.Y(n_313)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_203),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_183),
.B(n_193),
.Y(n_182)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_183),
.Y(n_243)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_187),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_187),
.Y(n_466)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_188),
.Y(n_192)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_188),
.Y(n_463)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_193),
.A2(n_204),
.B1(n_455),
.B2(n_458),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_193),
.A2(n_204),
.B1(n_405),
.B2(n_458),
.Y(n_478)
);

OAI21xp5_ASAP7_75t_L g545 ( 
.A1(n_193),
.A2(n_204),
.B(n_546),
.Y(n_545)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_194),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_194),
.A2(n_243),
.B1(n_244),
.B2(n_245),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_194),
.B(n_256),
.Y(n_353)
);

BUFx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_195),
.B(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_195),
.Y(n_265)
);

OA22x2_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_199),
.B1(n_201),
.B2(n_202),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_198),
.Y(n_440)
);

INVx8_ASAP7_75t_L g209 ( 
.A(n_199),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_202),
.Y(n_449)
);

INVxp33_ASAP7_75t_L g354 ( 
.A(n_203),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_204),
.B(n_216),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_204),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_204),
.A2(n_353),
.B(n_426),
.Y(n_425)
);

OAI22xp33_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_209),
.B1(n_210),
.B2(n_214),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_207),
.Y(n_258)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx6_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_214),
.Y(n_415)
);

BUFx12f_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_215),
.Y(n_391)
);

INVx4_ASAP7_75t_L g457 ( 
.A(n_215),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_216),
.B(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_225),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g538 ( 
.A1(n_223),
.A2(n_539),
.B(n_543),
.Y(n_538)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_226),
.Y(n_548)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_227),
.Y(n_320)
);

INVx6_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_231),
.Y(n_421)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_232),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_233),
.B(n_242),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_233),
.B(n_242),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_234),
.B(n_241),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g476 ( 
.A(n_234),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_238),
.Y(n_234)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_238),
.Y(n_402)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_244),
.A2(n_256),
.B(n_264),
.Y(n_255)
);

OA21x2_ASAP7_75t_L g315 ( 
.A1(n_244),
.A2(n_245),
.B(n_264),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_244),
.A2(n_404),
.B1(n_410),
.B2(n_416),
.Y(n_403)
);

BUFx2_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx4_ASAP7_75t_L g407 ( 
.A(n_248),
.Y(n_407)
);

INVx6_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_249),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_254),
.C(n_283),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_252),
.B(n_303),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_254),
.B(n_283),
.Y(n_303)
);

MAJx2_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_266),
.C(n_274),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_255),
.B(n_274),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g546 ( 
.A(n_256),
.Y(n_546)
);

OAI32xp33_ASAP7_75t_L g435 ( 
.A1(n_257),
.A2(n_436),
.A3(n_441),
.B1(n_445),
.B2(n_448),
.Y(n_435)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_262),
.Y(n_413)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_265),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_266),
.B(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_278),
.Y(n_296)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_279),
.Y(n_297)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_302),
.Y(n_284)
);

OR2x2_ASAP7_75t_L g373 ( 
.A(n_285),
.B(n_302),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_288),
.C(n_291),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g523 ( 
.A(n_286),
.B(n_524),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_SL g524 ( 
.A1(n_288),
.A2(n_289),
.B1(n_291),
.B2(n_525),
.Y(n_524)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_291),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_298),
.C(n_300),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_SL g428 ( 
.A(n_292),
.B(n_429),
.Y(n_428)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_299),
.B(n_300),
.Y(n_429)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_304),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_306),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_305),
.B(n_306),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_331),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_317),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_308),
.B(n_317),
.C(n_336),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_309),
.A2(n_314),
.B1(n_315),
.B2(n_316),
.Y(n_308)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_309),
.Y(n_316)
);

NOR2x1_ASAP7_75t_R g357 ( 
.A(n_309),
.B(n_315),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_309),
.A2(n_316),
.B1(n_359),
.B2(n_365),
.Y(n_358)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

AOI21xp33_ASAP7_75t_L g553 ( 
.A1(n_316),
.A2(n_365),
.B(n_554),
.Y(n_553)
);

XNOR2x1_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_330),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_326),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g339 ( 
.A(n_319),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_321),
.Y(n_343)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_326),
.B(n_330),
.C(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_328),
.Y(n_360)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_331),
.Y(n_336)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

NOR3xp33_ASAP7_75t_L g370 ( 
.A(n_334),
.B(n_371),
.C(n_374),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_337),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_335),
.B(n_337),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_340),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_338),
.B(n_356),
.C(n_367),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_341),
.A2(n_356),
.B1(n_366),
.B2(n_367),
.Y(n_340)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_341),
.Y(n_367)
);

OAI21xp33_ASAP7_75t_L g341 ( 
.A1(n_342),
.A2(n_352),
.B(n_355),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_342),
.B(n_352),
.Y(n_355)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

HB1xp67_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_354),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g535 ( 
.A1(n_355),
.A2(n_536),
.B1(n_550),
.B2(n_551),
.Y(n_535)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_355),
.Y(n_550)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_356),
.Y(n_366)
);

XNOR2x1_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_358),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g554 ( 
.A(n_357),
.Y(n_554)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_359),
.Y(n_365)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_363),
.Y(n_542)
);

INVx8_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_375),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_372),
.B(n_373),
.Y(n_371)
);

OAI21x1_ASAP7_75t_L g375 ( 
.A1(n_376),
.A2(n_522),
.B(n_527),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g376 ( 
.A1(n_377),
.A2(n_431),
.B(n_521),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_422),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_SL g521 ( 
.A(n_378),
.B(n_422),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_403),
.C(n_417),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g517 ( 
.A(n_379),
.B(n_518),
.Y(n_517)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_401),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_380),
.B(n_401),
.Y(n_424)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

BUFx3_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_396),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

HB1xp67_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g518 ( 
.A(n_403),
.B(n_417),
.Y(n_518)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx4_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_410),
.Y(n_426)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

INVx8_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_423),
.A2(n_427),
.B1(n_428),
.B2(n_430),
.Y(n_422)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_423),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_425),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_424),
.B(n_425),
.C(n_427),
.Y(n_526)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_L g431 ( 
.A1(n_432),
.A2(n_516),
.B(n_520),
.Y(n_431)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_433),
.A2(n_480),
.B(n_515),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_434),
.B(n_467),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_434),
.B(n_467),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_435),
.B(n_453),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_435),
.A2(n_453),
.B1(n_454),
.B2(n_492),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_435),
.Y(n_492)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

BUFx2_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

BUFx2_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

INVx3_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

INVx8_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_449),
.B(n_450),
.Y(n_448)
);

BUFx2_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

BUFx2_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_468),
.B(n_477),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_468),
.B(n_478),
.C(n_479),
.Y(n_519)
);

INVxp67_ASAP7_75t_L g490 ( 
.A(n_469),
.Y(n_490)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_478),
.B(n_479),
.Y(n_477)
);

OAI21xp5_ASAP7_75t_SL g480 ( 
.A1(n_481),
.A2(n_493),
.B(n_514),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_482),
.B(n_491),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_482),
.B(n_491),
.Y(n_514)
);

INVxp67_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

INVx1_ASAP7_75t_SL g485 ( 
.A(n_486),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

BUFx2_ASAP7_75t_L g489 ( 
.A(n_487),
.Y(n_489)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

AOI21xp5_ASAP7_75t_L g493 ( 
.A1(n_494),
.A2(n_508),
.B(n_513),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_495),
.B(n_503),
.Y(n_494)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_499),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_504),
.B(n_506),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

INVx5_ASAP7_75t_L g511 ( 
.A(n_507),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_509),
.B(n_512),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_509),
.B(n_512),
.Y(n_513)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

NOR2xp67_ASAP7_75t_SL g516 ( 
.A(n_517),
.B(n_519),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_517),
.B(n_519),
.Y(n_520)
);

NOR2xp67_ASAP7_75t_SL g522 ( 
.A(n_523),
.B(n_526),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_523),
.B(n_526),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_529),
.B(n_555),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_530),
.Y(n_529)
);

HB1xp67_ASAP7_75t_L g530 ( 
.A(n_531),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_532),
.B(n_533),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_532),
.B(n_533),
.Y(n_555)
);

OAI22xp5_ASAP7_75t_SL g533 ( 
.A1(n_534),
.A2(n_535),
.B1(n_552),
.B2(n_553),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_535),
.Y(n_534)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_536),
.Y(n_551)
);

AOI22xp5_ASAP7_75t_L g536 ( 
.A1(n_537),
.A2(n_538),
.B1(n_544),
.B2(n_549),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_538),
.Y(n_537)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_541),
.Y(n_540)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_544),
.Y(n_549)
);

XNOR2xp5_ASAP7_75t_L g544 ( 
.A(n_545),
.B(n_547),
.Y(n_544)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_553),
.Y(n_552)
);


endmodule