module fake_netlist_1_12610_n_734 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_107, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_106, n_15, n_61, n_21, n_99, n_93, n_51, n_96, n_39, n_734);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_107;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_106;
input n_15;
input n_61;
input n_21;
input n_99;
input n_93;
input n_51;
input n_96;
input n_39;
output n_734;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_732;
wire n_199;
wire n_351;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_724;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_623;
wire n_167;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_711;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_699;
wire n_519;
wire n_729;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_649;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_107), .Y(n_108) );
BUFx6f_ASAP7_75t_L g109 ( .A(n_61), .Y(n_109) );
NOR2xp33_ASAP7_75t_L g110 ( .A(n_14), .B(n_62), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_105), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_41), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_73), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_17), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_22), .Y(n_115) );
BUFx3_ASAP7_75t_L g116 ( .A(n_8), .Y(n_116) );
INVx1_ASAP7_75t_SL g117 ( .A(n_17), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_40), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_5), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_21), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_103), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_7), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_85), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_87), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_11), .Y(n_125) );
BUFx3_ASAP7_75t_L g126 ( .A(n_57), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_90), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_10), .Y(n_128) );
INVx1_ASAP7_75t_SL g129 ( .A(n_46), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_79), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_74), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_44), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g133 ( .A(n_9), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_5), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_63), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_52), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_9), .Y(n_137) );
INVx1_ASAP7_75t_SL g138 ( .A(n_88), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_29), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_32), .Y(n_140) );
BUFx2_ASAP7_75t_L g141 ( .A(n_37), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_24), .Y(n_142) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_25), .Y(n_143) );
INVxp33_ASAP7_75t_L g144 ( .A(n_99), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_10), .Y(n_145) );
INVxp67_ASAP7_75t_L g146 ( .A(n_72), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_70), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_0), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_80), .Y(n_149) );
CKINVDCx16_ASAP7_75t_R g150 ( .A(n_101), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_49), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_14), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_141), .B(n_0), .Y(n_153) );
AOI22xp5_ASAP7_75t_L g154 ( .A1(n_114), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_154) );
AND2x2_ASAP7_75t_L g155 ( .A(n_141), .B(n_1), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_109), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_109), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_109), .Y(n_158) );
BUFx3_ASAP7_75t_L g159 ( .A(n_126), .Y(n_159) );
HB1xp67_ASAP7_75t_L g160 ( .A(n_116), .Y(n_160) );
INVxp67_ASAP7_75t_L g161 ( .A(n_116), .Y(n_161) );
AND2x4_ASAP7_75t_L g162 ( .A(n_119), .B(n_2), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_109), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_109), .Y(n_164) );
OA21x2_ASAP7_75t_L g165 ( .A1(n_118), .A2(n_53), .B(n_104), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_118), .Y(n_166) );
AND2x4_ASAP7_75t_L g167 ( .A(n_119), .B(n_3), .Y(n_167) );
NAND2xp5_ASAP7_75t_SL g168 ( .A(n_143), .B(n_4), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_121), .Y(n_169) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_143), .Y(n_170) );
AND2x2_ASAP7_75t_L g171 ( .A(n_144), .B(n_4), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_121), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g173 ( .A(n_161), .B(n_146), .Y(n_173) );
BUFx3_ASAP7_75t_L g174 ( .A(n_159), .Y(n_174) );
CKINVDCx5p33_ASAP7_75t_R g175 ( .A(n_155), .Y(n_175) );
AOI22xp5_ASAP7_75t_L g176 ( .A1(n_155), .A2(n_114), .B1(n_125), .B2(n_122), .Y(n_176) );
OAI22xp33_ASAP7_75t_L g177 ( .A1(n_154), .A2(n_133), .B1(n_122), .B2(n_125), .Y(n_177) );
BUFx2_ASAP7_75t_L g178 ( .A(n_155), .Y(n_178) );
AND2x4_ASAP7_75t_L g179 ( .A(n_162), .B(n_145), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_162), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_170), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g182 ( .A(n_161), .B(n_111), .Y(n_182) );
INVx3_ASAP7_75t_L g183 ( .A(n_162), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_170), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_166), .B(n_169), .Y(n_185) );
NAND2xp33_ASAP7_75t_L g186 ( .A(n_166), .B(n_143), .Y(n_186) );
AND2x2_ASAP7_75t_L g187 ( .A(n_160), .B(n_150), .Y(n_187) );
BUFx3_ASAP7_75t_L g188 ( .A(n_159), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_162), .Y(n_189) );
BUFx3_ASAP7_75t_L g190 ( .A(n_159), .Y(n_190) );
INVx3_ASAP7_75t_L g191 ( .A(n_167), .Y(n_191) );
AND2x2_ASAP7_75t_L g192 ( .A(n_160), .B(n_145), .Y(n_192) );
AOI22xp5_ASAP7_75t_L g193 ( .A1(n_167), .A2(n_120), .B1(n_130), .B2(n_137), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_169), .B(n_147), .Y(n_194) );
BUFx4f_ASAP7_75t_L g195 ( .A(n_167), .Y(n_195) );
CKINVDCx11_ASAP7_75t_R g196 ( .A(n_167), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_172), .Y(n_197) );
BUFx3_ASAP7_75t_L g198 ( .A(n_165), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_170), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_183), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_178), .B(n_171), .Y(n_201) );
AND2x4_ASAP7_75t_L g202 ( .A(n_178), .B(n_153), .Y(n_202) );
HB1xp67_ASAP7_75t_L g203 ( .A(n_178), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_173), .B(n_171), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_183), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_195), .B(n_153), .Y(n_206) );
O2A1O1Ixp33_ASAP7_75t_L g207 ( .A1(n_192), .A2(n_172), .B(n_168), .C(n_115), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g208 ( .A(n_187), .B(n_108), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_183), .Y(n_209) );
AND2x2_ASAP7_75t_L g210 ( .A(n_187), .B(n_120), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_173), .B(n_108), .Y(n_211) );
INVx1_ASAP7_75t_SL g212 ( .A(n_196), .Y(n_212) );
INVx4_ASAP7_75t_L g213 ( .A(n_195), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_183), .Y(n_214) );
NAND3xp33_ASAP7_75t_SL g215 ( .A(n_193), .B(n_154), .C(n_123), .Y(n_215) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_195), .B(n_123), .Y(n_216) );
NAND2xp33_ASAP7_75t_L g217 ( .A(n_180), .B(n_127), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_183), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_191), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g220 ( .A(n_187), .B(n_127), .Y(n_220) );
INVx2_ASAP7_75t_SL g221 ( .A(n_195), .Y(n_221) );
CKINVDCx20_ASAP7_75t_R g222 ( .A(n_176), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_185), .B(n_131), .Y(n_223) );
A2O1A1Ixp33_ASAP7_75t_L g224 ( .A1(n_195), .A2(n_147), .B(n_134), .C(n_142), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_191), .Y(n_225) );
AOI22xp5_ASAP7_75t_L g226 ( .A1(n_175), .A2(n_152), .B1(n_148), .B2(n_128), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_185), .B(n_131), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_182), .B(n_136), .Y(n_228) );
AOI22xp33_ASAP7_75t_L g229 ( .A1(n_179), .A2(n_139), .B1(n_135), .B2(n_112), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_191), .Y(n_230) );
AND2x4_ASAP7_75t_L g231 ( .A(n_179), .B(n_117), .Y(n_231) );
INVx3_ASAP7_75t_L g232 ( .A(n_191), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_191), .Y(n_233) );
INVx2_ASAP7_75t_L g234 ( .A(n_198), .Y(n_234) );
NAND2xp5_ASAP7_75t_SL g235 ( .A(n_179), .B(n_136), .Y(n_235) );
AOI22xp5_ASAP7_75t_L g236 ( .A1(n_210), .A2(n_196), .B1(n_193), .B2(n_176), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_232), .Y(n_237) );
BUFx2_ASAP7_75t_L g238 ( .A(n_203), .Y(n_238) );
NOR3xp33_ASAP7_75t_SL g239 ( .A(n_215), .B(n_177), .C(n_182), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_206), .A2(n_189), .B(n_180), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_200), .A2(n_189), .B(n_198), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_202), .B(n_192), .Y(n_242) );
A2O1A1Ixp33_ASAP7_75t_L g243 ( .A1(n_207), .A2(n_197), .B(n_179), .C(n_198), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_202), .B(n_192), .Y(n_244) );
A2O1A1Ixp33_ASAP7_75t_L g245 ( .A1(n_200), .A2(n_197), .B(n_179), .C(n_198), .Y(n_245) );
INVx3_ASAP7_75t_L g246 ( .A(n_213), .Y(n_246) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_205), .A2(n_209), .B(n_225), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_232), .Y(n_248) );
NAND2xp5_ASAP7_75t_SL g249 ( .A(n_213), .B(n_174), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_205), .A2(n_174), .B(n_190), .Y(n_250) );
INVx2_ASAP7_75t_SL g251 ( .A(n_231), .Y(n_251) );
AOI22xp33_ASAP7_75t_L g252 ( .A1(n_202), .A2(n_177), .B1(n_194), .B2(n_190), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_202), .B(n_194), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_201), .B(n_174), .Y(n_254) );
OAI21xp33_ASAP7_75t_L g255 ( .A1(n_210), .A2(n_190), .B(n_188), .Y(n_255) );
OAI22xp5_ASAP7_75t_L g256 ( .A1(n_213), .A2(n_174), .B1(n_190), .B2(n_188), .Y(n_256) );
NAND2xp5_ASAP7_75t_SL g257 ( .A(n_213), .B(n_188), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_218), .Y(n_258) );
BUFx6f_ASAP7_75t_L g259 ( .A(n_234), .Y(n_259) );
NOR2xp33_ASAP7_75t_SL g260 ( .A(n_212), .B(n_188), .Y(n_260) );
BUFx2_ASAP7_75t_L g261 ( .A(n_231), .Y(n_261) );
AOI22xp5_ASAP7_75t_L g262 ( .A1(n_208), .A2(n_110), .B1(n_151), .B2(n_149), .Y(n_262) );
A2O1A1Ixp33_ASAP7_75t_L g263 ( .A1(n_209), .A2(n_113), .B(n_124), .C(n_132), .Y(n_263) );
AO22x1_ASAP7_75t_L g264 ( .A1(n_212), .A2(n_129), .B1(n_138), .B2(n_140), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_232), .Y(n_265) );
BUFx2_ASAP7_75t_L g266 ( .A(n_231), .Y(n_266) );
INVx2_ASAP7_75t_SL g267 ( .A(n_231), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_242), .B(n_220), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_258), .Y(n_269) );
AOI21xp5_ASAP7_75t_L g270 ( .A1(n_241), .A2(n_234), .B(n_225), .Y(n_270) );
BUFx6f_ASAP7_75t_L g271 ( .A(n_259), .Y(n_271) );
AO31x2_ASAP7_75t_L g272 ( .A1(n_245), .A2(n_224), .A3(n_234), .B(n_156), .Y(n_272) );
AOI22xp33_ASAP7_75t_L g273 ( .A1(n_238), .A2(n_222), .B1(n_221), .B2(n_235), .Y(n_273) );
NOR2xp33_ASAP7_75t_L g274 ( .A(n_236), .B(n_242), .Y(n_274) );
CKINVDCx5p33_ASAP7_75t_R g275 ( .A(n_264), .Y(n_275) );
O2A1O1Ixp33_ASAP7_75t_L g276 ( .A1(n_263), .A2(n_204), .B(n_223), .C(n_227), .Y(n_276) );
CKINVDCx5p33_ASAP7_75t_R g277 ( .A(n_261), .Y(n_277) );
NOR2xp33_ASAP7_75t_SL g278 ( .A(n_259), .B(n_221), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_244), .B(n_226), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_258), .Y(n_280) );
AND2x2_ASAP7_75t_L g281 ( .A(n_266), .B(n_226), .Y(n_281) );
AOI22xp33_ASAP7_75t_L g282 ( .A1(n_251), .A2(n_217), .B1(n_232), .B2(n_228), .Y(n_282) );
AOI21xp5_ASAP7_75t_L g283 ( .A1(n_245), .A2(n_247), .B(n_240), .Y(n_283) );
AOI21xp5_ASAP7_75t_L g284 ( .A1(n_249), .A2(n_230), .B(n_214), .Y(n_284) );
O2A1O1Ixp33_ASAP7_75t_SL g285 ( .A1(n_243), .A2(n_214), .B(n_230), .C(n_219), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_239), .B(n_229), .Y(n_286) );
A2O1A1Ixp33_ASAP7_75t_L g287 ( .A1(n_243), .A2(n_219), .B(n_233), .C(n_218), .Y(n_287) );
A2O1A1Ixp33_ASAP7_75t_L g288 ( .A1(n_255), .A2(n_233), .B(n_218), .C(n_211), .Y(n_288) );
INVx1_ASAP7_75t_SL g289 ( .A(n_246), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_252), .B(n_233), .Y(n_290) );
OA21x2_ASAP7_75t_L g291 ( .A1(n_263), .A2(n_164), .B(n_158), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_280), .Y(n_292) );
AND2x4_ASAP7_75t_L g293 ( .A(n_280), .B(n_246), .Y(n_293) );
AOI21xp5_ASAP7_75t_L g294 ( .A1(n_285), .A2(n_283), .B(n_276), .Y(n_294) );
INVx2_ASAP7_75t_SL g295 ( .A(n_269), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_279), .B(n_253), .Y(n_296) );
OAI221xp5_ASAP7_75t_L g297 ( .A1(n_274), .A2(n_262), .B1(n_267), .B2(n_254), .C(n_260), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_268), .B(n_286), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_269), .Y(n_299) );
AND2x2_ASAP7_75t_L g300 ( .A(n_281), .B(n_246), .Y(n_300) );
AO221x2_ASAP7_75t_L g301 ( .A1(n_275), .A2(n_256), .B1(n_7), .B2(n_8), .C(n_11), .Y(n_301) );
AOI21xp33_ASAP7_75t_L g302 ( .A1(n_290), .A2(n_249), .B(n_257), .Y(n_302) );
AO21x2_ASAP7_75t_L g303 ( .A1(n_287), .A2(n_257), .B(n_250), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_281), .B(n_237), .Y(n_304) );
OAI22xp33_ASAP7_75t_L g305 ( .A1(n_275), .A2(n_265), .B1(n_248), .B2(n_259), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_269), .Y(n_306) );
AND2x2_ASAP7_75t_L g307 ( .A(n_272), .B(n_259), .Y(n_307) );
INVx3_ASAP7_75t_L g308 ( .A(n_271), .Y(n_308) );
AND2x2_ASAP7_75t_L g309 ( .A(n_272), .B(n_291), .Y(n_309) );
NAND3xp33_ASAP7_75t_L g310 ( .A(n_291), .B(n_170), .C(n_165), .Y(n_310) );
AO31x2_ASAP7_75t_L g311 ( .A1(n_288), .A2(n_163), .A3(n_164), .B(n_156), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_271), .Y(n_312) );
CKINVDCx6p67_ASAP7_75t_R g313 ( .A(n_289), .Y(n_313) );
BUFx2_ASAP7_75t_L g314 ( .A(n_307), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_292), .Y(n_315) );
HB1xp67_ASAP7_75t_L g316 ( .A(n_295), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_292), .Y(n_317) );
OA21x2_ASAP7_75t_L g318 ( .A1(n_294), .A2(n_270), .B(n_284), .Y(n_318) );
BUFx3_ASAP7_75t_L g319 ( .A(n_313), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_299), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_299), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_306), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_296), .B(n_306), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_309), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_309), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_307), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_312), .Y(n_327) );
AND2x2_ASAP7_75t_L g328 ( .A(n_295), .B(n_272), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_312), .Y(n_329) );
NAND4xp25_ASAP7_75t_L g330 ( .A(n_298), .B(n_273), .C(n_282), .D(n_126), .Y(n_330) );
AND2x2_ASAP7_75t_L g331 ( .A(n_300), .B(n_272), .Y(n_331) );
AO21x2_ASAP7_75t_L g332 ( .A1(n_294), .A2(n_158), .B(n_156), .Y(n_332) );
OAI21xp5_ASAP7_75t_L g333 ( .A1(n_298), .A2(n_291), .B(n_289), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_300), .B(n_272), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_301), .B(n_272), .Y(n_335) );
OA21x2_ASAP7_75t_L g336 ( .A1(n_310), .A2(n_157), .B(n_158), .Y(n_336) );
INVx3_ASAP7_75t_L g337 ( .A(n_308), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_304), .Y(n_338) );
NAND2xp5_ASAP7_75t_SL g339 ( .A(n_305), .B(n_308), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_312), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_311), .Y(n_341) );
AND2x2_ASAP7_75t_L g342 ( .A(n_324), .B(n_311), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_338), .B(n_296), .Y(n_343) );
HB1xp67_ASAP7_75t_L g344 ( .A(n_316), .Y(n_344) );
AND2x4_ASAP7_75t_L g345 ( .A(n_324), .B(n_308), .Y(n_345) );
OR2x2_ASAP7_75t_L g346 ( .A(n_314), .B(n_304), .Y(n_346) );
INVx3_ASAP7_75t_L g347 ( .A(n_337), .Y(n_347) );
CKINVDCx20_ASAP7_75t_R g348 ( .A(n_319), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_322), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_324), .B(n_325), .Y(n_350) );
AND2x2_ASAP7_75t_L g351 ( .A(n_324), .B(n_311), .Y(n_351) );
NOR2x1_ASAP7_75t_SL g352 ( .A(n_319), .B(n_271), .Y(n_352) );
AND2x2_ASAP7_75t_L g353 ( .A(n_325), .B(n_311), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_322), .Y(n_354) );
AND2x2_ASAP7_75t_L g355 ( .A(n_325), .B(n_311), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_322), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_327), .Y(n_357) );
NOR3xp33_ASAP7_75t_SL g358 ( .A(n_330), .B(n_297), .C(n_277), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_325), .B(n_311), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_315), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_315), .Y(n_361) );
BUFx2_ASAP7_75t_L g362 ( .A(n_316), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_338), .B(n_301), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_327), .Y(n_364) );
INVx4_ASAP7_75t_L g365 ( .A(n_319), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_317), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_326), .B(n_291), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_327), .Y(n_368) );
OR2x2_ASAP7_75t_L g369 ( .A(n_314), .B(n_301), .Y(n_369) );
HB1xp67_ASAP7_75t_L g370 ( .A(n_327), .Y(n_370) );
INVxp67_ASAP7_75t_SL g371 ( .A(n_329), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_329), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_317), .B(n_301), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_320), .Y(n_374) );
BUFx2_ASAP7_75t_L g375 ( .A(n_319), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_320), .Y(n_376) );
HB1xp67_ASAP7_75t_L g377 ( .A(n_329), .Y(n_377) );
HB1xp67_ASAP7_75t_L g378 ( .A(n_329), .Y(n_378) );
BUFx3_ASAP7_75t_L g379 ( .A(n_337), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_321), .Y(n_380) );
HB1xp67_ASAP7_75t_L g381 ( .A(n_340), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_326), .B(n_301), .Y(n_382) );
OR2x2_ASAP7_75t_L g383 ( .A(n_314), .B(n_313), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_321), .Y(n_384) );
OR2x2_ASAP7_75t_L g385 ( .A(n_326), .B(n_313), .Y(n_385) );
HB1xp67_ASAP7_75t_L g386 ( .A(n_340), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_350), .B(n_331), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_349), .Y(n_388) );
AND2x4_ASAP7_75t_L g389 ( .A(n_350), .B(n_328), .Y(n_389) );
NAND4xp25_ASAP7_75t_L g390 ( .A(n_369), .B(n_330), .C(n_335), .D(n_297), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_349), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_354), .Y(n_392) );
NAND4xp25_ASAP7_75t_L g393 ( .A(n_369), .B(n_335), .C(n_331), .D(n_334), .Y(n_393) );
OR2x2_ASAP7_75t_L g394 ( .A(n_350), .B(n_331), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_357), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_367), .B(n_334), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_357), .Y(n_397) );
HB1xp67_ASAP7_75t_L g398 ( .A(n_362), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_357), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_354), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_367), .B(n_334), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_356), .Y(n_402) );
OR2x2_ASAP7_75t_L g403 ( .A(n_346), .B(n_328), .Y(n_403) );
OR2x2_ASAP7_75t_L g404 ( .A(n_346), .B(n_328), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_356), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_367), .B(n_335), .Y(n_406) );
INVx1_ASAP7_75t_SL g407 ( .A(n_375), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_343), .B(n_323), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_364), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_360), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_360), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_342), .B(n_341), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_342), .B(n_341), .Y(n_413) );
OR2x2_ASAP7_75t_L g414 ( .A(n_362), .B(n_341), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_342), .B(n_340), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_361), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_351), .B(n_340), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_343), .B(n_323), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_351), .B(n_333), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_351), .B(n_333), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_353), .B(n_332), .Y(n_421) );
CKINVDCx5p33_ASAP7_75t_R g422 ( .A(n_348), .Y(n_422) );
OR2x2_ASAP7_75t_L g423 ( .A(n_344), .B(n_332), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_353), .B(n_332), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_353), .B(n_332), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_361), .B(n_337), .Y(n_426) );
HB1xp67_ASAP7_75t_L g427 ( .A(n_344), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_364), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_355), .B(n_332), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_366), .B(n_337), .Y(n_430) );
AOI21xp33_ASAP7_75t_L g431 ( .A1(n_373), .A2(n_339), .B(n_337), .Y(n_431) );
OR2x6_ASAP7_75t_L g432 ( .A(n_365), .B(n_339), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_355), .B(n_336), .Y(n_433) );
NOR2xp33_ASAP7_75t_L g434 ( .A(n_363), .B(n_277), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_364), .Y(n_435) );
NAND2xp5_ASAP7_75t_SL g436 ( .A(n_365), .B(n_293), .Y(n_436) );
HB1xp67_ASAP7_75t_L g437 ( .A(n_383), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_355), .B(n_336), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_366), .Y(n_439) );
INVx2_ASAP7_75t_SL g440 ( .A(n_365), .Y(n_440) );
OR2x2_ASAP7_75t_L g441 ( .A(n_383), .B(n_318), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_359), .B(n_336), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_359), .B(n_336), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_359), .B(n_336), .Y(n_444) );
NOR4xp25_ASAP7_75t_SL g445 ( .A(n_375), .B(n_302), .C(n_336), .D(n_13), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_382), .B(n_318), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_382), .B(n_318), .Y(n_447) );
OR2x2_ASAP7_75t_L g448 ( .A(n_370), .B(n_318), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_382), .B(n_293), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_370), .B(n_318), .Y(n_450) );
BUFx2_ASAP7_75t_L g451 ( .A(n_365), .Y(n_451) );
INVxp67_ASAP7_75t_L g452 ( .A(n_385), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_377), .B(n_318), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_374), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_374), .Y(n_455) );
INVx2_ASAP7_75t_SL g456 ( .A(n_451), .Y(n_456) );
NAND4xp75_ASAP7_75t_L g457 ( .A(n_440), .B(n_358), .C(n_363), .D(n_373), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_387), .B(n_376), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_410), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_446), .B(n_377), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_410), .Y(n_461) );
OR2x2_ASAP7_75t_L g462 ( .A(n_394), .B(n_378), .Y(n_462) );
HB1xp67_ASAP7_75t_L g463 ( .A(n_427), .Y(n_463) );
INVxp67_ASAP7_75t_L g464 ( .A(n_451), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_395), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_387), .B(n_376), .Y(n_466) );
OR2x2_ASAP7_75t_L g467 ( .A(n_394), .B(n_378), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_446), .B(n_381), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_411), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_447), .B(n_381), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_411), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_395), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_412), .B(n_380), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_416), .Y(n_474) );
OR2x2_ASAP7_75t_L g475 ( .A(n_403), .B(n_386), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_416), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_389), .B(n_345), .Y(n_477) );
INVxp67_ASAP7_75t_L g478 ( .A(n_398), .Y(n_478) );
NAND2xp5_ASAP7_75t_SL g479 ( .A(n_440), .B(n_358), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_395), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_439), .Y(n_481) );
OR2x2_ASAP7_75t_L g482 ( .A(n_403), .B(n_386), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_447), .B(n_345), .Y(n_483) );
NAND2x1_ASAP7_75t_L g484 ( .A(n_432), .B(n_380), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_439), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_389), .B(n_412), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_413), .B(n_384), .Y(n_487) );
NOR2xp33_ASAP7_75t_L g488 ( .A(n_390), .B(n_384), .Y(n_488) );
NAND2xp5_ASAP7_75t_SL g489 ( .A(n_407), .B(n_385), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_454), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_454), .Y(n_491) );
INVxp67_ASAP7_75t_L g492 ( .A(n_437), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_389), .B(n_345), .Y(n_493) );
INVxp67_ASAP7_75t_SL g494 ( .A(n_448), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_455), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_455), .Y(n_496) );
AND3x2_ASAP7_75t_L g497 ( .A(n_452), .B(n_371), .C(n_345), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_413), .B(n_371), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_389), .B(n_345), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_388), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_388), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_397), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_406), .B(n_368), .Y(n_503) );
NAND2xp5_ASAP7_75t_SL g504 ( .A(n_407), .B(n_368), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_406), .B(n_368), .Y(n_505) );
HB1xp67_ASAP7_75t_L g506 ( .A(n_448), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_391), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_408), .B(n_372), .Y(n_508) );
INVx2_ASAP7_75t_L g509 ( .A(n_397), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_391), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_396), .B(n_379), .Y(n_511) );
OAI21xp33_ASAP7_75t_SL g512 ( .A1(n_390), .A2(n_347), .B(n_372), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_418), .B(n_372), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_396), .B(n_347), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_401), .B(n_379), .Y(n_515) );
NAND2x1p5_ASAP7_75t_L g516 ( .A(n_436), .B(n_379), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_392), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_401), .B(n_347), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_397), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_415), .B(n_347), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g521 ( .A(n_434), .B(n_6), .Y(n_521) );
OR2x2_ASAP7_75t_L g522 ( .A(n_404), .B(n_6), .Y(n_522) );
OR2x2_ASAP7_75t_L g523 ( .A(n_404), .B(n_12), .Y(n_523) );
AND2x4_ASAP7_75t_L g524 ( .A(n_432), .B(n_352), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_392), .Y(n_525) );
OR2x2_ASAP7_75t_L g526 ( .A(n_414), .B(n_12), .Y(n_526) );
INVx2_ASAP7_75t_L g527 ( .A(n_399), .Y(n_527) );
INVx2_ASAP7_75t_SL g528 ( .A(n_432), .Y(n_528) );
OR2x2_ASAP7_75t_L g529 ( .A(n_414), .B(n_13), .Y(n_529) );
CKINVDCx5p33_ASAP7_75t_R g530 ( .A(n_422), .Y(n_530) );
INVx2_ASAP7_75t_L g531 ( .A(n_399), .Y(n_531) );
INVx2_ASAP7_75t_L g532 ( .A(n_399), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_400), .Y(n_533) );
OR2x2_ASAP7_75t_L g534 ( .A(n_393), .B(n_415), .Y(n_534) );
INVxp67_ASAP7_75t_SL g535 ( .A(n_441), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_400), .Y(n_536) );
INVx2_ASAP7_75t_L g537 ( .A(n_409), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_402), .Y(n_538) );
HB1xp67_ASAP7_75t_L g539 ( .A(n_409), .Y(n_539) );
HB1xp67_ASAP7_75t_L g540 ( .A(n_409), .Y(n_540) );
OR2x2_ASAP7_75t_L g541 ( .A(n_462), .B(n_441), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_486), .B(n_421), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_463), .Y(n_543) );
OAI21xp5_ASAP7_75t_L g544 ( .A1(n_479), .A2(n_432), .B(n_423), .Y(n_544) );
BUFx3_ASAP7_75t_L g545 ( .A(n_456), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_486), .B(n_421), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_483), .B(n_424), .Y(n_547) );
OA22x2_ASAP7_75t_L g548 ( .A1(n_497), .A2(n_432), .B1(n_449), .B2(n_405), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_463), .Y(n_549) );
AOI22xp5_ASAP7_75t_L g550 ( .A1(n_488), .A2(n_393), .B1(n_424), .B2(n_425), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_459), .Y(n_551) );
INVx1_ASAP7_75t_SL g552 ( .A(n_530), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_488), .B(n_425), .Y(n_553) );
INVx2_ASAP7_75t_L g554 ( .A(n_465), .Y(n_554) );
INVxp67_ASAP7_75t_L g555 ( .A(n_456), .Y(n_555) );
NOR2xp33_ASAP7_75t_L g556 ( .A(n_492), .B(n_431), .Y(n_556) );
OAI32xp33_ASAP7_75t_L g557 ( .A1(n_512), .A2(n_423), .A3(n_402), .B1(n_405), .B2(n_453), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_499), .B(n_429), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_483), .B(n_429), .Y(n_559) );
INVx2_ASAP7_75t_L g560 ( .A(n_465), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_535), .B(n_419), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_460), .B(n_417), .Y(n_562) );
BUFx3_ASAP7_75t_L g563 ( .A(n_516), .Y(n_563) );
OAI21xp5_ASAP7_75t_L g564 ( .A1(n_479), .A2(n_453), .B(n_450), .Y(n_564) );
AOI21xp33_ASAP7_75t_L g565 ( .A1(n_521), .A2(n_529), .B(n_526), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_460), .B(n_417), .Y(n_566) );
NOR2xp33_ASAP7_75t_L g567 ( .A(n_478), .B(n_426), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_499), .B(n_419), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_477), .B(n_420), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_461), .Y(n_570) );
XNOR2xp5_ASAP7_75t_L g571 ( .A(n_530), .B(n_420), .Y(n_571) );
OR2x2_ASAP7_75t_L g572 ( .A(n_467), .B(n_433), .Y(n_572) );
INVxp67_ASAP7_75t_L g573 ( .A(n_506), .Y(n_573) );
OAI22xp33_ASAP7_75t_L g574 ( .A1(n_534), .A2(n_430), .B1(n_442), .B2(n_444), .Y(n_574) );
AND2x4_ASAP7_75t_L g575 ( .A(n_524), .B(n_528), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_493), .B(n_433), .Y(n_576) );
OR2x2_ASAP7_75t_L g577 ( .A(n_475), .B(n_438), .Y(n_577) );
OR2x2_ASAP7_75t_L g578 ( .A(n_482), .B(n_438), .Y(n_578) );
INVx1_ASAP7_75t_SL g579 ( .A(n_511), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_494), .B(n_450), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_469), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_515), .B(n_442), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_503), .B(n_443), .Y(n_583) );
INVx1_ASAP7_75t_SL g584 ( .A(n_498), .Y(n_584) );
AND2x2_ASAP7_75t_L g585 ( .A(n_503), .B(n_443), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_468), .B(n_444), .Y(n_586) );
INVx2_ASAP7_75t_L g587 ( .A(n_472), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_468), .B(n_428), .Y(n_588) );
AND2x2_ASAP7_75t_L g589 ( .A(n_470), .B(n_428), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_506), .B(n_428), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g591 ( .A(n_457), .B(n_435), .Y(n_591) );
AND2x4_ASAP7_75t_L g592 ( .A(n_524), .B(n_435), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_458), .B(n_435), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_466), .B(n_445), .Y(n_594) );
NAND2xp5_ASAP7_75t_SL g595 ( .A(n_524), .B(n_308), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_471), .Y(n_596) );
INVx2_ASAP7_75t_L g597 ( .A(n_472), .Y(n_597) );
OAI31xp33_ASAP7_75t_L g598 ( .A1(n_521), .A2(n_293), .A3(n_310), .B(n_302), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_470), .B(n_445), .Y(n_599) );
OAI21xp5_ASAP7_75t_L g600 ( .A1(n_489), .A2(n_157), .B(n_163), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_505), .B(n_352), .Y(n_601) );
AND2x2_ASAP7_75t_L g602 ( .A(n_505), .B(n_170), .Y(n_602) );
AND2x2_ASAP7_75t_L g603 ( .A(n_520), .B(n_170), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_473), .B(n_143), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_514), .B(n_518), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_487), .B(n_143), .Y(n_606) );
OR2x2_ASAP7_75t_L g607 ( .A(n_508), .B(n_157), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_474), .Y(n_608) );
NOR2xp33_ASAP7_75t_L g609 ( .A(n_522), .B(n_523), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_476), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_481), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_485), .Y(n_612) );
AND2x2_ASAP7_75t_L g613 ( .A(n_539), .B(n_170), .Y(n_613) );
AOI22xp5_ASAP7_75t_L g614 ( .A1(n_489), .A2(n_293), .B1(n_303), .B2(n_165), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_513), .B(n_303), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_490), .B(n_303), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_491), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_495), .B(n_303), .Y(n_618) );
OR2x2_ASAP7_75t_L g619 ( .A(n_541), .B(n_464), .Y(n_619) );
OAI211xp5_ASAP7_75t_SL g620 ( .A1(n_565), .A2(n_528), .B(n_504), .C(n_496), .Y(n_620) );
NOR2xp33_ASAP7_75t_L g621 ( .A(n_552), .B(n_500), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_543), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_553), .B(n_501), .Y(n_623) );
AOI22xp33_ASAP7_75t_L g624 ( .A1(n_550), .A2(n_484), .B1(n_516), .B2(n_538), .Y(n_624) );
OAI221xp5_ASAP7_75t_L g625 ( .A1(n_564), .A2(n_510), .B1(n_507), .B2(n_536), .C(n_533), .Y(n_625) );
OR2x2_ASAP7_75t_L g626 ( .A(n_580), .B(n_539), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_549), .Y(n_627) );
OA21x2_ASAP7_75t_SL g628 ( .A1(n_579), .A2(n_504), .B(n_16), .Y(n_628) );
AOI22xp33_ASAP7_75t_L g629 ( .A1(n_574), .A2(n_517), .B1(n_525), .B2(n_540), .Y(n_629) );
OAI211xp5_ASAP7_75t_SL g630 ( .A1(n_598), .A2(n_163), .B(n_164), .C(n_532), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_551), .Y(n_631) );
AOI22xp5_ASAP7_75t_L g632 ( .A1(n_574), .A2(n_540), .B1(n_537), .B2(n_532), .Y(n_632) );
AOI222xp33_ASAP7_75t_L g633 ( .A1(n_544), .A2(n_609), .B1(n_599), .B2(n_594), .C1(n_571), .C2(n_591), .Y(n_633) );
NOR2xp33_ASAP7_75t_L g634 ( .A(n_584), .B(n_480), .Y(n_634) );
INVx1_ASAP7_75t_SL g635 ( .A(n_545), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_573), .B(n_480), .Y(n_636) );
AND2x2_ASAP7_75t_L g637 ( .A(n_547), .B(n_502), .Y(n_637) );
INVxp67_ASAP7_75t_L g638 ( .A(n_556), .Y(n_638) );
INVx2_ASAP7_75t_L g639 ( .A(n_613), .Y(n_639) );
AOI221xp5_ASAP7_75t_L g640 ( .A1(n_556), .A2(n_537), .B1(n_531), .B2(n_527), .C(n_519), .Y(n_640) );
INVx2_ASAP7_75t_L g641 ( .A(n_613), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_570), .Y(n_642) );
NAND2x1p5_ASAP7_75t_L g643 ( .A(n_563), .B(n_502), .Y(n_643) );
INVx3_ASAP7_75t_L g644 ( .A(n_575), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_602), .B(n_509), .Y(n_645) );
OAI21xp33_ASAP7_75t_L g646 ( .A1(n_548), .A2(n_531), .B(n_527), .Y(n_646) );
AOI32xp33_ASAP7_75t_L g647 ( .A1(n_545), .A2(n_519), .A3(n_509), .B1(n_278), .B2(n_19), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_602), .B(n_15), .Y(n_648) );
AOI221xp5_ASAP7_75t_L g649 ( .A1(n_609), .A2(n_216), .B1(n_16), .B2(n_18), .C(n_19), .Y(n_649) );
AOI22xp5_ASAP7_75t_L g650 ( .A1(n_591), .A2(n_165), .B1(n_278), .B2(n_271), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_546), .B(n_15), .Y(n_651) );
INVxp67_ASAP7_75t_SL g652 ( .A(n_590), .Y(n_652) );
NOR3xp33_ASAP7_75t_L g653 ( .A(n_604), .B(n_181), .C(n_184), .Y(n_653) );
AOI221xp5_ASAP7_75t_L g654 ( .A1(n_557), .A2(n_18), .B1(n_20), .B2(n_21), .C(n_22), .Y(n_654) );
AOI22x1_ASAP7_75t_L g655 ( .A1(n_555), .A2(n_20), .B1(n_23), .B2(n_24), .Y(n_655) );
AOI221xp5_ASAP7_75t_L g656 ( .A1(n_567), .A2(n_23), .B1(n_199), .B2(n_184), .C(n_181), .Y(n_656) );
XNOR2xp5_ASAP7_75t_L g657 ( .A(n_601), .B(n_26), .Y(n_657) );
AND2x2_ASAP7_75t_L g658 ( .A(n_547), .B(n_165), .Y(n_658) );
AOI22xp5_ASAP7_75t_L g659 ( .A1(n_567), .A2(n_271), .B1(n_199), .B2(n_184), .Y(n_659) );
INVxp67_ASAP7_75t_SL g660 ( .A(n_606), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_581), .Y(n_661) );
NOR2x1_ASAP7_75t_L g662 ( .A(n_563), .B(n_27), .Y(n_662) );
INVx2_ASAP7_75t_SL g663 ( .A(n_601), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_546), .B(n_28), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_596), .Y(n_665) );
AO22x1_ASAP7_75t_L g666 ( .A1(n_575), .A2(n_30), .B1(n_31), .B2(n_33), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_608), .B(n_34), .Y(n_667) );
AOI22xp5_ASAP7_75t_L g668 ( .A1(n_548), .A2(n_199), .B1(n_181), .B2(n_186), .Y(n_668) );
INVxp67_ASAP7_75t_L g669 ( .A(n_603), .Y(n_669) );
OAI32xp33_ASAP7_75t_L g670 ( .A1(n_635), .A2(n_561), .A3(n_572), .B1(n_577), .B2(n_578), .Y(n_670) );
AOI211x1_ASAP7_75t_SL g671 ( .A1(n_628), .A2(n_600), .B(n_615), .C(n_593), .Y(n_671) );
AOI221xp5_ASAP7_75t_SL g672 ( .A1(n_638), .A2(n_605), .B1(n_559), .B2(n_586), .C(n_542), .Y(n_672) );
OAI21xp5_ASAP7_75t_L g673 ( .A1(n_633), .A2(n_603), .B(n_595), .Y(n_673) );
OAI211xp5_ASAP7_75t_L g674 ( .A1(n_633), .A2(n_595), .B(n_614), .C(n_607), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_631), .Y(n_675) );
AOI21xp33_ASAP7_75t_L g676 ( .A1(n_660), .A2(n_618), .B(n_616), .Y(n_676) );
OAI31xp33_ASAP7_75t_L g677 ( .A1(n_646), .A2(n_575), .A3(n_592), .B(n_586), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_642), .Y(n_678) );
AOI221x1_ASAP7_75t_L g679 ( .A1(n_620), .A2(n_617), .B1(n_612), .B2(n_611), .C(n_610), .Y(n_679) );
AOI21xp33_ASAP7_75t_L g680 ( .A1(n_668), .A2(n_592), .B(n_597), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_652), .B(n_605), .Y(n_681) );
O2A1O1Ixp33_ASAP7_75t_L g682 ( .A1(n_651), .A2(n_597), .B(n_560), .C(n_587), .Y(n_682) );
OAI221xp5_ASAP7_75t_L g683 ( .A1(n_629), .A2(n_559), .B1(n_587), .B2(n_560), .C(n_554), .Y(n_683) );
OAI21xp5_ASAP7_75t_L g684 ( .A1(n_654), .A2(n_592), .B(n_562), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_669), .B(n_558), .Y(n_685) );
OAI21xp5_ASAP7_75t_L g686 ( .A1(n_635), .A2(n_566), .B(n_562), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_661), .Y(n_687) );
OAI22xp33_ASAP7_75t_SL g688 ( .A1(n_644), .A2(n_554), .B1(n_566), .B2(n_582), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_665), .Y(n_689) );
A2O1A1Ixp33_ASAP7_75t_SL g690 ( .A1(n_647), .A2(n_630), .B(n_624), .C(n_648), .Y(n_690) );
NAND4xp25_ASAP7_75t_SL g691 ( .A(n_632), .B(n_585), .C(n_583), .D(n_589), .Y(n_691) );
AOI22xp5_ASAP7_75t_L g692 ( .A1(n_621), .A2(n_589), .B1(n_588), .B2(n_568), .Y(n_692) );
NAND2x1_ASAP7_75t_SL g693 ( .A(n_662), .B(n_588), .Y(n_693) );
OAI22xp33_ASAP7_75t_L g694 ( .A1(n_644), .A2(n_576), .B1(n_569), .B2(n_38), .Y(n_694) );
OAI22xp33_ASAP7_75t_L g695 ( .A1(n_625), .A2(n_35), .B1(n_36), .B2(n_39), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_640), .B(n_42), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_622), .Y(n_697) );
AOI221xp5_ASAP7_75t_L g698 ( .A1(n_673), .A2(n_623), .B1(n_627), .B2(n_634), .C(n_649), .Y(n_698) );
OAI221xp5_ASAP7_75t_L g699 ( .A1(n_671), .A2(n_655), .B1(n_657), .B2(n_643), .C(n_663), .Y(n_699) );
AOI221xp5_ASAP7_75t_L g700 ( .A1(n_670), .A2(n_636), .B1(n_645), .B2(n_641), .C(n_639), .Y(n_700) );
AOI21xp5_ASAP7_75t_L g701 ( .A1(n_688), .A2(n_666), .B(n_643), .Y(n_701) );
OA22x2_ASAP7_75t_L g702 ( .A1(n_679), .A2(n_637), .B1(n_664), .B2(n_658), .Y(n_702) );
AOI211xp5_ASAP7_75t_L g703 ( .A1(n_674), .A2(n_656), .B(n_619), .C(n_626), .Y(n_703) );
AOI21xp5_ASAP7_75t_L g704 ( .A1(n_682), .A2(n_667), .B(n_653), .Y(n_704) );
NOR2xp33_ASAP7_75t_SL g705 ( .A(n_694), .B(n_667), .Y(n_705) );
AOI21xp5_ASAP7_75t_L g706 ( .A1(n_682), .A2(n_659), .B(n_650), .Y(n_706) );
NAND4xp75_ASAP7_75t_L g707 ( .A(n_677), .B(n_43), .C(n_45), .D(n_47), .Y(n_707) );
AOI221xp5_ASAP7_75t_L g708 ( .A1(n_672), .A2(n_186), .B1(n_50), .B2(n_51), .C(n_54), .Y(n_708) );
AOI211x1_ASAP7_75t_L g709 ( .A1(n_691), .A2(n_48), .B(n_55), .C(n_56), .Y(n_709) );
AOI221xp5_ASAP7_75t_L g710 ( .A1(n_683), .A2(n_58), .B1(n_59), .B2(n_60), .C(n_64), .Y(n_710) );
AOI22xp5_ASAP7_75t_L g711 ( .A1(n_684), .A2(n_65), .B1(n_66), .B2(n_67), .Y(n_711) );
AOI221xp5_ASAP7_75t_L g712 ( .A1(n_698), .A2(n_676), .B1(n_680), .B2(n_690), .C(n_686), .Y(n_712) );
AOI211xp5_ASAP7_75t_L g713 ( .A1(n_699), .A2(n_695), .B(n_696), .C(n_681), .Y(n_713) );
NOR3xp33_ASAP7_75t_L g714 ( .A(n_708), .B(n_695), .C(n_689), .Y(n_714) );
AOI22xp5_ASAP7_75t_L g715 ( .A1(n_702), .A2(n_687), .B1(n_678), .B2(n_675), .Y(n_715) );
NOR2xp33_ASAP7_75t_L g716 ( .A(n_705), .B(n_697), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_703), .B(n_704), .Y(n_717) );
NAND2xp5_ASAP7_75t_SL g718 ( .A(n_701), .B(n_692), .Y(n_718) );
AND2x4_ASAP7_75t_L g719 ( .A(n_718), .B(n_685), .Y(n_719) );
NAND5xp2_ASAP7_75t_L g720 ( .A(n_717), .B(n_711), .C(n_710), .D(n_700), .E(n_706), .Y(n_720) );
NAND5xp2_ASAP7_75t_L g721 ( .A(n_712), .B(n_707), .C(n_709), .D(n_693), .E(n_75), .Y(n_721) );
AOI211x1_ASAP7_75t_L g722 ( .A1(n_715), .A2(n_68), .B(n_69), .C(n_71), .Y(n_722) );
AND4x1_ASAP7_75t_L g723 ( .A(n_720), .B(n_713), .C(n_716), .D(n_714), .Y(n_723) );
NOR3x1_ASAP7_75t_L g724 ( .A(n_721), .B(n_76), .C(n_77), .Y(n_724) );
XNOR2xp5_ASAP7_75t_L g725 ( .A(n_719), .B(n_78), .Y(n_725) );
AND2x4_ASAP7_75t_L g726 ( .A(n_723), .B(n_719), .Y(n_726) );
AO221x2_ASAP7_75t_L g727 ( .A1(n_724), .A2(n_722), .B1(n_82), .B2(n_83), .C(n_84), .Y(n_727) );
OAI22xp5_ASAP7_75t_L g728 ( .A1(n_726), .A2(n_725), .B1(n_86), .B2(n_89), .Y(n_728) );
INVx1_ASAP7_75t_L g729 ( .A(n_727), .Y(n_729) );
OAI22xp5_ASAP7_75t_L g730 ( .A1(n_729), .A2(n_81), .B1(n_91), .B2(n_92), .Y(n_730) );
OAI21xp33_ASAP7_75t_L g731 ( .A1(n_728), .A2(n_93), .B(n_94), .Y(n_731) );
AOI22xp5_ASAP7_75t_L g732 ( .A1(n_731), .A2(n_95), .B1(n_96), .B2(n_97), .Y(n_732) );
AO21x2_ASAP7_75t_L g733 ( .A1(n_732), .A2(n_730), .B(n_100), .Y(n_733) );
AOI22xp5_ASAP7_75t_L g734 ( .A1(n_733), .A2(n_98), .B1(n_102), .B2(n_106), .Y(n_734) );
endmodule