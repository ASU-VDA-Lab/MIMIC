module fake_jpeg_7130_n_241 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_241);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_241;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

INVx13_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_34),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g35 ( 
.A(n_23),
.B(n_0),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_35),
.B(n_41),
.Y(n_85)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_36),
.A2(n_31),
.B1(n_16),
.B2(n_17),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_40),
.Y(n_62)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_15),
.B(n_1),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_48),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_15),
.B(n_1),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_49),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_46),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_23),
.Y(n_49)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_51),
.B(n_70),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_32),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_53),
.B(n_30),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_55),
.Y(n_118)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_56),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_58),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_59),
.Y(n_104)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_61),
.Y(n_103)
);

INVx3_ASAP7_75t_SL g63 ( 
.A(n_45),
.Y(n_63)
);

INVxp33_ASAP7_75t_L g101 ( 
.A(n_63),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_40),
.A2(n_31),
.B1(n_32),
.B2(n_29),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_66),
.A2(n_65),
.B1(n_63),
.B2(n_60),
.Y(n_113)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_68),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_38),
.A2(n_31),
.B1(n_25),
.B2(n_29),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_69),
.A2(n_73),
.B1(n_75),
.B2(n_80),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_41),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_71),
.B(n_72),
.Y(n_110)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_34),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_38),
.A2(n_27),
.B1(n_26),
.B2(n_25),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_39),
.A2(n_36),
.B1(n_27),
.B2(n_26),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_74),
.A2(n_77),
.B1(n_30),
.B2(n_22),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_36),
.A2(n_28),
.B1(n_18),
.B2(n_17),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_76),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_45),
.A2(n_28),
.B1(n_18),
.B2(n_16),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_35),
.B(n_15),
.Y(n_78)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_78),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_SL g79 ( 
.A(n_47),
.Y(n_79)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_79),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_35),
.A2(n_30),
.B1(n_22),
.B2(n_19),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_37),
.B(n_2),
.Y(n_82)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_82),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_37),
.B(n_3),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_83),
.B(n_87),
.Y(n_107)
);

INVx2_ASAP7_75t_SL g86 ( 
.A(n_37),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_86),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_43),
.B(n_3),
.Y(n_87)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_43),
.Y(n_88)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_88),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_89),
.A2(n_22),
.B1(n_5),
.B2(n_7),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_35),
.B(n_4),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_90),
.B(n_91),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_94),
.B(n_99),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_85),
.B(n_30),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_105),
.Y(n_123)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_96),
.Y(n_120)
);

A2O1A1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_85),
.A2(n_64),
.B(n_53),
.C(n_80),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_75),
.B(n_30),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_69),
.A2(n_22),
.B1(n_5),
.B2(n_6),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_106),
.A2(n_111),
.B1(n_4),
.B2(n_9),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g108 ( 
.A(n_73),
.B(n_84),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_108),
.B(n_4),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_74),
.A2(n_22),
.B1(n_5),
.B2(n_7),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_113),
.A2(n_65),
.B1(n_60),
.B2(n_57),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_117),
.Y(n_122)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_110),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_121),
.B(n_127),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_112),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_124),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_105),
.A2(n_62),
.B(n_67),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_125),
.A2(n_132),
.B(n_141),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_112),
.B(n_61),
.Y(n_126)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_126),
.Y(n_167)
);

BUFx2_ASAP7_75t_L g127 ( 
.A(n_115),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_98),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_128),
.B(n_131),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_95),
.B(n_55),
.C(n_86),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_129),
.B(n_54),
.C(n_118),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_101),
.B(n_68),
.Y(n_130)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_130),
.Y(n_169)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_111),
.Y(n_131)
);

AND2x4_ASAP7_75t_L g132 ( 
.A(n_108),
.B(n_79),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_97),
.B(n_56),
.Y(n_133)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_133),
.Y(n_156)
);

NOR3xp33_ASAP7_75t_SL g135 ( 
.A(n_99),
.B(n_77),
.C(n_81),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_135),
.B(n_146),
.Y(n_154)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_94),
.B(n_59),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_136),
.B(n_140),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_97),
.B(n_81),
.Y(n_137)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_137),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_138),
.A2(n_145),
.B1(n_115),
.B2(n_102),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_SL g139 ( 
.A(n_92),
.B(n_55),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_139),
.B(n_123),
.Y(n_168)
);

OAI21xp33_ASAP7_75t_SL g141 ( 
.A1(n_93),
.A2(n_91),
.B(n_50),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_109),
.A2(n_91),
.B1(n_7),
.B2(n_8),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_142),
.Y(n_161)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_96),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_143),
.B(n_144),
.Y(n_150)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_94),
.Y(n_144)
);

AND2x2_ASAP7_75t_SL g146 ( 
.A(n_109),
.B(n_52),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_114),
.B(n_9),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_147),
.B(n_114),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_134),
.A2(n_104),
.B(n_92),
.Y(n_149)
);

AOI221xp5_ASAP7_75t_L g179 ( 
.A1(n_149),
.A2(n_132),
.B1(n_140),
.B2(n_135),
.C(n_145),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_152),
.B(n_164),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_131),
.A2(n_104),
.B1(n_106),
.B2(n_100),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_155),
.B(n_168),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_132),
.A2(n_116),
.B1(n_103),
.B2(n_119),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_157),
.A2(n_171),
.B1(n_122),
.B2(n_136),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_128),
.B(n_147),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_158),
.B(n_170),
.Y(n_187)
);

MAJx2_ASAP7_75t_L g162 ( 
.A(n_139),
.B(n_107),
.C(n_119),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_162),
.B(n_172),
.C(n_124),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_120),
.A2(n_116),
.B1(n_103),
.B2(n_102),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_163),
.A2(n_166),
.B1(n_143),
.B2(n_120),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_123),
.B(n_125),
.Y(n_164)
);

AO22x1_ASAP7_75t_L g166 ( 
.A1(n_132),
.A2(n_57),
.B1(n_54),
.B2(n_89),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g170 ( 
.A(n_146),
.Y(n_170)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_163),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_173),
.B(n_178),
.Y(n_193)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_150),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_174),
.Y(n_194)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_175),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_177),
.A2(n_180),
.B1(n_188),
.B2(n_161),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_164),
.B(n_144),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_179),
.B(n_154),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_149),
.A2(n_129),
.B1(n_122),
.B2(n_146),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_160),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_181),
.B(n_182),
.Y(n_200)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_151),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_152),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_183),
.B(n_184),
.Y(n_198)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_171),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_185),
.B(n_165),
.C(n_172),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_166),
.A2(n_121),
.B1(n_127),
.B2(n_12),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_153),
.B(n_118),
.Y(n_189)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_189),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_168),
.B(n_10),
.Y(n_190)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_190),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_192),
.B(n_195),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_186),
.B(n_165),
.C(n_154),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_175),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_196),
.B(n_205),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_197),
.B(n_190),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_173),
.A2(n_166),
.B1(n_169),
.B2(n_155),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_199),
.A2(n_204),
.B1(n_184),
.B2(n_188),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_186),
.B(n_162),
.C(n_148),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_203),
.B(n_185),
.Y(n_215)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_187),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_198),
.A2(n_176),
.B(n_148),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_206),
.B(n_208),
.C(n_209),
.Y(n_218)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_207),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_198),
.A2(n_176),
.B(n_148),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_191),
.A2(n_183),
.B(n_182),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_211),
.B(n_215),
.C(n_203),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_193),
.B(n_178),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_212),
.B(n_214),
.Y(n_216)
);

NOR3xp33_ASAP7_75t_SL g214 ( 
.A(n_197),
.B(n_180),
.C(n_174),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_210),
.A2(n_196),
.B1(n_191),
.B2(n_204),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_219),
.B(n_221),
.Y(n_227)
);

MAJx2_ASAP7_75t_L g228 ( 
.A(n_220),
.B(n_202),
.C(n_159),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_212),
.B(n_181),
.Y(n_221)
);

XOR2x2_ASAP7_75t_L g222 ( 
.A(n_213),
.B(n_195),
.Y(n_222)
);

AOI21x1_ASAP7_75t_L g224 ( 
.A1(n_222),
.A2(n_220),
.B(n_223),
.Y(n_224)
);

A2O1A1Ixp33_ASAP7_75t_SL g223 ( 
.A1(n_215),
.A2(n_161),
.B(n_192),
.C(n_194),
.Y(n_223)
);

INVxp67_ASAP7_75t_SL g229 ( 
.A(n_223),
.Y(n_229)
);

AOI221xp5_ASAP7_75t_L g230 ( 
.A1(n_224),
.A2(n_226),
.B1(n_228),
.B2(n_216),
.C(n_223),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_218),
.B(n_201),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_225),
.B(n_159),
.Y(n_231)
);

OAI31xp33_ASAP7_75t_L g226 ( 
.A1(n_222),
.A2(n_200),
.A3(n_202),
.B(n_167),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_230),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_231),
.B(n_232),
.Y(n_235)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_227),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_229),
.B(n_156),
.Y(n_233)
);

OAI321xp33_ASAP7_75t_L g236 ( 
.A1(n_233),
.A2(n_234),
.A3(n_217),
.B1(n_11),
.B2(n_14),
.C(n_10),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_229),
.B(n_156),
.Y(n_234)
);

NAND3xp33_ASAP7_75t_L g238 ( 
.A(n_236),
.B(n_10),
.C(n_11),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_238),
.B(n_239),
.C(n_237),
.Y(n_240)
);

INVxp33_ASAP7_75t_SL g239 ( 
.A(n_235),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_240),
.B(n_232),
.Y(n_241)
);


endmodule