module fake_jpeg_13600_n_374 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_374);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_374;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_35),
.Y(n_84)
);

INVx6_ASAP7_75t_SL g36 ( 
.A(n_20),
.Y(n_36)
);

INVx5_ASAP7_75t_SL g72 ( 
.A(n_36),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_37),
.B(n_59),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_21),
.B(n_13),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_39),
.B(n_43),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx3_ASAP7_75t_SL g74 ( 
.A(n_40),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_21),
.B(n_13),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_20),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_44),
.B(n_58),
.Y(n_90)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

BUFx12_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_25),
.B(n_0),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_51),
.B(n_60),
.Y(n_81)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_53),
.Y(n_87)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_57),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_21),
.B(n_13),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_32),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_24),
.B(n_0),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_45),
.A2(n_34),
.B1(n_26),
.B2(n_29),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_63),
.A2(n_70),
.B1(n_89),
.B2(n_91),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_60),
.A2(n_24),
.B1(n_33),
.B2(n_17),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_64),
.A2(n_78),
.B1(n_82),
.B2(n_27),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_37),
.B(n_18),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_65),
.B(n_71),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_54),
.A2(n_34),
.B1(n_26),
.B2(n_30),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_18),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_42),
.A2(n_24),
.B1(n_33),
.B2(n_17),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_52),
.A2(n_17),
.B1(n_33),
.B2(n_18),
.Y(n_82)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_35),
.Y(n_88)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_88),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_55),
.A2(n_34),
.B1(n_26),
.B2(n_30),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_58),
.A2(n_34),
.B1(n_23),
.B2(n_30),
.Y(n_91)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_93),
.B(n_48),
.Y(n_97)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_35),
.Y(n_94)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_94),
.Y(n_125)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_38),
.Y(n_95)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_95),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_56),
.A2(n_30),
.B1(n_23),
.B2(n_32),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_96),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_97),
.Y(n_144)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_98),
.Y(n_137)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_69),
.Y(n_99)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_99),
.Y(n_143)
);

O2A1O1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_81),
.A2(n_36),
.B(n_49),
.C(n_51),
.Y(n_101)
);

A2O1A1Ixp33_ASAP7_75t_L g168 ( 
.A1(n_101),
.A2(n_46),
.B(n_22),
.C(n_50),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_75),
.B(n_16),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_102),
.B(n_103),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_62),
.B(n_59),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_16),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_104),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_62),
.B(n_48),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_105),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_84),
.Y(n_106)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_106),
.Y(n_148)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_61),
.Y(n_107)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_107),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_65),
.B(n_44),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_108),
.B(n_116),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_81),
.B(n_25),
.Y(n_109)
);

NOR3xp33_ASAP7_75t_L g139 ( 
.A(n_109),
.B(n_118),
.C(n_133),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_81),
.B(n_48),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_110),
.B(n_112),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_71),
.B(n_28),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_111),
.B(n_119),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_72),
.B(n_46),
.Y(n_112)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_87),
.Y(n_113)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_113),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_61),
.B(n_66),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_114),
.B(n_76),
.C(n_27),
.Y(n_156)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_72),
.B(n_28),
.Y(n_116)
);

INVx5_ASAP7_75t_SL g117 ( 
.A(n_83),
.Y(n_117)
);

INVx13_ASAP7_75t_L g142 ( 
.A(n_117),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_66),
.B(n_28),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_86),
.B(n_27),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_120),
.B(n_130),
.Y(n_141)
);

BUFx16f_ASAP7_75t_L g122 ( 
.A(n_83),
.Y(n_122)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_122),
.Y(n_145)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_87),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_123),
.Y(n_135)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_84),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_124),
.B(n_127),
.Y(n_164)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_73),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_126),
.B(n_129),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_76),
.B(n_46),
.Y(n_127)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_79),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_73),
.Y(n_130)
);

INVx11_ASAP7_75t_L g131 ( 
.A(n_68),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_131),
.Y(n_163)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_86),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_85),
.Y(n_134)
);

AOI21xp33_ASAP7_75t_L g153 ( 
.A1(n_134),
.A2(n_32),
.B(n_22),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_121),
.A2(n_95),
.B1(n_94),
.B2(n_88),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_136),
.A2(n_151),
.B1(n_152),
.B2(n_155),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_128),
.A2(n_89),
.B1(n_57),
.B2(n_47),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_147),
.A2(n_150),
.B1(n_154),
.B2(n_161),
.Y(n_172)
);

FAx1_ASAP7_75t_SL g149 ( 
.A(n_100),
.B(n_32),
.CI(n_77),
.CON(n_149),
.SN(n_149)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_149),
.B(n_116),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_128),
.A2(n_74),
.B1(n_67),
.B2(n_38),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_121),
.A2(n_67),
.B1(n_85),
.B2(n_77),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_101),
.A2(n_74),
.B1(n_40),
.B2(n_47),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_153),
.B(n_165),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_103),
.A2(n_108),
.B1(n_100),
.B2(n_111),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_119),
.A2(n_57),
.B1(n_41),
.B2(n_40),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_156),
.B(n_159),
.C(n_117),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_99),
.B(n_41),
.C(n_92),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_120),
.A2(n_23),
.B1(n_30),
.B2(n_68),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_98),
.A2(n_23),
.B1(n_79),
.B2(n_92),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_168),
.B(n_169),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_114),
.A2(n_50),
.B1(n_22),
.B2(n_19),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_170),
.B(n_169),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_154),
.B(n_116),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_173),
.B(n_176),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_147),
.A2(n_114),
.B1(n_107),
.B2(n_124),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_174),
.A2(n_142),
.B1(n_148),
.B2(n_3),
.Y(n_240)
);

OR2x2_ASAP7_75t_L g231 ( 
.A(n_175),
.B(n_182),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_138),
.B(n_122),
.Y(n_176)
);

BUFx24_ASAP7_75t_SL g177 ( 
.A(n_158),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_177),
.B(n_183),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_140),
.B(n_115),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_178),
.B(n_180),
.Y(n_212)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_145),
.Y(n_179)
);

INVx5_ASAP7_75t_L g210 ( 
.A(n_179),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_140),
.B(n_115),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_167),
.A2(n_117),
.B1(n_129),
.B2(n_123),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_181),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_158),
.B(n_113),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_135),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_137),
.Y(n_184)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_184),
.Y(n_216)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_137),
.Y(n_185)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_185),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_144),
.B(n_134),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_186),
.B(n_200),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_146),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_187),
.B(n_193),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_141),
.B(n_133),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_188),
.B(n_198),
.Y(n_214)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_143),
.Y(n_189)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_189),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_144),
.A2(n_130),
.B1(n_126),
.B2(n_131),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_190),
.Y(n_241)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_148),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_191),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_167),
.B(n_132),
.C(n_125),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_192),
.B(n_199),
.C(n_205),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_146),
.Y(n_193)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_143),
.Y(n_195)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_195),
.Y(n_232)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_166),
.Y(n_196)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_196),
.Y(n_238)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_166),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_197),
.B(n_157),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_141),
.B(n_132),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_162),
.B(n_125),
.C(n_106),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_160),
.B(n_164),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_160),
.B(n_106),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_202),
.B(n_203),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_145),
.B(n_122),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_156),
.B(n_19),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g235 ( 
.A(n_204),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_159),
.B(n_50),
.C(n_22),
.Y(n_205)
);

BUFx24_ASAP7_75t_SL g206 ( 
.A(n_149),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_206),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_149),
.B(n_1),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_207),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_194),
.A2(n_150),
.B1(n_161),
.B2(n_139),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_209),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_269)
);

AO21x1_ASAP7_75t_L g213 ( 
.A1(n_171),
.A2(n_168),
.B(n_152),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_213),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_178),
.B(n_163),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_217),
.B(n_222),
.Y(n_252)
);

AOI322xp5_ASAP7_75t_L g219 ( 
.A1(n_200),
.A2(n_175),
.A3(n_193),
.B1(n_187),
.B2(n_182),
.C1(n_172),
.C2(n_201),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_219),
.B(n_4),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_180),
.B(n_163),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_188),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_225),
.B(n_226),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_198),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_172),
.A2(n_155),
.B1(n_136),
.B2(n_165),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_227),
.A2(n_240),
.B1(n_201),
.B2(n_185),
.Y(n_243)
);

OAI21xp33_ASAP7_75t_L g230 ( 
.A1(n_171),
.A2(n_146),
.B(n_142),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_230),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_170),
.B(n_157),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_234),
.B(n_236),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_236),
.B(n_199),
.C(n_205),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_237),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_194),
.B(n_192),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_239),
.B(n_189),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_243),
.A2(n_251),
.B1(n_254),
.B2(n_258),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_244),
.B(n_256),
.C(n_261),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_217),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_245),
.B(n_259),
.Y(n_273)
);

OAI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_231),
.A2(n_174),
.B1(n_181),
.B2(n_194),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_247),
.A2(n_266),
.B1(n_269),
.B2(n_240),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_222),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_248),
.B(n_212),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_250),
.B(n_220),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_227),
.A2(n_184),
.B1(n_195),
.B2(n_183),
.Y(n_251)
);

AOI32xp33_ASAP7_75t_L g254 ( 
.A1(n_211),
.A2(n_197),
.A3(n_142),
.B1(n_196),
.B2(n_179),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_233),
.A2(n_191),
.B1(n_2),
.B2(n_3),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_255),
.A2(n_221),
.B(n_208),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_239),
.B(n_1),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_225),
.A2(n_12),
.B1(n_4),
.B2(n_5),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_226),
.B(n_3),
.Y(n_260)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_260),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_234),
.B(n_4),
.C(n_5),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_216),
.Y(n_262)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_262),
.Y(n_296)
);

NAND3xp33_ASAP7_75t_L g284 ( 
.A(n_263),
.B(n_215),
.C(n_228),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_220),
.B(n_4),
.C(n_5),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_264),
.B(n_238),
.C(n_224),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_214),
.B(n_6),
.Y(n_265)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_265),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_209),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_216),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_267),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_237),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_268),
.B(n_257),
.Y(n_291)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_223),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_270),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_SL g271 ( 
.A(n_229),
.B(n_7),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_271),
.B(n_223),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_249),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_272),
.B(n_289),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_257),
.A2(n_213),
.B1(n_212),
.B2(n_214),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_275),
.A2(n_252),
.B1(n_266),
.B2(n_260),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_276),
.B(n_280),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_253),
.A2(n_241),
.B1(n_233),
.B2(n_208),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_278),
.A2(n_286),
.B1(n_288),
.B2(n_255),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_259),
.B(n_231),
.Y(n_280)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_281),
.Y(n_305)
);

OR2x2_ASAP7_75t_L g283 ( 
.A(n_251),
.B(n_218),
.Y(n_283)
);

OAI22xp33_ASAP7_75t_SL g314 ( 
.A1(n_283),
.A2(n_262),
.B1(n_232),
.B2(n_238),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_284),
.B(n_287),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_243),
.A2(n_211),
.B1(n_213),
.B2(n_241),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_291),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_250),
.B(n_235),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_292),
.B(n_295),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_293),
.B(n_280),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_253),
.A2(n_237),
.B(n_224),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_294),
.A2(n_268),
.B(n_245),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_244),
.B(n_232),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g326 ( 
.A(n_298),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_299),
.A2(n_315),
.B(n_290),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_295),
.B(n_256),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_300),
.B(n_311),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_304),
.A2(n_308),
.B1(n_290),
.B2(n_288),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_276),
.B(n_264),
.C(n_261),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_306),
.B(n_282),
.C(n_289),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_283),
.A2(n_252),
.B1(n_265),
.B2(n_258),
.Y(n_307)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_307),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_277),
.A2(n_246),
.B1(n_270),
.B2(n_267),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_273),
.Y(n_309)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_309),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_291),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_312),
.B(n_316),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_292),
.B(n_271),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_313),
.B(n_293),
.Y(n_332)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_314),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_273),
.Y(n_315)
);

FAx1_ASAP7_75t_SL g316 ( 
.A(n_275),
.B(n_242),
.CI(n_210),
.CON(n_316),
.SN(n_316)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_317),
.B(n_274),
.C(n_297),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_299),
.A2(n_294),
.B(n_287),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_318),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_319),
.B(n_324),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_322),
.A2(n_327),
.B1(n_309),
.B2(n_315),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_SL g324 ( 
.A(n_302),
.B(n_282),
.Y(n_324)
);

CKINVDCx14_ASAP7_75t_R g327 ( 
.A(n_310),
.Y(n_327)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_305),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_329),
.B(n_330),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_302),
.B(n_279),
.C(n_285),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_303),
.B(n_279),
.C(n_285),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_331),
.B(n_313),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_332),
.B(n_300),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_335),
.B(n_343),
.Y(n_346)
);

BUFx24_ASAP7_75t_SL g336 ( 
.A(n_320),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_SL g351 ( 
.A(n_336),
.B(n_344),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_317),
.B(n_303),
.C(n_306),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_337),
.B(n_338),
.Y(n_355)
);

CKINVDCx16_ASAP7_75t_R g338 ( 
.A(n_318),
.Y(n_338)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_339),
.Y(n_349)
);

NAND4xp25_ASAP7_75t_SL g341 ( 
.A(n_319),
.B(n_210),
.C(n_305),
.D(n_308),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_341),
.B(n_342),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_330),
.B(n_301),
.C(n_304),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_324),
.B(n_328),
.C(n_331),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_345),
.B(n_328),
.C(n_332),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_334),
.A2(n_325),
.B1(n_326),
.B2(n_321),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_347),
.A2(n_274),
.B1(n_341),
.B2(n_316),
.Y(n_359)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_348),
.B(n_352),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_337),
.B(n_322),
.C(n_323),
.Y(n_350)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_350),
.A2(n_353),
.B(n_335),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_342),
.B(n_316),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_334),
.A2(n_340),
.B(n_333),
.Y(n_353)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_354),
.Y(n_357)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_357),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_SL g358 ( 
.A(n_355),
.B(n_333),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_358),
.B(n_346),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_359),
.B(n_352),
.Y(n_365)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_360),
.A2(n_361),
.B(n_362),
.Y(n_363)
);

OAI21x1_ASAP7_75t_L g361 ( 
.A1(n_351),
.A2(n_296),
.B(n_8),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_SL g362 ( 
.A1(n_348),
.A2(n_7),
.B(n_8),
.Y(n_362)
);

HB1xp67_ASAP7_75t_L g369 ( 
.A(n_364),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_365),
.B(n_366),
.C(n_367),
.Y(n_368)
);

AOI21xp5_ASAP7_75t_L g366 ( 
.A1(n_356),
.A2(n_346),
.B(n_350),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_368),
.B(n_363),
.C(n_349),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_370),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_371),
.B(n_369),
.C(n_9),
.Y(n_372)
);

AOI221xp5_ASAP7_75t_L g373 ( 
.A1(n_372),
.A2(n_9),
.B1(n_10),
.B2(n_272),
.C(n_327),
.Y(n_373)
);

OAI21x1_ASAP7_75t_SL g374 ( 
.A1(n_373),
.A2(n_9),
.B(n_10),
.Y(n_374)
);


endmodule