module fake_jpeg_19123_n_33 (n_3, n_2, n_1, n_0, n_4, n_5, n_33);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_33;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx12f_ASAP7_75t_L g6 ( 
.A(n_5),
.Y(n_6)
);

AND2x2_ASAP7_75t_SL g7 ( 
.A(n_5),
.B(n_2),
.Y(n_7)
);

NOR2xp33_ASAP7_75t_L g8 ( 
.A(n_2),
.B(n_0),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_0),
.B(n_3),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_SL g12 ( 
.A(n_8),
.B(n_1),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_12),
.B(n_17),
.Y(n_20)
);

A2O1A1Ixp33_ASAP7_75t_L g13 ( 
.A1(n_7),
.A2(n_1),
.B(n_2),
.C(n_3),
.Y(n_13)
);

OA21x2_ASAP7_75t_L g19 ( 
.A1(n_13),
.A2(n_14),
.B(n_15),
.Y(n_19)
);

AOI21xp33_ASAP7_75t_L g14 ( 
.A1(n_11),
.A2(n_1),
.B(n_3),
.Y(n_14)
);

AOI32xp33_ASAP7_75t_L g15 ( 
.A1(n_7),
.A2(n_4),
.A3(n_9),
.B1(n_6),
.B2(n_10),
.Y(n_15)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g17 ( 
.A(n_7),
.B(n_4),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_17),
.B(n_6),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_18),
.B(n_22),
.Y(n_25)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_21),
.Y(n_23)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_18),
.B(n_17),
.C(n_16),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_24),
.B(n_19),
.C(n_25),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_26),
.B(n_28),
.C(n_19),
.Y(n_30)
);

NOR4xp25_ASAP7_75t_L g28 ( 
.A(n_24),
.B(n_19),
.C(n_15),
.D(n_13),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_27),
.Y(n_29)
);

O2A1O1Ixp33_ASAP7_75t_SL g31 ( 
.A1(n_29),
.A2(n_30),
.B(n_20),
.C(n_12),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_31),
.B(n_6),
.Y(n_32)
);

OAI221xp5_ASAP7_75t_L g33 ( 
.A1(n_32),
.A2(n_9),
.B1(n_16),
.B2(n_10),
.C(n_4),
.Y(n_33)
);


endmodule