module fake_jpeg_20184_n_78 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_78);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_78;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_48;
wire n_35;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_4),
.B(n_18),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_17),
.B(n_21),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_5),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_3),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_15),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_48),
.Y(n_57)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx3_ASAP7_75t_SL g49 ( 
.A(n_27),
.Y(n_49)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_45),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_50),
.A2(n_51),
.B1(n_52),
.B2(n_53),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_33),
.A2(n_16),
.B1(n_28),
.B2(n_34),
.Y(n_51)
);

BUFx16f_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_22),
.B(n_35),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_30),
.B(n_36),
.Y(n_54)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_57),
.B(n_54),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_59),
.B(n_60),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_57),
.B(n_47),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_59),
.A2(n_56),
.B1(n_55),
.B2(n_39),
.Y(n_61)
);

AND2x6_ASAP7_75t_L g63 ( 
.A(n_61),
.B(n_56),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_63),
.B(n_61),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_SL g66 ( 
.A1(n_64),
.A2(n_26),
.B(n_40),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_63),
.B(n_62),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_65),
.B(n_52),
.C(n_42),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_66),
.B(n_67),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_66),
.A2(n_55),
.B1(n_29),
.B2(n_24),
.Y(n_68)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_68),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_69),
.B(n_31),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_71),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g73 ( 
.A1(n_70),
.A2(n_68),
.B(n_25),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g75 ( 
.A(n_73),
.B(n_40),
.Y(n_75)
);

AOI322xp5_ASAP7_75t_L g74 ( 
.A1(n_72),
.A2(n_23),
.A3(n_46),
.B1(n_38),
.B2(n_37),
.C1(n_44),
.C2(n_43),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_74),
.B(n_75),
.C(n_58),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_76),
.A2(n_43),
.B1(n_58),
.B2(n_49),
.Y(n_77)
);

FAx1_ASAP7_75t_SL g78 ( 
.A(n_77),
.B(n_32),
.CI(n_58),
.CON(n_78),
.SN(n_78)
);


endmodule