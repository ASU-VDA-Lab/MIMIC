module fake_jpeg_11772_n_179 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_179);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_179;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_11),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx4f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx16f_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_17),
.B(n_7),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_36),
.B(n_37),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_7),
.Y(n_37)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_8),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_39),
.B(n_47),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_42),
.Y(n_94)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

INVx6_ASAP7_75t_SL g44 ( 
.A(n_35),
.Y(n_44)
);

NAND2x1_ASAP7_75t_SL g73 ( 
.A(n_44),
.B(n_56),
.Y(n_73)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_14),
.B(n_0),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_46),
.B(n_60),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_14),
.B(n_9),
.Y(n_47)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_48),
.Y(n_89)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_16),
.B(n_9),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_50),
.B(n_51),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_16),
.B(n_10),
.Y(n_51)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

INVx3_ASAP7_75t_SL g53 ( 
.A(n_19),
.Y(n_53)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_53),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_20),
.B(n_4),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_54),
.B(n_57),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

INVxp67_ASAP7_75t_SL g56 ( 
.A(n_26),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_59),
.Y(n_77)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_18),
.A2(n_33),
.B1(n_27),
.B2(n_34),
.Y(n_61)
);

OA22x2_ASAP7_75t_L g99 ( 
.A1(n_61),
.A2(n_67),
.B1(n_69),
.B2(n_38),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_31),
.B(n_4),
.C(n_1),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_62),
.B(n_63),
.Y(n_92)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_27),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_63),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_15),
.B(n_1),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_64),
.B(n_65),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_20),
.B(n_33),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_25),
.B(n_2),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_66),
.B(n_69),
.Y(n_87)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_15),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_25),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_22),
.B(n_23),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_23),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_80),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_81),
.B(n_88),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_45),
.A2(n_24),
.B1(n_53),
.B2(n_55),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_83),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_61),
.B(n_24),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_92),
.B(n_74),
.Y(n_120)
);

AO22x2_ASAP7_75t_L g95 ( 
.A1(n_48),
.A2(n_40),
.B1(n_58),
.B2(n_52),
.Y(n_95)
);

AO22x1_ASAP7_75t_L g107 ( 
.A1(n_95),
.A2(n_98),
.B1(n_100),
.B2(n_73),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_57),
.B(n_69),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_101),
.Y(n_117)
);

A2O1A1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_56),
.A2(n_57),
.B(n_41),
.C(n_38),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_98),
.Y(n_116)
);

OR2x2_ASAP7_75t_SL g100 ( 
.A(n_41),
.B(n_63),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_65),
.B(n_64),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_65),
.B(n_64),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_102),
.B(n_84),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_71),
.A2(n_99),
.B1(n_77),
.B2(n_95),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_103),
.A2(n_104),
.B1(n_109),
.B2(n_116),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_99),
.A2(n_77),
.B1(n_95),
.B2(n_79),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_97),
.Y(n_105)
);

INVx2_ASAP7_75t_SL g133 ( 
.A(n_105),
.Y(n_133)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_82),
.Y(n_106)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_106),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_107),
.A2(n_116),
.B(n_103),
.Y(n_139)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_80),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_108),
.B(n_111),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_95),
.A2(n_72),
.B1(n_87),
.B2(n_82),
.Y(n_109)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_76),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_112),
.B(n_114),
.Y(n_142)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_76),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_86),
.B(n_93),
.C(n_100),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_115),
.B(n_120),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_75),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_118),
.B(n_123),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_119),
.B(n_121),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_85),
.B(n_75),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_89),
.A2(n_91),
.B1(n_90),
.B2(n_78),
.Y(n_122)
);

XNOR2x1_ASAP7_75t_L g136 ( 
.A(n_122),
.B(n_124),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_73),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_90),
.B(n_78),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_89),
.B(n_70),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_125),
.B(n_128),
.Y(n_132)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_70),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_92),
.B(n_71),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_124),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_135),
.B(n_138),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_117),
.B(n_128),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_139),
.A2(n_140),
.B(n_134),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_107),
.A2(n_116),
.B(n_104),
.Y(n_140)
);

HB1xp67_ASAP7_75t_L g143 ( 
.A(n_137),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_143),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_129),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_144),
.B(n_146),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_139),
.A2(n_115),
.B(n_113),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_130),
.B(n_110),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_147),
.B(n_151),
.Y(n_158)
);

A2O1A1O1Ixp25_ASAP7_75t_L g153 ( 
.A1(n_148),
.A2(n_149),
.B(n_131),
.C(n_141),
.D(n_136),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_132),
.A2(n_113),
.B(n_126),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_130),
.B(n_109),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_150),
.B(n_131),
.Y(n_159)
);

HB1xp67_ASAP7_75t_L g151 ( 
.A(n_137),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_140),
.A2(n_127),
.B(n_118),
.Y(n_152)
);

NAND2xp33_ASAP7_75t_SL g157 ( 
.A(n_152),
.B(n_122),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_153),
.B(n_156),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_144),
.A2(n_134),
.B1(n_135),
.B2(n_136),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_157),
.A2(n_152),
.B(n_150),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_159),
.B(n_158),
.C(n_147),
.Y(n_165)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_155),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_160),
.A2(n_161),
.B1(n_164),
.B2(n_133),
.Y(n_167)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_154),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_162),
.A2(n_165),
.B(n_159),
.Y(n_166)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_158),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_166),
.B(n_165),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_167),
.B(n_168),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_163),
.Y(n_168)
);

BUFx12f_ASAP7_75t_L g169 ( 
.A(n_162),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_169),
.B(n_145),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_171),
.A2(n_142),
.B(n_133),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_172),
.B(n_153),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_173),
.B(n_174),
.C(n_175),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_170),
.A2(n_141),
.B1(n_169),
.B2(n_157),
.Y(n_174)
);

BUFx24_ASAP7_75t_SL g177 ( 
.A(n_175),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_172),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_178),
.B(n_176),
.Y(n_179)
);


endmodule