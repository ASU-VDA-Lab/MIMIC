module real_aes_7722_n_271 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_271);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_271;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_285;
wire n_624;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_766;
wire n_329;
wire n_852;
wire n_857;
wire n_461;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_560;
wire n_660;
wire n_814;
wire n_594;
wire n_856;
wire n_767;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_815;
wire n_519;
wire n_638;
wire n_564;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_352;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_281;
wire n_496;
wire n_693;
wire n_468;
wire n_746;
wire n_284;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_671;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_807;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_848;
wire n_392;
wire n_562;
wire n_404;
wire n_288;
wire n_598;
wire n_756;
wire n_735;
wire n_713;
wire n_728;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_692;
wire n_544;
wire n_789;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_472;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_314;
wire n_283;
wire n_753;
wire n_741;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_456;
wire n_717;
wire n_359;
wire n_312;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_639;
wire n_546;
wire n_587;
wire n_811;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_836;
wire n_793;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_686;
wire n_279;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_652;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_804;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_842;
wire n_849;
wire n_475;
wire n_554;
wire n_855;
wire n_798;
wire n_797;
wire n_668;
wire n_862;
AOI22xp5_ASAP7_75t_SL g698 ( .A1(n_0), .A2(n_222), .B1(n_651), .B2(n_686), .Y(n_698) );
AOI22xp33_ASAP7_75t_L g680 ( .A1(n_1), .A2(n_257), .B1(n_681), .B2(n_682), .Y(n_680) );
CKINVDCx20_ASAP7_75t_R g837 ( .A(n_2), .Y(n_837) );
AOI22xp33_ASAP7_75t_L g343 ( .A1(n_3), .A2(n_233), .B1(n_344), .B2(n_347), .Y(n_343) );
AOI22xp33_ASAP7_75t_L g444 ( .A1(n_4), .A2(n_216), .B1(n_421), .B2(n_445), .Y(n_444) );
AOI22xp5_ASAP7_75t_L g470 ( .A1(n_5), .A2(n_108), .B1(n_314), .B2(n_471), .Y(n_470) );
AOI22xp33_ASAP7_75t_SL g473 ( .A1(n_6), .A2(n_21), .B1(n_474), .B2(n_475), .Y(n_473) );
AOI22xp5_ASAP7_75t_L g549 ( .A1(n_7), .A2(n_60), .B1(n_307), .B2(n_332), .Y(n_549) );
CKINVDCx20_ASAP7_75t_R g653 ( .A(n_8), .Y(n_653) );
AOI22xp33_ASAP7_75t_L g587 ( .A1(n_9), .A2(n_115), .B1(n_559), .B2(n_588), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g352 ( .A1(n_10), .A2(n_69), .B1(n_353), .B2(n_355), .Y(n_352) );
INVx1_ASAP7_75t_L g665 ( .A(n_11), .Y(n_665) );
CKINVDCx20_ASAP7_75t_R g657 ( .A(n_12), .Y(n_657) );
AOI22xp33_ASAP7_75t_L g380 ( .A1(n_13), .A2(n_117), .B1(n_381), .B2(n_382), .Y(n_380) );
AOI22xp33_ASAP7_75t_L g318 ( .A1(n_14), .A2(n_249), .B1(n_319), .B2(n_326), .Y(n_318) );
AOI22xp33_ASAP7_75t_L g805 ( .A1(n_15), .A2(n_158), .B1(n_337), .B2(n_679), .Y(n_805) );
AOI22xp5_ASAP7_75t_L g562 ( .A1(n_16), .A2(n_135), .B1(n_395), .B2(n_563), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_17), .A2(n_53), .B1(n_360), .B2(n_534), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g329 ( .A1(n_18), .A2(n_106), .B1(n_330), .B2(n_335), .Y(n_329) );
AOI22xp33_ASAP7_75t_SL g678 ( .A1(n_19), .A2(n_146), .B1(n_335), .B2(n_679), .Y(n_678) );
AOI22xp33_ASAP7_75t_L g844 ( .A1(n_20), .A2(n_165), .B1(n_384), .B2(n_692), .Y(n_844) );
AOI22xp33_ASAP7_75t_L g458 ( .A1(n_22), .A2(n_128), .B1(n_459), .B2(n_460), .Y(n_458) );
INVx1_ASAP7_75t_L g830 ( .A(n_23), .Y(n_830) );
CKINVDCx20_ASAP7_75t_R g505 ( .A(n_24), .Y(n_505) );
CKINVDCx20_ASAP7_75t_R g702 ( .A(n_25), .Y(n_702) );
CKINVDCx20_ASAP7_75t_R g649 ( .A(n_26), .Y(n_649) );
AOI22xp33_ASAP7_75t_SL g422 ( .A1(n_27), .A2(n_154), .B1(n_423), .B2(n_424), .Y(n_422) );
AOI22xp5_ASAP7_75t_L g536 ( .A1(n_28), .A2(n_261), .B1(n_427), .B2(n_442), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g835 ( .A1(n_29), .A2(n_223), .B1(n_314), .B2(n_553), .Y(n_835) );
CKINVDCx20_ASAP7_75t_R g642 ( .A(n_30), .Y(n_642) );
NAND2xp5_ASAP7_75t_SL g416 ( .A(n_31), .B(n_417), .Y(n_416) );
AO22x2_ASAP7_75t_L g293 ( .A1(n_32), .A2(n_83), .B1(n_294), .B2(n_295), .Y(n_293) );
INVx1_ASAP7_75t_L g823 ( .A(n_32), .Y(n_823) );
AOI22xp5_ASAP7_75t_L g626 ( .A1(n_33), .A2(n_133), .B1(n_399), .B2(n_449), .Y(n_626) );
AOI22xp33_ASAP7_75t_SL g706 ( .A1(n_34), .A2(n_199), .B1(n_404), .B2(n_475), .Y(n_706) );
AOI22xp5_ASAP7_75t_L g847 ( .A1(n_35), .A2(n_151), .B1(n_400), .B2(n_730), .Y(n_847) );
AOI22xp5_ASAP7_75t_L g761 ( .A1(n_36), .A2(n_149), .B1(n_429), .B2(n_561), .Y(n_761) );
AOI22xp5_ASAP7_75t_L g555 ( .A1(n_37), .A2(n_243), .B1(n_386), .B2(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g572 ( .A(n_38), .Y(n_572) );
CKINVDCx20_ASAP7_75t_R g574 ( .A(n_39), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g359 ( .A1(n_40), .A2(n_113), .B1(n_360), .B2(n_363), .Y(n_359) );
AOI222xp33_ASAP7_75t_L g462 ( .A1(n_41), .A2(n_181), .B1(n_236), .B2(n_402), .C1(n_463), .C2(n_464), .Y(n_462) );
CKINVDCx20_ASAP7_75t_R g582 ( .A(n_42), .Y(n_582) );
CKINVDCx20_ASAP7_75t_R g792 ( .A(n_43), .Y(n_792) );
CKINVDCx20_ASAP7_75t_R g859 ( .A(n_44), .Y(n_859) );
CKINVDCx20_ASAP7_75t_R g725 ( .A(n_45), .Y(n_725) );
INVx1_ASAP7_75t_L g551 ( .A(n_46), .Y(n_551) );
AOI22xp33_ASAP7_75t_SL g418 ( .A1(n_47), .A2(n_162), .B1(n_332), .B2(n_392), .Y(n_418) );
AO22x2_ASAP7_75t_L g297 ( .A1(n_48), .A2(n_86), .B1(n_294), .B2(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g824 ( .A(n_48), .Y(n_824) );
AOI22xp5_ASAP7_75t_L g639 ( .A1(n_49), .A2(n_123), .B1(n_315), .B2(n_338), .Y(n_639) );
INVx1_ASAP7_75t_L g610 ( .A(n_50), .Y(n_610) );
CKINVDCx20_ASAP7_75t_R g738 ( .A(n_51), .Y(n_738) );
AOI22xp33_ASAP7_75t_L g476 ( .A1(n_52), .A2(n_255), .B1(n_389), .B2(n_477), .Y(n_476) );
AOI22xp33_ASAP7_75t_L g699 ( .A1(n_54), .A2(n_148), .B1(n_397), .B2(n_561), .Y(n_699) );
CKINVDCx20_ASAP7_75t_R g580 ( .A(n_55), .Y(n_580) );
CKINVDCx20_ASAP7_75t_R g412 ( .A(n_56), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g675 ( .A1(n_57), .A2(n_240), .B1(n_464), .B2(n_676), .Y(n_675) );
AOI22xp33_ASAP7_75t_L g782 ( .A1(n_58), .A2(n_114), .B1(n_783), .B2(n_784), .Y(n_782) );
AOI222xp33_ASAP7_75t_L g401 ( .A1(n_59), .A2(n_175), .B1(n_244), .B2(n_402), .C1(n_404), .C2(n_405), .Y(n_401) );
AOI22xp5_ASAP7_75t_SL g696 ( .A1(n_61), .A2(n_142), .B1(n_429), .B2(n_448), .Y(n_696) );
AOI22xp33_ASAP7_75t_SL g846 ( .A1(n_62), .A2(n_241), .B1(n_360), .B2(n_556), .Y(n_846) );
AOI22xp5_ASAP7_75t_L g305 ( .A1(n_63), .A2(n_252), .B1(n_306), .B2(n_313), .Y(n_305) );
CKINVDCx20_ASAP7_75t_R g734 ( .A(n_64), .Y(n_734) );
CKINVDCx20_ASAP7_75t_R g747 ( .A(n_65), .Y(n_747) );
CKINVDCx20_ASAP7_75t_R g756 ( .A(n_66), .Y(n_756) );
AOI22xp33_ASAP7_75t_L g763 ( .A1(n_67), .A2(n_265), .B1(n_421), .B2(n_764), .Y(n_763) );
AOI22xp33_ASAP7_75t_L g732 ( .A1(n_68), .A2(n_182), .B1(n_370), .B2(n_423), .Y(n_732) );
AOI22xp33_ASAP7_75t_L g394 ( .A1(n_70), .A2(n_170), .B1(n_395), .B2(n_397), .Y(n_394) );
AOI22xp33_ASAP7_75t_SL g420 ( .A1(n_71), .A2(n_186), .B1(n_395), .B2(n_421), .Y(n_420) );
AOI22xp5_ASAP7_75t_SL g695 ( .A1(n_72), .A2(n_129), .B1(n_384), .B2(n_556), .Y(n_695) );
AOI22xp33_ASAP7_75t_L g707 ( .A1(n_73), .A2(n_211), .B1(n_327), .B2(n_477), .Y(n_707) );
CKINVDCx20_ASAP7_75t_R g752 ( .A(n_74), .Y(n_752) );
AO22x2_ASAP7_75t_L g743 ( .A1(n_75), .A2(n_744), .B1(n_767), .B2(n_768), .Y(n_743) );
CKINVDCx20_ASAP7_75t_R g768 ( .A(n_75), .Y(n_768) );
AOI22xp33_ASAP7_75t_L g762 ( .A1(n_76), .A2(n_219), .B1(n_399), .B2(n_424), .Y(n_762) );
AOI22xp33_ASAP7_75t_SL g798 ( .A1(n_77), .A2(n_150), .B1(n_799), .B2(n_800), .Y(n_798) );
CKINVDCx20_ASAP7_75t_R g718 ( .A(n_78), .Y(n_718) );
AOI211xp5_ASAP7_75t_L g716 ( .A1(n_79), .A2(n_576), .B(n_717), .C(n_723), .Y(n_716) );
AOI22xp33_ASAP7_75t_L g778 ( .A1(n_80), .A2(n_226), .B1(n_779), .B2(n_780), .Y(n_778) );
AOI22xp33_ASAP7_75t_L g480 ( .A1(n_81), .A2(n_136), .B1(n_381), .B2(n_427), .Y(n_480) );
INVx1_ASAP7_75t_L g564 ( .A(n_82), .Y(n_564) );
CKINVDCx20_ASAP7_75t_R g646 ( .A(n_84), .Y(n_646) );
AOI22xp33_ASAP7_75t_L g447 ( .A1(n_85), .A2(n_260), .B1(n_448), .B2(n_449), .Y(n_447) );
CKINVDCx20_ASAP7_75t_R g669 ( .A(n_87), .Y(n_669) );
AOI22xp33_ASAP7_75t_L g486 ( .A1(n_88), .A2(n_192), .B1(n_364), .B2(n_400), .Y(n_486) );
AOI22xp5_ASAP7_75t_L g491 ( .A1(n_89), .A2(n_492), .B1(n_537), .B2(n_538), .Y(n_491) );
INVx1_ASAP7_75t_L g537 ( .A(n_89), .Y(n_537) );
CKINVDCx20_ASAP7_75t_R g407 ( .A(n_90), .Y(n_407) );
INVx1_ASAP7_75t_L g279 ( .A(n_91), .Y(n_279) );
AOI22xp5_ASAP7_75t_L g286 ( .A1(n_92), .A2(n_287), .B1(n_372), .B2(n_373), .Y(n_286) );
INVx1_ASAP7_75t_L g373 ( .A(n_92), .Y(n_373) );
AOI22xp5_ASAP7_75t_SL g566 ( .A1(n_93), .A2(n_567), .B1(n_596), .B2(n_597), .Y(n_566) );
INVx1_ASAP7_75t_L g597 ( .A(n_93), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g452 ( .A1(n_94), .A2(n_250), .B1(n_453), .B2(n_456), .Y(n_452) );
AOI22xp5_ASAP7_75t_L g481 ( .A1(n_95), .A2(n_191), .B1(n_395), .B2(n_482), .Y(n_481) );
AOI22xp33_ASAP7_75t_L g729 ( .A1(n_96), .A2(n_194), .B1(n_563), .B2(n_730), .Y(n_729) );
CKINVDCx20_ASAP7_75t_R g786 ( .A(n_97), .Y(n_786) );
INVx1_ASAP7_75t_L g275 ( .A(n_98), .Y(n_275) );
AOI22xp33_ASAP7_75t_SL g413 ( .A1(n_99), .A2(n_134), .B1(n_315), .B2(n_404), .Y(n_413) );
AOI22xp33_ASAP7_75t_SL g484 ( .A1(n_100), .A2(n_155), .B1(n_367), .B2(n_485), .Y(n_484) );
CKINVDCx20_ASAP7_75t_R g517 ( .A(n_101), .Y(n_517) );
XOR2x2_ASAP7_75t_L g437 ( .A(n_102), .B(n_438), .Y(n_437) );
AOI22xp33_ASAP7_75t_SL g689 ( .A1(n_103), .A2(n_224), .B1(n_386), .B2(n_690), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_104), .B(n_389), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_105), .A2(n_213), .B1(n_526), .B2(n_528), .Y(n_525) );
INVx1_ASAP7_75t_L g641 ( .A(n_107), .Y(n_641) );
AOI22xp33_ASAP7_75t_L g390 ( .A1(n_109), .A2(n_141), .B1(n_391), .B2(n_392), .Y(n_390) );
CKINVDCx20_ASAP7_75t_R g708 ( .A(n_110), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g365 ( .A1(n_111), .A2(n_140), .B1(n_366), .B2(n_370), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_112), .B(n_804), .Y(n_803) );
AOI22xp33_ASAP7_75t_SL g685 ( .A1(n_116), .A2(n_210), .B1(n_586), .B2(n_686), .Y(n_685) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_118), .A2(n_193), .B1(n_534), .B2(n_535), .Y(n_533) );
INVx1_ASAP7_75t_L g666 ( .A(n_119), .Y(n_666) );
CKINVDCx20_ASAP7_75t_R g797 ( .A(n_120), .Y(n_797) );
NAND2xp5_ASAP7_75t_L g802 ( .A(n_121), .B(n_389), .Y(n_802) );
AOI22xp33_ASAP7_75t_L g461 ( .A1(n_122), .A2(n_225), .B1(n_330), .B2(n_337), .Y(n_461) );
AOI22xp33_ASAP7_75t_SL g623 ( .A1(n_124), .A2(n_264), .B1(n_482), .B2(n_594), .Y(n_623) );
AOI22xp5_ASAP7_75t_L g704 ( .A1(n_125), .A2(n_171), .B1(n_314), .B2(n_338), .Y(n_704) );
AOI22xp33_ASAP7_75t_L g722 ( .A1(n_126), .A2(n_201), .B1(n_335), .B2(n_679), .Y(n_722) );
CKINVDCx20_ASAP7_75t_R g508 ( .A(n_127), .Y(n_508) );
CKINVDCx20_ASAP7_75t_R g788 ( .A(n_130), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_131), .B(n_319), .Y(n_721) );
AND2x2_ASAP7_75t_L g278 ( .A(n_132), .B(n_279), .Y(n_278) );
INVx1_ASAP7_75t_L g618 ( .A(n_137), .Y(n_618) );
AOI22xp33_ASAP7_75t_SL g687 ( .A1(n_138), .A2(n_168), .B1(n_370), .B2(n_453), .Y(n_687) );
CKINVDCx20_ASAP7_75t_R g724 ( .A(n_139), .Y(n_724) );
AND2x6_ASAP7_75t_L g274 ( .A(n_143), .B(n_275), .Y(n_274) );
HB1xp67_ASAP7_75t_L g817 ( .A(n_143), .Y(n_817) );
AO22x2_ASAP7_75t_L g301 ( .A1(n_144), .A2(n_217), .B1(n_294), .B2(n_298), .Y(n_301) );
INVx1_ASAP7_75t_L g620 ( .A(n_145), .Y(n_620) );
CKINVDCx16_ASAP7_75t_R g714 ( .A(n_147), .Y(n_714) );
CKINVDCx20_ASAP7_75t_R g500 ( .A(n_152), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g383 ( .A1(n_153), .A2(n_190), .B1(n_384), .B2(n_386), .Y(n_383) );
CKINVDCx20_ASAP7_75t_R g644 ( .A(n_156), .Y(n_644) );
CKINVDCx20_ASAP7_75t_R g654 ( .A(n_157), .Y(n_654) );
CKINVDCx20_ASAP7_75t_R g495 ( .A(n_159), .Y(n_495) );
AOI22xp33_ASAP7_75t_SL g560 ( .A1(n_160), .A2(n_245), .B1(n_482), .B2(n_561), .Y(n_560) );
OA22x2_ASAP7_75t_L g604 ( .A1(n_161), .A2(n_605), .B1(n_606), .B2(n_607), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_161), .Y(n_605) );
CKINVDCx20_ASAP7_75t_R g513 ( .A(n_163), .Y(n_513) );
AOI22xp33_ASAP7_75t_SL g627 ( .A1(n_164), .A2(n_268), .B1(n_421), .B2(n_628), .Y(n_627) );
AOI22xp33_ASAP7_75t_L g577 ( .A1(n_166), .A2(n_174), .B1(n_306), .B2(n_578), .Y(n_577) );
CKINVDCx20_ASAP7_75t_R g487 ( .A(n_167), .Y(n_487) );
AOI22xp33_ASAP7_75t_L g585 ( .A1(n_169), .A2(n_204), .B1(n_347), .B2(n_586), .Y(n_585) );
AOI22xp33_ASAP7_75t_L g765 ( .A1(n_172), .A2(n_247), .B1(n_382), .B2(n_766), .Y(n_765) );
AOI22xp33_ASAP7_75t_SL g426 ( .A1(n_173), .A2(n_237), .B1(n_381), .B2(n_427), .Y(n_426) );
CKINVDCx20_ASAP7_75t_R g430 ( .A(n_176), .Y(n_430) );
AOI22xp33_ASAP7_75t_L g616 ( .A1(n_177), .A2(n_206), .B1(n_337), .B2(n_464), .Y(n_616) );
AO22x2_ASAP7_75t_L g303 ( .A1(n_178), .A2(n_234), .B1(n_294), .B2(n_295), .Y(n_303) );
AOI22xp33_ASAP7_75t_L g624 ( .A1(n_179), .A2(n_208), .B1(n_353), .B2(n_445), .Y(n_624) );
CKINVDCx20_ASAP7_75t_R g839 ( .A(n_180), .Y(n_839) );
AOI22xp33_ASAP7_75t_L g591 ( .A1(n_183), .A2(n_207), .B1(n_592), .B2(n_594), .Y(n_591) );
AOI22xp33_ASAP7_75t_L g753 ( .A1(n_184), .A2(n_239), .B1(n_405), .B2(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g740 ( .A(n_185), .Y(n_740) );
INVx1_ASAP7_75t_L g638 ( .A(n_187), .Y(n_638) );
CKINVDCx20_ASAP7_75t_R g794 ( .A(n_188), .Y(n_794) );
CKINVDCx20_ASAP7_75t_R g674 ( .A(n_189), .Y(n_674) );
AOI22xp5_ASAP7_75t_L g552 ( .A1(n_195), .A2(n_266), .B1(n_510), .B2(n_553), .Y(n_552) );
INVx1_ASAP7_75t_L g570 ( .A(n_196), .Y(n_570) );
INVx1_ASAP7_75t_L g662 ( .A(n_197), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_198), .B(n_459), .Y(n_547) );
AOI22xp33_ASAP7_75t_SL g428 ( .A1(n_200), .A2(n_238), .B1(n_384), .B2(n_429), .Y(n_428) );
NAND2xp5_ASAP7_75t_SL g650 ( .A(n_202), .B(n_651), .Y(n_650) );
CKINVDCx20_ASAP7_75t_R g304 ( .A(n_203), .Y(n_304) );
AOI22xp33_ASAP7_75t_L g398 ( .A1(n_205), .A2(n_235), .B1(n_399), .B2(n_400), .Y(n_398) );
AOI22xp33_ASAP7_75t_L g842 ( .A1(n_209), .A2(n_258), .B1(n_594), .B2(n_843), .Y(n_842) );
CKINVDCx20_ASAP7_75t_R g759 ( .A(n_212), .Y(n_759) );
CKINVDCx20_ASAP7_75t_R g736 ( .A(n_214), .Y(n_736) );
AOI22xp33_ASAP7_75t_SL g557 ( .A1(n_215), .A2(n_221), .B1(n_558), .B2(n_559), .Y(n_557) );
NOR2xp33_ASAP7_75t_L g821 ( .A(n_217), .B(n_822), .Y(n_821) );
NAND2xp5_ASAP7_75t_SL g415 ( .A(n_218), .B(n_389), .Y(n_415) );
INVx1_ASAP7_75t_L g615 ( .A(n_220), .Y(n_615) );
CKINVDCx20_ASAP7_75t_R g659 ( .A(n_227), .Y(n_659) );
AOI22xp33_ASAP7_75t_L g388 ( .A1(n_228), .A2(n_242), .B1(n_319), .B2(n_389), .Y(n_388) );
CKINVDCx20_ASAP7_75t_R g748 ( .A(n_229), .Y(n_748) );
AOI22xp5_ASAP7_75t_L g826 ( .A1(n_230), .A2(n_827), .B1(n_848), .B2(n_849), .Y(n_826) );
CKINVDCx20_ASAP7_75t_R g848 ( .A(n_230), .Y(n_848) );
OAI22xp5_ASAP7_75t_L g773 ( .A1(n_231), .A2(n_774), .B1(n_775), .B2(n_806), .Y(n_773) );
INVx1_ASAP7_75t_L g806 ( .A(n_231), .Y(n_806) );
INVx1_ASAP7_75t_L g612 ( .A(n_232), .Y(n_612) );
INVx1_ASAP7_75t_L g820 ( .A(n_234), .Y(n_820) );
AOI22xp33_ASAP7_75t_SL g691 ( .A1(n_246), .A2(n_270), .B1(n_594), .B2(n_692), .Y(n_691) );
CKINVDCx20_ASAP7_75t_R g834 ( .A(n_248), .Y(n_834) );
AOI22xp33_ASAP7_75t_L g440 ( .A1(n_251), .A2(n_256), .B1(n_441), .B2(n_442), .Y(n_440) );
CKINVDCx20_ASAP7_75t_R g511 ( .A(n_253), .Y(n_511) );
INVx1_ASAP7_75t_L g294 ( .A(n_254), .Y(n_294) );
INVx1_ASAP7_75t_L g296 ( .A(n_254), .Y(n_296) );
AOI211xp5_ASAP7_75t_L g271 ( .A1(n_259), .A2(n_272), .B(n_280), .C(n_825), .Y(n_271) );
INVx1_ASAP7_75t_L g832 ( .A(n_262), .Y(n_832) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_263), .A2(n_269), .B1(n_366), .B2(n_531), .Y(n_530) );
CKINVDCx20_ASAP7_75t_R g469 ( .A(n_267), .Y(n_469) );
INVx1_ASAP7_75t_SL g272 ( .A(n_273), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_274), .B(n_276), .Y(n_273) );
HB1xp67_ASAP7_75t_L g816 ( .A(n_275), .Y(n_816) );
OAI21xp5_ASAP7_75t_L g857 ( .A1(n_276), .A2(n_815), .B(n_858), .Y(n_857) );
CKINVDCx20_ASAP7_75t_R g276 ( .A(n_277), .Y(n_276) );
INVxp67_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
AOI221xp5_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_603), .B1(n_810), .B2(n_811), .C(n_812), .Y(n_280) );
INVx1_ASAP7_75t_L g810 ( .A(n_281), .Y(n_810) );
AOI22xp5_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_283), .B1(n_432), .B2(n_602), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AOI22xp5_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_285), .B1(n_374), .B2(n_375), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
HB1xp67_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
INVx2_ASAP7_75t_SL g372 ( .A(n_287), .Y(n_372) );
AND2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_341), .Y(n_287) );
NOR2xp33_ASAP7_75t_L g288 ( .A(n_289), .B(n_317), .Y(n_288) );
OAI21xp5_ASAP7_75t_SL g289 ( .A1(n_290), .A2(n_304), .B(n_305), .Y(n_289) );
OAI21xp5_ASAP7_75t_SL g411 ( .A1(n_290), .A2(n_412), .B(n_413), .Y(n_411) );
OAI21xp5_ASAP7_75t_L g468 ( .A1(n_290), .A2(n_469), .B(n_470), .Y(n_468) );
OAI21xp5_ASAP7_75t_L g550 ( .A1(n_290), .A2(n_551), .B(n_552), .Y(n_550) );
INVx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx4_ASAP7_75t_L g403 ( .A(n_291), .Y(n_403) );
BUFx6f_ASAP7_75t_L g507 ( .A(n_291), .Y(n_507) );
BUFx3_ASAP7_75t_L g576 ( .A(n_291), .Y(n_576) );
INVx2_ASAP7_75t_SL g645 ( .A(n_291), .Y(n_645) );
INVx2_ASAP7_75t_L g703 ( .A(n_291), .Y(n_703) );
AND2x6_ASAP7_75t_L g291 ( .A(n_292), .B(n_299), .Y(n_291) );
AND2x4_ASAP7_75t_L g338 ( .A(n_292), .B(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g521 ( .A(n_292), .Y(n_521) );
AND2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_297), .Y(n_292) );
AND2x2_ASAP7_75t_L g312 ( .A(n_293), .B(n_301), .Y(n_312) );
INVx2_ASAP7_75t_L g325 ( .A(n_293), .Y(n_325) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g298 ( .A(n_296), .Y(n_298) );
INVx2_ASAP7_75t_L g311 ( .A(n_297), .Y(n_311) );
OR2x2_ASAP7_75t_L g324 ( .A(n_297), .B(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g328 ( .A(n_297), .B(n_325), .Y(n_328) );
INVx1_ASAP7_75t_L g334 ( .A(n_297), .Y(n_334) );
AND2x6_ASAP7_75t_L g346 ( .A(n_299), .B(n_323), .Y(n_346) );
AND2x2_ASAP7_75t_L g354 ( .A(n_299), .B(n_351), .Y(n_354) );
AND2x4_ASAP7_75t_L g362 ( .A(n_299), .B(n_328), .Y(n_362) );
AND2x2_ASAP7_75t_L g299 ( .A(n_300), .B(n_302), .Y(n_299) );
AND2x2_ASAP7_75t_L g322 ( .A(n_300), .B(n_303), .Y(n_322) );
INVx2_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_301), .B(n_303), .Y(n_350) );
AND2x2_ASAP7_75t_L g357 ( .A(n_301), .B(n_340), .Y(n_357) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g310 ( .A(n_303), .Y(n_310) );
INVx1_ASAP7_75t_L g340 ( .A(n_303), .Y(n_340) );
BUFx6f_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g619 ( .A(n_307), .Y(n_619) );
BUFx6f_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
BUFx6f_ASAP7_75t_L g404 ( .A(n_308), .Y(n_404) );
BUFx6f_ASAP7_75t_L g463 ( .A(n_308), .Y(n_463) );
BUFx4f_ASAP7_75t_SL g474 ( .A(n_308), .Y(n_474) );
BUFx2_ASAP7_75t_L g754 ( .A(n_308), .Y(n_754) );
AND2x4_ASAP7_75t_L g308 ( .A(n_309), .B(n_312), .Y(n_308) );
AND2x2_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
INVx1_ASAP7_75t_L g316 ( .A(n_310), .Y(n_316) );
AND2x2_ASAP7_75t_L g351 ( .A(n_311), .B(n_325), .Y(n_351) );
INVx1_ASAP7_75t_L g516 ( .A(n_311), .Y(n_516) );
AND2x4_ASAP7_75t_L g315 ( .A(n_312), .B(n_316), .Y(n_315) );
AND2x4_ASAP7_75t_L g332 ( .A(n_312), .B(n_333), .Y(n_332) );
NAND2x1p5_ASAP7_75t_L g515 ( .A(n_312), .B(n_516), .Y(n_515) );
BUFx4f_ASAP7_75t_SL g313 ( .A(n_314), .Y(n_313) );
INVx2_ASAP7_75t_L g406 ( .A(n_314), .Y(n_406) );
BUFx12f_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
BUFx6f_ASAP7_75t_L g464 ( .A(n_315), .Y(n_464) );
BUFx6f_ASAP7_75t_L g510 ( .A(n_315), .Y(n_510) );
NAND2xp5_ASAP7_75t_SL g317 ( .A(n_318), .B(n_329), .Y(n_317) );
INVx2_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx2_ASAP7_75t_L g417 ( .A(n_320), .Y(n_417) );
INVx2_ASAP7_75t_L g459 ( .A(n_320), .Y(n_459) );
INVx5_ASAP7_75t_L g477 ( .A(n_320), .Y(n_477) );
INVx4_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
AND2x4_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
AND2x6_ASAP7_75t_L g327 ( .A(n_322), .B(n_328), .Y(n_327) );
AND2x4_ASAP7_75t_L g364 ( .A(n_322), .B(n_351), .Y(n_364) );
INVx1_ASAP7_75t_L g499 ( .A(n_322), .Y(n_499) );
NAND2x1p5_ASAP7_75t_L g502 ( .A(n_322), .B(n_328), .Y(n_502) );
INVx2_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
OR2x2_ASAP7_75t_L g498 ( .A(n_324), .B(n_499), .Y(n_498) );
BUFx2_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
BUFx4f_ASAP7_75t_L g389 ( .A(n_327), .Y(n_389) );
BUFx2_ASAP7_75t_L g460 ( .A(n_327), .Y(n_460) );
INVx1_ASAP7_75t_SL g683 ( .A(n_327), .Y(n_683) );
AND2x2_ASAP7_75t_L g369 ( .A(n_328), .B(n_357), .Y(n_369) );
NAND2xp5_ASAP7_75t_SL g660 ( .A(n_328), .B(n_357), .Y(n_660) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
BUFx2_ASAP7_75t_L g391 ( .A(n_332), .Y(n_391) );
BUFx3_ASAP7_75t_L g475 ( .A(n_332), .Y(n_475) );
BUFx2_ASAP7_75t_L g679 ( .A(n_332), .Y(n_679) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
OR2x6_ASAP7_75t_L g371 ( .A(n_334), .B(n_350), .Y(n_371) );
INVx2_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_SL g336 ( .A(n_337), .Y(n_336) );
BUFx6f_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
BUFx3_ASAP7_75t_L g392 ( .A(n_338), .Y(n_392) );
BUFx2_ASAP7_75t_SL g471 ( .A(n_338), .Y(n_471) );
BUFx2_ASAP7_75t_SL g553 ( .A(n_338), .Y(n_553) );
INVx1_ASAP7_75t_L g522 ( .A(n_339), .Y(n_522) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
NOR2xp33_ASAP7_75t_L g341 ( .A(n_342), .B(n_358), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_343), .B(n_352), .Y(n_342) );
INVx2_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx5_ASAP7_75t_SL g482 ( .A(n_345), .Y(n_482) );
NOR2xp33_ASAP7_75t_L g664 ( .A(n_345), .B(n_665), .Y(n_664) );
INVx2_ASAP7_75t_SL g766 ( .A(n_345), .Y(n_766) );
INVx11_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx11_ASAP7_75t_L g385 ( .A(n_346), .Y(n_385) );
BUFx2_ASAP7_75t_SL g347 ( .A(n_348), .Y(n_347) );
BUFx3_ASAP7_75t_L g382 ( .A(n_348), .Y(n_382) );
BUFx3_ASAP7_75t_L g427 ( .A(n_348), .Y(n_427) );
BUFx3_ASAP7_75t_L g445 ( .A(n_348), .Y(n_445) );
BUFx2_ASAP7_75t_L g563 ( .A(n_348), .Y(n_563) );
INVx1_ASAP7_75t_L g658 ( .A(n_348), .Y(n_658) );
BUFx3_ASAP7_75t_L g686 ( .A(n_348), .Y(n_686) );
BUFx2_ASAP7_75t_SL g843 ( .A(n_348), .Y(n_843) );
AND2x4_ASAP7_75t_L g348 ( .A(n_349), .B(n_351), .Y(n_348) );
AND2x2_ASAP7_75t_L g651 ( .A(n_349), .B(n_516), .Y(n_651) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g356 ( .A(n_351), .B(n_357), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_351), .B(n_357), .Y(n_663) );
INVx1_ASAP7_75t_L g793 ( .A(n_353), .Y(n_793) );
BUFx2_ASAP7_75t_SL g353 ( .A(n_354), .Y(n_353) );
INVx2_ASAP7_75t_L g396 ( .A(n_354), .Y(n_396) );
BUFx2_ASAP7_75t_SL g448 ( .A(n_354), .Y(n_448) );
BUFx6f_ASAP7_75t_L g527 ( .A(n_354), .Y(n_527) );
INVx1_ASAP7_75t_L g443 ( .A(n_355), .Y(n_443) );
BUFx3_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
BUFx3_ASAP7_75t_L g381 ( .A(n_356), .Y(n_381) );
BUFx3_ASAP7_75t_L g561 ( .A(n_356), .Y(n_561) );
BUFx3_ASAP7_75t_L g595 ( .A(n_356), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_359), .B(n_365), .Y(n_358) );
INVx2_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx2_ASAP7_75t_L g386 ( .A(n_361), .Y(n_386) );
INVx3_ASAP7_75t_L g485 ( .A(n_361), .Y(n_485) );
INVx2_ASAP7_75t_L g535 ( .A(n_361), .Y(n_535) );
OAI22xp5_ASAP7_75t_SL g652 ( .A1(n_361), .A2(n_396), .B1(n_653), .B2(n_654), .Y(n_652) );
OAI22xp5_ASAP7_75t_L g733 ( .A1(n_361), .A2(n_734), .B1(n_735), .B2(n_736), .Y(n_733) );
INVx6_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
BUFx3_ASAP7_75t_L g429 ( .A(n_362), .Y(n_429) );
BUFx3_ASAP7_75t_L g451 ( .A(n_362), .Y(n_451) );
BUFx3_ASAP7_75t_L g790 ( .A(n_362), .Y(n_790) );
INVx4_ASAP7_75t_L g731 ( .A(n_363), .Y(n_731) );
BUFx6f_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
BUFx3_ASAP7_75t_L g397 ( .A(n_364), .Y(n_397) );
BUFx3_ASAP7_75t_L g421 ( .A(n_364), .Y(n_421) );
INVx2_ASAP7_75t_L g529 ( .A(n_364), .Y(n_529) );
BUFx3_ASAP7_75t_L g558 ( .A(n_364), .Y(n_558) );
BUFx6f_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx5_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx2_ASAP7_75t_L g399 ( .A(n_368), .Y(n_399) );
INVx1_ASAP7_75t_L g423 ( .A(n_368), .Y(n_423) );
INVx4_ASAP7_75t_L g455 ( .A(n_368), .Y(n_455) );
INVx3_ASAP7_75t_L g556 ( .A(n_368), .Y(n_556) );
BUFx3_ASAP7_75t_L g589 ( .A(n_368), .Y(n_589) );
INVx8_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_SL g370 ( .A(n_371), .Y(n_370) );
INVx6_ASAP7_75t_SL g400 ( .A(n_371), .Y(n_400) );
INVx1_ASAP7_75t_SL g559 ( .A(n_371), .Y(n_559) );
INVx1_ASAP7_75t_L g628 ( .A(n_371), .Y(n_628) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AO22x2_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_377), .B1(n_408), .B2(n_431), .Y(n_375) );
INVx2_ASAP7_75t_SL g376 ( .A(n_377), .Y(n_376) );
XOR2x2_ASAP7_75t_L g377 ( .A(n_378), .B(n_407), .Y(n_377) );
NAND4xp75_ASAP7_75t_L g378 ( .A(n_379), .B(n_387), .C(n_393), .D(n_401), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_380), .B(n_383), .Y(n_379) );
INVx1_ASAP7_75t_L g735 ( .A(n_384), .Y(n_735) );
INVx3_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx4_ASAP7_75t_L g441 ( .A(n_385), .Y(n_441) );
INVx2_ASAP7_75t_SL g534 ( .A(n_385), .Y(n_534) );
INVx4_ASAP7_75t_L g690 ( .A(n_385), .Y(n_690) );
AND2x2_ASAP7_75t_SL g387 ( .A(n_388), .B(n_390), .Y(n_387) );
AND2x2_ASAP7_75t_L g393 ( .A(n_394), .B(n_398), .Y(n_393) );
INVx3_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx3_ASAP7_75t_L g764 ( .A(n_396), .Y(n_764) );
BUFx2_ASAP7_75t_L g424 ( .A(n_400), .Y(n_424) );
BUFx2_ASAP7_75t_L g456 ( .A(n_400), .Y(n_456) );
BUFx4f_ASAP7_75t_SL g531 ( .A(n_400), .Y(n_531) );
BUFx2_ASAP7_75t_L g784 ( .A(n_400), .Y(n_784) );
INVx4_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
OAI21xp5_ASAP7_75t_SL g796 ( .A1(n_403), .A2(n_797), .B(n_798), .Y(n_796) );
INVx4_ASAP7_75t_L g504 ( .A(n_404), .Y(n_504) );
BUFx2_ASAP7_75t_L g676 ( .A(n_404), .Y(n_676) );
INVx1_ASAP7_75t_L g726 ( .A(n_405), .Y(n_726) );
INVx3_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx4_ASAP7_75t_SL g431 ( .A(n_408), .Y(n_431) );
XOR2x2_ASAP7_75t_L g408 ( .A(n_409), .B(n_430), .Y(n_408) );
NAND3x1_ASAP7_75t_L g409 ( .A(n_410), .B(n_419), .C(n_425), .Y(n_409) );
NOR2xp33_ASAP7_75t_L g410 ( .A(n_411), .B(n_414), .Y(n_410) );
NAND3xp33_ASAP7_75t_L g414 ( .A(n_415), .B(n_416), .C(n_418), .Y(n_414) );
AND2x2_ASAP7_75t_L g419 ( .A(n_420), .B(n_422), .Y(n_419) );
AND2x2_ASAP7_75t_L g425 ( .A(n_426), .B(n_428), .Y(n_425) );
INVx1_ASAP7_75t_L g602 ( .A(n_432), .Y(n_602) );
AOI22xp5_ASAP7_75t_L g432 ( .A1(n_433), .A2(n_434), .B1(n_490), .B2(n_601), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
HB1xp67_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
AO22x1_ASAP7_75t_SL g436 ( .A1(n_437), .A2(n_465), .B1(n_488), .B2(n_489), .Y(n_436) );
INVx1_ASAP7_75t_L g488 ( .A(n_437), .Y(n_488) );
NAND4xp75_ASAP7_75t_L g438 ( .A(n_439), .B(n_446), .C(n_457), .D(n_462), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_440), .B(n_444), .Y(n_439) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx2_ASAP7_75t_L g781 ( .A(n_445), .Y(n_781) );
AND2x2_ASAP7_75t_L g446 ( .A(n_447), .B(n_452), .Y(n_446) );
INVx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx3_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx3_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
BUFx6f_ASAP7_75t_L g783 ( .A(n_455), .Y(n_783) );
AND2x2_ASAP7_75t_SL g457 ( .A(n_458), .B(n_461), .Y(n_457) );
BUFx4f_ASAP7_75t_L g800 ( .A(n_464), .Y(n_800) );
INVx3_ASAP7_75t_SL g489 ( .A(n_465), .Y(n_489) );
AOI22xp5_ASAP7_75t_L g539 ( .A1(n_465), .A2(n_489), .B1(n_540), .B2(n_598), .Y(n_539) );
XOR2x2_ASAP7_75t_L g465 ( .A(n_466), .B(n_487), .Y(n_465) );
NAND2xp5_ASAP7_75t_SL g466 ( .A(n_467), .B(n_478), .Y(n_466) );
NOR2xp33_ASAP7_75t_L g467 ( .A(n_468), .B(n_472), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_473), .B(n_476), .Y(n_472) );
INVx1_ASAP7_75t_L g838 ( .A(n_474), .Y(n_838) );
BUFx6f_ASAP7_75t_L g681 ( .A(n_477), .Y(n_681) );
HB1xp67_ASAP7_75t_L g804 ( .A(n_477), .Y(n_804) );
NOR2xp33_ASAP7_75t_L g478 ( .A(n_479), .B(n_483), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_480), .B(n_481), .Y(n_479) );
INVx1_ASAP7_75t_L g787 ( .A(n_482), .Y(n_787) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_484), .B(n_486), .Y(n_483) );
INVx1_ASAP7_75t_L g601 ( .A(n_490), .Y(n_601) );
AOI22xp5_ASAP7_75t_L g490 ( .A1(n_491), .A2(n_539), .B1(n_599), .B2(n_600), .Y(n_490) );
INVx1_ASAP7_75t_L g599 ( .A(n_491), .Y(n_599) );
INVx1_ASAP7_75t_L g538 ( .A(n_492), .Y(n_538) );
AND2x2_ASAP7_75t_L g492 ( .A(n_493), .B(n_523), .Y(n_492) );
NOR3xp33_ASAP7_75t_L g493 ( .A(n_494), .B(n_503), .C(n_512), .Y(n_493) );
OAI22xp5_ASAP7_75t_L g494 ( .A1(n_495), .A2(n_496), .B1(n_500), .B2(n_501), .Y(n_494) );
OAI22xp5_ASAP7_75t_L g746 ( .A1(n_496), .A2(n_747), .B1(n_748), .B2(n_749), .Y(n_746) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx2_ASAP7_75t_L g571 ( .A(n_497), .Y(n_571) );
INVx1_ASAP7_75t_SL g831 ( .A(n_497), .Y(n_831) );
INVx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
BUFx6f_ASAP7_75t_L g611 ( .A(n_498), .Y(n_611) );
OAI21xp5_ASAP7_75t_L g637 ( .A1(n_498), .A2(n_638), .B(n_639), .Y(n_637) );
OAI22xp5_ASAP7_75t_L g569 ( .A1(n_501), .A2(n_570), .B1(n_571), .B2(n_572), .Y(n_569) );
BUFx3_ASAP7_75t_L g613 ( .A(n_501), .Y(n_613) );
OAI22xp5_ASAP7_75t_L g640 ( .A1(n_501), .A2(n_515), .B1(n_641), .B2(n_642), .Y(n_640) );
INVx2_ASAP7_75t_L g720 ( .A(n_501), .Y(n_720) );
OAI22xp5_ASAP7_75t_L g829 ( .A1(n_501), .A2(n_830), .B1(n_831), .B2(n_832), .Y(n_829) );
BUFx3_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx1_ASAP7_75t_L g750 ( .A(n_502), .Y(n_750) );
OAI222xp33_ASAP7_75t_L g503 ( .A1(n_504), .A2(n_505), .B1(n_506), .B2(n_508), .C1(n_509), .C2(n_511), .Y(n_503) );
OAI22xp5_ASAP7_75t_L g643 ( .A1(n_504), .A2(n_644), .B1(n_645), .B2(n_646), .Y(n_643) );
INVx3_ASAP7_75t_L g799 ( .A(n_504), .Y(n_799) );
OAI21xp33_ASAP7_75t_L g614 ( .A1(n_506), .A2(n_615), .B(n_616), .Y(n_614) );
OAI21xp33_ASAP7_75t_L g833 ( .A1(n_506), .A2(n_834), .B(n_835), .Y(n_833) );
INVx2_ASAP7_75t_SL g506 ( .A(n_507), .Y(n_506) );
INVx2_ASAP7_75t_L g673 ( .A(n_507), .Y(n_673) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
BUFx3_ASAP7_75t_L g578 ( .A(n_510), .Y(n_578) );
OAI22xp5_ASAP7_75t_L g512 ( .A1(n_513), .A2(n_514), .B1(n_517), .B2(n_518), .Y(n_512) );
OAI22xp5_ASAP7_75t_L g836 ( .A1(n_514), .A2(n_837), .B1(n_838), .B2(n_839), .Y(n_836) );
HB1xp67_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
BUFx3_ASAP7_75t_L g581 ( .A(n_515), .Y(n_581) );
OAI22xp5_ASAP7_75t_L g617 ( .A1(n_515), .A2(n_618), .B1(n_619), .B2(n_620), .Y(n_617) );
INVx4_ASAP7_75t_L g758 ( .A(n_515), .Y(n_758) );
INVx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx2_ASAP7_75t_L g583 ( .A(n_519), .Y(n_583) );
CKINVDCx16_ASAP7_75t_R g519 ( .A(n_520), .Y(n_519) );
OAI22xp5_ASAP7_75t_L g755 ( .A1(n_520), .A2(n_756), .B1(n_757), .B2(n_759), .Y(n_755) );
OR2x6_ASAP7_75t_L g520 ( .A(n_521), .B(n_522), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g523 ( .A(n_524), .B(n_532), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_525), .B(n_530), .Y(n_524) );
BUFx3_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx3_ASAP7_75t_L g593 ( .A(n_527), .Y(n_593) );
BUFx6f_ASAP7_75t_L g692 ( .A(n_527), .Y(n_692) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx2_ASAP7_75t_L g586 ( .A(n_529), .Y(n_586) );
OAI21xp5_ASAP7_75t_SL g648 ( .A1(n_529), .A2(n_649), .B(n_650), .Y(n_648) );
NAND2xp5_ASAP7_75t_SL g532 ( .A(n_533), .B(n_536), .Y(n_532) );
INVx1_ASAP7_75t_L g600 ( .A(n_539), .Y(n_600) );
INVx1_ASAP7_75t_L g598 ( .A(n_540), .Y(n_598) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
OAI22xp5_ASAP7_75t_SL g541 ( .A1(n_542), .A2(n_543), .B1(n_565), .B2(n_566), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
XOR2x2_ASAP7_75t_L g543 ( .A(n_544), .B(n_564), .Y(n_543) );
NAND4xp75_ASAP7_75t_SL g544 ( .A(n_545), .B(n_554), .C(n_560), .D(n_562), .Y(n_544) );
NOR2xp67_ASAP7_75t_SL g545 ( .A(n_546), .B(n_550), .Y(n_545) );
NAND3xp33_ASAP7_75t_L g546 ( .A(n_547), .B(n_548), .C(n_549), .Y(n_546) );
AND2x2_ASAP7_75t_L g554 ( .A(n_555), .B(n_557), .Y(n_554) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx2_ASAP7_75t_SL g596 ( .A(n_567), .Y(n_596) );
AND2x2_ASAP7_75t_SL g567 ( .A(n_568), .B(n_584), .Y(n_567) );
NOR3xp33_ASAP7_75t_L g568 ( .A(n_569), .B(n_573), .C(n_579), .Y(n_568) );
OAI21xp33_ASAP7_75t_L g573 ( .A1(n_574), .A2(n_575), .B(n_577), .Y(n_573) );
OAI21xp33_ASAP7_75t_L g751 ( .A1(n_575), .A2(n_752), .B(n_753), .Y(n_751) );
INVx3_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
OAI22xp5_ASAP7_75t_L g579 ( .A1(n_580), .A2(n_581), .B1(n_582), .B2(n_583), .Y(n_579) );
AND4x1_ASAP7_75t_L g584 ( .A(n_585), .B(n_587), .C(n_590), .D(n_591), .Y(n_584) );
INVx3_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx2_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
BUFx4f_ASAP7_75t_SL g594 ( .A(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g811 ( .A(n_603), .Y(n_811) );
AOI22xp5_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_629), .B1(n_808), .B2(n_809), .Y(n_603) );
INVx1_ASAP7_75t_L g808 ( .A(n_604), .Y(n_808) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g607 ( .A(n_608), .B(n_621), .Y(n_607) );
NOR3xp33_ASAP7_75t_L g608 ( .A(n_609), .B(n_614), .C(n_617), .Y(n_608) );
OAI22xp5_ASAP7_75t_L g609 ( .A1(n_610), .A2(n_611), .B1(n_612), .B2(n_613), .Y(n_609) );
OAI22xp5_ASAP7_75t_L g723 ( .A1(n_619), .A2(n_724), .B1(n_725), .B2(n_726), .Y(n_723) );
NOR2xp33_ASAP7_75t_L g621 ( .A(n_622), .B(n_625), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_623), .B(n_624), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_626), .B(n_627), .Y(n_625) );
INVx1_ASAP7_75t_L g809 ( .A(n_629), .Y(n_809) );
AOI22xp5_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_709), .B1(n_710), .B2(n_807), .Y(n_629) );
INVx1_ASAP7_75t_SL g807 ( .A(n_630), .Y(n_807) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
XNOR2xp5_ASAP7_75t_L g632 ( .A(n_633), .B(n_667), .Y(n_632) );
BUFx2_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
XNOR2x1_ASAP7_75t_L g634 ( .A(n_635), .B(n_666), .Y(n_634) );
AND3x2_ASAP7_75t_L g635 ( .A(n_636), .B(n_647), .C(n_655), .Y(n_635) );
NOR3xp33_ASAP7_75t_L g636 ( .A(n_637), .B(n_640), .C(n_643), .Y(n_636) );
NOR2xp33_ASAP7_75t_L g647 ( .A(n_648), .B(n_652), .Y(n_647) );
NOR3xp33_ASAP7_75t_L g655 ( .A(n_656), .B(n_661), .C(n_664), .Y(n_655) );
OAI22xp5_ASAP7_75t_L g656 ( .A1(n_657), .A2(n_658), .B1(n_659), .B2(n_660), .Y(n_656) );
NOR2xp33_ASAP7_75t_L g661 ( .A(n_662), .B(n_663), .Y(n_661) );
INVx1_ASAP7_75t_L g742 ( .A(n_663), .Y(n_742) );
XOR2x2_ASAP7_75t_L g667 ( .A(n_668), .B(n_693), .Y(n_667) );
XNOR2xp5_ASAP7_75t_L g668 ( .A(n_669), .B(n_670), .Y(n_668) );
NAND3xp33_ASAP7_75t_L g670 ( .A(n_671), .B(n_684), .C(n_688), .Y(n_670) );
NOR2xp33_ASAP7_75t_L g671 ( .A(n_672), .B(n_677), .Y(n_671) );
OAI21xp5_ASAP7_75t_SL g672 ( .A1(n_673), .A2(n_674), .B(n_675), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_678), .B(n_680), .Y(n_677) );
INVx1_ASAP7_75t_SL g682 ( .A(n_683), .Y(n_682) );
AND2x2_ASAP7_75t_L g684 ( .A(n_685), .B(n_687), .Y(n_684) );
AND2x2_ASAP7_75t_L g688 ( .A(n_689), .B(n_691), .Y(n_688) );
INVx1_ASAP7_75t_SL g739 ( .A(n_692), .Y(n_739) );
XOR2x2_ASAP7_75t_L g693 ( .A(n_694), .B(n_708), .Y(n_693) );
NAND4xp75_ASAP7_75t_SL g694 ( .A(n_695), .B(n_696), .C(n_697), .D(n_700), .Y(n_694) );
AND2x2_ASAP7_75t_L g697 ( .A(n_698), .B(n_699), .Y(n_697) );
NOR2xp33_ASAP7_75t_L g700 ( .A(n_701), .B(n_705), .Y(n_700) );
OAI21xp5_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_703), .B(n_704), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_706), .B(n_707), .Y(n_705) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
XNOR2xp5_ASAP7_75t_SL g710 ( .A(n_711), .B(n_771), .Y(n_710) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
AOI22xp5_ASAP7_75t_L g712 ( .A1(n_713), .A2(n_743), .B1(n_769), .B2(n_770), .Y(n_712) );
INVx2_ASAP7_75t_L g769 ( .A(n_713), .Y(n_769) );
XNOR2xp5_ASAP7_75t_L g713 ( .A(n_714), .B(n_715), .Y(n_713) );
AND2x2_ASAP7_75t_L g715 ( .A(n_716), .B(n_727), .Y(n_715) );
OAI211xp5_ASAP7_75t_L g717 ( .A1(n_718), .A2(n_719), .B(n_721), .C(n_722), .Y(n_717) );
INVx2_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
NOR3xp33_ASAP7_75t_L g727 ( .A(n_728), .B(n_733), .C(n_737), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_729), .B(n_732), .Y(n_728) );
INVx3_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx4_ASAP7_75t_L g779 ( .A(n_731), .Y(n_779) );
OAI22xp5_ASAP7_75t_L g737 ( .A1(n_738), .A2(n_739), .B1(n_740), .B2(n_741), .Y(n_737) );
OAI22xp5_ASAP7_75t_L g791 ( .A1(n_741), .A2(n_792), .B1(n_793), .B2(n_794), .Y(n_791) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx2_ASAP7_75t_L g770 ( .A(n_743), .Y(n_770) );
XNOR2xp5_ASAP7_75t_L g772 ( .A(n_743), .B(n_773), .Y(n_772) );
INVx1_ASAP7_75t_SL g767 ( .A(n_744), .Y(n_767) );
AND2x2_ASAP7_75t_SL g744 ( .A(n_745), .B(n_760), .Y(n_744) );
NOR3xp33_ASAP7_75t_L g745 ( .A(n_746), .B(n_751), .C(n_755), .Y(n_745) );
INVx2_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx2_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
AND4x1_ASAP7_75t_L g760 ( .A(n_761), .B(n_762), .C(n_763), .D(n_765), .Y(n_760) );
HB1xp67_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
INVx1_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
AND2x2_ASAP7_75t_SL g775 ( .A(n_776), .B(n_795), .Y(n_775) );
NOR3xp33_ASAP7_75t_L g776 ( .A(n_777), .B(n_785), .C(n_791), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g777 ( .A(n_778), .B(n_782), .Y(n_777) );
INVx2_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
OAI22xp5_ASAP7_75t_L g785 ( .A1(n_786), .A2(n_787), .B1(n_788), .B2(n_789), .Y(n_785) );
INVx1_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
NOR2xp33_ASAP7_75t_L g795 ( .A(n_796), .B(n_801), .Y(n_795) );
NAND3xp33_ASAP7_75t_L g801 ( .A(n_802), .B(n_803), .C(n_805), .Y(n_801) );
INVx2_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
NOR2x1_ASAP7_75t_L g813 ( .A(n_814), .B(n_818), .Y(n_813) );
OR2x2_ASAP7_75t_SL g863 ( .A(n_814), .B(n_819), .Y(n_863) );
NAND2xp5_ASAP7_75t_L g814 ( .A(n_815), .B(n_817), .Y(n_814) );
CKINVDCx20_ASAP7_75t_R g851 ( .A(n_815), .Y(n_851) );
INVx1_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
NAND2xp5_ASAP7_75t_L g858 ( .A(n_816), .B(n_855), .Y(n_858) );
CKINVDCx16_ASAP7_75t_R g855 ( .A(n_817), .Y(n_855) );
CKINVDCx20_ASAP7_75t_R g818 ( .A(n_819), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g819 ( .A(n_820), .B(n_821), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g822 ( .A(n_823), .B(n_824), .Y(n_822) );
OAI322xp33_ASAP7_75t_L g825 ( .A1(n_826), .A2(n_850), .A3(n_852), .B1(n_856), .B2(n_859), .C1(n_860), .C2(n_861), .Y(n_825) );
INVx1_ASAP7_75t_L g849 ( .A(n_827), .Y(n_849) );
XNOR2x1_ASAP7_75t_L g860 ( .A(n_827), .B(n_859), .Y(n_860) );
AND2x2_ASAP7_75t_L g827 ( .A(n_828), .B(n_840), .Y(n_827) );
NOR3xp33_ASAP7_75t_L g828 ( .A(n_829), .B(n_833), .C(n_836), .Y(n_828) );
NOR2xp33_ASAP7_75t_L g840 ( .A(n_841), .B(n_845), .Y(n_840) );
NAND2xp5_ASAP7_75t_L g841 ( .A(n_842), .B(n_844), .Y(n_841) );
NAND2xp5_ASAP7_75t_L g845 ( .A(n_846), .B(n_847), .Y(n_845) );
HB1xp67_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
HB1xp67_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
HB1xp67_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
INVx1_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
CKINVDCx16_ASAP7_75t_R g856 ( .A(n_857), .Y(n_856) );
CKINVDCx20_ASAP7_75t_R g861 ( .A(n_862), .Y(n_861) );
CKINVDCx20_ASAP7_75t_R g862 ( .A(n_863), .Y(n_862) );
endmodule