module fake_jpeg_17506_n_390 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_390);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_390;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_1),
.Y(n_14)
);

INVx4_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_3),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_2),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_38),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_39),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_40),
.Y(n_87)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_41),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_30),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_42),
.B(n_46),
.Y(n_90)
);

AOI21xp33_ASAP7_75t_L g43 ( 
.A1(n_22),
.A2(n_7),
.B(n_12),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_43),
.B(n_53),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_22),
.B(n_27),
.Y(n_47)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_48),
.B(n_50),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_49),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g50 ( 
.A(n_26),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_16),
.B(n_7),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

BUFx4f_ASAP7_75t_SL g96 ( 
.A(n_54),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_55),
.Y(n_97)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_56),
.Y(n_120)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_57),
.B(n_59),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_27),
.B(n_7),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_16),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_30),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_60),
.Y(n_101)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_61),
.B(n_23),
.Y(n_109)
);

BUFx8_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g83 ( 
.A(n_62),
.Y(n_83)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_63),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_21),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_64),
.Y(n_82)
);

BUFx16f_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

CKINVDCx6p67_ASAP7_75t_R g92 ( 
.A(n_65),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_18),
.Y(n_66)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_66),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_18),
.Y(n_67)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_67),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_18),
.Y(n_68)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_68),
.Y(n_114)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_69),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_43),
.A2(n_31),
.B1(n_15),
.B2(n_25),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_70),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_72),
.B(n_76),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_56),
.A2(n_31),
.B1(n_15),
.B2(n_25),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_74),
.A2(n_75),
.B1(n_107),
.B2(n_115),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_48),
.A2(n_16),
.B1(n_34),
.B2(n_17),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_53),
.B(n_37),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_77),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_60),
.A2(n_37),
.B1(n_36),
.B2(n_14),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_80),
.A2(n_13),
.B1(n_12),
.B2(n_11),
.Y(n_137)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_85),
.Y(n_163)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_86),
.Y(n_160)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_67),
.Y(n_94)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_94),
.Y(n_129)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_95),
.B(n_102),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_42),
.B(n_59),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_99),
.B(n_105),
.Y(n_145)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_39),
.Y(n_100)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_100),
.Y(n_142)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_54),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_103),
.B(n_108),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_63),
.B(n_36),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_61),
.B(n_33),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_106),
.B(n_32),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_45),
.A2(n_34),
.B1(n_17),
.B2(n_14),
.Y(n_107)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_64),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_109),
.B(n_119),
.Y(n_140)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_64),
.Y(n_111)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_111),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_57),
.A2(n_17),
.B1(n_34),
.B2(n_33),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_64),
.Y(n_116)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_116),
.Y(n_127)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_41),
.Y(n_117)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_117),
.Y(n_151)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_40),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_118),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_49),
.B(n_23),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_79),
.B(n_19),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_121),
.B(n_124),
.Y(n_175)
);

INVx5_ASAP7_75t_SL g123 ( 
.A(n_92),
.Y(n_123)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_123),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_79),
.B(n_90),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_81),
.Y(n_125)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_125),
.Y(n_185)
);

BUFx12f_ASAP7_75t_L g126 ( 
.A(n_81),
.Y(n_126)
);

BUFx24_ASAP7_75t_L g204 ( 
.A(n_126),
.Y(n_204)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_87),
.Y(n_132)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_132),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_98),
.B(n_19),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_133),
.B(n_143),
.Y(n_177)
);

AND2x2_ASAP7_75t_SL g135 ( 
.A(n_84),
.B(n_65),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_135),
.B(n_170),
.C(n_121),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_137),
.B(n_165),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_78),
.A2(n_65),
.B1(n_20),
.B2(n_13),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_138),
.A2(n_146),
.B(n_161),
.Y(n_194)
);

A2O1A1Ixp33_ASAP7_75t_L g139 ( 
.A1(n_93),
.A2(n_62),
.B(n_20),
.C(n_23),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_139),
.B(n_153),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_101),
.B(n_19),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_114),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_144),
.B(n_155),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_120),
.A2(n_62),
.B(n_32),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_96),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_147),
.B(n_148),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_89),
.B(n_23),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_87),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_149),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_104),
.B(n_19),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_150),
.B(n_167),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_74),
.A2(n_44),
.B1(n_51),
.B2(n_52),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_154),
.A2(n_5),
.B1(n_9),
.B2(n_8),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_113),
.B(n_23),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_83),
.B(n_62),
.Y(n_156)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_156),
.Y(n_195)
);

AO22x1_ASAP7_75t_L g157 ( 
.A1(n_78),
.A2(n_55),
.B1(n_29),
.B2(n_32),
.Y(n_157)
);

AO22x1_ASAP7_75t_SL g173 ( 
.A1(n_157),
.A2(n_88),
.B1(n_97),
.B2(n_91),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_88),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_158),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_83),
.A2(n_91),
.B1(n_111),
.B2(n_71),
.Y(n_161)
);

O2A1O1Ixp33_ASAP7_75t_L g162 ( 
.A1(n_115),
.A2(n_19),
.B(n_32),
.C(n_28),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_162),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_73),
.A2(n_7),
.B1(n_12),
.B2(n_10),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_164),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_192)
);

NAND2x1p5_ASAP7_75t_L g165 ( 
.A(n_75),
.B(n_29),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_77),
.B(n_29),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_166),
.B(n_168),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_96),
.B(n_29),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_82),
.B(n_29),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_96),
.B(n_29),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_169),
.B(n_103),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_82),
.B(n_28),
.C(n_5),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_172),
.B(n_157),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_173),
.A2(n_192),
.B1(n_208),
.B2(n_210),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_128),
.A2(n_112),
.B1(n_110),
.B2(n_85),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_176),
.A2(n_182),
.B1(n_184),
.B2(n_190),
.Y(n_217)
);

AOI32xp33_ASAP7_75t_L g179 ( 
.A1(n_128),
.A2(n_92),
.A3(n_86),
.B1(n_102),
.B2(n_95),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_179),
.B(n_194),
.Y(n_247)
);

NAND2xp33_ASAP7_75t_SL g180 ( 
.A(n_165),
.B(n_108),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_180),
.A2(n_203),
.B(n_130),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_181),
.B(n_183),
.Y(n_233)
);

NAND3xp33_ASAP7_75t_L g183 ( 
.A(n_124),
.B(n_92),
.C(n_5),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_141),
.A2(n_5),
.B1(n_9),
.B2(n_8),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_153),
.B(n_28),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_186),
.B(n_140),
.Y(n_216)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_151),
.Y(n_187)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_187),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_165),
.B(n_6),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_189),
.B(n_212),
.C(n_136),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_162),
.A2(n_6),
.B1(n_8),
.B2(n_2),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_135),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_193),
.A2(n_196),
.B1(n_202),
.B2(n_209),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_143),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g202 ( 
.A1(n_142),
.A2(n_4),
.B1(n_132),
.B2(n_129),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_146),
.A2(n_4),
.B(n_139),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_145),
.B(n_147),
.Y(n_205)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_205),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_152),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_206),
.B(n_211),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_164),
.A2(n_4),
.B1(n_137),
.B2(n_122),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_135),
.A2(n_4),
.B1(n_150),
.B2(n_152),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_122),
.A2(n_4),
.B1(n_166),
.B2(n_151),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_159),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_167),
.B(n_169),
.C(n_133),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_142),
.A2(n_129),
.B1(n_157),
.B2(n_170),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_213),
.A2(n_163),
.B1(n_134),
.B2(n_144),
.Y(n_230)
);

INVx13_ASAP7_75t_L g214 ( 
.A(n_123),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_214),
.B(n_160),
.Y(n_223)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_159),
.Y(n_215)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_215),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_216),
.B(n_232),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_178),
.B(n_145),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_218),
.B(n_234),
.Y(n_267)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_187),
.Y(n_219)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_219),
.Y(n_262)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_185),
.Y(n_220)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_220),
.Y(n_278)
);

INVx6_ASAP7_75t_L g222 ( 
.A(n_214),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_222),
.A2(n_227),
.B1(n_237),
.B2(n_249),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_223),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_191),
.B(n_127),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_226),
.B(n_236),
.Y(n_272)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_174),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_228),
.B(n_235),
.C(n_241),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_230),
.B(n_247),
.Y(n_256)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_204),
.Y(n_231)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_231),
.Y(n_280)
);

OR2x2_ASAP7_75t_L g232 ( 
.A(n_175),
.B(n_163),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_178),
.B(n_131),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_174),
.B(n_127),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_200),
.A2(n_134),
.B1(n_160),
.B2(n_125),
.Y(n_237)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_204),
.Y(n_239)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_239),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_215),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_240),
.B(n_243),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_172),
.B(n_126),
.C(n_149),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_181),
.Y(n_242)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_242),
.Y(n_286)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_188),
.Y(n_243)
);

HAxp5_ASAP7_75t_SL g261 ( 
.A(n_244),
.B(n_194),
.CON(n_261),
.SN(n_261)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_212),
.B(n_126),
.C(n_158),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_245),
.B(n_176),
.C(n_190),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_207),
.Y(n_246)
);

NOR3xp33_ASAP7_75t_L g268 ( 
.A(n_246),
.B(n_195),
.C(n_192),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_177),
.B(n_130),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_248),
.B(n_255),
.Y(n_270)
);

INVx1_ASAP7_75t_SL g249 ( 
.A(n_197),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_200),
.A2(n_126),
.B1(n_180),
.B2(n_197),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_250),
.A2(n_251),
.B1(n_171),
.B2(n_184),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_197),
.A2(n_208),
.B1(n_175),
.B2(n_177),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_201),
.B(n_206),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_252),
.Y(n_271)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_188),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_253),
.B(n_199),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_186),
.B(n_210),
.Y(n_255)
);

NAND3xp33_ASAP7_75t_SL g257 ( 
.A(n_251),
.B(n_209),
.C(n_203),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_257),
.B(n_268),
.Y(n_290)
);

OR2x2_ASAP7_75t_L g258 ( 
.A(n_242),
.B(n_211),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_258),
.B(n_263),
.Y(n_317)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_259),
.Y(n_296)
);

MAJx2_ASAP7_75t_L g260 ( 
.A(n_249),
.B(n_189),
.C(n_171),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_260),
.B(n_281),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_261),
.A2(n_230),
.B1(n_227),
.B2(n_238),
.Y(n_291)
);

OR2x2_ASAP7_75t_L g263 ( 
.A(n_255),
.B(n_193),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_264),
.A2(n_221),
.B1(n_243),
.B2(n_253),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_229),
.A2(n_182),
.B1(n_173),
.B2(n_179),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_265),
.A2(n_284),
.B1(n_217),
.B2(n_225),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_218),
.B(n_196),
.Y(n_269)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_269),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_234),
.B(n_248),
.Y(n_273)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_273),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_216),
.B(n_173),
.Y(n_275)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_275),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_276),
.B(n_279),
.C(n_287),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_228),
.B(n_204),
.C(n_198),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_224),
.B(n_173),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_232),
.B(n_198),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_282),
.B(n_267),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_229),
.A2(n_199),
.B1(n_185),
.B2(n_204),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_235),
.B(n_241),
.C(n_245),
.Y(n_287)
);

OAI32xp33_ASAP7_75t_L g289 ( 
.A1(n_247),
.A2(n_250),
.A3(n_244),
.B1(n_225),
.B2(n_217),
.Y(n_289)
);

XNOR2x2_ASAP7_75t_SL g306 ( 
.A(n_289),
.B(n_260),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_291),
.A2(n_306),
.B(n_315),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_292),
.A2(n_300),
.B1(n_302),
.B2(n_303),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_256),
.A2(n_233),
.B1(n_238),
.B2(n_254),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_294),
.A2(n_312),
.B1(n_315),
.B2(n_270),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_288),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_295),
.B(n_301),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_274),
.B(n_287),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_299),
.B(n_316),
.C(n_298),
.Y(n_335)
);

OAI22x1_ASAP7_75t_L g300 ( 
.A1(n_285),
.A2(n_222),
.B1(n_239),
.B2(n_231),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_288),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_256),
.A2(n_221),
.B1(n_220),
.B2(n_219),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_281),
.A2(n_275),
.B1(n_276),
.B2(n_271),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_304),
.A2(n_308),
.B1(n_266),
.B2(n_277),
.Y(n_325)
);

OA22x2_ASAP7_75t_L g308 ( 
.A1(n_284),
.A2(n_265),
.B1(n_282),
.B2(n_263),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_262),
.Y(n_309)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_309),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_262),
.Y(n_310)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_310),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_259),
.Y(n_311)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_311),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_264),
.A2(n_270),
.B1(n_289),
.B2(n_279),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_272),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_313),
.B(n_314),
.Y(n_326)
);

OAI22x1_ASAP7_75t_L g315 ( 
.A1(n_260),
.A2(n_258),
.B1(n_263),
.B2(n_266),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_274),
.B(n_267),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_318),
.B(n_321),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_307),
.A2(n_273),
.B1(n_286),
.B2(n_269),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_320),
.A2(n_323),
.B1(n_325),
.B2(n_331),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_316),
.B(n_272),
.Y(n_321)
);

INVx1_ASAP7_75t_SL g322 ( 
.A(n_291),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_322),
.A2(n_333),
.B1(n_317),
.B2(n_308),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_312),
.A2(n_286),
.B1(n_271),
.B2(n_258),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_296),
.Y(n_324)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_324),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_299),
.B(n_280),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_327),
.B(n_338),
.Y(n_346)
);

INVx3_ASAP7_75t_SL g330 ( 
.A(n_300),
.Y(n_330)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_330),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_293),
.A2(n_280),
.B1(n_283),
.B2(n_278),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_296),
.Y(n_332)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_332),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_302),
.A2(n_278),
.B1(n_283),
.B2(n_317),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g351 ( 
.A1(n_334),
.A2(n_290),
.B(n_308),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_335),
.B(n_339),
.C(n_294),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_298),
.B(n_305),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_305),
.B(n_314),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_319),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_340),
.B(n_353),
.Y(n_358)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_341),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_342),
.B(n_343),
.C(n_348),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_335),
.B(n_303),
.C(n_297),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_338),
.B(n_327),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_347),
.B(n_352),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_321),
.B(n_297),
.C(n_292),
.Y(n_348)
);

AOI32xp33_ASAP7_75t_L g366 ( 
.A1(n_351),
.A2(n_356),
.A3(n_355),
.B1(n_345),
.B2(n_352),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_339),
.B(n_306),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_326),
.B(n_308),
.C(n_313),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_326),
.B(n_318),
.C(n_324),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_354),
.B(n_356),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_325),
.B(n_334),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_L g357 ( 
.A1(n_351),
.A2(n_322),
.B(n_332),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_357),
.A2(n_368),
.B1(n_361),
.B2(n_366),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_344),
.B(n_329),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_359),
.B(n_358),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_349),
.A2(n_330),
.B1(n_336),
.B2(n_337),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_362),
.A2(n_363),
.B1(n_364),
.B2(n_346),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_353),
.A2(n_323),
.B1(n_333),
.B2(n_331),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_354),
.A2(n_320),
.B1(n_328),
.B2(n_348),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_366),
.B(n_346),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_343),
.A2(n_350),
.B1(n_345),
.B2(n_342),
.Y(n_368)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_369),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_370),
.B(n_371),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_368),
.B(n_347),
.Y(n_371)
);

OR2x2_ASAP7_75t_L g377 ( 
.A(n_372),
.B(n_373),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_SL g373 ( 
.A(n_359),
.B(n_364),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_360),
.B(n_367),
.C(n_363),
.Y(n_374)
);

OAI21xp33_ASAP7_75t_L g376 ( 
.A1(n_374),
.A2(n_375),
.B(n_361),
.Y(n_376)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_376),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_378),
.B(n_374),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_380),
.B(n_382),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_377),
.B(n_379),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_L g383 ( 
.A1(n_381),
.A2(n_376),
.B(n_370),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_383),
.B(n_369),
.C(n_371),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_385),
.Y(n_386)
);

NAND3xp33_ASAP7_75t_L g387 ( 
.A(n_386),
.B(n_384),
.C(n_380),
.Y(n_387)
);

AOI22xp33_ASAP7_75t_L g388 ( 
.A1(n_387),
.A2(n_360),
.B1(n_362),
.B2(n_357),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_SL g389 ( 
.A(n_388),
.B(n_365),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_389),
.B(n_365),
.Y(n_390)
);


endmodule