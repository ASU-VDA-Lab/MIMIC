module fake_jpeg_19270_n_330 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_330);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_330;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx14_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx24_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx6_ASAP7_75t_SL g39 ( 
.A(n_17),
.Y(n_39)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx4_ASAP7_75t_SL g41 ( 
.A(n_17),
.Y(n_41)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_47),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_33),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_53),
.B(n_57),
.Y(n_72)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_43),
.B(n_25),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_45),
.A2(n_31),
.B1(n_25),
.B2(n_33),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_60),
.A2(n_63),
.B1(n_41),
.B2(n_39),
.Y(n_73)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_41),
.A2(n_31),
.B1(n_29),
.B2(n_35),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_64),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_18),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_67),
.B(n_32),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_66),
.A2(n_31),
.B1(n_41),
.B2(n_39),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_68),
.A2(n_73),
.B1(n_87),
.B2(n_99),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_69),
.B(n_83),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g70 ( 
.A(n_66),
.Y(n_70)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_70),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_71),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_62),
.A2(n_41),
.B1(n_22),
.B2(n_37),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_75),
.A2(n_94),
.B1(n_98),
.B2(n_103),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_47),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_76),
.B(n_88),
.Y(n_126)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g132 ( 
.A(n_77),
.Y(n_132)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g137 ( 
.A(n_78),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_58),
.B(n_46),
.C(n_37),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_79),
.B(n_38),
.Y(n_122)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_80),
.Y(n_115)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_81),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_56),
.B(n_20),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_59),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_84),
.B(n_85),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_59),
.B(n_19),
.Y(n_85)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_86),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_50),
.A2(n_20),
.B1(n_18),
.B2(n_32),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_48),
.B(n_26),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_56),
.B(n_37),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_89),
.A2(n_91),
.B1(n_38),
.B2(n_42),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_65),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_90),
.B(n_92),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_48),
.B(n_46),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_62),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_93),
.B(n_100),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_50),
.A2(n_22),
.B1(n_36),
.B2(n_26),
.Y(n_94)
);

INVx2_ASAP7_75t_SL g96 ( 
.A(n_52),
.Y(n_96)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_96),
.Y(n_127)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_52),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_51),
.A2(n_39),
.B1(n_36),
.B2(n_16),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_51),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_53),
.B(n_19),
.Y(n_101)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_101),
.Y(n_128)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_47),
.Y(n_102)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_102),
.Y(n_129)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_67),
.Y(n_103)
);

INVxp33_ASAP7_75t_SL g104 ( 
.A(n_53),
.Y(n_104)
);

NOR2x1_ASAP7_75t_L g139 ( 
.A(n_104),
.B(n_27),
.Y(n_139)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_105),
.A2(n_107),
.B1(n_108),
.B2(n_23),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_52),
.Y(n_106)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_106),
.Y(n_110)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_49),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_47),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_69),
.A2(n_22),
.B1(n_35),
.B2(n_36),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_113),
.A2(n_124),
.B1(n_139),
.B2(n_96),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_72),
.A2(n_35),
.B1(n_30),
.B2(n_28),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_118),
.A2(n_119),
.B1(n_105),
.B2(n_98),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_91),
.A2(n_28),
.B1(n_30),
.B2(n_16),
.Y(n_119)
);

O2A1O1Ixp33_ASAP7_75t_SL g120 ( 
.A1(n_89),
.A2(n_38),
.B(n_42),
.C(n_44),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_120),
.A2(n_133),
.B(n_27),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_122),
.B(n_74),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_83),
.B(n_82),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_123),
.B(n_118),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_79),
.A2(n_38),
.B1(n_44),
.B2(n_42),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_89),
.A2(n_27),
.B(n_21),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_130),
.A2(n_133),
.B(n_120),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_131),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_91),
.A2(n_44),
.B(n_1),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_135),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_122),
.B(n_95),
.C(n_81),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_140),
.B(n_148),
.C(n_115),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_129),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_141),
.B(n_145),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_112),
.B(n_108),
.Y(n_142)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_142),
.Y(n_191)
);

O2A1O1Ixp33_ASAP7_75t_L g143 ( 
.A1(n_113),
.A2(n_86),
.B(n_80),
.C(n_107),
.Y(n_143)
);

O2A1O1Ixp33_ASAP7_75t_L g196 ( 
.A1(n_143),
.A2(n_0),
.B(n_1),
.C(n_3),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_144),
.A2(n_116),
.B1(n_134),
.B2(n_137),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_126),
.B(n_109),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_146),
.B(n_154),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_147),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_131),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_149),
.B(n_158),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_128),
.B(n_97),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_150),
.B(n_156),
.Y(n_181)
);

AND2x4_ASAP7_75t_L g151 ( 
.A(n_120),
.B(n_74),
.Y(n_151)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_151),
.Y(n_193)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_116),
.Y(n_152)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_152),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_139),
.A2(n_78),
.B1(n_77),
.B2(n_102),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_153),
.A2(n_134),
.B1(n_137),
.B2(n_71),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_123),
.B(n_97),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_129),
.Y(n_155)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_155),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_128),
.B(n_27),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_157),
.A2(n_169),
.B1(n_171),
.B2(n_143),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g158 ( 
.A(n_115),
.Y(n_158)
);

INVx5_ASAP7_75t_SL g159 ( 
.A(n_132),
.Y(n_159)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_159),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_160),
.A2(n_124),
.B(n_138),
.Y(n_173)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_110),
.Y(n_161)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_161),
.Y(n_199)
);

FAx1_ASAP7_75t_SL g162 ( 
.A(n_130),
.B(n_27),
.CI(n_24),
.CON(n_162),
.SN(n_162)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_162),
.B(n_163),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_139),
.B(n_24),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_163),
.B(n_165),
.Y(n_194)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_132),
.Y(n_164)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_164),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_121),
.A2(n_100),
.B1(n_24),
.B2(n_34),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_132),
.Y(n_166)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_166),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_114),
.A2(n_106),
.B1(n_34),
.B2(n_2),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_127),
.Y(n_170)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_170),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_114),
.A2(n_34),
.B1(n_1),
.B2(n_2),
.Y(n_171)
);

OA22x2_ASAP7_75t_L g172 ( 
.A1(n_151),
.A2(n_149),
.B1(n_144),
.B2(n_153),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_172),
.A2(n_173),
.B(n_180),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_170),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_174),
.B(n_197),
.Y(n_219)
);

AOI322xp5_ASAP7_75t_L g176 ( 
.A1(n_151),
.A2(n_125),
.A3(n_136),
.B1(n_111),
.B2(n_119),
.C1(n_127),
.C2(n_117),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_176),
.Y(n_212)
);

BUFx10_ASAP7_75t_L g179 ( 
.A(n_151),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_179),
.B(n_202),
.Y(n_230)
);

OA22x2_ASAP7_75t_L g180 ( 
.A1(n_160),
.A2(n_111),
.B1(n_110),
.B2(n_117),
.Y(n_180)
);

BUFx12f_ASAP7_75t_L g182 ( 
.A(n_152),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_182),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_183),
.B(n_10),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_184),
.A2(n_196),
.B(n_10),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_185),
.B(n_187),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_148),
.B(n_137),
.C(n_15),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_190),
.B(n_140),
.C(n_162),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_195),
.A2(n_165),
.B1(n_167),
.B2(n_147),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_166),
.Y(n_197)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_161),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_168),
.A2(n_146),
.B1(n_154),
.B2(n_167),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_203),
.B(n_204),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_168),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_207),
.B(n_194),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_189),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_208),
.B(n_181),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_210),
.A2(n_217),
.B1(n_218),
.B2(n_222),
.Y(n_247)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_175),
.Y(n_211)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_211),
.Y(n_233)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_201),
.Y(n_213)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_213),
.Y(n_237)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_192),
.Y(n_214)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_214),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_200),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_215),
.B(n_216),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_178),
.B(n_142),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_193),
.A2(n_157),
.B1(n_162),
.B2(n_158),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_193),
.A2(n_142),
.B1(n_159),
.B2(n_4),
.Y(n_218)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_187),
.Y(n_220)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_220),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_195),
.A2(n_173),
.B1(n_177),
.B2(n_178),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_177),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_223),
.A2(n_186),
.B1(n_172),
.B2(n_180),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_172),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_224),
.B(n_225),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_190),
.B(n_0),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_226),
.A2(n_228),
.B(n_196),
.Y(n_236)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_180),
.Y(n_227)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_227),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_180),
.A2(n_3),
.B(n_5),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_229),
.B(n_232),
.C(n_194),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_198),
.A2(n_202),
.B1(n_199),
.B2(n_191),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_231),
.A2(n_199),
.B1(n_198),
.B2(n_186),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_183),
.B(n_10),
.C(n_6),
.Y(n_232)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_235),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_236),
.A2(n_241),
.B(n_255),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_238),
.B(n_229),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_240),
.A2(n_205),
.B1(n_215),
.B2(n_224),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_221),
.A2(n_227),
.B(n_222),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_221),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_242),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_206),
.A2(n_188),
.B1(n_191),
.B2(n_172),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_245),
.A2(n_251),
.B1(n_205),
.B2(n_220),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_248),
.B(n_250),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_207),
.B(n_179),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_249),
.B(n_238),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_219),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_232),
.B(n_179),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_252),
.B(n_253),
.Y(n_263)
);

BUFx8_ASAP7_75t_L g253 ( 
.A(n_209),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_206),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_254),
.B(n_250),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_228),
.A2(n_179),
.B(n_182),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_256),
.B(n_259),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_257),
.A2(n_237),
.B1(n_243),
.B2(n_233),
.Y(n_279)
);

BUFx12f_ASAP7_75t_SL g260 ( 
.A(n_249),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_260),
.A2(n_269),
.B(n_9),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_248),
.B(n_210),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g282 ( 
.A(n_264),
.B(n_266),
.Y(n_282)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_265),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_247),
.B(n_216),
.Y(n_266)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_267),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_247),
.B(n_217),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_268),
.B(n_253),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_241),
.A2(n_226),
.B(n_230),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_251),
.A2(n_212),
.B1(n_218),
.B2(n_223),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_270),
.B(n_274),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_239),
.A2(n_208),
.B1(n_219),
.B2(n_225),
.Y(n_271)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_271),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_234),
.B(n_213),
.C(n_214),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_273),
.B(n_255),
.C(n_237),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_246),
.A2(n_244),
.B1(n_239),
.B2(n_234),
.Y(n_274)
);

FAx1_ASAP7_75t_SL g275 ( 
.A(n_236),
.B(n_211),
.CI(n_182),
.CON(n_275),
.SN(n_275)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_275),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_276),
.B(n_277),
.C(n_280),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_262),
.B(n_244),
.C(n_246),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_279),
.B(n_285),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_264),
.B(n_243),
.C(n_233),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_284),
.B(n_256),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_272),
.B(n_209),
.Y(n_285)
);

O2A1O1Ixp33_ASAP7_75t_L g288 ( 
.A1(n_261),
.A2(n_253),
.B(n_209),
.C(n_7),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_288),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_290),
.A2(n_269),
.B(n_261),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_273),
.B(n_5),
.C(n_6),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_291),
.B(n_263),
.C(n_275),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_291),
.B(n_258),
.Y(n_292)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_292),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_294),
.B(n_296),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_295),
.A2(n_283),
.B(n_267),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_280),
.B(n_260),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_297),
.B(n_298),
.Y(n_305)
);

HB1xp67_ASAP7_75t_L g298 ( 
.A(n_277),
.Y(n_298)
);

FAx1_ASAP7_75t_SL g300 ( 
.A(n_282),
.B(n_266),
.CI(n_268),
.CON(n_300),
.SN(n_300)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_300),
.B(n_286),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_276),
.B(n_259),
.C(n_274),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_301),
.B(n_287),
.C(n_281),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_282),
.B(n_270),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_303),
.B(n_284),
.C(n_289),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_307),
.B(n_309),
.C(n_293),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_302),
.A2(n_288),
.B(n_278),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_308),
.A2(n_312),
.B(n_299),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_297),
.B(n_279),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_310),
.B(n_311),
.Y(n_318)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_313),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_314),
.B(n_315),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_305),
.B(n_293),
.C(n_301),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_309),
.B(n_296),
.C(n_303),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_316),
.B(n_317),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_310),
.A2(n_304),
.B1(n_300),
.B2(n_306),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_318),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_319),
.B(n_300),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_306),
.C(n_294),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_323),
.B(n_324),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_325),
.Y(n_326)
);

NAND3xp33_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_320),
.C(n_321),
.Y(n_327)
);

BUFx24_ASAP7_75t_SL g328 ( 
.A(n_327),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_328),
.B(n_286),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_5),
.Y(n_330)
);


endmodule