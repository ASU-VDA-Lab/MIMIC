module real_jpeg_4488_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx8_ASAP7_75t_L g130 ( 
.A(n_0),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_1),
.A2(n_95),
.B1(n_96),
.B2(n_97),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_1),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_1),
.A2(n_95),
.B1(n_145),
.B2(n_146),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_1),
.A2(n_95),
.B1(n_203),
.B2(n_208),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g322 ( 
.A1(n_1),
.A2(n_70),
.B1(n_95),
.B2(n_323),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_2),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g293 ( 
.A1(n_2),
.A2(n_41),
.B1(n_204),
.B2(n_294),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_2),
.B(n_303),
.C(n_307),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_2),
.B(n_123),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_2),
.B(n_67),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_2),
.B(n_179),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_2),
.B(n_376),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_3),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_3),
.Y(n_64)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_3),
.Y(n_169)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_4),
.Y(n_117)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_5),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_5),
.Y(n_321)
);

BUFx5_ASAP7_75t_L g346 ( 
.A(n_5),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_5),
.Y(n_383)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_6),
.A2(n_70),
.B1(n_72),
.B2(n_73),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_6),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_6),
.A2(n_72),
.B1(n_131),
.B2(n_185),
.Y(n_245)
);

OAI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_7),
.A2(n_190),
.B1(n_194),
.B2(n_195),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_7),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_8),
.A2(n_155),
.B1(n_174),
.B2(n_177),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_8),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_8),
.A2(n_177),
.B1(n_232),
.B2(n_233),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_L g271 ( 
.A1(n_8),
.A2(n_177),
.B1(n_272),
.B2(n_276),
.Y(n_271)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_9),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_9),
.Y(n_104)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_11),
.A2(n_79),
.B1(n_81),
.B2(n_82),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_11),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_11),
.A2(n_25),
.B1(n_81),
.B2(n_221),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_L g327 ( 
.A1(n_11),
.A2(n_81),
.B1(n_185),
.B2(n_328),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_11),
.A2(n_81),
.B1(n_343),
.B2(n_344),
.Y(n_342)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_12),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_12),
.Y(n_96)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_12),
.Y(n_99)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_12),
.Y(n_107)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_12),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_12),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_12),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_13),
.A2(n_137),
.B1(n_139),
.B2(n_140),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_13),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_13),
.A2(n_139),
.B1(n_238),
.B2(n_240),
.Y(n_237)
);

OAI22xp33_ASAP7_75t_SL g312 ( 
.A1(n_13),
.A2(n_139),
.B1(n_313),
.B2(n_317),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_SL g364 ( 
.A1(n_13),
.A2(n_139),
.B1(n_204),
.B2(n_365),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_14),
.A2(n_249),
.B1(n_250),
.B2(n_251),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_14),
.Y(n_249)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_15),
.Y(n_158)
);

BUFx5_ASAP7_75t_L g160 ( 
.A(n_15),
.Y(n_160)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_15),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_15),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_16),
.A2(n_59),
.B1(n_60),
.B2(n_65),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_16),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_16),
.A2(n_65),
.B1(n_182),
.B2(n_185),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_257),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_256),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2x1_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_222),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_21),
.B(n_222),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_148),
.C(n_199),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_22),
.B(n_284),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_75),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_23),
.B(n_76),
.C(n_112),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_46),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_24),
.A2(n_46),
.B1(n_47),
.B2(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_24),
.Y(n_266)
);

OAI32xp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_28),
.A3(n_30),
.B1(n_34),
.B2(n_40),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_26),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_26),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_26),
.Y(n_122)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_26),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_26),
.Y(n_373)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_27),
.Y(n_90)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_27),
.Y(n_138)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_27),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g377 ( 
.A(n_27),
.Y(n_377)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_32),
.A2(n_88),
.B1(n_90),
.B2(n_91),
.Y(n_87)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_37),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_36),
.Y(n_110)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_38),
.Y(n_37)
);

INVx6_ASAP7_75t_SL g38 ( 
.A(n_39),
.Y(n_38)
);

OAI21xp33_ASAP7_75t_SL g213 ( 
.A1(n_40),
.A2(n_41),
.B(n_214),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_42),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_41),
.B(n_87),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_41),
.A2(n_48),
.B(n_319),
.Y(n_339)
);

OAI21xp33_ASAP7_75t_SL g370 ( 
.A1(n_41),
.A2(n_371),
.B(n_374),
.Y(n_370)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_57),
.B1(n_66),
.B2(n_68),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_48),
.A2(n_189),
.B1(n_247),
.B2(n_248),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_48),
.A2(n_312),
.B(n_319),
.Y(n_311)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_49),
.A2(n_69),
.B1(n_188),
.B2(n_197),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_49),
.A2(n_58),
.B1(n_271),
.B2(n_280),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_49),
.B(n_322),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_49),
.A2(n_320),
.B1(n_352),
.B2(n_353),
.Y(n_351)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_53),
.Y(n_49)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_52),
.Y(n_198)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_52),
.Y(n_281)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_56),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_56),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_56),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_56),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx8_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_66),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx3_ASAP7_75t_L g337 ( 
.A(n_74),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_76),
.A2(n_77),
.B1(n_111),
.B2(n_112),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_85),
.B(n_93),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_78),
.A2(n_87),
.B1(n_236),
.B2(n_237),
.Y(n_235)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_86),
.B(n_94),
.Y(n_218)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_101),
.Y(n_100)
);

INVx4_ASAP7_75t_SL g146 ( 
.A(n_88),
.Y(n_146)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_90),
.Y(n_145)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_100),
.Y(n_93)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx8_ASAP7_75t_L g240 ( 
.A(n_99),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_100),
.A2(n_213),
.B(n_217),
.Y(n_212)
);

INVx2_ASAP7_75t_SL g236 ( 
.A(n_100),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_105),
.B1(n_108),
.B2(n_110),
.Y(n_101)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_135),
.B(n_143),
.Y(n_112)
);

AOI22x1_ASAP7_75t_L g228 ( 
.A1(n_113),
.A2(n_123),
.B1(n_229),
.B2(n_230),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_113),
.B(n_229),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g369 ( 
.A1(n_113),
.A2(n_143),
.B(n_370),
.Y(n_369)
);

INVx2_ASAP7_75t_SL g113 ( 
.A(n_114),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_114),
.A2(n_136),
.B1(n_147),
.B2(n_220),
.Y(n_219)
);

OR2x2_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_123),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_118),
.B1(n_120),
.B2(n_121),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_117),
.Y(n_120)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_117),
.Y(n_126)
);

INVx3_ASAP7_75t_L g389 ( 
.A(n_117),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx5_ASAP7_75t_L g232 ( 
.A(n_119),
.Y(n_232)
);

INVx6_ASAP7_75t_L g392 ( 
.A(n_120),
.Y(n_392)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_123),
.Y(n_147)
);

AO22x2_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_127),
.B1(n_131),
.B2(n_133),
.Y(n_123)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_126),
.Y(n_134)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_129),
.Y(n_367)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_130),
.Y(n_132)
);

INVx11_ASAP7_75t_L g156 ( 
.A(n_130),
.Y(n_156)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_130),
.Y(n_162)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_130),
.Y(n_184)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_130),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_130),
.Y(n_386)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_147),
.Y(n_143)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_144),
.Y(n_229)
);

INVx4_ASAP7_75t_L g385 ( 
.A(n_145),
.Y(n_385)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_146),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_147),
.A2(n_220),
.B(n_269),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_148),
.A2(n_149),
.B1(n_199),
.B2(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_187),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_150),
.B(n_187),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_151),
.A2(n_173),
.B1(n_178),
.B2(n_180),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_151),
.A2(n_293),
.B(n_296),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_151),
.A2(n_178),
.B1(n_327),
.B2(n_364),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_SL g399 ( 
.A1(n_151),
.A2(n_296),
.B(n_364),
.Y(n_399)
);

INVx2_ASAP7_75t_SL g151 ( 
.A(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_152),
.B(n_202),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_152),
.A2(n_179),
.B1(n_181),
.B2(n_245),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_163),
.Y(n_152)
);

OAI22xp33_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_157),
.B1(n_159),
.B2(n_161),
.Y(n_153)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_156),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_156),
.Y(n_186)
);

INVx6_ASAP7_75t_L g210 ( 
.A(n_156),
.Y(n_210)
);

INVx6_ASAP7_75t_L g329 ( 
.A(n_156),
.Y(n_329)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx5_ASAP7_75t_L g306 ( 
.A(n_158),
.Y(n_306)
);

INVx4_ASAP7_75t_SL g159 ( 
.A(n_160),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_163),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_163),
.A2(n_201),
.B(n_327),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_167),
.B1(n_170),
.B2(n_171),
.Y(n_163)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_168),
.Y(n_275)
);

INVx5_ASAP7_75t_L g279 ( 
.A(n_168),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_169),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_169),
.Y(n_253)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_173),
.A2(n_178),
.B(n_201),
.Y(n_200)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx5_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

BUFx2_ASAP7_75t_L g295 ( 
.A(n_176),
.Y(n_295)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_179),
.B(n_202),
.Y(n_296)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx4_ASAP7_75t_SL g182 ( 
.A(n_183),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx11_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_192),
.Y(n_191)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_193),
.Y(n_316)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_195),
.Y(n_343)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_199),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_211),
.C(n_219),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_200),
.B(n_219),
.Y(n_262)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx5_ASAP7_75t_SL g204 ( 
.A(n_205),
.Y(n_204)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx6_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_210),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_211),
.A2(n_212),
.B1(n_262),
.B2(n_263),
.Y(n_261)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_225),
.A2(n_243),
.B1(n_254),
.B2(n_255),
.Y(n_224)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_225),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_228),
.A2(n_235),
.B1(n_241),
.B2(n_242),
.Y(n_227)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_228),
.Y(n_241)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_235),
.Y(n_242)
);

INVx8_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_243),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_246),
.Y(n_243)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx4_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx4_ASAP7_75t_L g318 ( 
.A(n_253),
.Y(n_318)
);

INVx8_ASAP7_75t_L g345 ( 
.A(n_253),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_258),
.A2(n_286),
.B(n_411),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

OR2x2_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_283),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_260),
.B(n_283),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_264),
.C(n_267),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_261),
.B(n_408),
.Y(n_407)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_262),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_264),
.A2(n_265),
.B1(n_267),
.B2(n_409),
.Y(n_408)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_267),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_270),
.C(n_282),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g401 ( 
.A(n_268),
.B(n_402),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_270),
.B(n_282),
.Y(n_402)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_271),
.Y(n_380)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx4_ASAP7_75t_SL g273 ( 
.A(n_274),
.Y(n_273)
);

INVx4_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_279),
.Y(n_309)
);

INVx4_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_287),
.A2(n_405),
.B(n_410),
.Y(n_286)
);

AO21x1_ASAP7_75t_SL g287 ( 
.A1(n_288),
.A2(n_394),
.B(n_404),
.Y(n_287)
);

OAI21x1_ASAP7_75t_L g288 ( 
.A1(n_289),
.A2(n_358),
.B(n_393),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_290),
.A2(n_332),
.B(n_357),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_310),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_291),
.B(n_310),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_292),
.B(n_297),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_292),
.A2(n_297),
.B1(n_298),
.B2(n_355),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_292),
.Y(n_355)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_302),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx3_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_324),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_311),
.B(n_325),
.C(n_331),
.Y(n_359)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_312),
.Y(n_353)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx6_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx4_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx4_ASAP7_75t_L g323 ( 
.A(n_316),
.Y(n_323)
);

INVx4_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_322),
.Y(n_319)
);

INVx4_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_325),
.A2(n_326),
.B1(n_330),
.B2(n_331),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

NAND2xp33_ASAP7_75t_SL g390 ( 
.A(n_328),
.B(n_391),
.Y(n_390)
);

INVx8_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_333),
.A2(n_350),
.B(n_356),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_334),
.A2(n_340),
.B(n_349),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_339),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_338),
.Y(n_335)
);

INVx1_ASAP7_75t_SL g336 ( 
.A(n_337),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_341),
.B(n_348),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_341),
.B(n_348),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_342),
.A2(n_346),
.B(n_347),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_342),
.Y(n_352)
);

INVx4_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g379 ( 
.A1(n_347),
.A2(n_380),
.B(n_381),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_354),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_351),
.B(n_354),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_360),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_359),
.B(n_360),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_378),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_362),
.A2(n_363),
.B1(n_368),
.B2(n_369),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_363),
.B(n_368),
.C(n_378),
.Y(n_395)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx6_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx6_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVxp33_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

AOI32xp33_ASAP7_75t_L g384 ( 
.A1(n_375),
.A2(n_385),
.A3(n_386),
.B1(n_387),
.B2(n_390),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_384),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_379),
.B(n_384),
.Y(n_400)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx3_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx4_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx4_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_396),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_SL g404 ( 
.A(n_395),
.B(n_396),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_397),
.A2(n_398),
.B1(n_401),
.B2(n_403),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_SL g398 ( 
.A(n_399),
.B(n_400),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_399),
.B(n_400),
.C(n_403),
.Y(n_406)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_401),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_407),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_SL g410 ( 
.A(n_406),
.B(n_407),
.Y(n_410)
);


endmodule