module real_aes_17018_n_312 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_19, n_40, n_239, n_100, n_54, n_112, n_35, n_42, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_232, n_6, n_69, n_73, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_292, n_116, n_94, n_289, n_280, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_304, n_311, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_89, n_277, n_93, n_182, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_195, n_300, n_252, n_283, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_183, n_266, n_205, n_177, n_22, n_140, n_219, n_180, n_212, n_210, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_14, n_194, n_137, n_225, n_16, n_39, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_312);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_19;
input n_40;
input n_239;
input n_100;
input n_54;
input n_112;
input n_35;
input n_42;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_232;
input n_6;
input n_69;
input n_73;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_304;
input n_311;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_89;
input n_277;
input n_93;
input n_182;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_195;
input n_300;
input n_252;
input n_283;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_183;
input n_266;
input n_205;
input n_177;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_312;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1328;
wire n_1034;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_553;
wire n_1367;
wire n_744;
wire n_1325;
wire n_1382;
wire n_1225;
wire n_875;
wire n_1199;
wire n_951;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_1537;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1639;
wire n_1224;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_368;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1383;
wire n_1346;
wire n_1675;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_1600;
wire n_619;
wire n_1284;
wire n_1095;
wire n_1250;
wire n_360;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_488;
wire n_1380;
wire n_1658;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_1301;
wire n_728;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_1003;
wire n_346;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_1351;
wire n_972;
wire n_1628;
wire n_1587;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_1397;
wire n_765;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1615;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1666;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1495;
wire n_1510;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1648;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_1488;
wire n_337;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_667;
wire n_991;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1417;
wire n_1370;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_1260;
wire n_328;
wire n_355;
wire n_1606;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1594;
wire n_537;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_948;
wire n_399;
wire n_700;
wire n_1499;
wire n_1269;
wire n_677;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_1338;
wire n_981;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1189;
wire n_1070;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_1145;
wire n_645;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_985;
wire n_777;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_1179;
wire n_334;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_720;
wire n_354;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_1403;
wire n_643;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_1409;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1133;
wire n_1593;
wire n_313;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_325;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1172;
wire n_459;
wire n_998;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_967;
wire n_1159;
wire n_474;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_1185;
wire n_661;
wire n_1102;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_1377;
wire n_800;
wire n_1170;
wire n_1175;
wire n_778;
wire n_522;
wire n_1475;
wire n_943;
wire n_977;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1268;
wire n_1113;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_1644;
wire n_594;
wire n_856;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_370;
wire n_1663;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_316;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1411;
wire n_1263;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1671;
wire n_1414;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1670;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1331;
wire n_714;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_1592;
wire n_1605;
wire n_663;
wire n_588;
wire n_1682;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_1378;
wire n_524;
wire n_1496;
wire n_1191;
wire n_705;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_1617;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1143;
wire n_929;
wire n_1190;
wire n_543;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1466;
wire n_1396;
wire n_921;
wire n_1176;
wire n_640;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_1679;
wire n_317;
wire n_1595;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_578;
wire n_372;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_559;
wire n_466;
wire n_1049;
wire n_1277;
wire n_1584;
wire n_984;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_924;
wire n_1264;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1290;
wire n_1318;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_1100;
wire n_398;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_331;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1647;
wire n_1252;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1573;
wire n_1130;
wire n_794;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_1300;
wire n_575;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_1630;
wire n_1352;
wire n_729;
wire n_394;
wire n_1323;
wire n_1280;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
NOR2xp33_ASAP7_75t_L g337 ( .A(n_0), .B(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g366 ( .A(n_0), .Y(n_366) );
AND2x2_ASAP7_75t_L g564 ( .A(n_0), .B(n_227), .Y(n_564) );
AND2x2_ASAP7_75t_L g582 ( .A(n_0), .B(n_467), .Y(n_582) );
AOI22xp33_ASAP7_75t_SL g1129 ( .A1(n_1), .A2(n_280), .B1(n_844), .B2(n_1078), .Y(n_1129) );
AOI221xp5_ASAP7_75t_L g1144 ( .A1(n_1), .A2(n_3), .B1(n_585), .B2(n_592), .C(n_1145), .Y(n_1144) );
AOI22xp33_ASAP7_75t_SL g524 ( .A1(n_2), .A2(n_39), .B1(n_525), .B2(n_529), .Y(n_524) );
INVxp67_ASAP7_75t_SL g620 ( .A(n_2), .Y(n_620) );
AOI22xp33_ASAP7_75t_SL g1135 ( .A1(n_3), .A2(n_7), .B1(n_541), .B2(n_1039), .Y(n_1135) );
AOI22xp33_ASAP7_75t_SL g1075 ( .A1(n_4), .A2(n_279), .B1(n_1076), .B2(n_1078), .Y(n_1075) );
AOI221xp5_ASAP7_75t_L g1098 ( .A1(n_4), .A2(n_232), .B1(n_1003), .B2(n_1099), .C(n_1100), .Y(n_1098) );
INVx1_ASAP7_75t_L g1234 ( .A(n_5), .Y(n_1234) );
XOR2x2_ASAP7_75t_L g317 ( .A(n_6), .B(n_318), .Y(n_317) );
AOI22xp5_ASAP7_75t_L g1459 ( .A1(n_6), .A2(n_50), .B1(n_1434), .B2(n_1440), .Y(n_1459) );
A2O1A1Ixp33_ASAP7_75t_L g1153 ( .A1(n_7), .A2(n_1154), .B(n_1155), .C(n_1160), .Y(n_1153) );
OAI22xp5_ASAP7_75t_L g1299 ( .A1(n_8), .A2(n_199), .B1(n_908), .B2(n_1300), .Y(n_1299) );
INVxp67_ASAP7_75t_SL g1167 ( .A(n_9), .Y(n_1167) );
AND4x1_ASAP7_75t_L g1207 ( .A(n_9), .B(n_1169), .C(n_1172), .D(n_1192), .Y(n_1207) );
AOI22xp33_ASAP7_75t_L g801 ( .A1(n_10), .A2(n_290), .B1(n_802), .B2(n_803), .Y(n_801) );
INVx1_ASAP7_75t_L g824 ( .A(n_10), .Y(n_824) );
INVx2_ASAP7_75t_L g376 ( .A(n_11), .Y(n_376) );
OAI22xp5_ASAP7_75t_SL g994 ( .A1(n_12), .A2(n_253), .B1(n_836), .B2(n_995), .Y(n_994) );
OAI221xp5_ASAP7_75t_L g1010 ( .A1(n_12), .A2(n_253), .B1(n_610), .B2(n_612), .C(n_1011), .Y(n_1010) );
XNOR2x1_ASAP7_75t_L g972 ( .A(n_13), .B(n_973), .Y(n_972) );
INVx1_ASAP7_75t_L g1280 ( .A(n_14), .Y(n_1280) );
INVx1_ASAP7_75t_L g903 ( .A(n_15), .Y(n_903) );
INVx1_ASAP7_75t_L g1278 ( .A(n_16), .Y(n_1278) );
AOI22xp33_ASAP7_75t_L g1289 ( .A1(n_16), .A2(n_62), .B1(n_1290), .B2(n_1291), .Y(n_1289) );
OAI22xp5_ASAP7_75t_L g1171 ( .A1(n_17), .A2(n_152), .B1(n_569), .B2(n_573), .Y(n_1171) );
OAI211xp5_ASAP7_75t_L g1173 ( .A1(n_17), .A2(n_950), .B(n_1174), .C(n_1177), .Y(n_1173) );
AOI22xp5_ASAP7_75t_L g1473 ( .A1(n_18), .A2(n_200), .B1(n_1430), .B2(n_1437), .Y(n_1473) );
AOI22xp33_ASAP7_75t_L g1182 ( .A1(n_19), .A2(n_83), .B1(n_1110), .B2(n_1183), .Y(n_1182) );
AOI22xp33_ASAP7_75t_L g1201 ( .A1(n_19), .A2(n_29), .B1(n_534), .B2(n_1200), .Y(n_1201) );
INVx1_ASAP7_75t_L g1381 ( .A(n_20), .Y(n_1381) );
AOI221xp5_ASAP7_75t_L g1402 ( .A1(n_20), .A2(n_134), .B1(n_534), .B2(n_1403), .C(n_1405), .Y(n_1402) );
INVx1_ASAP7_75t_L g1009 ( .A(n_21), .Y(n_1009) );
HB1xp67_ASAP7_75t_L g1422 ( .A(n_22), .Y(n_1422) );
AND2x2_ASAP7_75t_L g1431 ( .A(n_22), .B(n_1420), .Y(n_1431) );
AOI22xp5_ASAP7_75t_L g1458 ( .A1(n_23), .A2(n_178), .B1(n_1430), .B2(n_1437), .Y(n_1458) );
OAI22xp5_ASAP7_75t_SL g866 ( .A1(n_24), .A2(n_260), .B1(n_323), .B2(n_349), .Y(n_866) );
INVxp67_ASAP7_75t_SL g906 ( .A(n_24), .Y(n_906) );
INVx1_ASAP7_75t_L g922 ( .A(n_25), .Y(n_922) );
OAI211xp5_ASAP7_75t_L g931 ( .A1(n_25), .A2(n_932), .B(n_933), .C(n_940), .Y(n_931) );
INVxp67_ASAP7_75t_L g1066 ( .A(n_26), .Y(n_1066) );
CKINVDCx5p33_ASAP7_75t_R g1170 ( .A(n_27), .Y(n_1170) );
AOI22xp5_ASAP7_75t_L g1464 ( .A1(n_28), .A2(n_245), .B1(n_1430), .B2(n_1437), .Y(n_1464) );
AOI221xp5_ASAP7_75t_L g1190 ( .A1(n_29), .A2(n_294), .B1(n_630), .B2(n_939), .C(n_1191), .Y(n_1190) );
AOI22xp33_ASAP7_75t_L g767 ( .A1(n_30), .A2(n_45), .B1(n_535), .B2(n_705), .Y(n_767) );
INVx1_ASAP7_75t_L g780 ( .A(n_30), .Y(n_780) );
INVx1_ASAP7_75t_L g1390 ( .A(n_31), .Y(n_1390) );
OAI22xp33_ASAP7_75t_L g1399 ( .A1(n_31), .A2(n_46), .B1(n_718), .B2(n_720), .Y(n_1399) );
INVx1_ASAP7_75t_L g677 ( .A(n_32), .Y(n_677) );
AOI22xp5_ASAP7_75t_L g641 ( .A1(n_33), .A2(n_43), .B1(n_642), .B2(n_643), .Y(n_641) );
AOI22xp33_ASAP7_75t_L g703 ( .A1(n_33), .A2(n_150), .B1(n_704), .B2(n_706), .Y(n_703) );
AOI22xp33_ASAP7_75t_L g1130 ( .A1(n_34), .A2(n_91), .B1(n_1072), .B2(n_1131), .Y(n_1130) );
AOI221xp5_ASAP7_75t_L g1156 ( .A1(n_34), .A2(n_182), .B1(n_1022), .B2(n_1100), .C(n_1157), .Y(n_1156) );
AOI221xp5_ASAP7_75t_L g946 ( .A1(n_35), .A2(n_276), .B1(n_625), .B2(n_876), .C(n_939), .Y(n_946) );
INVxp67_ASAP7_75t_SL g958 ( .A(n_35), .Y(n_958) );
AOI22xp5_ASAP7_75t_L g1453 ( .A1(n_36), .A2(n_117), .B1(n_1430), .B2(n_1437), .Y(n_1453) );
INVx1_ASAP7_75t_L g928 ( .A(n_37), .Y(n_928) );
OAI22xp5_ASAP7_75t_L g947 ( .A1(n_37), .A2(n_192), .B1(n_948), .B2(n_950), .Y(n_947) );
AOI221xp5_ASAP7_75t_L g756 ( .A1(n_38), .A2(n_304), .B1(n_432), .B2(n_757), .C(n_758), .Y(n_756) );
AOI221xp5_ASAP7_75t_L g778 ( .A1(n_38), .A2(n_118), .B1(n_771), .B2(n_772), .C(n_779), .Y(n_778) );
AOI221xp5_ASAP7_75t_L g584 ( .A1(n_39), .A2(n_96), .B1(n_585), .B2(n_587), .C(n_591), .Y(n_584) );
INVx1_ASAP7_75t_L g806 ( .A(n_40), .Y(n_806) );
NAND5xp2_ASAP7_75t_L g1307 ( .A(n_41), .B(n_1308), .C(n_1325), .D(n_1336), .E(n_1340), .Y(n_1307) );
INVx1_ASAP7_75t_L g1346 ( .A(n_41), .Y(n_1346) );
AOI22xp5_ASAP7_75t_L g1451 ( .A1(n_41), .A2(n_159), .B1(n_1440), .B2(n_1452), .Y(n_1451) );
XNOR2xp5_ASAP7_75t_L g1638 ( .A(n_42), .B(n_1639), .Y(n_1638) );
AOI22xp33_ASAP7_75t_SL g690 ( .A1(n_43), .A2(n_161), .B1(n_691), .B2(n_693), .Y(n_690) );
INVx1_ASAP7_75t_L g805 ( .A(n_44), .Y(n_805) );
INVx1_ASAP7_75t_L g774 ( .A(n_45), .Y(n_774) );
OAI221xp5_ASAP7_75t_L g1384 ( .A1(n_46), .A2(n_273), .B1(n_658), .B2(n_659), .C(n_1385), .Y(n_1384) );
INVxp67_ASAP7_75t_SL g945 ( .A(n_47), .Y(n_945) );
AOI22xp33_ASAP7_75t_L g967 ( .A1(n_47), .A2(n_131), .B1(n_968), .B2(n_969), .Y(n_967) );
BUFx6f_ASAP7_75t_L g325 ( .A(n_48), .Y(n_325) );
INVx1_ASAP7_75t_L g1175 ( .A(n_49), .Y(n_1175) );
OAI22xp33_ASAP7_75t_L g1194 ( .A1(n_49), .A2(n_98), .B1(n_543), .B2(n_1195), .Y(n_1194) );
CKINVDCx5p33_ASAP7_75t_R g1376 ( .A(n_51), .Y(n_1376) );
INVx1_ASAP7_75t_L g1008 ( .A(n_52), .Y(n_1008) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_53), .A2(n_233), .B1(n_531), .B2(n_534), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_53), .A2(n_133), .B1(n_594), .B2(n_596), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g1531 ( .A1(n_54), .A2(n_218), .B1(n_1434), .B2(n_1440), .Y(n_1531) );
AOI221xp5_ASAP7_75t_L g1313 ( .A1(n_55), .A2(n_158), .B1(n_483), .B2(n_876), .C(n_939), .Y(n_1313) );
AOI22xp33_ASAP7_75t_L g1329 ( .A1(n_55), .A2(n_212), .B1(n_404), .B2(n_706), .Y(n_1329) );
CKINVDCx5p33_ASAP7_75t_R g1139 ( .A(n_56), .Y(n_1139) );
AOI22xp33_ASAP7_75t_L g1314 ( .A1(n_57), .A2(n_212), .B1(n_803), .B2(n_1183), .Y(n_1314) );
AOI22xp33_ASAP7_75t_L g1328 ( .A1(n_57), .A2(n_158), .B1(n_706), .B2(n_1042), .Y(n_1328) );
INVxp67_ASAP7_75t_SL g1388 ( .A(n_58), .Y(n_1388) );
OAI22xp5_ASAP7_75t_L g1408 ( .A1(n_58), .A2(n_729), .B1(n_1409), .B2(n_1411), .Y(n_1408) );
INVx1_ASAP7_75t_L g346 ( .A(n_59), .Y(n_346) );
AOI22xp33_ASAP7_75t_L g1083 ( .A1(n_60), .A2(n_147), .B1(n_1071), .B2(n_1084), .Y(n_1083) );
AOI21xp33_ASAP7_75t_L g1111 ( .A1(n_60), .A2(n_630), .B(n_1112), .Y(n_1111) );
AOI221xp5_ASAP7_75t_L g1178 ( .A1(n_61), .A2(n_293), .B1(n_1112), .B2(n_1179), .C(n_1181), .Y(n_1178) );
AOI22xp33_ASAP7_75t_SL g1202 ( .A1(n_61), .A2(n_268), .B1(n_704), .B2(n_1203), .Y(n_1202) );
INVx1_ASAP7_75t_L g1268 ( .A(n_62), .Y(n_1268) );
INVx1_ASAP7_75t_L g1126 ( .A(n_63), .Y(n_1126) );
AOI221xp5_ASAP7_75t_L g645 ( .A1(n_64), .A2(n_291), .B1(n_646), .B2(n_648), .C(n_650), .Y(n_645) );
AOI221xp5_ASAP7_75t_L g696 ( .A1(n_64), .A2(n_262), .B1(n_697), .B2(n_699), .C(n_702), .Y(n_696) );
OAI211xp5_ASAP7_75t_SL g747 ( .A1(n_65), .A2(n_715), .B(n_722), .C(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g783 ( .A(n_65), .Y(n_783) );
OAI22xp5_ASAP7_75t_L g420 ( .A1(n_66), .A2(n_226), .B1(n_421), .B2(n_425), .Y(n_420) );
OAI22xp5_ASAP7_75t_L g470 ( .A1(n_66), .A2(n_226), .B1(n_471), .B2(n_473), .Y(n_470) );
CKINVDCx5p33_ASAP7_75t_R g1088 ( .A(n_67), .Y(n_1088) );
OAI21xp5_ASAP7_75t_SL g1117 ( .A1(n_68), .A2(n_569), .B(n_1118), .Y(n_1117) );
CKINVDCx5p33_ASAP7_75t_R g1320 ( .A(n_69), .Y(n_1320) );
AOI22xp33_ASAP7_75t_L g1225 ( .A1(n_70), .A2(n_210), .B1(n_529), .B2(n_1226), .Y(n_1225) );
AOI22xp33_ASAP7_75t_SL g1253 ( .A1(n_70), .A2(n_258), .B1(n_802), .B2(n_1110), .Y(n_1253) );
INVxp67_ASAP7_75t_SL g683 ( .A(n_71), .Y(n_683) );
OAI22xp5_ASAP7_75t_L g707 ( .A1(n_71), .A2(n_299), .B1(n_708), .B2(n_711), .Y(n_707) );
INVx1_ASAP7_75t_L g1392 ( .A(n_72), .Y(n_1392) );
OAI222xp33_ASAP7_75t_L g1395 ( .A1(n_72), .A2(n_259), .B1(n_273), .B2(n_692), .C1(n_962), .C2(n_1396), .Y(n_1395) );
AOI22xp33_ASAP7_75t_SL g1080 ( .A1(n_73), .A2(n_232), .B1(n_541), .B2(n_1081), .Y(n_1080) );
AOI22xp33_ASAP7_75t_L g1108 ( .A1(n_73), .A2(n_279), .B1(n_1109), .B2(n_1110), .Y(n_1108) );
AOI22xp33_ASAP7_75t_L g538 ( .A1(n_74), .A2(n_96), .B1(n_529), .B2(n_539), .Y(n_538) );
INVxp67_ASAP7_75t_SL g623 ( .A(n_74), .Y(n_623) );
OR2x2_ASAP7_75t_L g926 ( .A(n_75), .B(n_559), .Y(n_926) );
OAI221xp5_ASAP7_75t_L g941 ( .A1(n_76), .A2(n_191), .B1(n_612), .B2(n_942), .C(n_943), .Y(n_941) );
OAI322xp33_ASAP7_75t_L g956 ( .A1(n_76), .A2(n_407), .A3(n_550), .B1(n_890), .B2(n_957), .C1(n_960), .C2(n_963), .Y(n_956) );
AOI22xp33_ASAP7_75t_L g1436 ( .A1(n_77), .A2(n_160), .B1(n_1437), .B2(n_1440), .Y(n_1436) );
AOI22xp33_ASAP7_75t_SL g1041 ( .A1(n_78), .A2(n_186), .B1(n_706), .B2(n_1042), .Y(n_1041) );
AOI22xp33_ASAP7_75t_L g1054 ( .A1(n_78), .A2(n_88), .B1(n_597), .B2(n_802), .Y(n_1054) );
AOI22xp33_ASAP7_75t_SL g1224 ( .A1(n_79), .A2(n_204), .B1(n_693), .B2(n_1222), .Y(n_1224) );
INVx1_ASAP7_75t_L g1248 ( .A(n_79), .Y(n_1248) );
AOI22xp33_ASAP7_75t_SL g869 ( .A1(n_80), .A2(n_149), .B1(n_580), .B2(n_870), .Y(n_869) );
INVxp67_ASAP7_75t_SL g899 ( .A(n_80), .Y(n_899) );
INVx1_ASAP7_75t_L g976 ( .A(n_81), .Y(n_976) );
AOI22xp33_ASAP7_75t_SL g984 ( .A1(n_82), .A2(n_255), .B1(n_901), .B2(n_985), .Y(n_984) );
AOI221xp5_ASAP7_75t_L g1001 ( .A1(n_82), .A2(n_90), .B1(n_872), .B2(n_1002), .C(n_1003), .Y(n_1001) );
AOI22xp33_ASAP7_75t_L g1199 ( .A1(n_83), .A2(n_294), .B1(n_534), .B2(n_1200), .Y(n_1199) );
AOI22xp33_ASAP7_75t_L g1429 ( .A1(n_84), .A2(n_269), .B1(n_1430), .B2(n_1434), .Y(n_1429) );
AOI22xp33_ASAP7_75t_L g1655 ( .A1(n_85), .A2(n_243), .B1(n_525), .B2(n_985), .Y(n_1655) );
AOI221xp5_ASAP7_75t_L g1660 ( .A1(n_85), .A2(n_238), .B1(n_586), .B2(n_592), .C(n_772), .Y(n_1660) );
AOI22xp5_ASAP7_75t_L g1476 ( .A1(n_86), .A2(n_144), .B1(n_1440), .B2(n_1449), .Y(n_1476) );
INVx1_ASAP7_75t_L g978 ( .A(n_87), .Y(n_978) );
AOI22xp33_ASAP7_75t_SL g1045 ( .A1(n_88), .A2(n_257), .B1(n_706), .B2(n_1042), .Y(n_1045) );
INVx1_ASAP7_75t_L g1648 ( .A(n_89), .Y(n_1648) );
AOI22xp33_ASAP7_75t_L g1661 ( .A1(n_89), .A2(n_266), .B1(n_597), .B2(n_1109), .Y(n_1661) );
AOI22xp33_ASAP7_75t_L g993 ( .A1(n_90), .A2(n_175), .B1(n_697), .B2(n_968), .Y(n_993) );
AOI22xp33_ASAP7_75t_SL g1147 ( .A1(n_91), .A2(n_130), .B1(n_596), .B2(n_802), .Y(n_1147) );
INVx1_ASAP7_75t_L g340 ( .A(n_92), .Y(n_340) );
INVx1_ASAP7_75t_L g1277 ( .A(n_93), .Y(n_1277) );
AOI221xp5_ASAP7_75t_L g1285 ( .A1(n_93), .A2(n_205), .B1(n_625), .B2(n_630), .C(n_1099), .Y(n_1285) );
CKINVDCx5p33_ASAP7_75t_R g1036 ( .A(n_94), .Y(n_1036) );
CKINVDCx5p33_ASAP7_75t_R g1096 ( .A(n_95), .Y(n_1096) );
XNOR2xp5_ASAP7_75t_L g793 ( .A(n_97), .B(n_794), .Y(n_793) );
INVx1_ASAP7_75t_L g1176 ( .A(n_98), .Y(n_1176) );
OAI211xp5_ASAP7_75t_L g1317 ( .A1(n_99), .A2(n_1249), .B(n_1318), .C(n_1319), .Y(n_1317) );
INVx1_ASAP7_75t_L g1342 ( .A(n_99), .Y(n_1342) );
INVx1_ASAP7_75t_L g944 ( .A(n_100), .Y(n_944) );
AOI22xp33_ASAP7_75t_L g1532 ( .A1(n_101), .A2(n_289), .B1(n_1430), .B2(n_1437), .Y(n_1532) );
CKINVDCx5p33_ASAP7_75t_R g1091 ( .A(n_102), .Y(n_1091) );
OAI22xp5_ASAP7_75t_L g1114 ( .A1(n_102), .A2(n_121), .B1(n_1115), .B2(n_1116), .Y(n_1114) );
CKINVDCx5p33_ASAP7_75t_R g1378 ( .A(n_103), .Y(n_1378) );
AOI22xp33_ASAP7_75t_L g877 ( .A1(n_104), .A2(n_211), .B1(n_580), .B2(n_878), .Y(n_877) );
AOI22xp33_ASAP7_75t_L g895 ( .A1(n_104), .A2(n_230), .B1(n_529), .B2(n_541), .Y(n_895) );
INVx1_ASAP7_75t_L g369 ( .A(n_105), .Y(n_369) );
AOI21xp33_ASAP7_75t_L g814 ( .A1(n_106), .A2(n_772), .B(n_815), .Y(n_814) );
INVx1_ASAP7_75t_L g823 ( .A(n_106), .Y(n_823) );
INVx1_ASAP7_75t_L g851 ( .A(n_107), .Y(n_851) );
INVx1_ASAP7_75t_L g1642 ( .A(n_108), .Y(n_1642) );
CKINVDCx5p33_ASAP7_75t_R g1382 ( .A(n_109), .Y(n_1382) );
OAI221xp5_ASAP7_75t_L g1184 ( .A1(n_110), .A2(n_240), .B1(n_608), .B2(n_1185), .C(n_1186), .Y(n_1184) );
INVx1_ASAP7_75t_L g1206 ( .A(n_110), .Y(n_1206) );
INVx1_ASAP7_75t_L g1420 ( .A(n_111), .Y(n_1420) );
AOI221xp5_ASAP7_75t_L g798 ( .A1(n_112), .A2(n_228), .B1(n_592), .B2(n_771), .C(n_799), .Y(n_798) );
AOI22xp33_ASAP7_75t_L g828 ( .A1(n_112), .A2(n_164), .B1(n_525), .B2(n_556), .Y(n_828) );
INVx1_ASAP7_75t_L g1031 ( .A(n_113), .Y(n_1031) );
INVx1_ASAP7_75t_L g1030 ( .A(n_114), .Y(n_1030) );
INVx1_ASAP7_75t_L g1389 ( .A(n_115), .Y(n_1389) );
AOI221xp5_ASAP7_75t_L g1038 ( .A1(n_116), .A2(n_256), .B1(n_968), .B2(n_1039), .C(n_1040), .Y(n_1038) );
AOI221xp5_ASAP7_75t_L g1053 ( .A1(n_116), .A2(n_208), .B1(n_586), .B2(n_588), .C(n_1003), .Y(n_1053) );
INVx1_ASAP7_75t_L g763 ( .A(n_118), .Y(n_763) );
OAI22xp33_ASAP7_75t_L g1265 ( .A1(n_119), .A2(n_271), .B1(n_543), .B2(n_1195), .Y(n_1265) );
INVx1_ASAP7_75t_L g1294 ( .A(n_119), .Y(n_1294) );
INVx1_ASAP7_75t_L g515 ( .A(n_120), .Y(n_515) );
OAI221xp5_ASAP7_75t_L g607 ( .A1(n_120), .A2(n_122), .B1(n_608), .B2(n_612), .C(n_616), .Y(n_607) );
CKINVDCx5p33_ASAP7_75t_R g1090 ( .A(n_121), .Y(n_1090) );
INVx1_ASAP7_75t_L g506 ( .A(n_122), .Y(n_506) );
OAI211xp5_ASAP7_75t_L g855 ( .A1(n_123), .A2(n_856), .B(n_857), .C(n_859), .Y(n_855) );
INVxp33_ASAP7_75t_SL g885 ( .A(n_123), .Y(n_885) );
CKINVDCx5p33_ASAP7_75t_R g1653 ( .A(n_124), .Y(n_1653) );
OAI22xp33_ASAP7_75t_L g725 ( .A1(n_125), .A2(n_156), .B1(n_726), .B2(n_729), .Y(n_725) );
INVxp67_ASAP7_75t_SL g734 ( .A(n_125), .Y(n_734) );
INVx1_ASAP7_75t_L g1269 ( .A(n_126), .Y(n_1269) );
AOI221xp5_ASAP7_75t_L g1288 ( .A1(n_126), .A2(n_249), .B1(n_591), .B2(n_625), .C(n_1157), .Y(n_1288) );
AOI22xp33_ASAP7_75t_SL g1463 ( .A1(n_127), .A2(n_195), .B1(n_1434), .B2(n_1440), .Y(n_1463) );
INVx1_ASAP7_75t_L g1647 ( .A(n_128), .Y(n_1647) );
AOI21xp33_ASAP7_75t_L g1668 ( .A1(n_128), .A2(n_630), .B(n_772), .Y(n_1668) );
OAI22xp5_ASAP7_75t_L g1643 ( .A1(n_129), .A2(n_155), .B1(n_573), .B2(n_841), .Y(n_1643) );
OAI211xp5_ASAP7_75t_L g1658 ( .A1(n_129), .A2(n_578), .B(n_1659), .C(n_1662), .Y(n_1658) );
AOI22xp33_ASAP7_75t_L g1133 ( .A1(n_130), .A2(n_182), .B1(n_1072), .B2(n_1134), .Y(n_1133) );
AOI221xp5_ASAP7_75t_L g938 ( .A1(n_131), .A2(n_201), .B1(n_592), .B2(n_872), .C(n_939), .Y(n_938) );
OAI22xp33_ASAP7_75t_L g746 ( .A1(n_132), .A2(n_309), .B1(n_726), .B2(n_729), .Y(n_746) );
INVxp33_ASAP7_75t_SL g787 ( .A(n_132), .Y(n_787) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_133), .A2(n_162), .B1(n_531), .B2(n_534), .Y(n_536) );
INVx1_ASAP7_75t_L g1363 ( .A(n_134), .Y(n_1363) );
INVx1_ASAP7_75t_L g1215 ( .A(n_135), .Y(n_1215) );
OAI221xp5_ASAP7_75t_L g1246 ( .A1(n_135), .A2(n_136), .B1(n_808), .B2(n_809), .C(n_1247), .Y(n_1246) );
INVx1_ASAP7_75t_L g1216 ( .A(n_136), .Y(n_1216) );
CKINVDCx5p33_ASAP7_75t_R g749 ( .A(n_137), .Y(n_749) );
OA21x2_ASAP7_75t_L g974 ( .A1(n_138), .A2(n_559), .B(n_975), .Y(n_974) );
INVx1_ASAP7_75t_L g753 ( .A(n_139), .Y(n_753) );
AOI221xp5_ASAP7_75t_L g770 ( .A1(n_139), .A2(n_221), .B1(n_771), .B2(n_772), .C(n_773), .Y(n_770) );
AOI221xp5_ASAP7_75t_L g661 ( .A1(n_140), .A2(n_150), .B1(n_643), .B2(n_662), .C(n_664), .Y(n_661) );
AOI221xp5_ASAP7_75t_L g694 ( .A1(n_140), .A2(n_291), .B1(n_525), .B2(n_529), .C(n_695), .Y(n_694) );
OAI22xp33_ASAP7_75t_L g542 ( .A1(n_141), .A2(n_251), .B1(n_543), .B2(n_550), .Y(n_542) );
INVx1_ASAP7_75t_L g604 ( .A(n_141), .Y(n_604) );
OAI22xp33_ASAP7_75t_L g445 ( .A1(n_142), .A2(n_151), .B1(n_446), .B2(n_449), .Y(n_445) );
OAI22xp33_ASAP7_75t_L g457 ( .A1(n_142), .A2(n_151), .B1(n_458), .B2(n_464), .Y(n_457) );
OAI221xp5_ASAP7_75t_L g807 ( .A1(n_143), .A2(n_301), .B1(n_808), .B2(n_809), .C(n_810), .Y(n_807) );
OAI22xp33_ASAP7_75t_L g835 ( .A1(n_143), .A2(n_301), .B1(n_508), .B2(n_836), .Y(n_835) );
AO22x1_ASAP7_75t_L g1070 ( .A1(n_145), .A2(n_181), .B1(n_1071), .B2(n_1072), .Y(n_1070) );
NAND2xp5_ASAP7_75t_L g1105 ( .A(n_145), .B(n_1106), .Y(n_1105) );
INVx1_ASAP7_75t_L g1339 ( .A(n_146), .Y(n_1339) );
AOI22xp33_ASAP7_75t_SL g1102 ( .A1(n_147), .A2(n_181), .B1(n_594), .B2(n_1103), .Y(n_1102) );
INVx1_ASAP7_75t_L g435 ( .A(n_148), .Y(n_435) );
INVx1_ASAP7_75t_L g894 ( .A(n_149), .Y(n_894) );
INVx1_ASAP7_75t_L g356 ( .A(n_153), .Y(n_356) );
CKINVDCx5p33_ASAP7_75t_R g862 ( .A(n_154), .Y(n_862) );
INVxp67_ASAP7_75t_SL g671 ( .A(n_156), .Y(n_671) );
OAI22xp5_ASAP7_75t_L g568 ( .A1(n_157), .A2(n_173), .B1(n_569), .B2(n_573), .Y(n_568) );
OAI211xp5_ASAP7_75t_L g577 ( .A1(n_157), .A2(n_578), .B(n_583), .C(n_599), .Y(n_577) );
INVx1_ASAP7_75t_L g665 ( .A(n_161), .Y(n_665) );
AOI221xp5_ASAP7_75t_L g624 ( .A1(n_162), .A2(n_233), .B1(n_625), .B2(n_626), .C(n_630), .Y(n_624) );
CKINVDCx5p33_ASAP7_75t_R g860 ( .A(n_163), .Y(n_860) );
AOI22xp33_ASAP7_75t_SL g816 ( .A1(n_164), .A2(n_278), .B1(n_580), .B2(n_594), .Y(n_816) );
OAI211xp5_ASAP7_75t_L g796 ( .A1(n_165), .A2(n_578), .B(n_797), .C(n_804), .Y(n_796) );
OAI22xp5_ASAP7_75t_L g840 ( .A1(n_165), .A2(n_292), .B1(n_573), .B2(n_841), .Y(n_840) );
INVx1_ASAP7_75t_L g874 ( .A(n_166), .Y(n_874) );
AOI22xp33_ASAP7_75t_SL g1221 ( .A1(n_167), .A2(n_263), .B1(n_693), .B2(n_1222), .Y(n_1221) );
AOI22xp33_ASAP7_75t_L g1241 ( .A1(n_167), .A2(n_204), .B1(n_597), .B2(n_1242), .Y(n_1241) );
INVx1_ASAP7_75t_L g983 ( .A(n_168), .Y(n_983) );
AOI221xp5_ASAP7_75t_L g1017 ( .A1(n_168), .A2(n_203), .B1(n_588), .B2(n_1018), .C(n_1022), .Y(n_1017) );
OAI211xp5_ASAP7_75t_L g1309 ( .A1(n_169), .A2(n_1310), .B(n_1311), .C(n_1316), .Y(n_1309) );
NOR2xp33_ASAP7_75t_L g1324 ( .A(n_169), .B(n_908), .Y(n_1324) );
AOI221xp5_ASAP7_75t_L g1043 ( .A1(n_170), .A2(n_208), .B1(n_697), .B2(n_968), .C(n_1044), .Y(n_1043) );
AOI22xp33_ASAP7_75t_L g1056 ( .A1(n_170), .A2(n_256), .B1(n_597), .B2(n_870), .Y(n_1056) );
AND2x2_ASAP7_75t_L g1432 ( .A(n_171), .B(n_1433), .Y(n_1432) );
AND2x2_ASAP7_75t_L g1435 ( .A(n_171), .B(n_267), .Y(n_1435) );
INVx2_ASAP7_75t_L g1439 ( .A(n_171), .Y(n_1439) );
CKINVDCx5p33_ASAP7_75t_R g955 ( .A(n_172), .Y(n_955) );
INVx1_ASAP7_75t_L g1664 ( .A(n_174), .Y(n_1664) );
INVx1_ASAP7_75t_L g1016 ( .A(n_175), .Y(n_1016) );
OAI22xp5_ASAP7_75t_L g1140 ( .A1(n_176), .A2(n_254), .B1(n_569), .B2(n_908), .Y(n_1140) );
OAI211xp5_ASAP7_75t_L g1142 ( .A1(n_176), .A2(n_950), .B(n_1143), .C(n_1148), .Y(n_1142) );
AOI22xp5_ASAP7_75t_L g1447 ( .A1(n_177), .A2(n_224), .B1(n_1430), .B2(n_1440), .Y(n_1447) );
CKINVDCx5p33_ASAP7_75t_R g1095 ( .A(n_179), .Y(n_1095) );
XOR2x2_ASAP7_75t_L g501 ( .A(n_180), .B(n_502), .Y(n_501) );
AOI22xp33_ASAP7_75t_L g1448 ( .A1(n_183), .A2(n_188), .B1(n_1437), .B2(n_1449), .Y(n_1448) );
AOI22xp33_ASAP7_75t_L g1312 ( .A1(n_184), .A2(n_248), .B1(n_803), .B2(n_878), .Y(n_1312) );
AOI22xp33_ASAP7_75t_SL g1330 ( .A1(n_184), .A2(n_265), .B1(n_525), .B2(n_1331), .Y(n_1330) );
AOI22xp33_ASAP7_75t_SL g1649 ( .A1(n_185), .A2(n_238), .B1(n_525), .B2(n_985), .Y(n_1649) );
AOI22xp33_ASAP7_75t_SL g1669 ( .A1(n_185), .A2(n_243), .B1(n_594), .B2(n_1110), .Y(n_1669) );
AOI221xp5_ASAP7_75t_L g1057 ( .A1(n_186), .A2(n_257), .B1(n_588), .B2(n_630), .C(n_771), .Y(n_1057) );
INVx1_ASAP7_75t_L g1273 ( .A(n_187), .Y(n_1273) );
INVx1_ASAP7_75t_L g992 ( .A(n_189), .Y(n_992) );
AOI22xp33_ASAP7_75t_L g1004 ( .A1(n_189), .A2(n_242), .B1(n_803), .B2(n_1005), .Y(n_1004) );
OAI211xp5_ASAP7_75t_L g429 ( .A1(n_190), .A2(n_405), .B(n_430), .C(n_434), .Y(n_429) );
INVx1_ASAP7_75t_L g489 ( .A(n_190), .Y(n_489) );
INVx1_ASAP7_75t_L g920 ( .A(n_191), .Y(n_920) );
INVx1_ASAP7_75t_L g924 ( .A(n_192), .Y(n_924) );
CKINVDCx5p33_ASAP7_75t_R g811 ( .A(n_193), .Y(n_811) );
OAI22xp5_ASAP7_75t_L g1235 ( .A1(n_194), .A2(n_307), .B1(n_550), .B2(n_1236), .Y(n_1235) );
INVx1_ASAP7_75t_L g1244 ( .A(n_194), .Y(n_1244) );
INVx1_ASAP7_75t_L g970 ( .A(n_195), .Y(n_970) );
CKINVDCx5p33_ASAP7_75t_R g1321 ( .A(n_196), .Y(n_1321) );
INVx2_ASAP7_75t_L g375 ( .A(n_197), .Y(n_375) );
INVx1_ASAP7_75t_L g414 ( .A(n_197), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_197), .B(n_376), .Y(n_549) );
AOI22xp5_ASAP7_75t_L g1477 ( .A1(n_198), .A2(n_300), .B1(n_1430), .B2(n_1437), .Y(n_1477) );
OAI211xp5_ASAP7_75t_L g1286 ( .A1(n_199), .A2(n_578), .B(n_1287), .C(n_1293), .Y(n_1286) );
INVx1_ASAP7_75t_L g1357 ( .A(n_200), .Y(n_1357) );
AO22x1_ASAP7_75t_L g1633 ( .A1(n_200), .A2(n_1634), .B1(n_1637), .B2(n_1671), .Y(n_1633) );
INVx1_ASAP7_75t_L g961 ( .A(n_201), .Y(n_961) );
INVx1_ASAP7_75t_L g368 ( .A(n_202), .Y(n_368) );
INVx1_ASAP7_75t_L g991 ( .A(n_203), .Y(n_991) );
INVx1_ASAP7_75t_L g1274 ( .A(n_205), .Y(n_1274) );
INVx1_ASAP7_75t_L g937 ( .A(n_206), .Y(n_937) );
OAI22xp5_ASAP7_75t_L g1322 ( .A1(n_207), .A2(n_272), .B1(n_1318), .B2(n_1323), .Y(n_1322) );
INVx1_ASAP7_75t_L g1341 ( .A(n_207), .Y(n_1341) );
BUFx3_ASAP7_75t_L g381 ( .A(n_209), .Y(n_381) );
AOI221xp5_ASAP7_75t_L g1240 ( .A1(n_210), .A2(n_216), .B1(n_586), .B2(n_592), .C(n_772), .Y(n_1240) );
AOI22xp33_ASAP7_75t_L g900 ( .A1(n_211), .A2(n_244), .B1(n_529), .B2(n_901), .Y(n_900) );
INVx1_ASAP7_75t_L g1051 ( .A(n_213), .Y(n_1051) );
CKINVDCx5p33_ASAP7_75t_R g750 ( .A(n_214), .Y(n_750) );
OAI22xp5_ASAP7_75t_L g1262 ( .A1(n_215), .A2(n_217), .B1(n_508), .B2(n_1263), .Y(n_1262) );
OAI221xp5_ASAP7_75t_L g1283 ( .A1(n_215), .A2(n_217), .B1(n_608), .B2(n_1185), .C(n_1284), .Y(n_1283) );
AOI22xp33_ASAP7_75t_SL g1220 ( .A1(n_216), .A2(n_258), .B1(n_529), .B2(n_1076), .Y(n_1220) );
AOI21xp33_ASAP7_75t_L g875 ( .A1(n_219), .A2(n_772), .B(n_876), .Y(n_875) );
INVx1_ASAP7_75t_L g893 ( .A(n_219), .Y(n_893) );
AOI22xp5_ASAP7_75t_L g1258 ( .A1(n_220), .A2(n_1259), .B1(n_1260), .B2(n_1301), .Y(n_1258) );
INVx1_ASAP7_75t_L g1301 ( .A(n_220), .Y(n_1301) );
AOI21xp33_ASAP7_75t_L g766 ( .A1(n_221), .A2(n_701), .B(n_702), .Y(n_766) );
XOR2x2_ASAP7_75t_L g846 ( .A(n_222), .B(n_847), .Y(n_846) );
CKINVDCx5p33_ASAP7_75t_R g1371 ( .A(n_223), .Y(n_1371) );
NAND2xp5_ASAP7_75t_L g1210 ( .A(n_224), .B(n_1211), .Y(n_1210) );
AOI22xp5_ASAP7_75t_L g1230 ( .A1(n_224), .A2(n_1231), .B1(n_1232), .B2(n_1254), .Y(n_1230) );
INVx1_ASAP7_75t_L g1256 ( .A(n_224), .Y(n_1256) );
OAI22xp33_ASAP7_75t_L g1136 ( .A1(n_225), .A2(n_237), .B1(n_543), .B2(n_550), .Y(n_1136) );
INVx1_ASAP7_75t_L g1149 ( .A(n_225), .Y(n_1149) );
BUFx3_ASAP7_75t_L g338 ( .A(n_227), .Y(n_338) );
INVx1_ASAP7_75t_L g467 ( .A(n_227), .Y(n_467) );
AOI22xp33_ASAP7_75t_L g834 ( .A1(n_228), .A2(n_278), .B1(n_525), .B2(n_697), .Y(n_834) );
XNOR2x1_ASAP7_75t_L g1027 ( .A(n_229), .B(n_1028), .Y(n_1027) );
NAND2xp5_ASAP7_75t_SL g868 ( .A(n_230), .B(n_772), .Y(n_868) );
CKINVDCx5p33_ASAP7_75t_R g755 ( .A(n_231), .Y(n_755) );
INVx1_ASAP7_75t_L g1050 ( .A(n_234), .Y(n_1050) );
CKINVDCx5p33_ASAP7_75t_R g1229 ( .A(n_235), .Y(n_1229) );
INVx1_ASAP7_75t_L g1127 ( .A(n_236), .Y(n_1127) );
INVx1_ASAP7_75t_L g1150 ( .A(n_237), .Y(n_1150) );
INVx1_ASAP7_75t_L g934 ( .A(n_239), .Y(n_934) );
INVx1_ASAP7_75t_L g1205 ( .A(n_240), .Y(n_1205) );
INVx1_ASAP7_75t_L g1663 ( .A(n_241), .Y(n_1663) );
NAND2xp33_ASAP7_75t_SL g986 ( .A(n_242), .B(n_987), .Y(n_986) );
NAND2xp5_ASAP7_75t_SL g871 ( .A(n_244), .B(n_872), .Y(n_871) );
INVx1_ASAP7_75t_L g737 ( .A(n_246), .Y(n_737) );
XNOR2x2_ASAP7_75t_L g1121 ( .A(n_247), .B(n_1122), .Y(n_1121) );
AOI22xp33_ASAP7_75t_SL g1327 ( .A1(n_248), .A2(n_311), .B1(n_525), .B2(n_985), .Y(n_1327) );
INVx1_ASAP7_75t_L g1281 ( .A(n_249), .Y(n_1281) );
INVx1_ASAP7_75t_L g383 ( .A(n_250), .Y(n_383) );
INVx1_ASAP7_75t_L g390 ( .A(n_250), .Y(n_390) );
INVx1_ASAP7_75t_L g600 ( .A(n_251), .Y(n_600) );
CKINVDCx5p33_ASAP7_75t_R g1367 ( .A(n_252), .Y(n_1367) );
INVx1_ASAP7_75t_L g1013 ( .A(n_255), .Y(n_1013) );
INVx1_ASAP7_75t_L g1414 ( .A(n_259), .Y(n_1414) );
OAI21xp33_ASAP7_75t_L g880 ( .A1(n_260), .A2(n_881), .B(n_884), .Y(n_880) );
AOI22xp5_ASAP7_75t_SL g1472 ( .A1(n_261), .A2(n_308), .B1(n_1440), .B2(n_1449), .Y(n_1472) );
INVx1_ASAP7_75t_L g666 ( .A(n_262), .Y(n_666) );
AOI21xp33_ASAP7_75t_L g1250 ( .A1(n_263), .A2(n_630), .B(n_1251), .Y(n_1250) );
CKINVDCx5p33_ASAP7_75t_R g1034 ( .A(n_264), .Y(n_1034) );
AOI221xp5_ASAP7_75t_SL g1315 ( .A1(n_265), .A2(n_311), .B1(n_483), .B2(n_628), .C(n_1003), .Y(n_1315) );
INVx1_ASAP7_75t_L g1654 ( .A(n_266), .Y(n_1654) );
INVx1_ASAP7_75t_L g1433 ( .A(n_267), .Y(n_1433) );
AND2x2_ASAP7_75t_L g1441 ( .A(n_267), .B(n_1439), .Y(n_1441) );
INVxp67_ASAP7_75t_SL g1189 ( .A(n_268), .Y(n_1189) );
INVx1_ASAP7_75t_L g441 ( .A(n_270), .Y(n_441) );
OAI211xp5_ASAP7_75t_L g479 ( .A1(n_270), .A2(n_330), .B(n_480), .C(n_485), .Y(n_479) );
INVx1_ASAP7_75t_L g1295 ( .A(n_271), .Y(n_1295) );
INVx1_ASAP7_75t_L g1335 ( .A(n_272), .Y(n_1335) );
XNOR2xp5_ASAP7_75t_L g738 ( .A(n_274), .B(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g322 ( .A(n_275), .Y(n_322) );
INVxp67_ASAP7_75t_SL g965 ( .A(n_276), .Y(n_965) );
INVxp67_ASAP7_75t_SL g1218 ( .A(n_277), .Y(n_1218) );
OAI211xp5_ASAP7_75t_L g1238 ( .A1(n_277), .A2(n_578), .B(n_1239), .C(n_1243), .Y(n_1238) );
NAND2xp5_ASAP7_75t_L g1158 ( .A(n_280), .B(n_1159), .Y(n_1158) );
INVx1_ASAP7_75t_L g741 ( .A(n_281), .Y(n_741) );
OAI21xp5_ASAP7_75t_SL g1059 ( .A1(n_282), .A2(n_841), .B(n_1060), .Y(n_1059) );
INVx1_ASAP7_75t_L g761 ( .A(n_283), .Y(n_761) );
INVx1_ASAP7_75t_L g355 ( .A(n_284), .Y(n_355) );
INVx1_ASAP7_75t_L g328 ( .A(n_285), .Y(n_328) );
CKINVDCx5p33_ASAP7_75t_R g1120 ( .A(n_286), .Y(n_1120) );
INVxp67_ASAP7_75t_SL g1187 ( .A(n_287), .Y(n_1187) );
AOI22xp33_ASAP7_75t_SL g1197 ( .A1(n_287), .A2(n_293), .B1(n_541), .B2(n_1198), .Y(n_1197) );
BUFx6f_ASAP7_75t_L g327 ( .A(n_288), .Y(n_327) );
INVx1_ASAP7_75t_L g833 ( .A(n_290), .Y(n_833) );
INVxp67_ASAP7_75t_SL g681 ( .A(n_295), .Y(n_681) );
OAI221xp5_ASAP7_75t_L g717 ( .A1(n_295), .A2(n_298), .B1(n_718), .B2(n_720), .C(n_722), .Y(n_717) );
INVx1_ASAP7_75t_L g839 ( .A(n_296), .Y(n_839) );
CKINVDCx5p33_ASAP7_75t_R g1365 ( .A(n_297), .Y(n_1365) );
OAI221xp5_ASAP7_75t_L g652 ( .A1(n_298), .A2(n_299), .B1(n_653), .B2(n_658), .C(n_659), .Y(n_652) );
INVx2_ASAP7_75t_L g336 ( .A(n_302), .Y(n_336) );
INVx1_ASAP7_75t_L g364 ( .A(n_302), .Y(n_364) );
INVx1_ASAP7_75t_L g413 ( .A(n_302), .Y(n_413) );
CKINVDCx5p33_ASAP7_75t_R g567 ( .A(n_303), .Y(n_567) );
INVx1_ASAP7_75t_L g775 ( .A(n_304), .Y(n_775) );
CKINVDCx5p33_ASAP7_75t_R g1298 ( .A(n_305), .Y(n_1298) );
OAI22xp33_ASAP7_75t_SL g1656 ( .A1(n_306), .A2(n_310), .B1(n_508), .B2(n_836), .Y(n_1656) );
OAI221xp5_ASAP7_75t_L g1665 ( .A1(n_306), .A2(n_310), .B1(n_608), .B2(n_809), .C(n_1666), .Y(n_1665) );
INVx1_ASAP7_75t_L g1245 ( .A(n_307), .Y(n_1245) );
INVxp67_ASAP7_75t_SL g744 ( .A(n_309), .Y(n_744) );
A2O1A1Ixp33_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_911), .B(n_1352), .C(n_1677), .Y(n_312) );
OAI21xp33_ASAP7_75t_L g1352 ( .A1(n_313), .A2(n_911), .B(n_1353), .Y(n_1352) );
AOI22xp33_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_790), .B1(n_791), .B2(n_910), .Y(n_313) );
INVx1_ASAP7_75t_L g910 ( .A(n_314), .Y(n_910) );
AOI22xp5_ASAP7_75t_L g314 ( .A1(n_315), .A2(n_316), .B1(n_634), .B2(n_789), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
OA22x2_ASAP7_75t_L g316 ( .A1(n_317), .A2(n_500), .B1(n_501), .B2(n_633), .Y(n_316) );
INVx1_ASAP7_75t_L g633 ( .A(n_317), .Y(n_633) );
NAND3xp33_ASAP7_75t_L g318 ( .A(n_319), .B(n_419), .C(n_456), .Y(n_318) );
NOR2xp33_ASAP7_75t_L g319 ( .A(n_320), .B(n_370), .Y(n_319) );
OAI33xp33_ASAP7_75t_L g320 ( .A1(n_321), .A2(n_333), .A3(n_339), .B1(n_354), .B2(n_357), .B3(n_367), .Y(n_320) );
OAI22xp5_ASAP7_75t_L g321 ( .A1(n_322), .A2(n_323), .B1(n_328), .B2(n_329), .Y(n_321) );
OAI22xp5_ASAP7_75t_L g392 ( .A1(n_322), .A2(n_355), .B1(n_393), .B2(n_398), .Y(n_392) );
OAI22xp5_ASAP7_75t_L g367 ( .A1(n_323), .A2(n_347), .B1(n_368), .B2(n_369), .Y(n_367) );
BUFx2_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
BUFx3_ASAP7_75t_L g647 ( .A(n_324), .Y(n_647) );
BUFx2_ASAP7_75t_L g1370 ( .A(n_324), .Y(n_1370) );
INVx2_ASAP7_75t_L g1375 ( .A(n_324), .Y(n_1375) );
OR2x2_ASAP7_75t_L g324 ( .A(n_325), .B(n_326), .Y(n_324) );
NAND2x1_ASAP7_75t_L g332 ( .A(n_325), .B(n_327), .Y(n_332) );
OR2x2_ASAP7_75t_L g345 ( .A(n_325), .B(n_327), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_325), .B(n_353), .Y(n_352) );
INVx2_ASAP7_75t_L g469 ( .A(n_325), .Y(n_469) );
AND2x2_ASAP7_75t_L g484 ( .A(n_325), .B(n_327), .Y(n_484) );
BUFx2_ASAP7_75t_L g488 ( .A(n_325), .Y(n_488) );
INVx1_ASAP7_75t_L g566 ( .A(n_325), .Y(n_566) );
AND2x2_ASAP7_75t_L g581 ( .A(n_325), .B(n_353), .Y(n_581) );
AND2x2_ASAP7_75t_L g565 ( .A(n_326), .B(n_566), .Y(n_565) );
HB1xp67_ASAP7_75t_L g864 ( .A(n_326), .Y(n_864) );
INVx2_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx2_ASAP7_75t_L g353 ( .A(n_327), .Y(n_353) );
AND2x2_ASAP7_75t_L g468 ( .A(n_327), .B(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g494 ( .A(n_327), .Y(n_494) );
OAI22xp5_ASAP7_75t_L g402 ( .A1(n_328), .A2(n_356), .B1(n_403), .B2(n_405), .Y(n_402) );
HB1xp67_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
OAI22xp33_ASAP7_75t_L g354 ( .A1(n_330), .A2(n_341), .B1(n_355), .B2(n_356), .Y(n_354) );
BUFx6f_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
BUFx4f_ASAP7_75t_L g649 ( .A(n_331), .Y(n_649) );
OR2x6_ASAP7_75t_L g659 ( .A(n_331), .B(n_660), .Y(n_659) );
INVx4_ASAP7_75t_L g858 ( .A(n_331), .Y(n_858) );
BUFx4f_ASAP7_75t_L g1323 ( .A(n_331), .Y(n_1323) );
BUFx6f_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
BUFx3_ASAP7_75t_L g680 ( .A(n_332), .Y(n_680) );
OAI33xp33_ASAP7_75t_L g1361 ( .A1(n_333), .A2(n_1362), .A3(n_1366), .B1(n_1372), .B2(n_1379), .B3(n_1383), .Y(n_1361) );
INVx2_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
OAI221xp5_ASAP7_75t_L g664 ( .A1(n_334), .A2(n_647), .B1(n_649), .B2(n_665), .C(n_666), .Y(n_664) );
HB1xp67_ASAP7_75t_L g777 ( .A(n_334), .Y(n_777) );
AND2x4_ASAP7_75t_L g334 ( .A(n_335), .B(n_337), .Y(n_334) );
INVx1_ASAP7_75t_L g952 ( .A(n_335), .Y(n_952) );
OR2x2_ASAP7_75t_L g1040 ( .A(n_335), .B(n_695), .Y(n_1040) );
OR2x6_ASAP7_75t_L g1333 ( .A(n_335), .B(n_695), .Y(n_1333) );
BUFx2_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx2_ASAP7_75t_L g523 ( .A(n_336), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_336), .B(n_564), .Y(n_655) );
AND2x4_ASAP7_75t_L g365 ( .A(n_338), .B(n_366), .Y(n_365) );
INVx2_ASAP7_75t_L g463 ( .A(n_338), .Y(n_463) );
BUFx2_ASAP7_75t_L g478 ( .A(n_338), .Y(n_478) );
AND2x4_ASAP7_75t_L g492 ( .A(n_338), .B(n_493), .Y(n_492) );
OAI22xp5_ASAP7_75t_L g339 ( .A1(n_340), .A2(n_341), .B1(n_346), .B2(n_347), .Y(n_339) );
OAI22xp33_ASAP7_75t_L g377 ( .A1(n_340), .A2(n_368), .B1(n_378), .B2(n_384), .Y(n_377) );
OAI221xp5_ASAP7_75t_L g1186 ( .A1(n_341), .A2(n_1187), .B1(n_1188), .B2(n_1189), .C(n_1190), .Y(n_1186) );
INVx2_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx2_ASAP7_75t_SL g342 ( .A(n_343), .Y(n_342) );
BUFx6f_ASAP7_75t_L g644 ( .A(n_343), .Y(n_644) );
OAI22xp5_ASAP7_75t_L g773 ( .A1(n_343), .A2(n_774), .B1(n_775), .B2(n_776), .Y(n_773) );
OAI22x1_ASAP7_75t_SL g779 ( .A1(n_343), .A2(n_755), .B1(n_776), .B2(n_780), .Y(n_779) );
BUFx3_ASAP7_75t_L g1012 ( .A(n_343), .Y(n_1012) );
INVx3_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx2_ASAP7_75t_L g461 ( .A(n_344), .Y(n_461) );
BUFx4f_ASAP7_75t_L g619 ( .A(n_344), .Y(n_619) );
INVx3_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
OAI22xp5_ASAP7_75t_L g415 ( .A1(n_346), .A2(n_369), .B1(n_416), .B2(n_418), .Y(n_415) );
INVx2_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx4_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx2_ASAP7_75t_L g622 ( .A(n_350), .Y(n_622) );
INVx2_ASAP7_75t_L g776 ( .A(n_350), .Y(n_776) );
INVx2_ASAP7_75t_SL g936 ( .A(n_350), .Y(n_936) );
INVx1_ASAP7_75t_L g1015 ( .A(n_350), .Y(n_1015) );
BUFx6f_ASAP7_75t_L g1154 ( .A(n_350), .Y(n_1154) );
INVx8_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
OR2x2_ASAP7_75t_L g477 ( .A(n_351), .B(n_478), .Y(n_477) );
BUFx2_ASAP7_75t_L g663 ( .A(n_351), .Y(n_663) );
BUFx6f_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx2_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_360), .B(n_365), .Y(n_359) );
AND2x4_ASAP7_75t_L g781 ( .A(n_360), .B(n_365), .Y(n_781) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
OR2x2_ASAP7_75t_L g373 ( .A(n_362), .B(n_374), .Y(n_373) );
HB1xp67_ASAP7_75t_L g455 ( .A(n_362), .Y(n_455) );
OR2x2_ASAP7_75t_L g548 ( .A(n_362), .B(n_549), .Y(n_548) );
AND2x2_ASAP7_75t_SL g651 ( .A(n_362), .B(n_365), .Y(n_651) );
INVx2_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
BUFx2_ASAP7_75t_L g499 ( .A(n_363), .Y(n_499) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx4_ASAP7_75t_L g592 ( .A(n_365), .Y(n_592) );
NAND4xp25_ASAP7_75t_L g867 ( .A(n_365), .B(n_868), .C(n_869), .D(n_871), .Y(n_867) );
INVx4_ASAP7_75t_L g1003 ( .A(n_365), .Y(n_1003) );
INVx1_ASAP7_75t_SL g1181 ( .A(n_365), .Y(n_1181) );
INVx1_ASAP7_75t_L g497 ( .A(n_366), .Y(n_497) );
AND2x4_ASAP7_75t_L g631 ( .A(n_366), .B(n_463), .Y(n_631) );
OAI33xp33_ASAP7_75t_L g370 ( .A1(n_371), .A2(n_377), .A3(n_392), .B1(n_402), .B2(n_407), .B3(n_415), .Y(n_370) );
BUFx3_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
OAI22xp5_ASAP7_75t_SL g1645 ( .A1(n_372), .A2(n_1646), .B1(n_1650), .B2(n_1651), .Y(n_1645) );
BUFx4f_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
BUFx8_ASAP7_75t_L g820 ( .A(n_373), .Y(n_820) );
BUFx2_ASAP7_75t_L g890 ( .A(n_373), .Y(n_890) );
BUFx4f_ASAP7_75t_L g981 ( .A(n_373), .Y(n_981) );
BUFx2_ASAP7_75t_L g702 ( .A(n_374), .Y(n_702) );
NAND2xp33_ASAP7_75t_SL g374 ( .A(n_375), .B(n_376), .Y(n_374) );
HB1xp67_ASAP7_75t_L g453 ( .A(n_375), .Y(n_453) );
INVx1_ASAP7_75t_L g514 ( .A(n_375), .Y(n_514) );
AND3x4_ASAP7_75t_L g522 ( .A(n_375), .B(n_439), .C(n_523), .Y(n_522) );
AND2x2_ASAP7_75t_L g1407 ( .A(n_375), .B(n_439), .Y(n_1407) );
INVx3_ASAP7_75t_L g411 ( .A(n_376), .Y(n_411) );
BUFx3_ASAP7_75t_L g439 ( .A(n_376), .Y(n_439) );
HB1xp67_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g417 ( .A(n_379), .Y(n_417) );
BUFx4f_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
OR2x4_ASAP7_75t_L g423 ( .A(n_380), .B(n_424), .Y(n_423) );
OR2x4_ASAP7_75t_L g448 ( .A(n_380), .B(n_411), .Y(n_448) );
INVx2_ASAP7_75t_L g545 ( .A(n_380), .Y(n_545) );
BUFx3_ASAP7_75t_L g1396 ( .A(n_380), .Y(n_1396) );
BUFx3_ASAP7_75t_L g1410 ( .A(n_380), .Y(n_1410) );
OR2x2_ASAP7_75t_L g380 ( .A(n_381), .B(n_382), .Y(n_380) );
BUFx6f_ASAP7_75t_L g391 ( .A(n_381), .Y(n_391) );
INVx2_ASAP7_75t_L g397 ( .A(n_381), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_381), .B(n_390), .Y(n_401) );
AND2x4_ASAP7_75t_L g432 ( .A(n_381), .B(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g528 ( .A(n_382), .Y(n_528) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVxp67_ASAP7_75t_L g396 ( .A(n_383), .Y(n_396) );
INVx2_ASAP7_75t_SL g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
BUFx6f_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
OR2x2_ASAP7_75t_L g572 ( .A(n_387), .B(n_548), .Y(n_572) );
INVx3_ASAP7_75t_L g765 ( .A(n_387), .Y(n_765) );
BUFx6f_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
BUFx3_ASAP7_75t_L g406 ( .A(n_388), .Y(n_406) );
BUFx2_ASAP7_75t_L g723 ( .A(n_388), .Y(n_723) );
NAND2x1p5_ASAP7_75t_L g388 ( .A(n_389), .B(n_391), .Y(n_388) );
BUFx2_ASAP7_75t_L g444 ( .A(n_389), .Y(n_444) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx2_ASAP7_75t_L g433 ( .A(n_390), .Y(n_433) );
BUFx2_ASAP7_75t_L g440 ( .A(n_391), .Y(n_440) );
INVx2_ASAP7_75t_L g510 ( .A(n_391), .Y(n_510) );
AND2x4_ASAP7_75t_L g535 ( .A(n_391), .B(n_520), .Y(n_535) );
INVx1_ASAP7_75t_L g1200 ( .A(n_393), .Y(n_1200) );
INVx2_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
BUFx6f_ASAP7_75t_L g404 ( .A(n_394), .Y(n_404) );
AND2x4_ASAP7_75t_L g450 ( .A(n_394), .B(n_424), .Y(n_450) );
INVx2_ASAP7_75t_L g959 ( .A(n_394), .Y(n_959) );
BUFx6f_ASAP7_75t_L g1042 ( .A(n_394), .Y(n_1042) );
INVx2_ASAP7_75t_L g1652 ( .A(n_394), .Y(n_1652) );
BUFx6f_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
BUFx8_ASAP7_75t_L g533 ( .A(n_395), .Y(n_533) );
INVx2_ASAP7_75t_L g692 ( .A(n_395), .Y(n_692) );
BUFx6f_ASAP7_75t_L g701 ( .A(n_395), .Y(n_701) );
AND2x4_ASAP7_75t_L g395 ( .A(n_396), .B(n_397), .Y(n_395) );
AND2x4_ASAP7_75t_L g527 ( .A(n_397), .B(n_528), .Y(n_527) );
OAI22xp33_ASAP7_75t_L g1267 ( .A1(n_398), .A2(n_962), .B1(n_1268), .B2(n_1269), .Y(n_1267) );
OAI22xp5_ASAP7_75t_L g1275 ( .A1(n_398), .A2(n_1276), .B1(n_1277), .B2(n_1278), .Y(n_1275) );
INVx3_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx3_ASAP7_75t_L g418 ( .A(n_399), .Y(n_418) );
CKINVDCx8_ASAP7_75t_R g832 ( .A(n_399), .Y(n_832) );
BUFx6f_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g561 ( .A(n_400), .Y(n_561) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
BUFx2_ASAP7_75t_L g428 ( .A(n_401), .Y(n_428) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
BUFx6f_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
OAI221xp5_ASAP7_75t_L g1405 ( .A1(n_406), .A2(n_1371), .B1(n_1376), .B2(n_1406), .C(n_1407), .Y(n_1405) );
OAI221xp5_ASAP7_75t_L g1409 ( .A1(n_406), .A2(n_759), .B1(n_1365), .B2(n_1378), .C(n_1410), .Y(n_1409) );
OAI33xp33_ASAP7_75t_L g1266 ( .A1(n_407), .A2(n_820), .A3(n_1267), .B1(n_1270), .B2(n_1275), .B3(n_1279), .Y(n_1266) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
NAND3xp33_ASAP7_75t_L g1079 ( .A(n_408), .B(n_1080), .C(n_1083), .Y(n_1079) );
AOI33xp33_ASAP7_75t_L g1196 ( .A1(n_408), .A2(n_522), .A3(n_1197), .B1(n_1199), .B2(n_1201), .B3(n_1202), .Y(n_1196) );
BUFx2_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
BUFx2_ASAP7_75t_L g537 ( .A(n_409), .Y(n_537) );
BUFx2_ASAP7_75t_L g1227 ( .A(n_409), .Y(n_1227) );
INVx3_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx3_ASAP7_75t_L g830 ( .A(n_410), .Y(n_830) );
NAND3x1_ASAP7_75t_L g410 ( .A(n_411), .B(n_412), .C(n_414), .Y(n_410) );
INVx1_ASAP7_75t_L g424 ( .A(n_411), .Y(n_424) );
OR2x6_ASAP7_75t_L g427 ( .A(n_411), .B(n_428), .Y(n_427) );
AND2x4_ASAP7_75t_L g431 ( .A(n_411), .B(n_432), .Y(n_431) );
AND2x4_ASAP7_75t_L g513 ( .A(n_411), .B(n_514), .Y(n_513) );
NAND2x1p5_ASAP7_75t_L g695 ( .A(n_411), .B(n_414), .Y(n_695) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g512 ( .A(n_413), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_413), .B(n_582), .Y(n_674) );
OAI22xp33_ASAP7_75t_L g960 ( .A1(n_416), .A2(n_944), .B1(n_961), .B2(n_962), .Y(n_960) );
INVx2_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
OAI221xp5_ASAP7_75t_L g891 ( .A1(n_418), .A2(n_892), .B1(n_893), .B2(n_894), .C(n_895), .Y(n_891) );
OAI22xp5_ASAP7_75t_L g957 ( .A1(n_418), .A2(n_934), .B1(n_958), .B2(n_959), .Y(n_957) );
OAI22xp5_ASAP7_75t_L g1411 ( .A1(n_418), .A2(n_1367), .B1(n_1382), .B2(n_1412), .Y(n_1411) );
OAI31xp33_ASAP7_75t_L g419 ( .A1(n_420), .A2(n_429), .A3(n_445), .B(n_451), .Y(n_419) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx2_ASAP7_75t_SL g422 ( .A(n_423), .Y(n_422) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g827 ( .A(n_428), .Y(n_827) );
BUFx3_ASAP7_75t_L g966 ( .A(n_428), .Y(n_966) );
CKINVDCx8_ASAP7_75t_R g430 ( .A(n_431), .Y(n_430) );
BUFx3_ASAP7_75t_L g529 ( .A(n_432), .Y(n_529) );
BUFx2_ASAP7_75t_L g556 ( .A(n_432), .Y(n_556) );
INVx2_ASAP7_75t_L g698 ( .A(n_432), .Y(n_698) );
AND2x2_ASAP7_75t_L g712 ( .A(n_432), .B(n_710), .Y(n_712) );
BUFx2_ASAP7_75t_L g985 ( .A(n_432), .Y(n_985) );
BUFx2_ASAP7_75t_L g1039 ( .A(n_432), .Y(n_1039) );
BUFx2_ASAP7_75t_L g1198 ( .A(n_432), .Y(n_1198) );
INVx1_ASAP7_75t_L g520 ( .A(n_433), .Y(n_520) );
AOI22xp33_ASAP7_75t_L g434 ( .A1(n_435), .A2(n_436), .B1(n_441), .B2(n_442), .Y(n_434) );
AOI22xp33_ASAP7_75t_L g485 ( .A1(n_435), .A2(n_486), .B1(n_489), .B2(n_490), .Y(n_485) );
BUFx3_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_438), .B(n_440), .Y(n_437) );
AND2x4_ASAP7_75t_L g443 ( .A(n_438), .B(n_444), .Y(n_443) );
INVx3_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
BUFx6f_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
AND2x2_ASAP7_75t_SL g451 ( .A(n_452), .B(n_454), .Y(n_451) );
INVx1_ASAP7_75t_SL g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
OAI31xp33_ASAP7_75t_SL g456 ( .A1(n_457), .A2(n_470), .A3(n_479), .B(n_495), .Y(n_456) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
AND2x4_ASAP7_75t_SL g1415 ( .A(n_459), .B(n_1416), .Y(n_1415) );
NAND2xp5_ASAP7_75t_L g1683 ( .A(n_459), .B(n_1684), .Y(n_1683) );
INVx3_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
OR2x6_ASAP7_75t_L g460 ( .A(n_461), .B(n_462), .Y(n_460) );
OR2x6_ASAP7_75t_L g472 ( .A(n_461), .B(n_466), .Y(n_472) );
INVxp67_ASAP7_75t_L g1159 ( .A(n_461), .Y(n_1159) );
BUFx4f_ASAP7_75t_L g1364 ( .A(n_461), .Y(n_1364) );
INVxp67_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g482 ( .A(n_463), .Y(n_482) );
INVx3_ASAP7_75t_SL g464 ( .A(n_465), .Y(n_464) );
AND2x4_ASAP7_75t_L g465 ( .A(n_466), .B(n_468), .Y(n_465) );
HB1xp67_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
BUFx6f_ASAP7_75t_L g590 ( .A(n_468), .Y(n_590) );
INVx2_ASAP7_75t_L g629 ( .A(n_468), .Y(n_629) );
BUFx3_ASAP7_75t_L g772 ( .A(n_468), .Y(n_772) );
HB1xp67_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx2_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
AND2x4_ASAP7_75t_L g487 ( .A(n_478), .B(n_488), .Y(n_487) );
INVx3_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_482), .B(n_483), .Y(n_481) );
BUFx6f_ASAP7_75t_L g586 ( .A(n_483), .Y(n_586) );
AND2x6_ASAP7_75t_L g598 ( .A(n_483), .B(n_564), .Y(n_598) );
AND2x4_ASAP7_75t_SL g611 ( .A(n_483), .B(n_582), .Y(n_611) );
BUFx3_ASAP7_75t_L g625 ( .A(n_483), .Y(n_625) );
BUFx3_ASAP7_75t_L g771 ( .A(n_483), .Y(n_771) );
BUFx3_ASAP7_75t_L g872 ( .A(n_483), .Y(n_872) );
INVx1_ASAP7_75t_L g1113 ( .A(n_483), .Y(n_1113) );
BUFx6f_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g1021 ( .A(n_484), .Y(n_1021) );
BUFx3_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g614 ( .A(n_488), .Y(n_614) );
INVx1_ASAP7_75t_L g657 ( .A(n_488), .Y(n_657) );
BUFx2_ASAP7_75t_L g861 ( .A(n_488), .Y(n_861) );
INVx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_493), .B(n_564), .Y(n_571) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
BUFx3_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
AND2x4_ASAP7_75t_L g496 ( .A(n_497), .B(n_498), .Y(n_496) );
NOR2xp33_ASAP7_75t_L g1416 ( .A(n_497), .B(n_1417), .Y(n_1416) );
INVx1_ASAP7_75t_L g1684 ( .A(n_497), .Y(n_1684) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
OR2x2_ASAP7_75t_L g570 ( .A(n_499), .B(n_571), .Y(n_570) );
INVxp67_ASAP7_75t_L g575 ( .A(n_499), .Y(n_575) );
OR2x2_ASAP7_75t_L g658 ( .A(n_499), .B(n_571), .Y(n_658) );
INVx1_ASAP7_75t_L g687 ( .A(n_499), .Y(n_687) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
NAND3xp33_ASAP7_75t_L g502 ( .A(n_503), .B(n_557), .C(n_576), .Y(n_502) );
NOR3xp33_ASAP7_75t_L g503 ( .A(n_504), .B(n_542), .C(n_553), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_505), .B(n_521), .Y(n_504) );
AOI22xp33_ASAP7_75t_L g505 ( .A1(n_506), .A2(n_507), .B1(n_515), .B2(n_516), .Y(n_505) );
AOI221x1_ASAP7_75t_L g888 ( .A1(n_507), .A2(n_516), .B1(n_851), .B2(n_860), .C(n_889), .Y(n_888) );
AOI22xp5_ASAP7_75t_L g1214 ( .A1(n_507), .A2(n_516), .B1(n_1215), .B2(n_1216), .Y(n_1214) );
INVx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
NAND2x1_ASAP7_75t_L g508 ( .A(n_509), .B(n_511), .Y(n_508) );
AND2x6_ASAP7_75t_L g719 ( .A(n_509), .B(n_513), .Y(n_719) );
AND2x2_ASAP7_75t_L g921 ( .A(n_509), .B(n_511), .Y(n_921) );
AND2x2_ASAP7_75t_L g996 ( .A(n_509), .B(n_511), .Y(n_996) );
AND2x4_ASAP7_75t_SL g1035 ( .A(n_509), .B(n_511), .Y(n_1035) );
INVx3_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
AND2x4_ASAP7_75t_L g516 ( .A(n_511), .B(n_517), .Y(n_516) );
AND2x4_ASAP7_75t_L g555 ( .A(n_511), .B(n_556), .Y(n_555) );
AND2x4_ASAP7_75t_SL g837 ( .A(n_511), .B(n_517), .Y(n_837) );
AND2x4_ASAP7_75t_L g511 ( .A(n_512), .B(n_513), .Y(n_511) );
OR2x2_ASAP7_75t_L g562 ( .A(n_512), .B(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g669 ( .A(n_512), .Y(n_669) );
NAND2x1p5_ASAP7_75t_L g574 ( .A(n_513), .B(n_527), .Y(n_574) );
AND2x2_ASAP7_75t_L g721 ( .A(n_513), .B(n_519), .Y(n_721) );
INVx1_ASAP7_75t_L g724 ( .A(n_513), .Y(n_724) );
AOI22xp33_ASAP7_75t_L g919 ( .A1(n_516), .A2(n_920), .B1(n_921), .B2(n_922), .Y(n_919) );
AOI22xp33_ASAP7_75t_L g1089 ( .A1(n_516), .A2(n_921), .B1(n_1090), .B2(n_1091), .Y(n_1089) );
AOI22xp33_ASAP7_75t_L g1125 ( .A1(n_516), .A2(n_921), .B1(n_1126), .B2(n_1127), .Y(n_1125) );
AOI22xp33_ASAP7_75t_L g1204 ( .A1(n_516), .A2(n_996), .B1(n_1205), .B2(n_1206), .Y(n_1204) );
HB1xp67_ASAP7_75t_L g1264 ( .A(n_516), .Y(n_1264) );
INVx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
AOI33xp33_ASAP7_75t_L g521 ( .A1(n_522), .A2(n_524), .A3(n_530), .B1(n_536), .B2(n_537), .B3(n_538), .Y(n_521) );
INVx1_ASAP7_75t_L g1044 ( .A(n_522), .Y(n_1044) );
BUFx3_ASAP7_75t_L g1074 ( .A(n_522), .Y(n_1074) );
AOI33xp33_ASAP7_75t_L g1219 ( .A1(n_522), .A2(n_1220), .A3(n_1221), .B1(n_1224), .B2(n_1225), .B3(n_1227), .Y(n_1219) );
AOI33xp33_ASAP7_75t_L g1326 ( .A1(n_522), .A2(n_1327), .A3(n_1328), .B1(n_1329), .B2(n_1330), .B3(n_1332), .Y(n_1326) );
INVx2_ASAP7_75t_SL g632 ( .A(n_523), .Y(n_632) );
INVx1_ASAP7_75t_L g732 ( .A(n_523), .Y(n_732) );
OAI31xp33_ASAP7_75t_SL g745 ( .A1(n_523), .A2(n_746), .A3(n_747), .B(n_751), .Y(n_745) );
INVx8_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
CKINVDCx5p33_ASAP7_75t_R g757 ( .A(n_526), .Y(n_757) );
INVx2_ASAP7_75t_L g844 ( .A(n_526), .Y(n_844) );
INVx2_ASAP7_75t_L g968 ( .A(n_526), .Y(n_968) );
INVx3_ASAP7_75t_L g1226 ( .A(n_526), .Y(n_1226) );
INVx8_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
BUFx3_ASAP7_75t_L g541 ( .A(n_527), .Y(n_541) );
BUFx3_ASAP7_75t_L g705 ( .A(n_527), .Y(n_705) );
AND2x2_ASAP7_75t_L g709 ( .A(n_527), .B(n_710), .Y(n_709) );
HB1xp67_ASAP7_75t_L g901 ( .A(n_527), .Y(n_901) );
INVx1_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx3_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
AND2x4_ASAP7_75t_L g551 ( .A(n_533), .B(n_552), .Y(n_551) );
INVx2_ASAP7_75t_SL g822 ( .A(n_533), .Y(n_822) );
HB1xp67_ASAP7_75t_L g1071 ( .A(n_533), .Y(n_1071) );
INVx2_ASAP7_75t_SL g1276 ( .A(n_533), .Y(n_1276) );
INVx3_ASAP7_75t_L g1412 ( .A(n_533), .Y(n_1412) );
BUFx3_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
BUFx2_ASAP7_75t_L g693 ( .A(n_535), .Y(n_693) );
BUFx12f_ASAP7_75t_L g706 ( .A(n_535), .Y(n_706) );
AND2x4_ASAP7_75t_L g730 ( .A(n_535), .B(n_728), .Y(n_730) );
INVx5_ASAP7_75t_L g988 ( .A(n_535), .Y(n_988) );
BUFx3_ASAP7_75t_L g1072 ( .A(n_535), .Y(n_1072) );
AOI33xp33_ASAP7_75t_L g1128 ( .A1(n_537), .A2(n_1074), .A3(n_1129), .B1(n_1130), .B2(n_1133), .B3(n_1135), .Y(n_1128) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx2_ASAP7_75t_SL g1077 ( .A(n_541), .Y(n_1077) );
NAND2xp5_ASAP7_75t_L g904 ( .A(n_543), .B(n_685), .Y(n_904) );
OR2x6_ASAP7_75t_L g543 ( .A(n_544), .B(n_546), .Y(n_543) );
OR2x2_ASAP7_75t_L g1236 ( .A(n_544), .B(n_546), .Y(n_1236) );
INVx2_ASAP7_75t_SL g1272 ( .A(n_544), .Y(n_1272) );
INVx2_ASAP7_75t_SL g544 ( .A(n_545), .Y(n_544) );
INVxp67_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g882 ( .A(n_547), .B(n_883), .Y(n_882) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g552 ( .A(n_548), .Y(n_552) );
OR2x2_ASAP7_75t_L g560 ( .A(n_548), .B(n_561), .Y(n_560) );
INVx1_ASAP7_75t_L g710 ( .A(n_549), .Y(n_710) );
INVx1_ASAP7_75t_L g728 ( .A(n_549), .Y(n_728) );
INVxp67_ASAP7_75t_L g1026 ( .A(n_550), .Y(n_1026) );
INVx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g842 ( .A1(n_551), .A2(n_805), .B1(n_806), .B2(n_843), .Y(n_842) );
AOI22xp33_ASAP7_75t_L g1118 ( .A1(n_551), .A2(n_843), .B1(n_1095), .B2(n_1096), .Y(n_1118) );
INVx2_ASAP7_75t_L g1195 ( .A(n_551), .Y(n_1195) );
AOI22xp33_ASAP7_75t_L g1670 ( .A1(n_551), .A2(n_843), .B1(n_1663), .B2(n_1664), .Y(n_1670) );
AND2x4_ASAP7_75t_L g843 ( .A(n_552), .B(n_844), .Y(n_843) );
AND2x4_ASAP7_75t_L g1061 ( .A(n_552), .B(n_844), .Y(n_1061) );
NOR4xp25_ASAP7_75t_L g1261 ( .A(n_553), .B(n_1262), .C(n_1265), .D(n_1266), .Y(n_1261) );
INVx2_ASAP7_75t_SL g553 ( .A(n_554), .Y(n_553) );
AND5x1_ASAP7_75t_L g847 ( .A(n_554), .B(n_848), .C(n_888), .D(n_902), .E(n_905), .Y(n_847) );
NAND5xp2_ASAP7_75t_L g918 ( .A(n_554), .B(n_919), .C(n_923), .D(n_926), .E(n_927), .Y(n_918) );
NAND3xp33_ASAP7_75t_SL g1032 ( .A(n_554), .B(n_1033), .C(n_1037), .Y(n_1032) );
AND4x1_ASAP7_75t_L g1192 ( .A(n_554), .B(n_1193), .C(n_1196), .D(n_1204), .Y(n_1192) );
INVx3_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
NOR3xp33_ASAP7_75t_L g818 ( .A(n_555), .B(n_819), .C(n_835), .Y(n_818) );
NOR3xp33_ASAP7_75t_SL g979 ( .A(n_555), .B(n_980), .C(n_994), .Y(n_979) );
INVx3_ASAP7_75t_L g1086 ( .A(n_555), .Y(n_1086) );
HB1xp67_ASAP7_75t_L g1137 ( .A(n_555), .Y(n_1137) );
AOI221xp5_ASAP7_75t_L g1334 ( .A1(n_555), .A2(n_837), .B1(n_1035), .B2(n_1320), .C(n_1335), .Y(n_1334) );
BUFx2_ASAP7_75t_L g1078 ( .A(n_556), .Y(n_1078) );
AOI21xp33_ASAP7_75t_SL g557 ( .A1(n_558), .A2(n_567), .B(n_568), .Y(n_557) );
AOI21xp5_ASAP7_75t_L g838 ( .A1(n_558), .A2(n_839), .B(n_840), .Y(n_838) );
AOI221xp5_ASAP7_75t_L g1029 ( .A1(n_558), .A2(n_925), .B1(n_1030), .B2(n_1031), .C(n_1032), .Y(n_1029) );
NAND2xp5_ASAP7_75t_L g1119 ( .A(n_558), .B(n_1120), .Y(n_1119) );
AOI21xp5_ASAP7_75t_L g1138 ( .A1(n_558), .A2(n_1139), .B(n_1140), .Y(n_1138) );
AOI21xp33_ASAP7_75t_L g1169 ( .A1(n_558), .A2(n_1170), .B(n_1171), .Y(n_1169) );
NAND2xp33_ASAP7_75t_L g1228 ( .A(n_558), .B(n_1229), .Y(n_1228) );
AOI21xp33_ASAP7_75t_L g1297 ( .A1(n_558), .A2(n_1298), .B(n_1299), .Y(n_1297) );
AOI21xp5_ASAP7_75t_L g1641 ( .A1(n_558), .A2(n_1642), .B(n_1643), .Y(n_1641) );
INVx8_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
AND2x4_ASAP7_75t_L g559 ( .A(n_560), .B(n_562), .Y(n_559) );
INVx1_ASAP7_75t_L g886 ( .A(n_560), .Y(n_886) );
BUFx3_ASAP7_75t_L g754 ( .A(n_561), .Y(n_754) );
INVx1_ASAP7_75t_L g670 ( .A(n_563), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .Y(n_563) );
INVx1_ASAP7_75t_L g615 ( .A(n_564), .Y(n_615) );
AND2x2_ASAP7_75t_L g1058 ( .A(n_564), .B(n_861), .Y(n_1058) );
INVx3_ASAP7_75t_L g595 ( .A(n_565), .Y(n_595) );
AND2x2_ASAP7_75t_L g603 ( .A(n_565), .B(n_582), .Y(n_603) );
BUFx6f_ASAP7_75t_L g878 ( .A(n_565), .Y(n_878) );
INVx2_ASAP7_75t_L g954 ( .A(n_569), .Y(n_954) );
HB1xp67_ASAP7_75t_L g1300 ( .A(n_569), .Y(n_1300) );
AND2x4_ASAP7_75t_L g569 ( .A(n_570), .B(n_572), .Y(n_569) );
INVx2_ASAP7_75t_SL g785 ( .A(n_570), .Y(n_785) );
AND2x4_ASAP7_75t_L g841 ( .A(n_570), .B(n_572), .Y(n_841) );
INVx2_ASAP7_75t_L g887 ( .A(n_572), .Y(n_887) );
OR2x2_ASAP7_75t_L g573 ( .A(n_574), .B(n_575), .Y(n_573) );
INVx2_ASAP7_75t_L g716 ( .A(n_574), .Y(n_716) );
OR2x6_ASAP7_75t_L g908 ( .A(n_574), .B(n_575), .Y(n_908) );
OAI21xp5_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_607), .B(n_632), .Y(n_576) );
INVx2_ASAP7_75t_SL g578 ( .A(n_579), .Y(n_578) );
INVx3_ASAP7_75t_L g950 ( .A(n_579), .Y(n_950) );
AOI221xp5_ASAP7_75t_SL g1097 ( .A1(n_579), .A2(n_598), .B1(n_1088), .B2(n_1098), .C(n_1102), .Y(n_1097) );
AND2x4_ASAP7_75t_L g579 ( .A(n_580), .B(n_582), .Y(n_579) );
BUFx2_ASAP7_75t_L g1103 ( .A(n_580), .Y(n_1103) );
BUFx6f_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
BUFx3_ASAP7_75t_L g597 ( .A(n_581), .Y(n_597) );
INVx2_ASAP7_75t_L g676 ( .A(n_581), .Y(n_676) );
BUFx3_ASAP7_75t_L g803 ( .A(n_581), .Y(n_803) );
AND2x4_ASAP7_75t_L g606 ( .A(n_582), .B(n_590), .Y(n_606) );
AND2x2_ASAP7_75t_L g736 ( .A(n_582), .B(n_590), .Y(n_736) );
BUFx2_ASAP7_75t_L g865 ( .A(n_582), .Y(n_865) );
AND2x2_ASAP7_75t_L g1000 ( .A(n_582), .B(n_675), .Y(n_1000) );
AOI21xp5_ASAP7_75t_SL g583 ( .A1(n_584), .A2(n_593), .B(n_598), .Y(n_583) );
BUFx2_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
HB1xp67_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g1146 ( .A(n_588), .Y(n_1146) );
INVx2_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx2_ASAP7_75t_L g1107 ( .A(n_589), .Y(n_1107) );
INVx2_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g800 ( .A(n_590), .Y(n_800) );
BUFx6f_ASAP7_75t_L g1002 ( .A(n_590), .Y(n_1002) );
HB1xp67_ASAP7_75t_SL g591 ( .A(n_592), .Y(n_591) );
INVx2_ASAP7_75t_SL g594 ( .A(n_595), .Y(n_594) );
INVx2_ASAP7_75t_L g802 ( .A(n_595), .Y(n_802) );
INVx1_ASAP7_75t_L g870 ( .A(n_595), .Y(n_870) );
INVx2_ASAP7_75t_L g1183 ( .A(n_595), .Y(n_1183) );
INVx1_ASAP7_75t_L g1290 ( .A(n_595), .Y(n_1290) );
BUFx3_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx1_ASAP7_75t_SL g1292 ( .A(n_597), .Y(n_1292) );
AOI21xp5_ASAP7_75t_L g797 ( .A1(n_598), .A2(n_798), .B(n_801), .Y(n_797) );
INVx1_ASAP7_75t_L g940 ( .A(n_598), .Y(n_940) );
AOI221xp5_ASAP7_75t_L g999 ( .A1(n_598), .A2(n_978), .B1(n_1000), .B2(n_1001), .C(n_1004), .Y(n_999) );
AOI221xp5_ASAP7_75t_L g1052 ( .A1(n_598), .A2(n_1000), .B1(n_1030), .B2(n_1053), .C(n_1054), .Y(n_1052) );
AOI21xp5_ASAP7_75t_L g1143 ( .A1(n_598), .A2(n_1144), .B(n_1147), .Y(n_1143) );
AOI21xp5_ASAP7_75t_L g1177 ( .A1(n_598), .A2(n_1178), .B(n_1182), .Y(n_1177) );
AOI21xp5_ASAP7_75t_L g1239 ( .A1(n_598), .A2(n_1240), .B(n_1241), .Y(n_1239) );
AOI21xp5_ASAP7_75t_L g1287 ( .A1(n_598), .A2(n_1288), .B(n_1289), .Y(n_1287) );
AOI21xp5_ASAP7_75t_L g1659 ( .A1(n_598), .A2(n_1660), .B(n_1661), .Y(n_1659) );
AOI22xp33_ASAP7_75t_L g599 ( .A1(n_600), .A2(n_601), .B1(n_604), .B2(n_605), .Y(n_599) );
AOI22xp33_ASAP7_75t_L g1148 ( .A1(n_601), .A2(n_1149), .B1(n_1150), .B2(n_1151), .Y(n_1148) );
AOI22xp33_ASAP7_75t_L g1293 ( .A1(n_601), .A2(n_1294), .B1(n_1295), .B2(n_1296), .Y(n_1293) );
INVx2_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
AND2x4_ASAP7_75t_L g686 ( .A(n_603), .B(n_687), .Y(n_686) );
AOI22xp33_ASAP7_75t_L g804 ( .A1(n_603), .A2(n_606), .B1(n_805), .B2(n_806), .Y(n_804) );
BUFx6f_ASAP7_75t_L g949 ( .A(n_603), .Y(n_949) );
INVxp67_ASAP7_75t_SL g942 ( .A(n_605), .Y(n_942) );
AOI22xp33_ASAP7_75t_L g1174 ( .A1(n_605), .A2(n_949), .B1(n_1175), .B2(n_1176), .Y(n_1174) );
BUFx6f_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
AOI22xp5_ASAP7_75t_L g1007 ( .A1(n_606), .A2(n_949), .B1(n_1008), .B2(n_1009), .Y(n_1007) );
AOI22xp5_ASAP7_75t_L g1049 ( .A1(n_606), .A2(n_949), .B1(n_1050), .B2(n_1051), .Y(n_1049) );
AOI22xp33_ASAP7_75t_L g1094 ( .A1(n_606), .A2(n_949), .B1(n_1095), .B2(n_1096), .Y(n_1094) );
INVx1_ASAP7_75t_L g1152 ( .A(n_606), .Y(n_1152) );
AOI22xp33_ASAP7_75t_L g1243 ( .A1(n_606), .A2(n_949), .B1(n_1244), .B2(n_1245), .Y(n_1243) );
HB1xp67_ASAP7_75t_L g1296 ( .A(n_606), .Y(n_1296) );
AOI22xp33_ASAP7_75t_L g1662 ( .A1(n_606), .A2(n_949), .B1(n_1663), .B2(n_1664), .Y(n_1662) );
INVx2_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx2_ASAP7_75t_L g808 ( .A(n_609), .Y(n_808) );
INVx1_ASAP7_75t_L g932 ( .A(n_609), .Y(n_932) );
AOI22xp33_ASAP7_75t_L g1160 ( .A1(n_609), .A2(n_613), .B1(n_1126), .B2(n_1127), .Y(n_1160) );
INVx4_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx2_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
BUFx3_ASAP7_75t_L g852 ( .A(n_611), .Y(n_852) );
INVx2_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx2_ASAP7_75t_L g809 ( .A(n_613), .Y(n_809) );
NOR2x1_ASAP7_75t_L g613 ( .A(n_614), .B(n_615), .Y(n_613) );
INVx1_ASAP7_75t_L g854 ( .A(n_615), .Y(n_854) );
OAI221xp5_ASAP7_75t_L g616 ( .A1(n_617), .A2(n_620), .B1(n_621), .B2(n_623), .C(n_624), .Y(n_616) );
INVx2_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
BUFx6f_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx4_ASAP7_75t_L g856 ( .A(n_619), .Y(n_856) );
INVx3_ASAP7_75t_L g1318 ( .A(n_619), .Y(n_1318) );
INVx1_ASAP7_75t_L g642 ( .A(n_621), .Y(n_642) );
BUFx2_ASAP7_75t_L g1188 ( .A(n_621), .Y(n_1188) );
BUFx6f_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx2_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx2_ASAP7_75t_L g1099 ( .A(n_627), .Y(n_1099) );
INVx2_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
HB1xp67_ASAP7_75t_L g1157 ( .A(n_628), .Y(n_1157) );
INVx1_ASAP7_75t_L g1180 ( .A(n_628), .Y(n_1180) );
INVx2_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx2_ASAP7_75t_L g939 ( .A(n_629), .Y(n_939) );
INVx2_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g815 ( .A(n_631), .Y(n_815) );
INVx3_ASAP7_75t_L g876 ( .A(n_631), .Y(n_876) );
INVx2_ASAP7_75t_L g1022 ( .A(n_631), .Y(n_1022) );
AOI21xp5_ASAP7_75t_SL g1092 ( .A1(n_632), .A2(n_1093), .B(n_1117), .Y(n_1092) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
BUFx2_ASAP7_75t_SL g789 ( .A(n_635), .Y(n_789) );
INVxp67_ASAP7_75t_SL g635 ( .A(n_636), .Y(n_635) );
XNOR2x1_ASAP7_75t_L g636 ( .A(n_637), .B(n_738), .Y(n_636) );
XNOR2x1_ASAP7_75t_L g637 ( .A(n_638), .B(n_737), .Y(n_637) );
OR2x2_ASAP7_75t_L g638 ( .A(n_639), .B(n_688), .Y(n_638) );
NAND3xp33_ASAP7_75t_SL g639 ( .A(n_640), .B(n_667), .C(n_682), .Y(n_639) );
AOI211xp5_ASAP7_75t_SL g640 ( .A1(n_641), .A2(n_645), .B(n_652), .C(n_661), .Y(n_640) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
OAI221xp5_ASAP7_75t_L g933 ( .A1(n_644), .A2(n_934), .B1(n_935), .B2(n_937), .C(n_938), .Y(n_933) );
OAI221xp5_ASAP7_75t_L g943 ( .A1(n_644), .A2(n_663), .B1(n_944), .B2(n_945), .C(n_946), .Y(n_943) );
OAI221xp5_ASAP7_75t_SL g1284 ( .A1(n_644), .A2(n_1188), .B1(n_1273), .B2(n_1280), .C(n_1285), .Y(n_1284) );
INVx2_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVxp67_ASAP7_75t_SL g648 ( .A(n_649), .Y(n_648) );
INVx2_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx2_ASAP7_75t_L g1383 ( .A(n_651), .Y(n_1383) );
INVx1_ASAP7_75t_L g784 ( .A(n_653), .Y(n_784) );
INVx2_ASAP7_75t_SL g1386 ( .A(n_653), .Y(n_1386) );
NAND2x2_ASAP7_75t_L g653 ( .A(n_654), .B(n_656), .Y(n_653) );
INVx1_ASAP7_75t_L g660 ( .A(n_654), .Y(n_660) );
INVx2_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx2_ASAP7_75t_SL g656 ( .A(n_657), .Y(n_656) );
CKINVDCx5p33_ASAP7_75t_R g788 ( .A(n_659), .Y(n_788) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
AOI222xp33_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_671), .B1(n_672), .B2(n_677), .C1(n_678), .C2(n_681), .Y(n_667) );
AOI21xp33_ASAP7_75t_SL g786 ( .A1(n_668), .A2(n_787), .B(n_788), .Y(n_786) );
AOI222xp33_ASAP7_75t_L g1387 ( .A1(n_668), .A2(n_672), .B1(n_678), .B2(n_1388), .C1(n_1389), .C2(n_1390), .Y(n_1387) );
AND2x4_ASAP7_75t_L g668 ( .A(n_669), .B(n_670), .Y(n_668) );
AOI222xp33_ASAP7_75t_L g782 ( .A1(n_672), .A2(n_749), .B1(n_761), .B2(n_783), .C1(n_784), .C2(n_785), .Y(n_782) );
AND2x4_ASAP7_75t_L g672 ( .A(n_673), .B(n_675), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
OR2x2_ASAP7_75t_L g679 ( .A(n_674), .B(n_680), .Y(n_679) );
INVx3_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g1110 ( .A(n_676), .Y(n_1110) );
AOI211xp5_ASAP7_75t_L g713 ( .A1(n_677), .A2(n_714), .B(n_717), .C(n_725), .Y(n_713) );
AOI222xp33_ASAP7_75t_L g769 ( .A1(n_678), .A2(n_750), .B1(n_770), .B2(n_777), .C1(n_778), .C2(n_781), .Y(n_769) );
INVx2_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx2_ASAP7_75t_SL g813 ( .A(n_680), .Y(n_813) );
BUFx3_ASAP7_75t_L g1377 ( .A(n_680), .Y(n_1377) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_683), .B(n_684), .Y(n_682) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx3_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
HB1xp67_ASAP7_75t_L g740 ( .A(n_686), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g1391 ( .A(n_686), .B(n_1392), .Y(n_1391) );
AND2x4_ASAP7_75t_L g735 ( .A(n_687), .B(n_736), .Y(n_735) );
A2O1A1Ixp33_ASAP7_75t_L g688 ( .A1(n_689), .A2(n_713), .B(n_731), .C(n_733), .Y(n_688) );
AOI221xp5_ASAP7_75t_L g689 ( .A1(n_690), .A2(n_694), .B1(n_696), .B2(n_703), .C(n_707), .Y(n_689) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
OR2x6_ASAP7_75t_SL g726 ( .A(n_692), .B(n_727), .Y(n_726) );
INVx3_ASAP7_75t_L g883 ( .A(n_692), .Y(n_883) );
BUFx2_ASAP7_75t_L g1132 ( .A(n_692), .Y(n_1132) );
OAI221xp5_ASAP7_75t_L g1646 ( .A1(n_692), .A2(n_825), .B1(n_1647), .B2(n_1648), .C(n_1649), .Y(n_1646) );
INVx3_ASAP7_75t_L g759 ( .A(n_695), .Y(n_759) );
INVx2_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g969 ( .A(n_698), .Y(n_969) );
INVx1_ASAP7_75t_L g1203 ( .A(n_698), .Y(n_1203) );
INVx2_ASAP7_75t_L g1331 ( .A(n_698), .Y(n_1331) );
INVx2_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
OAI221xp5_ASAP7_75t_L g752 ( .A1(n_700), .A2(n_753), .B1(n_754), .B2(n_755), .C(n_756), .Y(n_752) );
INVx3_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx2_ASAP7_75t_SL g892 ( .A(n_701), .Y(n_892) );
INVx5_ASAP7_75t_L g898 ( .A(n_701), .Y(n_898) );
INVx2_ASAP7_75t_SL g1223 ( .A(n_701), .Y(n_1223) );
BUFx2_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g1404 ( .A(n_705), .Y(n_1404) );
BUFx2_ASAP7_75t_L g1084 ( .A(n_706), .Y(n_1084) );
INVx2_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
AOI22xp5_ASAP7_75t_L g760 ( .A1(n_709), .A2(n_712), .B1(n_741), .B2(n_761), .Y(n_760) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx2_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
AOI221xp5_ASAP7_75t_L g1394 ( .A1(n_716), .A2(n_1389), .B1(n_1395), .B2(n_1397), .C(n_1399), .Y(n_1394) );
INVx4_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
AOI22xp33_ASAP7_75t_L g748 ( .A1(n_719), .A2(n_721), .B1(n_749), .B2(n_750), .Y(n_748) );
INVx2_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
CKINVDCx5p33_ASAP7_75t_R g1401 ( .A(n_722), .Y(n_1401) );
OR2x6_ASAP7_75t_L g722 ( .A(n_723), .B(n_724), .Y(n_722) );
INVx2_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
HB1xp67_ASAP7_75t_L g1398 ( .A(n_728), .Y(n_1398) );
INVx3_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
HB1xp67_ASAP7_75t_L g879 ( .A(n_731), .Y(n_879) );
INVx1_ASAP7_75t_L g1162 ( .A(n_731), .Y(n_1162) );
BUFx2_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
BUFx2_ASAP7_75t_L g817 ( .A(n_732), .Y(n_817) );
AOI21x1_ASAP7_75t_L g1308 ( .A1(n_732), .A2(n_1309), .B(n_1324), .Y(n_1308) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_734), .B(n_735), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_735), .B(n_744), .Y(n_743) );
INVx2_ASAP7_75t_L g1338 ( .A(n_735), .Y(n_1338) );
NAND2xp33_ASAP7_75t_SL g1413 ( .A(n_735), .B(n_1414), .Y(n_1413) );
AOI211x1_ASAP7_75t_L g739 ( .A1(n_740), .A2(n_741), .B(n_742), .C(n_768), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_743), .B(n_745), .Y(n_742) );
NAND3xp33_ASAP7_75t_L g751 ( .A(n_752), .B(n_760), .C(n_762), .Y(n_751) );
OAI221xp5_ASAP7_75t_L g897 ( .A1(n_754), .A2(n_874), .B1(n_898), .B2(n_899), .C(n_900), .Y(n_897) );
INVx3_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
OAI211xp5_ASAP7_75t_L g762 ( .A1(n_763), .A2(n_764), .B(n_766), .C(n_767), .Y(n_762) );
INVx3_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
INVx2_ASAP7_75t_L g962 ( .A(n_765), .Y(n_962) );
NAND3xp33_ASAP7_75t_L g768 ( .A(n_769), .B(n_782), .C(n_786), .Y(n_768) );
INVx1_ASAP7_75t_L g1252 ( .A(n_772), .Y(n_1252) );
INVx1_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
OA22x2_ASAP7_75t_L g791 ( .A1(n_792), .A2(n_845), .B1(n_846), .B2(n_909), .Y(n_791) );
INVx1_ASAP7_75t_L g909 ( .A(n_792), .Y(n_909) );
INVx1_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
AND4x1_ASAP7_75t_L g794 ( .A(n_795), .B(n_818), .C(n_838), .D(n_842), .Y(n_794) );
OAI21xp5_ASAP7_75t_L g795 ( .A1(n_796), .A2(n_807), .B(n_817), .Y(n_795) );
INVx2_ASAP7_75t_SL g799 ( .A(n_800), .Y(n_799) );
BUFx2_ASAP7_75t_L g1185 ( .A(n_809), .Y(n_1185) );
OAI211xp5_ASAP7_75t_L g810 ( .A1(n_811), .A2(n_812), .B(n_814), .C(n_816), .Y(n_810) );
OAI221xp5_ASAP7_75t_L g831 ( .A1(n_811), .A2(n_822), .B1(n_832), .B2(n_833), .C(n_834), .Y(n_831) );
OAI211xp5_ASAP7_75t_L g873 ( .A1(n_812), .A2(n_874), .B(n_875), .C(n_877), .Y(n_873) );
INVx5_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
OAI22xp5_ASAP7_75t_SL g819 ( .A1(n_820), .A2(n_821), .B1(n_829), .B2(n_831), .Y(n_819) );
OAI221xp5_ASAP7_75t_L g821 ( .A1(n_822), .A2(n_823), .B1(n_824), .B2(n_825), .C(n_828), .Y(n_821) );
INVx3_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
BUFx2_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
CKINVDCx5p33_ASAP7_75t_R g829 ( .A(n_830), .Y(n_829) );
INVx2_ASAP7_75t_L g896 ( .A(n_830), .Y(n_896) );
INVx2_ASAP7_75t_L g1650 ( .A(n_830), .Y(n_1650) );
OAI221xp5_ASAP7_75t_L g1651 ( .A1(n_832), .A2(n_1652), .B1(n_1653), .B2(n_1654), .C(n_1655), .Y(n_1651) );
INVx1_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
AOI22xp5_ASAP7_75t_L g1033 ( .A1(n_837), .A2(n_1034), .B1(n_1035), .B2(n_1036), .Y(n_1033) );
INVx1_ASAP7_75t_SL g977 ( .A(n_841), .Y(n_977) );
NAND2xp5_ASAP7_75t_L g927 ( .A(n_843), .B(n_928), .Y(n_927) );
AOI22xp5_ASAP7_75t_L g1025 ( .A1(n_843), .A2(n_1008), .B1(n_1009), .B2(n_1026), .Y(n_1025) );
INVx2_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
AOI21xp5_ASAP7_75t_L g848 ( .A1(n_849), .A2(n_879), .B(n_880), .Y(n_848) );
NAND4xp25_ASAP7_75t_L g849 ( .A(n_850), .B(n_853), .C(n_867), .D(n_873), .Y(n_849) );
NAND2xp5_ASAP7_75t_L g850 ( .A(n_851), .B(n_852), .Y(n_850) );
AOI222xp33_ASAP7_75t_L g1055 ( .A1(n_852), .A2(n_1034), .B1(n_1036), .B2(n_1056), .C1(n_1057), .C2(n_1058), .Y(n_1055) );
INVx1_ASAP7_75t_L g1115 ( .A(n_852), .Y(n_1115) );
AOI22xp5_ASAP7_75t_L g853 ( .A1(n_854), .A2(n_855), .B1(n_865), .B2(n_866), .Y(n_853) );
AOI22xp5_ASAP7_75t_L g1316 ( .A1(n_854), .A2(n_865), .B1(n_1317), .B2(n_1322), .Y(n_1316) );
OAI22xp5_ASAP7_75t_L g1366 ( .A1(n_857), .A2(n_1367), .B1(n_1368), .B2(n_1371), .Y(n_1366) );
INVx2_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
INVx2_ASAP7_75t_L g1249 ( .A(n_858), .Y(n_1249) );
INVx1_ASAP7_75t_L g1667 ( .A(n_858), .Y(n_1667) );
AOI22xp33_ASAP7_75t_L g859 ( .A1(n_860), .A2(n_861), .B1(n_862), .B2(n_863), .Y(n_859) );
AOI22xp5_ASAP7_75t_L g1319 ( .A1(n_861), .A2(n_863), .B1(n_1320), .B2(n_1321), .Y(n_1319) );
AOI22xp5_ASAP7_75t_L g884 ( .A1(n_862), .A2(n_885), .B1(n_886), .B2(n_887), .Y(n_884) );
INVx1_ASAP7_75t_L g863 ( .A(n_864), .Y(n_863) );
INVx3_ASAP7_75t_L g1006 ( .A(n_878), .Y(n_1006) );
BUFx6f_ASAP7_75t_L g1242 ( .A(n_878), .Y(n_1242) );
NAND2x1_ASAP7_75t_L g1337 ( .A(n_881), .B(n_1338), .Y(n_1337) );
INVx2_ASAP7_75t_SL g881 ( .A(n_882), .Y(n_881) );
AOI22xp33_ASAP7_75t_L g1060 ( .A1(n_882), .A2(n_1050), .B1(n_1051), .B2(n_1061), .Y(n_1060) );
INVx2_ASAP7_75t_L g990 ( .A(n_883), .Y(n_990) );
INVx2_ASAP7_75t_L g1406 ( .A(n_883), .Y(n_1406) );
AOI222xp33_ASAP7_75t_L g1340 ( .A1(n_886), .A2(n_887), .B1(n_1061), .B2(n_1321), .C1(n_1341), .C2(n_1342), .Y(n_1340) );
OAI22xp5_ASAP7_75t_SL g889 ( .A1(n_890), .A2(n_891), .B1(n_896), .B2(n_897), .Y(n_889) );
OAI211xp5_ASAP7_75t_L g982 ( .A1(n_892), .A2(n_983), .B(n_984), .C(n_986), .Y(n_982) );
OAI22xp5_ASAP7_75t_L g980 ( .A1(n_896), .A2(n_981), .B1(n_982), .B2(n_989), .Y(n_980) );
BUFx3_ASAP7_75t_L g964 ( .A(n_898), .Y(n_964) );
INVx8_ASAP7_75t_L g1134 ( .A(n_898), .Y(n_1134) );
NAND2xp5_ASAP7_75t_L g902 ( .A(n_903), .B(n_904), .Y(n_902) );
NAND2xp5_ASAP7_75t_L g905 ( .A(n_906), .B(n_907), .Y(n_905) );
NAND2xp5_ASAP7_75t_L g1217 ( .A(n_907), .B(n_1218), .Y(n_1217) );
INVx5_ASAP7_75t_L g907 ( .A(n_908), .Y(n_907) );
INVx3_ASAP7_75t_L g925 ( .A(n_908), .Y(n_925) );
OAI22xp5_ASAP7_75t_L g911 ( .A1(n_912), .A2(n_1302), .B1(n_1350), .B2(n_1351), .Y(n_911) );
INVx1_ASAP7_75t_L g1350 ( .A(n_912), .Y(n_1350) );
XOR2x2_ASAP7_75t_L g912 ( .A(n_913), .B(n_1164), .Y(n_912) );
XOR2xp5_ASAP7_75t_L g913 ( .A(n_914), .B(n_1063), .Y(n_913) );
AOI22xp5_ASAP7_75t_L g914 ( .A1(n_915), .A2(n_916), .B1(n_971), .B2(n_1062), .Y(n_914) );
INVx2_ASAP7_75t_L g915 ( .A(n_916), .Y(n_915) );
XNOR2x1_ASAP7_75t_L g916 ( .A(n_917), .B(n_970), .Y(n_916) );
NOR2x1_ASAP7_75t_L g917 ( .A(n_918), .B(n_929), .Y(n_917) );
NAND2xp5_ASAP7_75t_L g923 ( .A(n_924), .B(n_925), .Y(n_923) );
AOI22xp5_ASAP7_75t_L g975 ( .A1(n_925), .A2(n_976), .B1(n_977), .B2(n_978), .Y(n_975) );
NAND2xp5_ASAP7_75t_L g1087 ( .A(n_925), .B(n_1088), .Y(n_1087) );
NAND2xp5_ASAP7_75t_L g929 ( .A(n_930), .B(n_953), .Y(n_929) );
OAI31xp33_ASAP7_75t_L g930 ( .A1(n_931), .A2(n_941), .A3(n_947), .B(n_951), .Y(n_930) );
HB1xp67_ASAP7_75t_L g935 ( .A(n_936), .Y(n_935) );
OAI22xp5_ASAP7_75t_L g1362 ( .A1(n_936), .A2(n_1363), .B1(n_1364), .B2(n_1365), .Y(n_1362) );
OAI22xp5_ASAP7_75t_L g1379 ( .A1(n_936), .A2(n_1380), .B1(n_1381), .B2(n_1382), .Y(n_1379) );
OAI221xp5_ASAP7_75t_L g963 ( .A1(n_937), .A2(n_964), .B1(n_965), .B2(n_966), .C(n_967), .Y(n_963) );
INVx1_ASAP7_75t_L g948 ( .A(n_949), .Y(n_948) );
OAI21xp5_ASAP7_75t_L g1172 ( .A1(n_951), .A2(n_1173), .B(n_1184), .Y(n_1172) );
INVx1_ASAP7_75t_L g951 ( .A(n_952), .Y(n_951) );
BUFx2_ASAP7_75t_L g1024 ( .A(n_952), .Y(n_1024) );
AOI21xp5_ASAP7_75t_SL g953 ( .A1(n_954), .A2(n_955), .B(n_956), .Y(n_953) );
AOI21xp5_ASAP7_75t_L g1233 ( .A1(n_954), .A2(n_1234), .B(n_1235), .Y(n_1233) );
OAI22xp33_ASAP7_75t_L g1279 ( .A1(n_962), .A2(n_1271), .B1(n_1280), .B2(n_1281), .Y(n_1279) );
OAI22xp5_ASAP7_75t_L g1270 ( .A1(n_964), .A2(n_1271), .B1(n_1273), .B2(n_1274), .Y(n_1270) );
OAI221xp5_ASAP7_75t_L g989 ( .A1(n_966), .A2(n_990), .B1(n_991), .B2(n_992), .C(n_993), .Y(n_989) );
INVx1_ASAP7_75t_L g1062 ( .A(n_971), .Y(n_1062) );
XNOR2x1_ASAP7_75t_L g971 ( .A(n_972), .B(n_1027), .Y(n_971) );
NAND4xp75_ASAP7_75t_L g973 ( .A(n_974), .B(n_979), .C(n_997), .D(n_1025), .Y(n_973) );
INVx2_ASAP7_75t_L g987 ( .A(n_988), .Y(n_987) );
INVx1_ASAP7_75t_L g995 ( .A(n_996), .Y(n_995) );
OAI21xp5_ASAP7_75t_L g997 ( .A1(n_998), .A2(n_1010), .B(n_1023), .Y(n_997) );
NAND2xp5_ASAP7_75t_L g998 ( .A(n_999), .B(n_1007), .Y(n_998) );
INVx2_ASAP7_75t_L g1310 ( .A(n_1000), .Y(n_1310) );
INVx1_ASAP7_75t_L g1005 ( .A(n_1006), .Y(n_1005) );
INVx2_ASAP7_75t_SL g1109 ( .A(n_1006), .Y(n_1109) );
OAI221xp5_ASAP7_75t_L g1011 ( .A1(n_1012), .A2(n_1013), .B1(n_1014), .B2(n_1016), .C(n_1017), .Y(n_1011) );
BUFx3_ASAP7_75t_L g1014 ( .A(n_1015), .Y(n_1014) );
INVx2_ASAP7_75t_L g1018 ( .A(n_1019), .Y(n_1018) );
INVx1_ASAP7_75t_L g1019 ( .A(n_1020), .Y(n_1019) );
INVx1_ASAP7_75t_L g1020 ( .A(n_1021), .Y(n_1020) );
BUFx2_ASAP7_75t_L g1101 ( .A(n_1021), .Y(n_1101) );
INVx1_ASAP7_75t_L g1023 ( .A(n_1024), .Y(n_1023) );
INVx2_ASAP7_75t_L g1047 ( .A(n_1024), .Y(n_1047) );
AND2x2_ASAP7_75t_L g1028 ( .A(n_1029), .B(n_1046), .Y(n_1028) );
AOI22xp5_ASAP7_75t_L g1037 ( .A1(n_1038), .A2(n_1041), .B1(n_1043), .B2(n_1045), .Y(n_1037) );
INVx1_ASAP7_75t_L g1082 ( .A(n_1039), .Y(n_1082) );
AOI21xp5_ASAP7_75t_L g1046 ( .A1(n_1047), .A2(n_1048), .B(n_1059), .Y(n_1046) );
OAI21xp5_ASAP7_75t_L g1237 ( .A1(n_1047), .A2(n_1238), .B(n_1246), .Y(n_1237) );
A2O1A1Ixp33_ASAP7_75t_L g1393 ( .A1(n_1047), .A2(n_1394), .B(n_1400), .C(n_1413), .Y(n_1393) );
OAI21xp5_ASAP7_75t_L g1657 ( .A1(n_1047), .A2(n_1658), .B(n_1665), .Y(n_1657) );
NAND3xp33_ASAP7_75t_L g1048 ( .A(n_1049), .B(n_1052), .C(n_1055), .Y(n_1048) );
INVx1_ASAP7_75t_L g1116 ( .A(n_1058), .Y(n_1116) );
OAI22x1_ASAP7_75t_L g1063 ( .A1(n_1064), .A2(n_1065), .B1(n_1121), .B2(n_1163), .Y(n_1063) );
INVx2_ASAP7_75t_L g1064 ( .A(n_1065), .Y(n_1064) );
XNOR2x1_ASAP7_75t_L g1065 ( .A(n_1066), .B(n_1067), .Y(n_1065) );
AND3x2_ASAP7_75t_L g1067 ( .A(n_1068), .B(n_1092), .C(n_1119), .Y(n_1067) );
NOR2xp33_ASAP7_75t_SL g1068 ( .A(n_1069), .B(n_1085), .Y(n_1068) );
OAI21xp5_ASAP7_75t_SL g1069 ( .A1(n_1070), .A2(n_1073), .B(n_1079), .Y(n_1069) );
NAND2xp5_ASAP7_75t_L g1073 ( .A(n_1074), .B(n_1075), .Y(n_1073) );
INVx2_ASAP7_75t_L g1076 ( .A(n_1077), .Y(n_1076) );
INVx1_ASAP7_75t_L g1081 ( .A(n_1082), .Y(n_1081) );
NAND3xp33_ASAP7_75t_L g1085 ( .A(n_1086), .B(n_1087), .C(n_1089), .Y(n_1085) );
NAND4xp25_ASAP7_75t_SL g1213 ( .A(n_1086), .B(n_1214), .C(n_1217), .D(n_1219), .Y(n_1213) );
NAND3xp33_ASAP7_75t_L g1093 ( .A(n_1094), .B(n_1097), .C(n_1104), .Y(n_1093) );
INVx2_ASAP7_75t_L g1100 ( .A(n_1101), .Y(n_1100) );
AOI31xp33_ASAP7_75t_L g1104 ( .A1(n_1105), .A2(n_1108), .A3(n_1111), .B(n_1114), .Y(n_1104) );
BUFx2_ASAP7_75t_L g1106 ( .A(n_1107), .Y(n_1106) );
INVx1_ASAP7_75t_L g1112 ( .A(n_1113), .Y(n_1112) );
INVx1_ASAP7_75t_L g1191 ( .A(n_1113), .Y(n_1191) );
INVx1_ASAP7_75t_L g1163 ( .A(n_1121), .Y(n_1163) );
NAND3xp33_ASAP7_75t_L g1122 ( .A(n_1123), .B(n_1138), .C(n_1141), .Y(n_1122) );
NOR3xp33_ASAP7_75t_L g1123 ( .A(n_1124), .B(n_1136), .C(n_1137), .Y(n_1123) );
NAND2xp5_ASAP7_75t_L g1124 ( .A(n_1125), .B(n_1128), .Y(n_1124) );
INVx2_ASAP7_75t_L g1131 ( .A(n_1132), .Y(n_1131) );
NOR3xp33_ASAP7_75t_L g1644 ( .A(n_1137), .B(n_1645), .C(n_1656), .Y(n_1644) );
OAI21xp5_ASAP7_75t_L g1141 ( .A1(n_1142), .A2(n_1153), .B(n_1161), .Y(n_1141) );
INVx1_ASAP7_75t_L g1145 ( .A(n_1146), .Y(n_1145) );
INVx1_ASAP7_75t_L g1151 ( .A(n_1152), .Y(n_1151) );
NAND2xp5_ASAP7_75t_L g1155 ( .A(n_1156), .B(n_1158), .Y(n_1155) );
INVx1_ASAP7_75t_L g1380 ( .A(n_1159), .Y(n_1380) );
OAI21xp5_ASAP7_75t_L g1282 ( .A1(n_1161), .A2(n_1283), .B(n_1286), .Y(n_1282) );
INVx2_ASAP7_75t_L g1161 ( .A(n_1162), .Y(n_1161) );
XNOR2x1_ASAP7_75t_L g1164 ( .A(n_1165), .B(n_1258), .Y(n_1164) );
OAI22x1_ASAP7_75t_L g1165 ( .A1(n_1166), .A2(n_1208), .B1(n_1209), .B2(n_1257), .Y(n_1165) );
INVx2_ASAP7_75t_L g1257 ( .A(n_1166), .Y(n_1257) );
AO21x2_ASAP7_75t_L g1166 ( .A1(n_1167), .A2(n_1168), .B(n_1207), .Y(n_1166) );
NAND3xp33_ASAP7_75t_SL g1168 ( .A(n_1169), .B(n_1172), .C(n_1192), .Y(n_1168) );
INVx1_ASAP7_75t_L g1179 ( .A(n_1180), .Y(n_1179) );
INVx1_ASAP7_75t_L g1193 ( .A(n_1194), .Y(n_1193) );
INVx2_ASAP7_75t_L g1208 ( .A(n_1209), .Y(n_1208) );
NAND2x1p5_ASAP7_75t_L g1209 ( .A(n_1210), .B(n_1230), .Y(n_1209) );
NAND2xp5_ASAP7_75t_L g1211 ( .A(n_1212), .B(n_1228), .Y(n_1211) );
INVxp67_ASAP7_75t_L g1212 ( .A(n_1213), .Y(n_1212) );
NOR2xp33_ASAP7_75t_SL g1254 ( .A(n_1213), .B(n_1255), .Y(n_1254) );
INVx2_ASAP7_75t_L g1222 ( .A(n_1223), .Y(n_1222) );
NAND2xp5_ASAP7_75t_L g1255 ( .A(n_1228), .B(n_1256), .Y(n_1255) );
INVx1_ASAP7_75t_L g1231 ( .A(n_1232), .Y(n_1231) );
NAND2xp5_ASAP7_75t_L g1232 ( .A(n_1233), .B(n_1237), .Y(n_1232) );
OAI211xp5_ASAP7_75t_L g1247 ( .A1(n_1248), .A2(n_1249), .B(n_1250), .C(n_1253), .Y(n_1247) );
INVx1_ASAP7_75t_L g1251 ( .A(n_1252), .Y(n_1251) );
INVx1_ASAP7_75t_L g1259 ( .A(n_1260), .Y(n_1259) );
AND3x2_ASAP7_75t_L g1260 ( .A(n_1261), .B(n_1282), .C(n_1297), .Y(n_1260) );
INVx1_ASAP7_75t_L g1263 ( .A(n_1264), .Y(n_1263) );
INVx1_ASAP7_75t_L g1271 ( .A(n_1272), .Y(n_1271) );
INVx1_ASAP7_75t_SL g1291 ( .A(n_1292), .Y(n_1291) );
CKINVDCx14_ASAP7_75t_R g1351 ( .A(n_1302), .Y(n_1351) );
CKINVDCx6p67_ASAP7_75t_R g1302 ( .A(n_1303), .Y(n_1302) );
HB1xp67_ASAP7_75t_L g1303 ( .A(n_1304), .Y(n_1303) );
HB1xp67_ASAP7_75t_L g1304 ( .A(n_1305), .Y(n_1304) );
INVx1_ASAP7_75t_L g1305 ( .A(n_1306), .Y(n_1305) );
NAND3xp33_ASAP7_75t_L g1306 ( .A(n_1307), .B(n_1343), .C(n_1347), .Y(n_1306) );
INVx1_ASAP7_75t_L g1344 ( .A(n_1308), .Y(n_1344) );
AOI22xp5_ASAP7_75t_L g1311 ( .A1(n_1312), .A2(n_1313), .B1(n_1314), .B2(n_1315), .Y(n_1311) );
INVx1_ASAP7_75t_L g1345 ( .A(n_1325), .Y(n_1345) );
AND2x2_ASAP7_75t_L g1325 ( .A(n_1326), .B(n_1334), .Y(n_1325) );
INVx1_ASAP7_75t_L g1332 ( .A(n_1333), .Y(n_1332) );
INVx1_ASAP7_75t_L g1349 ( .A(n_1336), .Y(n_1349) );
NAND2xp5_ASAP7_75t_L g1336 ( .A(n_1337), .B(n_1339), .Y(n_1336) );
INVx1_ASAP7_75t_L g1348 ( .A(n_1340), .Y(n_1348) );
OAI21xp5_ASAP7_75t_L g1343 ( .A1(n_1344), .A2(n_1345), .B(n_1346), .Y(n_1343) );
OAI21xp33_ASAP7_75t_L g1347 ( .A1(n_1346), .A2(n_1348), .B(n_1349), .Y(n_1347) );
NAND2xp5_ASAP7_75t_SL g1677 ( .A(n_1353), .B(n_1678), .Y(n_1677) );
AOI221xp5_ASAP7_75t_L g1353 ( .A1(n_1354), .A2(n_1415), .B1(n_1423), .B2(n_1631), .C(n_1633), .Y(n_1353) );
INVx1_ASAP7_75t_L g1354 ( .A(n_1355), .Y(n_1354) );
INVx1_ASAP7_75t_L g1355 ( .A(n_1356), .Y(n_1355) );
XNOR2x1_ASAP7_75t_L g1356 ( .A(n_1357), .B(n_1358), .Y(n_1356) );
NOR2x1_ASAP7_75t_L g1358 ( .A(n_1359), .B(n_1393), .Y(n_1358) );
NAND3xp33_ASAP7_75t_L g1359 ( .A(n_1360), .B(n_1387), .C(n_1391), .Y(n_1359) );
NOR2xp33_ASAP7_75t_L g1360 ( .A(n_1361), .B(n_1384), .Y(n_1360) );
INVx4_ASAP7_75t_L g1368 ( .A(n_1369), .Y(n_1368) );
INVx4_ASAP7_75t_L g1369 ( .A(n_1370), .Y(n_1369) );
OAI22xp5_ASAP7_75t_L g1372 ( .A1(n_1373), .A2(n_1376), .B1(n_1377), .B2(n_1378), .Y(n_1372) );
INVx4_ASAP7_75t_L g1373 ( .A(n_1374), .Y(n_1373) );
BUFx2_ASAP7_75t_L g1374 ( .A(n_1375), .Y(n_1374) );
INVx2_ASAP7_75t_L g1385 ( .A(n_1386), .Y(n_1385) );
BUFx2_ASAP7_75t_L g1397 ( .A(n_1398), .Y(n_1397) );
NOR3xp33_ASAP7_75t_L g1400 ( .A(n_1401), .B(n_1402), .C(n_1408), .Y(n_1400) );
INVx1_ASAP7_75t_L g1403 ( .A(n_1404), .Y(n_1403) );
OR2x2_ASAP7_75t_L g1681 ( .A(n_1417), .B(n_1682), .Y(n_1681) );
INVx1_ASAP7_75t_L g1417 ( .A(n_1418), .Y(n_1417) );
NOR2xp33_ASAP7_75t_L g1418 ( .A(n_1419), .B(n_1421), .Y(n_1418) );
NOR2xp33_ASAP7_75t_L g1636 ( .A(n_1419), .B(n_1422), .Y(n_1636) );
INVx1_ASAP7_75t_L g1674 ( .A(n_1419), .Y(n_1674) );
HB1xp67_ASAP7_75t_L g1419 ( .A(n_1420), .Y(n_1419) );
INVx1_ASAP7_75t_L g1421 ( .A(n_1422), .Y(n_1421) );
NOR2xp33_ASAP7_75t_L g1676 ( .A(n_1422), .B(n_1674), .Y(n_1676) );
INVx1_ASAP7_75t_L g1423 ( .A(n_1424), .Y(n_1423) );
AOI211xp5_ASAP7_75t_L g1424 ( .A1(n_1425), .A2(n_1545), .B(n_1591), .C(n_1615), .Y(n_1424) );
OAI211xp5_ASAP7_75t_L g1425 ( .A1(n_1426), .A2(n_1442), .B(n_1487), .C(n_1533), .Y(n_1425) );
NAND2xp5_ASAP7_75t_L g1565 ( .A(n_1426), .B(n_1566), .Y(n_1565) );
OAI211xp5_ASAP7_75t_L g1615 ( .A1(n_1426), .A2(n_1616), .B(n_1618), .C(n_1624), .Y(n_1615) );
INVx2_ASAP7_75t_L g1426 ( .A(n_1427), .Y(n_1426) );
OAI221xp5_ASAP7_75t_L g1517 ( .A1(n_1427), .A2(n_1518), .B1(n_1524), .B2(n_1527), .C(n_1529), .Y(n_1517) );
OAI32xp33_ASAP7_75t_L g1583 ( .A1(n_1427), .A2(n_1488), .A3(n_1505), .B1(n_1540), .B2(n_1584), .Y(n_1583) );
OAI221xp5_ASAP7_75t_L g1591 ( .A1(n_1427), .A2(n_1516), .B1(n_1592), .B2(n_1599), .C(n_1601), .Y(n_1591) );
INVx3_ASAP7_75t_L g1427 ( .A(n_1428), .Y(n_1427) );
INVx3_ASAP7_75t_L g1511 ( .A(n_1428), .Y(n_1511) );
AND2x2_ASAP7_75t_L g1514 ( .A(n_1428), .B(n_1515), .Y(n_1514) );
AND2x2_ASAP7_75t_L g1528 ( .A(n_1428), .B(n_1461), .Y(n_1528) );
OR2x2_ASAP7_75t_L g1550 ( .A(n_1428), .B(n_1483), .Y(n_1550) );
AND2x2_ASAP7_75t_L g1595 ( .A(n_1428), .B(n_1474), .Y(n_1595) );
AND2x2_ASAP7_75t_L g1607 ( .A(n_1428), .B(n_1499), .Y(n_1607) );
NAND2xp5_ASAP7_75t_L g1614 ( .A(n_1428), .B(n_1483), .Y(n_1614) );
NOR2xp33_ASAP7_75t_L g1619 ( .A(n_1428), .B(n_1620), .Y(n_1619) );
AND2x4_ASAP7_75t_SL g1428 ( .A(n_1429), .B(n_1436), .Y(n_1428) );
INVx2_ASAP7_75t_L g1632 ( .A(n_1430), .Y(n_1632) );
AND2x6_ASAP7_75t_L g1430 ( .A(n_1431), .B(n_1432), .Y(n_1430) );
AND2x2_ASAP7_75t_L g1434 ( .A(n_1431), .B(n_1435), .Y(n_1434) );
AND2x4_ASAP7_75t_L g1437 ( .A(n_1431), .B(n_1438), .Y(n_1437) );
AND2x6_ASAP7_75t_L g1440 ( .A(n_1431), .B(n_1441), .Y(n_1440) );
AND2x2_ASAP7_75t_L g1449 ( .A(n_1431), .B(n_1435), .Y(n_1449) );
AND2x2_ASAP7_75t_L g1452 ( .A(n_1431), .B(n_1435), .Y(n_1452) );
HB1xp67_ASAP7_75t_L g1673 ( .A(n_1432), .Y(n_1673) );
AND2x2_ASAP7_75t_L g1438 ( .A(n_1433), .B(n_1439), .Y(n_1438) );
AOI221xp5_ASAP7_75t_L g1442 ( .A1(n_1443), .A2(n_1454), .B1(n_1465), .B2(n_1482), .C(n_1484), .Y(n_1442) );
A2O1A1Ixp33_ASAP7_75t_SL g1512 ( .A1(n_1443), .A2(n_1493), .B(n_1513), .C(n_1514), .Y(n_1512) );
INVx1_ASAP7_75t_L g1543 ( .A(n_1443), .Y(n_1543) );
AND2x2_ASAP7_75t_L g1443 ( .A(n_1444), .B(n_1450), .Y(n_1443) );
INVx1_ASAP7_75t_L g1444 ( .A(n_1445), .Y(n_1444) );
OR2x2_ASAP7_75t_L g1505 ( .A(n_1445), .B(n_1450), .Y(n_1505) );
INVx1_ASAP7_75t_L g1445 ( .A(n_1446), .Y(n_1445) );
OR2x2_ASAP7_75t_L g1469 ( .A(n_1446), .B(n_1470), .Y(n_1469) );
AND2x2_ASAP7_75t_L g1485 ( .A(n_1446), .B(n_1470), .Y(n_1485) );
AND2x2_ASAP7_75t_L g1496 ( .A(n_1446), .B(n_1471), .Y(n_1496) );
INVx1_ASAP7_75t_L g1508 ( .A(n_1446), .Y(n_1508) );
NOR2xp33_ASAP7_75t_L g1520 ( .A(n_1446), .B(n_1450), .Y(n_1520) );
NAND2xp5_ASAP7_75t_L g1446 ( .A(n_1447), .B(n_1448), .Y(n_1446) );
NOR2xp33_ASAP7_75t_L g1467 ( .A(n_1450), .B(n_1457), .Y(n_1467) );
CKINVDCx5p33_ASAP7_75t_R g1481 ( .A(n_1450), .Y(n_1481) );
AND2x2_ASAP7_75t_L g1486 ( .A(n_1450), .B(n_1457), .Y(n_1486) );
NAND2xp5_ASAP7_75t_L g1523 ( .A(n_1450), .B(n_1480), .Y(n_1523) );
AND2x2_ASAP7_75t_L g1564 ( .A(n_1450), .B(n_1496), .Y(n_1564) );
AND2x2_ASAP7_75t_L g1577 ( .A(n_1450), .B(n_1508), .Y(n_1577) );
NAND2xp5_ASAP7_75t_L g1597 ( .A(n_1450), .B(n_1598), .Y(n_1597) );
AND2x2_ASAP7_75t_L g1450 ( .A(n_1451), .B(n_1453), .Y(n_1450) );
AND2x2_ASAP7_75t_L g1526 ( .A(n_1451), .B(n_1453), .Y(n_1526) );
AND2x2_ASAP7_75t_L g1454 ( .A(n_1455), .B(n_1460), .Y(n_1454) );
AND2x2_ASAP7_75t_L g1513 ( .A(n_1455), .B(n_1507), .Y(n_1513) );
AND2x2_ASAP7_75t_L g1519 ( .A(n_1455), .B(n_1520), .Y(n_1519) );
OR2x2_ASAP7_75t_L g1560 ( .A(n_1455), .B(n_1523), .Y(n_1560) );
AND2x2_ASAP7_75t_L g1590 ( .A(n_1455), .B(n_1499), .Y(n_1590) );
AND2x2_ASAP7_75t_L g1625 ( .A(n_1455), .B(n_1488), .Y(n_1625) );
INVx1_ASAP7_75t_L g1455 ( .A(n_1456), .Y(n_1455) );
NAND2xp5_ASAP7_75t_L g1478 ( .A(n_1456), .B(n_1479), .Y(n_1478) );
AND2x2_ASAP7_75t_L g1534 ( .A(n_1456), .B(n_1485), .Y(n_1534) );
NOR2xp33_ASAP7_75t_L g1538 ( .A(n_1456), .B(n_1505), .Y(n_1538) );
NAND2xp5_ASAP7_75t_L g1544 ( .A(n_1456), .B(n_1488), .Y(n_1544) );
AND2x2_ASAP7_75t_L g1551 ( .A(n_1456), .B(n_1552), .Y(n_1551) );
NAND2xp5_ASAP7_75t_L g1555 ( .A(n_1456), .B(n_1495), .Y(n_1555) );
NAND2xp5_ASAP7_75t_L g1563 ( .A(n_1456), .B(n_1490), .Y(n_1563) );
INVx3_ASAP7_75t_L g1456 ( .A(n_1457), .Y(n_1456) );
INVx2_ASAP7_75t_L g1493 ( .A(n_1457), .Y(n_1493) );
NAND2xp5_ASAP7_75t_L g1578 ( .A(n_1457), .B(n_1461), .Y(n_1578) );
OR2x2_ASAP7_75t_L g1620 ( .A(n_1457), .B(n_1490), .Y(n_1620) );
AND2x2_ASAP7_75t_L g1457 ( .A(n_1458), .B(n_1459), .Y(n_1457) );
INVx1_ASAP7_75t_L g1460 ( .A(n_1461), .Y(n_1460) );
INVx1_ASAP7_75t_L g1535 ( .A(n_1461), .Y(n_1535) );
NAND2xp5_ASAP7_75t_L g1599 ( .A(n_1461), .B(n_1600), .Y(n_1599) );
INVx1_ASAP7_75t_L g1461 ( .A(n_1462), .Y(n_1461) );
OR2x2_ASAP7_75t_L g1482 ( .A(n_1462), .B(n_1483), .Y(n_1482) );
INVx1_ASAP7_75t_L g1490 ( .A(n_1462), .Y(n_1490) );
AND2x2_ASAP7_75t_L g1499 ( .A(n_1462), .B(n_1483), .Y(n_1499) );
INVx1_ASAP7_75t_L g1516 ( .A(n_1462), .Y(n_1516) );
NAND2xp5_ASAP7_75t_L g1462 ( .A(n_1463), .B(n_1464), .Y(n_1462) );
OAI32xp33_ASAP7_75t_L g1465 ( .A1(n_1466), .A2(n_1468), .A3(n_1474), .B1(n_1475), .B2(n_1478), .Y(n_1465) );
INVx1_ASAP7_75t_L g1466 ( .A(n_1467), .Y(n_1466) );
AND2x2_ASAP7_75t_L g1600 ( .A(n_1467), .B(n_1485), .Y(n_1600) );
AND2x2_ASAP7_75t_L g1525 ( .A(n_1468), .B(n_1526), .Y(n_1525) );
NAND2xp5_ASAP7_75t_SL g1540 ( .A(n_1468), .B(n_1493), .Y(n_1540) );
AND2x2_ASAP7_75t_L g1582 ( .A(n_1468), .B(n_1481), .Y(n_1582) );
OAI21xp5_ASAP7_75t_L g1587 ( .A1(n_1468), .A2(n_1588), .B(n_1590), .Y(n_1587) );
NAND2xp5_ASAP7_75t_L g1594 ( .A(n_1468), .B(n_1486), .Y(n_1594) );
INVx1_ASAP7_75t_L g1468 ( .A(n_1469), .Y(n_1468) );
INVx1_ASAP7_75t_L g1480 ( .A(n_1470), .Y(n_1480) );
AND2x2_ASAP7_75t_L g1507 ( .A(n_1470), .B(n_1508), .Y(n_1507) );
INVx1_ASAP7_75t_L g1470 ( .A(n_1471), .Y(n_1470) );
INVx1_ASAP7_75t_L g1598 ( .A(n_1471), .Y(n_1598) );
NAND2xp5_ASAP7_75t_L g1471 ( .A(n_1472), .B(n_1473), .Y(n_1471) );
OAI21xp33_ASAP7_75t_L g1536 ( .A1(n_1474), .A2(n_1537), .B(n_1539), .Y(n_1536) );
AOI221xp5_ASAP7_75t_L g1624 ( .A1(n_1474), .A2(n_1506), .B1(n_1625), .B2(n_1626), .C(n_1627), .Y(n_1624) );
INVx2_ASAP7_75t_L g1474 ( .A(n_1475), .Y(n_1474) );
AOI22xp33_ASAP7_75t_L g1518 ( .A1(n_1475), .A2(n_1519), .B1(n_1521), .B2(n_1522), .Y(n_1518) );
AND2x2_ASAP7_75t_L g1521 ( .A(n_1475), .B(n_1490), .Y(n_1521) );
CKINVDCx6p67_ASAP7_75t_R g1569 ( .A(n_1475), .Y(n_1569) );
AND2x4_ASAP7_75t_L g1475 ( .A(n_1476), .B(n_1477), .Y(n_1475) );
AND2x2_ASAP7_75t_L g1483 ( .A(n_1476), .B(n_1477), .Y(n_1483) );
AND2x2_ASAP7_75t_L g1479 ( .A(n_1480), .B(n_1481), .Y(n_1479) );
AND2x2_ASAP7_75t_L g1495 ( .A(n_1481), .B(n_1496), .Y(n_1495) );
OR2x2_ASAP7_75t_L g1500 ( .A(n_1481), .B(n_1501), .Y(n_1500) );
AND2x2_ASAP7_75t_L g1506 ( .A(n_1481), .B(n_1507), .Y(n_1506) );
OR2x2_ASAP7_75t_L g1539 ( .A(n_1481), .B(n_1540), .Y(n_1539) );
AND2x2_ASAP7_75t_L g1603 ( .A(n_1481), .B(n_1604), .Y(n_1603) );
OR2x2_ASAP7_75t_L g1510 ( .A(n_1482), .B(n_1511), .Y(n_1510) );
INVx1_ASAP7_75t_L g1585 ( .A(n_1482), .Y(n_1585) );
OR2x2_ASAP7_75t_L g1489 ( .A(n_1483), .B(n_1490), .Y(n_1489) );
AOI21xp33_ASAP7_75t_L g1558 ( .A1(n_1483), .A2(n_1529), .B(n_1559), .Y(n_1558) );
NAND2xp5_ASAP7_75t_SL g1574 ( .A(n_1483), .B(n_1575), .Y(n_1574) );
AND2x2_ASAP7_75t_L g1630 ( .A(n_1483), .B(n_1511), .Y(n_1630) );
INVx1_ASAP7_75t_L g1570 ( .A(n_1484), .Y(n_1570) );
AND2x2_ASAP7_75t_L g1617 ( .A(n_1484), .B(n_1515), .Y(n_1617) );
AND2x2_ASAP7_75t_L g1626 ( .A(n_1484), .B(n_1516), .Y(n_1626) );
AND2x2_ASAP7_75t_L g1484 ( .A(n_1485), .B(n_1486), .Y(n_1484) );
INVx1_ASAP7_75t_L g1501 ( .A(n_1485), .Y(n_1501) );
AOI211xp5_ASAP7_75t_L g1487 ( .A1(n_1488), .A2(n_1491), .B(n_1497), .C(n_1517), .Y(n_1487) );
INVx2_ASAP7_75t_SL g1488 ( .A(n_1489), .Y(n_1488) );
NOR2xp33_ASAP7_75t_L g1572 ( .A(n_1489), .B(n_1573), .Y(n_1572) );
INVx1_ASAP7_75t_L g1491 ( .A(n_1492), .Y(n_1491) );
OR2x2_ASAP7_75t_L g1492 ( .A(n_1493), .B(n_1494), .Y(n_1492) );
INVx2_ASAP7_75t_L g1504 ( .A(n_1493), .Y(n_1504) );
NAND2xp5_ASAP7_75t_SL g1557 ( .A(n_1493), .B(n_1521), .Y(n_1557) );
NAND2xp5_ASAP7_75t_L g1611 ( .A(n_1493), .B(n_1577), .Y(n_1611) );
INVx1_ASAP7_75t_L g1494 ( .A(n_1495), .Y(n_1494) );
INVx1_ASAP7_75t_L g1606 ( .A(n_1496), .Y(n_1606) );
OAI211xp5_ASAP7_75t_L g1497 ( .A1(n_1498), .A2(n_1500), .B(n_1502), .C(n_1512), .Y(n_1497) );
CKINVDCx14_ASAP7_75t_R g1498 ( .A(n_1499), .Y(n_1498) );
NOR2xp33_ASAP7_75t_L g1547 ( .A(n_1500), .B(n_1510), .Y(n_1547) );
OR2x2_ASAP7_75t_L g1589 ( .A(n_1501), .B(n_1526), .Y(n_1589) );
OAI21xp5_ASAP7_75t_L g1502 ( .A1(n_1503), .A2(n_1506), .B(n_1509), .Y(n_1502) );
NOR2xp33_ASAP7_75t_L g1503 ( .A(n_1504), .B(n_1505), .Y(n_1503) );
AOI311xp33_ASAP7_75t_L g1579 ( .A1(n_1504), .A2(n_1549), .A3(n_1580), .B(n_1583), .C(n_1586), .Y(n_1579) );
AND2x2_ASAP7_75t_L g1613 ( .A(n_1504), .B(n_1506), .Y(n_1613) );
INVx1_ASAP7_75t_L g1573 ( .A(n_1506), .Y(n_1573) );
AND2x2_ASAP7_75t_L g1552 ( .A(n_1507), .B(n_1526), .Y(n_1552) );
INVx1_ASAP7_75t_L g1605 ( .A(n_1507), .Y(n_1605) );
INVx1_ASAP7_75t_L g1509 ( .A(n_1510), .Y(n_1509) );
NAND2xp5_ASAP7_75t_L g1584 ( .A(n_1511), .B(n_1585), .Y(n_1584) );
AOI221xp5_ASAP7_75t_L g1553 ( .A1(n_1514), .A2(n_1554), .B1(n_1556), .B2(n_1565), .C(n_1567), .Y(n_1553) );
INVx1_ASAP7_75t_L g1541 ( .A(n_1515), .Y(n_1541) );
INVx1_ASAP7_75t_L g1515 ( .A(n_1516), .Y(n_1515) );
INVx1_ASAP7_75t_L g1522 ( .A(n_1523), .Y(n_1522) );
AOI21xp5_ASAP7_75t_L g1627 ( .A1(n_1524), .A2(n_1628), .B(n_1629), .Y(n_1627) );
CKINVDCx5p33_ASAP7_75t_R g1524 ( .A(n_1525), .Y(n_1524) );
AND2x2_ASAP7_75t_L g1602 ( .A(n_1526), .B(n_1534), .Y(n_1602) );
INVx1_ASAP7_75t_L g1527 ( .A(n_1528), .Y(n_1527) );
INVx1_ASAP7_75t_L g1566 ( .A(n_1529), .Y(n_1566) );
INVx1_ASAP7_75t_L g1529 ( .A(n_1530), .Y(n_1529) );
AND2x2_ASAP7_75t_L g1530 ( .A(n_1531), .B(n_1532), .Y(n_1530) );
AOI221xp5_ASAP7_75t_L g1533 ( .A1(n_1534), .A2(n_1535), .B1(n_1536), .B2(n_1541), .C(n_1542), .Y(n_1533) );
INVxp33_ASAP7_75t_SL g1537 ( .A(n_1538), .Y(n_1537) );
OAI31xp33_ASAP7_75t_L g1609 ( .A1(n_1541), .A2(n_1559), .A3(n_1588), .B(n_1610), .Y(n_1609) );
NOR2xp33_ASAP7_75t_L g1542 ( .A(n_1543), .B(n_1544), .Y(n_1542) );
OAI211xp5_ASAP7_75t_L g1556 ( .A1(n_1543), .A2(n_1557), .B(n_1558), .C(n_1561), .Y(n_1556) );
NAND2xp5_ASAP7_75t_L g1580 ( .A(n_1543), .B(n_1581), .Y(n_1580) );
INVx1_ASAP7_75t_L g1621 ( .A(n_1544), .Y(n_1621) );
NAND3xp33_ASAP7_75t_L g1545 ( .A(n_1546), .B(n_1553), .C(n_1579), .Y(n_1545) );
NOR2xp33_ASAP7_75t_L g1546 ( .A(n_1547), .B(n_1548), .Y(n_1546) );
AND2x2_ASAP7_75t_L g1548 ( .A(n_1549), .B(n_1551), .Y(n_1548) );
AOI22xp33_ASAP7_75t_SL g1592 ( .A1(n_1549), .A2(n_1593), .B1(n_1595), .B2(n_1596), .Y(n_1592) );
INVx1_ASAP7_75t_L g1549 ( .A(n_1550), .Y(n_1549) );
INVx1_ASAP7_75t_L g1623 ( .A(n_1552), .Y(n_1623) );
INVx1_ASAP7_75t_L g1554 ( .A(n_1555), .Y(n_1554) );
INVx1_ASAP7_75t_L g1559 ( .A(n_1560), .Y(n_1559) );
NAND2xp5_ASAP7_75t_L g1561 ( .A(n_1562), .B(n_1564), .Y(n_1561) );
INVx1_ASAP7_75t_L g1562 ( .A(n_1563), .Y(n_1562) );
OAI211xp5_ASAP7_75t_L g1567 ( .A1(n_1568), .A2(n_1570), .B(n_1571), .C(n_1574), .Y(n_1567) );
CKINVDCx6p67_ASAP7_75t_R g1568 ( .A(n_1569), .Y(n_1568) );
INVx1_ASAP7_75t_L g1571 ( .A(n_1572), .Y(n_1571) );
INVxp33_ASAP7_75t_SL g1628 ( .A(n_1575), .Y(n_1628) );
NOR2xp33_ASAP7_75t_L g1575 ( .A(n_1576), .B(n_1578), .Y(n_1575) );
CKINVDCx14_ASAP7_75t_R g1576 ( .A(n_1577), .Y(n_1576) );
INVx1_ASAP7_75t_L g1581 ( .A(n_1582), .Y(n_1581) );
INVxp67_ASAP7_75t_L g1586 ( .A(n_1587), .Y(n_1586) );
INVx1_ASAP7_75t_L g1588 ( .A(n_1589), .Y(n_1588) );
NAND2xp5_ASAP7_75t_L g1622 ( .A(n_1589), .B(n_1623), .Y(n_1622) );
INVx1_ASAP7_75t_L g1593 ( .A(n_1594), .Y(n_1593) );
INVx1_ASAP7_75t_L g1596 ( .A(n_1597), .Y(n_1596) );
O2A1O1Ixp33_ASAP7_75t_L g1601 ( .A1(n_1602), .A2(n_1603), .B(n_1607), .C(n_1608), .Y(n_1601) );
NAND2xp5_ASAP7_75t_L g1604 ( .A(n_1605), .B(n_1606), .Y(n_1604) );
AOI21xp5_ASAP7_75t_L g1608 ( .A1(n_1609), .A2(n_1612), .B(n_1614), .Y(n_1608) );
INVx1_ASAP7_75t_L g1610 ( .A(n_1611), .Y(n_1610) );
INVx1_ASAP7_75t_L g1612 ( .A(n_1613), .Y(n_1612) );
INVx1_ASAP7_75t_L g1616 ( .A(n_1617), .Y(n_1616) );
OAI21xp33_ASAP7_75t_L g1618 ( .A1(n_1619), .A2(n_1621), .B(n_1622), .Y(n_1618) );
INVx1_ASAP7_75t_L g1629 ( .A(n_1630), .Y(n_1629) );
CKINVDCx20_ASAP7_75t_R g1631 ( .A(n_1632), .Y(n_1631) );
BUFx2_ASAP7_75t_SL g1634 ( .A(n_1635), .Y(n_1634) );
BUFx3_ASAP7_75t_L g1635 ( .A(n_1636), .Y(n_1635) );
INVxp33_ASAP7_75t_L g1637 ( .A(n_1638), .Y(n_1637) );
HB1xp67_ASAP7_75t_L g1639 ( .A(n_1640), .Y(n_1639) );
AND4x1_ASAP7_75t_L g1640 ( .A(n_1641), .B(n_1644), .C(n_1657), .D(n_1670), .Y(n_1640) );
OAI211xp5_ASAP7_75t_L g1666 ( .A1(n_1653), .A2(n_1667), .B(n_1668), .C(n_1669), .Y(n_1666) );
HB1xp67_ASAP7_75t_L g1671 ( .A(n_1672), .Y(n_1671) );
OAI21xp5_ASAP7_75t_L g1672 ( .A1(n_1673), .A2(n_1674), .B(n_1675), .Y(n_1672) );
INVx1_ASAP7_75t_L g1675 ( .A(n_1676), .Y(n_1675) );
INVxp67_ASAP7_75t_L g1678 ( .A(n_1679), .Y(n_1678) );
BUFx3_ASAP7_75t_L g1679 ( .A(n_1680), .Y(n_1679) );
INVx3_ASAP7_75t_L g1680 ( .A(n_1681), .Y(n_1680) );
INVx1_ASAP7_75t_L g1682 ( .A(n_1683), .Y(n_1682) );
endmodule