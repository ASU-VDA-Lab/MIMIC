module fake_jpeg_29783_n_55 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_55);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_55;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_3),
.Y(n_7)
);

INVx6_ASAP7_75t_SL g8 ( 
.A(n_5),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_0),
.B(n_4),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

INVx4_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx5_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

AND2x2_ASAP7_75t_L g14 ( 
.A(n_6),
.B(n_3),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_15),
.B(n_16),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_14),
.B(n_9),
.Y(n_16)
);

AO22x2_ASAP7_75t_L g17 ( 
.A1(n_14),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g27 ( 
.A1(n_17),
.A2(n_18),
.B(n_1),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_SL g18 ( 
.A1(n_14),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_14),
.B(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_19),
.Y(n_29)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_10),
.A2(n_6),
.B1(n_1),
.B2(n_2),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_21),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_10),
.B(n_0),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_22),
.B(n_11),
.C(n_12),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_17),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_15),
.A2(n_16),
.B1(n_19),
.B2(n_18),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_24),
.A2(n_26),
.B1(n_27),
.B2(n_30),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_22),
.A2(n_7),
.B1(n_12),
.B2(n_11),
.Y(n_26)
);

XOR2xp5_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_21),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_32),
.C(n_36),
.Y(n_38)
);

CKINVDCx14_ASAP7_75t_R g33 ( 
.A(n_27),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_33),
.Y(n_37)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_35),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_29),
.A2(n_17),
.B1(n_20),
.B2(n_8),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_29),
.C(n_23),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_40),
.C(n_37),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_28),
.C(n_26),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_34),
.A2(n_30),
.B1(n_17),
.B2(n_7),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_32),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_38),
.B(n_35),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_43),
.B(n_44),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_42),
.B(n_36),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g48 ( 
.A1(n_45),
.A2(n_46),
.B(n_17),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_37),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_47),
.B(n_17),
.C(n_7),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_SL g53 ( 
.A1(n_48),
.A2(n_51),
.B(n_13),
.Y(n_53)
);

MAJx2_ASAP7_75t_L g52 ( 
.A(n_50),
.B(n_13),
.C(n_12),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_SL g51 ( 
.A1(n_44),
.A2(n_8),
.B(n_13),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_52),
.B(n_53),
.C(n_49),
.Y(n_54)
);

OAI21x1_ASAP7_75t_L g55 ( 
.A1(n_54),
.A2(n_12),
.B(n_2),
.Y(n_55)
);


endmodule