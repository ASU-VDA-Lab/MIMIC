module real_aes_8136_n_222 (n_17, n_28, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_165, n_51, n_195, n_176, n_27, n_163, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_84, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_16, n_116, n_94, n_39, n_5, n_45, n_60, n_38, n_155, n_118, n_143, n_139, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_107, n_184, n_53, n_36, n_222);
input n_17;
input n_28;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_84;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_16;
input n_116;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_107;
input n_184;
input n_53;
input n_36;
output n_222;
wire n_480;
wire n_476;
wire n_599;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_631;
wire n_357;
wire n_503;
wire n_287;
wire n_635;
wire n_673;
wire n_386;
wire n_518;
wire n_254;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_461;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_578;
wire n_372;
wire n_528;
wire n_495;
wire n_370;
wire n_384;
wire n_352;
wire n_467;
wire n_327;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_281;
wire n_496;
wire n_693;
wire n_468;
wire n_234;
wire n_284;
wire n_316;
wire n_656;
wire n_532;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_617;
wire n_552;
wire n_402;
wire n_602;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_246;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_392;
wire n_562;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_269;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_649;
wire n_663;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_498;
wire n_481;
wire n_691;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_472;
wire n_452;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_681;
wire n_359;
wire n_456;
wire n_717;
wire n_712;
wire n_266;
wire n_312;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_705;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_541;
wire n_224;
wire n_546;
wire n_587;
wire n_639;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_228;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_0), .A2(n_129), .B1(n_351), .B2(n_526), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g670 ( .A1(n_1), .A2(n_41), .B1(n_399), .B2(n_599), .Y(n_670) );
CKINVDCx20_ASAP7_75t_R g482 ( .A(n_2), .Y(n_482) );
CKINVDCx20_ASAP7_75t_R g654 ( .A(n_3), .Y(n_654) );
AOI22xp33_ASAP7_75t_SL g669 ( .A1(n_4), .A2(n_214), .B1(n_306), .B2(n_309), .Y(n_669) );
AOI22xp33_ASAP7_75t_SL g587 ( .A1(n_5), .A2(n_29), .B1(n_358), .B2(n_588), .Y(n_587) );
AOI22xp5_ASAP7_75t_L g698 ( .A1(n_6), .A2(n_102), .B1(n_347), .B2(n_399), .Y(n_698) );
CKINVDCx20_ASAP7_75t_R g534 ( .A(n_7), .Y(n_534) );
CKINVDCx20_ASAP7_75t_R g492 ( .A(n_8), .Y(n_492) );
AOI22xp33_ASAP7_75t_L g467 ( .A1(n_9), .A2(n_39), .B1(n_313), .B2(n_468), .Y(n_467) );
AOI22xp33_ASAP7_75t_SL g335 ( .A1(n_10), .A2(n_103), .B1(n_262), .B2(n_336), .Y(n_335) );
AOI22xp33_ASAP7_75t_SL g719 ( .A1(n_11), .A2(n_116), .B1(n_293), .B2(n_316), .Y(n_719) );
AOI22xp33_ASAP7_75t_L g354 ( .A1(n_12), .A2(n_219), .B1(n_315), .B2(n_355), .Y(n_354) );
CKINVDCx20_ASAP7_75t_R g377 ( .A(n_13), .Y(n_377) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_14), .A2(n_178), .B1(n_395), .B2(n_400), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g637 ( .A1(n_15), .A2(n_31), .B1(n_599), .B2(n_638), .Y(n_637) );
CKINVDCx20_ASAP7_75t_R g382 ( .A(n_16), .Y(n_382) );
CKINVDCx20_ASAP7_75t_R g371 ( .A(n_17), .Y(n_371) );
AOI22xp33_ASAP7_75t_L g627 ( .A1(n_18), .A2(n_108), .B1(n_520), .B2(n_552), .Y(n_627) );
CKINVDCx20_ASAP7_75t_R g655 ( .A(n_19), .Y(n_655) );
AOI22xp33_ASAP7_75t_L g388 ( .A1(n_20), .A2(n_165), .B1(n_242), .B2(n_389), .Y(n_388) );
AOI22x1_ASAP7_75t_L g408 ( .A1(n_21), .A2(n_409), .B1(n_457), .B2(n_458), .Y(n_408) );
INVx1_ASAP7_75t_L g457 ( .A(n_21), .Y(n_457) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_22), .A2(n_212), .B1(n_551), .B2(n_604), .Y(n_603) );
AO22x2_ASAP7_75t_L g245 ( .A1(n_23), .A2(n_77), .B1(n_246), .B2(n_247), .Y(n_245) );
INVx1_ASAP7_75t_L g686 ( .A(n_23), .Y(n_686) );
CKINVDCx20_ASAP7_75t_R g613 ( .A(n_24), .Y(n_613) );
AOI22xp33_ASAP7_75t_L g464 ( .A1(n_25), .A2(n_58), .B1(n_465), .B2(n_466), .Y(n_464) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_26), .A2(n_192), .B1(n_399), .B2(n_599), .Y(n_598) );
CKINVDCx20_ASAP7_75t_R g450 ( .A(n_27), .Y(n_450) );
CKINVDCx20_ASAP7_75t_R g329 ( .A(n_28), .Y(n_329) );
AOI22xp5_ASAP7_75t_L g697 ( .A1(n_30), .A2(n_208), .B1(n_358), .B2(n_391), .Y(n_697) );
AOI22xp33_ASAP7_75t_L g312 ( .A1(n_32), .A2(n_110), .B1(n_313), .B2(n_316), .Y(n_312) );
CKINVDCx20_ASAP7_75t_R g444 ( .A(n_33), .Y(n_444) );
AOI22xp33_ASAP7_75t_SL g582 ( .A1(n_34), .A2(n_151), .B1(n_349), .B2(n_583), .Y(n_582) );
CKINVDCx20_ASAP7_75t_R g601 ( .A(n_35), .Y(n_601) );
CKINVDCx20_ASAP7_75t_R g327 ( .A(n_36), .Y(n_327) );
AOI22xp33_ASAP7_75t_L g348 ( .A1(n_37), .A2(n_84), .B1(n_349), .B2(n_351), .Y(n_348) );
AOI22xp33_ASAP7_75t_L g729 ( .A1(n_38), .A2(n_215), .B1(n_280), .B2(n_284), .Y(n_729) );
AO22x2_ASAP7_75t_L g249 ( .A1(n_40), .A2(n_79), .B1(n_246), .B2(n_250), .Y(n_249) );
INVx1_ASAP7_75t_L g687 ( .A(n_40), .Y(n_687) );
AOI22xp33_ASAP7_75t_SL g584 ( .A1(n_42), .A2(n_83), .B1(n_399), .B2(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g479 ( .A(n_43), .Y(n_479) );
AOI22xp33_ASAP7_75t_SL g555 ( .A1(n_44), .A2(n_152), .B1(n_389), .B2(n_395), .Y(n_555) );
CKINVDCx20_ASAP7_75t_R g701 ( .A(n_45), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_46), .B(n_268), .Y(n_602) );
CKINVDCx20_ASAP7_75t_R g648 ( .A(n_47), .Y(n_648) );
AOI22xp5_ASAP7_75t_L g695 ( .A1(n_48), .A2(n_164), .B1(n_316), .B2(n_397), .Y(n_695) );
AOI22xp33_ASAP7_75t_L g720 ( .A1(n_49), .A2(n_221), .B1(n_638), .B2(n_721), .Y(n_720) );
CKINVDCx20_ASAP7_75t_R g415 ( .A(n_50), .Y(n_415) );
AOI22xp5_ASAP7_75t_L g666 ( .A1(n_51), .A2(n_76), .B1(n_292), .B2(n_389), .Y(n_666) );
CKINVDCx20_ASAP7_75t_R g623 ( .A(n_52), .Y(n_623) );
AOI22xp33_ASAP7_75t_L g297 ( .A1(n_53), .A2(n_91), .B1(n_298), .B2(n_300), .Y(n_297) );
AOI22xp5_ASAP7_75t_L g256 ( .A1(n_54), .A2(n_181), .B1(n_257), .B2(n_262), .Y(n_256) );
AOI22xp33_ASAP7_75t_SL g305 ( .A1(n_55), .A2(n_184), .B1(n_306), .B2(n_309), .Y(n_305) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_56), .A2(n_106), .B1(n_290), .B2(n_417), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_57), .A2(n_69), .B1(n_345), .B2(n_524), .Y(n_523) );
CKINVDCx20_ASAP7_75t_R g658 ( .A(n_59), .Y(n_658) );
CKINVDCx20_ASAP7_75t_R g663 ( .A(n_60), .Y(n_663) );
CKINVDCx20_ASAP7_75t_R g629 ( .A(n_61), .Y(n_629) );
CKINVDCx20_ASAP7_75t_R g544 ( .A(n_62), .Y(n_544) );
CKINVDCx20_ASAP7_75t_R g421 ( .A(n_63), .Y(n_421) );
CKINVDCx20_ASAP7_75t_R g333 ( .A(n_64), .Y(n_333) );
AOI22xp5_ASAP7_75t_L g705 ( .A1(n_65), .A2(n_111), .B1(n_443), .B2(n_520), .Y(n_705) );
AOI22xp33_ASAP7_75t_L g471 ( .A1(n_66), .A2(n_175), .B1(n_472), .B2(n_473), .Y(n_471) );
AOI22xp33_ASAP7_75t_L g337 ( .A1(n_67), .A2(n_173), .B1(n_338), .B2(n_340), .Y(n_337) );
CKINVDCx20_ASAP7_75t_R g436 ( .A(n_68), .Y(n_436) );
CKINVDCx20_ASAP7_75t_R g704 ( .A(n_70), .Y(n_704) );
AOI22xp5_ASAP7_75t_L g474 ( .A1(n_71), .A2(n_85), .B1(n_428), .B2(n_475), .Y(n_474) );
AOI222xp33_ASAP7_75t_L g609 ( .A1(n_72), .A2(n_130), .B1(n_135), .B2(n_262), .C1(n_610), .C2(n_612), .Y(n_609) );
CKINVDCx20_ASAP7_75t_R g642 ( .A(n_73), .Y(n_642) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_74), .A2(n_149), .B1(n_347), .B2(n_395), .Y(n_667) );
AOI22xp33_ASAP7_75t_L g702 ( .A1(n_75), .A2(n_121), .B1(n_284), .B2(n_513), .Y(n_702) );
CKINVDCx20_ASAP7_75t_R g713 ( .A(n_78), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_80), .B(n_508), .Y(n_507) );
AOI22xp33_ASAP7_75t_SL g580 ( .A1(n_81), .A2(n_205), .B1(n_326), .B2(n_379), .Y(n_580) );
AND2x2_ASAP7_75t_L g229 ( .A(n_82), .B(n_230), .Y(n_229) );
AOI22xp33_ASAP7_75t_L g426 ( .A1(n_86), .A2(n_150), .B1(n_427), .B2(n_428), .Y(n_426) );
CKINVDCx20_ASAP7_75t_R g592 ( .A(n_87), .Y(n_592) );
INVx1_ASAP7_75t_L g226 ( .A(n_88), .Y(n_226) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_89), .A2(n_138), .B1(n_389), .B2(n_607), .Y(n_606) );
AOI211xp5_ASAP7_75t_L g222 ( .A1(n_90), .A2(n_223), .B(n_231), .C(n_688), .Y(n_222) );
AOI22xp33_ASAP7_75t_L g356 ( .A1(n_92), .A2(n_120), .B1(n_308), .B2(n_357), .Y(n_356) );
AOI22xp33_ASAP7_75t_L g378 ( .A1(n_93), .A2(n_109), .B1(n_258), .B2(n_379), .Y(n_378) );
AOI22xp5_ASAP7_75t_L g659 ( .A1(n_94), .A2(n_210), .B1(n_258), .B2(n_552), .Y(n_659) );
AOI22xp5_ASAP7_75t_L g693 ( .A1(n_95), .A2(n_187), .B1(n_560), .B2(n_694), .Y(n_693) );
AOI22xp33_ASAP7_75t_SL g550 ( .A1(n_96), .A2(n_100), .B1(n_551), .B2(n_552), .Y(n_550) );
OA22x2_ASAP7_75t_L g538 ( .A1(n_97), .A2(n_539), .B1(n_540), .B2(n_563), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_97), .Y(n_539) );
CKINVDCx20_ASAP7_75t_R g531 ( .A(n_98), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_99), .B(n_276), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_101), .B(n_339), .Y(n_549) );
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_104), .A2(n_107), .B1(n_349), .B2(n_597), .Y(n_596) );
OA22x2_ASAP7_75t_L g362 ( .A1(n_105), .A2(n_363), .B1(n_364), .B2(n_401), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_105), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_112), .B(n_578), .Y(n_577) );
CKINVDCx20_ASAP7_75t_R g445 ( .A(n_113), .Y(n_445) );
CKINVDCx20_ASAP7_75t_R g700 ( .A(n_114), .Y(n_700) );
AOI22xp33_ASAP7_75t_L g344 ( .A1(n_115), .A2(n_186), .B1(n_345), .B2(n_347), .Y(n_344) );
INVx2_ASAP7_75t_L g230 ( .A(n_117), .Y(n_230) );
XOR2xp5_ASAP7_75t_L g689 ( .A(n_118), .B(n_690), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_119), .B(n_548), .Y(n_547) );
CKINVDCx20_ASAP7_75t_R g500 ( .A(n_122), .Y(n_500) );
CKINVDCx20_ASAP7_75t_R g412 ( .A(n_123), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_124), .B(n_509), .Y(n_727) );
CKINVDCx20_ASAP7_75t_R g486 ( .A(n_125), .Y(n_486) );
CKINVDCx20_ASAP7_75t_R g515 ( .A(n_126), .Y(n_515) );
AND2x6_ASAP7_75t_L g225 ( .A(n_127), .B(n_226), .Y(n_225) );
HB1xp67_ASAP7_75t_L g680 ( .A(n_127), .Y(n_680) );
AO22x2_ASAP7_75t_L g253 ( .A1(n_128), .A2(n_176), .B1(n_246), .B2(n_250), .Y(n_253) );
AOI22xp33_ASAP7_75t_L g725 ( .A1(n_131), .A2(n_204), .B1(n_332), .B2(n_513), .Y(n_725) );
AOI22xp33_ASAP7_75t_L g394 ( .A1(n_132), .A2(n_200), .B1(n_395), .B2(n_397), .Y(n_394) );
CKINVDCx20_ASAP7_75t_R g485 ( .A(n_133), .Y(n_485) );
CKINVDCx20_ASAP7_75t_R g240 ( .A(n_134), .Y(n_240) );
AOI22xp33_ASAP7_75t_L g390 ( .A1(n_136), .A2(n_161), .B1(n_391), .B2(n_392), .Y(n_390) );
AOI22xp33_ASAP7_75t_SL g562 ( .A1(n_137), .A2(n_206), .B1(n_315), .B2(n_347), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g279 ( .A1(n_139), .A2(n_146), .B1(n_280), .B2(n_284), .Y(n_279) );
AOI22xp5_ASAP7_75t_L g635 ( .A1(n_140), .A2(n_160), .B1(n_308), .B2(n_636), .Y(n_635) );
AOI22xp33_ASAP7_75t_SL g559 ( .A1(n_141), .A2(n_197), .B1(n_560), .B2(n_561), .Y(n_559) );
CKINVDCx20_ASAP7_75t_R g491 ( .A(n_142), .Y(n_491) );
AOI22xp33_ASAP7_75t_L g289 ( .A1(n_143), .A2(n_220), .B1(n_290), .B2(n_293), .Y(n_289) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_144), .A2(n_168), .B1(n_336), .B2(n_511), .Y(n_510) );
AO22x2_ASAP7_75t_L g255 ( .A1(n_145), .A2(n_194), .B1(n_246), .B2(n_247), .Y(n_255) );
AOI22xp33_ASAP7_75t_L g733 ( .A1(n_147), .A2(n_182), .B1(n_298), .B2(n_309), .Y(n_733) );
AOI22xp5_ASAP7_75t_L g460 ( .A1(n_148), .A2(n_461), .B1(n_493), .B2(n_494), .Y(n_460) );
INVx1_ASAP7_75t_L g493 ( .A(n_148), .Y(n_493) );
AOI22xp33_ASAP7_75t_SL g556 ( .A1(n_153), .A2(n_177), .B1(n_476), .B2(n_557), .Y(n_556) );
CKINVDCx20_ASAP7_75t_R g381 ( .A(n_154), .Y(n_381) );
CKINVDCx20_ASAP7_75t_R g626 ( .A(n_155), .Y(n_626) );
AOI22xp33_ASAP7_75t_SL g545 ( .A1(n_156), .A2(n_196), .B1(n_280), .B2(n_520), .Y(n_545) );
AOI22xp33_ASAP7_75t_SL g589 ( .A1(n_157), .A2(n_190), .B1(n_590), .B2(n_591), .Y(n_589) );
AOI22xp33_ASAP7_75t_SL g731 ( .A1(n_158), .A2(n_216), .B1(n_420), .B2(n_732), .Y(n_731) );
CKINVDCx20_ASAP7_75t_R g425 ( .A(n_159), .Y(n_425) );
CKINVDCx20_ASAP7_75t_R g529 ( .A(n_162), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_163), .B(n_277), .Y(n_728) );
CKINVDCx20_ASAP7_75t_R g505 ( .A(n_166), .Y(n_505) );
CKINVDCx20_ASAP7_75t_R g624 ( .A(n_167), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_169), .B(n_268), .Y(n_267) );
AOI22xp33_ASAP7_75t_SL g575 ( .A1(n_170), .A2(n_202), .B1(n_257), .B2(n_552), .Y(n_575) );
NAND2xp5_ASAP7_75t_SL g579 ( .A(n_171), .B(n_338), .Y(n_579) );
CKINVDCx20_ASAP7_75t_R g647 ( .A(n_172), .Y(n_647) );
CKINVDCx20_ASAP7_75t_R g367 ( .A(n_174), .Y(n_367) );
NOR2xp33_ASAP7_75t_L g684 ( .A(n_176), .B(n_685), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_179), .B(n_488), .Y(n_487) );
CKINVDCx20_ASAP7_75t_R g448 ( .A(n_180), .Y(n_448) );
CKINVDCx20_ASAP7_75t_R g724 ( .A(n_183), .Y(n_724) );
INVx1_ASAP7_75t_L g671 ( .A(n_185), .Y(n_671) );
CKINVDCx20_ASAP7_75t_R g318 ( .A(n_188), .Y(n_318) );
OA22x2_ASAP7_75t_L g320 ( .A1(n_189), .A2(n_321), .B1(n_322), .B2(n_359), .Y(n_320) );
CKINVDCx20_ASAP7_75t_R g321 ( .A(n_189), .Y(n_321) );
CKINVDCx20_ASAP7_75t_R g535 ( .A(n_191), .Y(n_535) );
CKINVDCx20_ASAP7_75t_R g432 ( .A(n_193), .Y(n_432) );
INVx1_ASAP7_75t_L g683 ( .A(n_194), .Y(n_683) );
AOI211xp5_ASAP7_75t_L g502 ( .A1(n_195), .A2(n_503), .B(n_504), .C(n_514), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g398 ( .A1(n_198), .A2(n_201), .B1(n_399), .B2(n_400), .Y(n_398) );
CKINVDCx20_ASAP7_75t_R g574 ( .A(n_199), .Y(n_574) );
CKINVDCx20_ASAP7_75t_R g640 ( .A(n_203), .Y(n_640) );
INVx1_ASAP7_75t_L g246 ( .A(n_207), .Y(n_246) );
INVx1_ASAP7_75t_L g248 ( .A(n_207), .Y(n_248) );
CKINVDCx20_ASAP7_75t_R g631 ( .A(n_209), .Y(n_631) );
CKINVDCx20_ASAP7_75t_R g516 ( .A(n_211), .Y(n_516) );
OA22x2_ASAP7_75t_L g616 ( .A1(n_213), .A2(n_617), .B1(n_618), .B2(n_619), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_213), .Y(n_617) );
CKINVDCx20_ASAP7_75t_R g454 ( .A(n_217), .Y(n_454) );
CKINVDCx20_ASAP7_75t_R g661 ( .A(n_218), .Y(n_661) );
INVx1_ASAP7_75t_SL g223 ( .A(n_224), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_225), .B(n_227), .Y(n_224) );
HB1xp67_ASAP7_75t_L g679 ( .A(n_226), .Y(n_679) );
OAI21xp5_ASAP7_75t_L g711 ( .A1(n_227), .A2(n_678), .B(n_712), .Y(n_711) );
CKINVDCx20_ASAP7_75t_R g227 ( .A(n_228), .Y(n_227) );
INVxp67_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
AOI221xp5_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_566), .B1(n_673), .B2(n_674), .C(n_675), .Y(n_231) );
INVx1_ASAP7_75t_L g673 ( .A(n_232), .Y(n_673) );
XOR2xp5_ASAP7_75t_L g232 ( .A(n_233), .B(n_405), .Y(n_232) );
AOI22xp5_ASAP7_75t_L g233 ( .A1(n_234), .A2(n_235), .B1(n_319), .B2(n_404), .Y(n_233) );
INVx2_ASAP7_75t_SL g234 ( .A(n_235), .Y(n_234) );
INVx3_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
XOR2x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_318), .Y(n_236) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_238), .B(n_287), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_239), .B(n_266), .Y(n_238) );
OAI21xp5_ASAP7_75t_L g239 ( .A1(n_240), .A2(n_241), .B(n_256), .Y(n_239) );
INVx2_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
INVx2_ASAP7_75t_SL g328 ( .A(n_242), .Y(n_328) );
BUFx6f_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
INVx2_ASAP7_75t_SL g484 ( .A(n_243), .Y(n_484) );
BUFx3_ASAP7_75t_L g503 ( .A(n_243), .Y(n_503) );
INVx2_ASAP7_75t_L g573 ( .A(n_243), .Y(n_573) );
INVx4_ASAP7_75t_L g611 ( .A(n_243), .Y(n_611) );
AND2x6_ASAP7_75t_L g243 ( .A(n_244), .B(n_251), .Y(n_243) );
AND2x4_ASAP7_75t_L g263 ( .A(n_244), .B(n_264), .Y(n_263) );
INVx1_ASAP7_75t_L g384 ( .A(n_244), .Y(n_384) );
AND2x2_ASAP7_75t_L g244 ( .A(n_245), .B(n_249), .Y(n_244) );
AND2x2_ASAP7_75t_L g261 ( .A(n_245), .B(n_253), .Y(n_261) );
INVx2_ASAP7_75t_L g274 ( .A(n_245), .Y(n_274) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
INVx1_ASAP7_75t_L g250 ( .A(n_248), .Y(n_250) );
OR2x2_ASAP7_75t_L g273 ( .A(n_249), .B(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g278 ( .A(n_249), .B(n_274), .Y(n_278) );
INVx2_ASAP7_75t_L g283 ( .A(n_249), .Y(n_283) );
INVx1_ASAP7_75t_L g286 ( .A(n_249), .Y(n_286) );
AND2x6_ASAP7_75t_L g292 ( .A(n_251), .B(n_272), .Y(n_292) );
AND2x2_ASAP7_75t_L g299 ( .A(n_251), .B(n_296), .Y(n_299) );
AND2x4_ASAP7_75t_L g308 ( .A(n_251), .B(n_278), .Y(n_308) );
AND2x2_ASAP7_75t_L g251 ( .A(n_252), .B(n_254), .Y(n_251) );
AND2x2_ASAP7_75t_L g271 ( .A(n_252), .B(n_255), .Y(n_271) );
INVx2_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g295 ( .A(n_253), .B(n_265), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_253), .B(n_255), .Y(n_303) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
INVx1_ASAP7_75t_L g260 ( .A(n_255), .Y(n_260) );
INVx1_ASAP7_75t_L g265 ( .A(n_255), .Y(n_265) );
BUFx3_ASAP7_75t_L g447 ( .A(n_257), .Y(n_447) );
INVx2_ASAP7_75t_L g489 ( .A(n_257), .Y(n_489) );
BUFx6f_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
BUFx6f_ASAP7_75t_L g332 ( .A(n_258), .Y(n_332) );
BUFx12f_ASAP7_75t_L g520 ( .A(n_258), .Y(n_520) );
AND2x4_ASAP7_75t_L g258 ( .A(n_259), .B(n_261), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g282 ( .A(n_260), .B(n_283), .Y(n_282) );
AND2x4_ASAP7_75t_L g281 ( .A(n_261), .B(n_282), .Y(n_281) );
AND2x4_ASAP7_75t_L g284 ( .A(n_261), .B(n_285), .Y(n_284) );
NAND2x1p5_ASAP7_75t_L g453 ( .A(n_261), .B(n_317), .Y(n_453) );
BUFx2_ASAP7_75t_SL g262 ( .A(n_263), .Y(n_262) );
BUFx6f_ASAP7_75t_L g513 ( .A(n_263), .Y(n_513) );
BUFx2_ASAP7_75t_SL g552 ( .A(n_263), .Y(n_552) );
INVx1_ASAP7_75t_L g385 ( .A(n_264), .Y(n_385) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
NAND3xp33_ASAP7_75t_L g266 ( .A(n_267), .B(n_275), .C(n_279), .Y(n_266) );
INVx2_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
INVx5_ASAP7_75t_L g339 ( .A(n_269), .Y(n_339) );
INVx2_ASAP7_75t_L g509 ( .A(n_269), .Y(n_509) );
INVx4_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
AND2x4_ASAP7_75t_L g270 ( .A(n_271), .B(n_272), .Y(n_270) );
AND2x6_ASAP7_75t_L g277 ( .A(n_271), .B(n_278), .Y(n_277) );
AND2x4_ASAP7_75t_L g315 ( .A(n_271), .B(n_296), .Y(n_315) );
INVx1_ASAP7_75t_L g370 ( .A(n_271), .Y(n_370) );
NAND2x1p5_ASAP7_75t_L g374 ( .A(n_271), .B(n_278), .Y(n_374) );
INVx2_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
OR2x2_ASAP7_75t_L g369 ( .A(n_273), .B(n_370), .Y(n_369) );
AND2x2_ASAP7_75t_L g296 ( .A(n_274), .B(n_283), .Y(n_296) );
BUFx4f_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
INVx1_ASAP7_75t_SL g341 ( .A(n_277), .Y(n_341) );
BUFx2_ASAP7_75t_L g578 ( .A(n_277), .Y(n_578) );
AND2x2_ASAP7_75t_L g311 ( .A(n_278), .B(n_295), .Y(n_311) );
BUFx4f_ASAP7_75t_SL g280 ( .A(n_281), .Y(n_280) );
BUFx6f_ASAP7_75t_L g326 ( .A(n_281), .Y(n_326) );
BUFx2_ASAP7_75t_L g392 ( .A(n_281), .Y(n_392) );
BUFx6f_ASAP7_75t_L g443 ( .A(n_281), .Y(n_443) );
BUFx6f_ASAP7_75t_L g604 ( .A(n_281), .Y(n_604) );
INVx1_ASAP7_75t_L g317 ( .A(n_283), .Y(n_317) );
BUFx2_ASAP7_75t_L g336 ( .A(n_284), .Y(n_336) );
BUFx2_ASAP7_75t_L g379 ( .A(n_284), .Y(n_379) );
BUFx3_ASAP7_75t_L g551 ( .A(n_284), .Y(n_551) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
OR2x6_ASAP7_75t_L g352 ( .A(n_286), .B(n_303), .Y(n_352) );
NOR2x1_ASAP7_75t_L g287 ( .A(n_288), .B(n_304), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_289), .B(n_297), .Y(n_288) );
INVx4_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx5_ASAP7_75t_SL g355 ( .A(n_291), .Y(n_355) );
INVx1_ASAP7_75t_L g607 ( .A(n_291), .Y(n_607) );
INVx2_ASAP7_75t_SL g732 ( .A(n_291), .Y(n_732) );
INVx11_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
INVx11_ASAP7_75t_L g376 ( .A(n_292), .Y(n_376) );
BUFx3_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
BUFx3_ASAP7_75t_L g358 ( .A(n_294), .Y(n_358) );
BUFx3_ASAP7_75t_L g389 ( .A(n_294), .Y(n_389) );
AND2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_295), .B(n_296), .Y(n_424) );
AND2x4_ASAP7_75t_L g301 ( .A(n_296), .B(n_302), .Y(n_301) );
INVx3_ASAP7_75t_L g346 ( .A(n_298), .Y(n_346) );
BUFx3_ASAP7_75t_L g472 ( .A(n_298), .Y(n_472) );
BUFx6f_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx2_ASAP7_75t_L g396 ( .A(n_299), .Y(n_396) );
BUFx2_ASAP7_75t_SL g590 ( .A(n_299), .Y(n_590) );
HB1xp67_ASAP7_75t_L g417 ( .A(n_300), .Y(n_417) );
BUFx3_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
BUFx2_ASAP7_75t_L g347 ( .A(n_301), .Y(n_347) );
BUFx3_ASAP7_75t_L g400 ( .A(n_301), .Y(n_400) );
BUFx3_ASAP7_75t_L g469 ( .A(n_301), .Y(n_469) );
BUFx2_ASAP7_75t_SL g591 ( .A(n_301), .Y(n_591) );
BUFx2_ASAP7_75t_SL g644 ( .A(n_301), .Y(n_644) );
BUFx3_ASAP7_75t_L g721 ( .A(n_301), .Y(n_721) );
AND2x2_ASAP7_75t_L g316 ( .A(n_302), .B(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_305), .B(n_312), .Y(n_304) );
INVxp67_ASAP7_75t_L g530 ( .A(n_306), .Y(n_530) );
INVx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx3_ASAP7_75t_L g561 ( .A(n_307), .Y(n_561) );
INVx2_ASAP7_75t_L g583 ( .A(n_307), .Y(n_583) );
INVx2_ASAP7_75t_L g597 ( .A(n_307), .Y(n_597) );
INVx6_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
BUFx3_ASAP7_75t_L g391 ( .A(n_308), .Y(n_391) );
BUFx3_ASAP7_75t_L g420 ( .A(n_308), .Y(n_420) );
BUFx3_ASAP7_75t_L g465 ( .A(n_308), .Y(n_465) );
INVx3_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
BUFx3_ASAP7_75t_L g350 ( .A(n_310), .Y(n_350) );
INVx5_ASAP7_75t_L g397 ( .A(n_310), .Y(n_397) );
INVx4_ASAP7_75t_L g476 ( .A(n_310), .Y(n_476) );
INVx1_ASAP7_75t_L g636 ( .A(n_310), .Y(n_636) );
INVx8_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx2_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
OAI22xp5_ASAP7_75t_L g533 ( .A1(n_314), .A2(n_534), .B1(n_535), .B2(n_536), .Y(n_533) );
INVx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
BUFx3_ASAP7_75t_L g399 ( .A(n_315), .Y(n_399) );
BUFx3_ASAP7_75t_L g638 ( .A(n_315), .Y(n_638) );
INVx1_ASAP7_75t_L g404 ( .A(n_319), .Y(n_404) );
AOI22xp5_ASAP7_75t_L g319 ( .A1(n_320), .A2(n_360), .B1(n_402), .B2(n_403), .Y(n_319) );
INVx1_ASAP7_75t_L g402 ( .A(n_320), .Y(n_402) );
INVx1_ASAP7_75t_SL g359 ( .A(n_322), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_323), .B(n_342), .Y(n_322) );
NOR2x1_ASAP7_75t_L g323 ( .A(n_324), .B(n_334), .Y(n_323) );
OAI222xp33_ASAP7_75t_L g324 ( .A1(n_325), .A2(n_327), .B1(n_328), .B2(n_329), .C1(n_330), .C2(n_333), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
OAI222xp33_ASAP7_75t_L g440 ( .A1(n_328), .A2(n_441), .B1(n_444), .B2(n_445), .C1(n_446), .C2(n_448), .Y(n_440) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
BUFx4f_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_335), .B(n_337), .Y(n_334) );
BUFx6f_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_SL g340 ( .A(n_341), .Y(n_340) );
INVx1_ASAP7_75t_SL g548 ( .A(n_341), .Y(n_548) );
NOR2xp33_ASAP7_75t_L g342 ( .A(n_343), .B(n_353), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_344), .B(n_348), .Y(n_343) );
INVx2_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
OAI221xp5_ASAP7_75t_SL g411 ( .A1(n_346), .A2(n_412), .B1(n_413), .B2(n_415), .C(n_416), .Y(n_411) );
INVx3_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_SL g351 ( .A(n_352), .Y(n_351) );
OAI22xp5_ASAP7_75t_L g380 ( .A1(n_352), .A2(n_381), .B1(n_382), .B2(n_383), .Y(n_380) );
INVx6_ASAP7_75t_SL g429 ( .A(n_352), .Y(n_429) );
INVx1_ASAP7_75t_SL g557 ( .A(n_352), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_354), .B(n_356), .Y(n_353) );
HB1xp67_ASAP7_75t_L g524 ( .A(n_355), .Y(n_524) );
BUFx3_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g403 ( .A(n_360), .Y(n_403) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx2_ASAP7_75t_L g401 ( .A(n_364), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_365), .B(n_386), .Y(n_364) );
NOR3xp33_ASAP7_75t_L g365 ( .A(n_366), .B(n_375), .C(n_380), .Y(n_365) );
OAI22xp5_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_368), .B1(n_371), .B2(n_372), .Y(n_366) );
OAI22xp5_ASAP7_75t_L g653 ( .A1(n_368), .A2(n_654), .B1(n_655), .B2(n_656), .Y(n_653) );
BUFx3_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
BUFx6f_ASAP7_75t_L g435 ( .A(n_369), .Y(n_435) );
INVx2_ASAP7_75t_L g481 ( .A(n_369), .Y(n_481) );
OAI221xp5_ASAP7_75t_L g699 ( .A1(n_369), .A2(n_439), .B1(n_700), .B2(n_701), .C(n_702), .Y(n_699) );
OAI22xp5_ASAP7_75t_L g478 ( .A1(n_372), .A2(n_479), .B1(n_480), .B2(n_482), .Y(n_478) );
OA211x2_ASAP7_75t_L g600 ( .A1(n_372), .A2(n_601), .B(n_602), .C(n_603), .Y(n_600) );
INVx1_ASAP7_75t_SL g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g656 ( .A(n_373), .Y(n_656) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
BUFx3_ASAP7_75t_L g439 ( .A(n_374), .Y(n_439) );
OAI21xp33_ASAP7_75t_SL g375 ( .A1(n_376), .A2(n_377), .B(n_378), .Y(n_375) );
INVx3_ASAP7_75t_L g473 ( .A(n_376), .Y(n_473) );
INVx4_ASAP7_75t_L g560 ( .A(n_376), .Y(n_560) );
INVx4_ASAP7_75t_L g588 ( .A(n_376), .Y(n_588) );
CKINVDCx16_ASAP7_75t_R g456 ( .A(n_383), .Y(n_456) );
OR2x6_ASAP7_75t_L g383 ( .A(n_384), .B(n_385), .Y(n_383) );
NOR2xp33_ASAP7_75t_L g386 ( .A(n_387), .B(n_393), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_388), .B(n_390), .Y(n_387) );
BUFx2_ASAP7_75t_L g466 ( .A(n_389), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_394), .B(n_398), .Y(n_393) );
INVx3_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx3_ASAP7_75t_L g694 ( .A(n_396), .Y(n_694) );
BUFx2_ASAP7_75t_L g427 ( .A(n_397), .Y(n_427) );
HB1xp67_ASAP7_75t_L g414 ( .A(n_399), .Y(n_414) );
OAI22xp5_ASAP7_75t_SL g405 ( .A1(n_406), .A2(n_407), .B1(n_497), .B2(n_498), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
AOI22xp5_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_459), .B1(n_495), .B2(n_496), .Y(n_407) );
INVx2_ASAP7_75t_L g495 ( .A(n_408), .Y(n_495) );
INVx1_ASAP7_75t_SL g458 ( .A(n_409), .Y(n_458) );
AND2x2_ASAP7_75t_SL g409 ( .A(n_410), .B(n_430), .Y(n_409) );
NOR2xp33_ASAP7_75t_L g410 ( .A(n_411), .B(n_418), .Y(n_410) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
OAI221xp5_ASAP7_75t_SL g418 ( .A1(n_419), .A2(n_421), .B1(n_422), .B2(n_425), .C(n_426), .Y(n_418) );
INVx3_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
OAI22xp5_ASAP7_75t_L g645 ( .A1(n_422), .A2(n_646), .B1(n_647), .B2(n_648), .Y(n_645) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g532 ( .A(n_423), .Y(n_532) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
BUFx4f_ASAP7_75t_SL g428 ( .A(n_429), .Y(n_428) );
BUFx2_ASAP7_75t_L g585 ( .A(n_429), .Y(n_585) );
BUFx2_ASAP7_75t_L g599 ( .A(n_429), .Y(n_599) );
NOR3xp33_ASAP7_75t_L g430 ( .A(n_431), .B(n_440), .C(n_449), .Y(n_430) );
OAI22xp5_ASAP7_75t_L g431 ( .A1(n_432), .A2(n_433), .B1(n_436), .B2(n_437), .Y(n_431) );
INVx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
OAI22xp5_ASAP7_75t_SL g621 ( .A1(n_437), .A2(n_622), .B1(n_623), .B2(n_624), .Y(n_621) );
INVx2_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
BUFx3_ASAP7_75t_L g506 ( .A(n_439), .Y(n_506) );
OAI221xp5_ASAP7_75t_L g483 ( .A1(n_441), .A2(n_484), .B1(n_485), .B2(n_486), .C(n_487), .Y(n_483) );
OAI22xp5_ASAP7_75t_L g514 ( .A1(n_441), .A2(n_515), .B1(n_516), .B2(n_517), .Y(n_514) );
INVx2_ASAP7_75t_SL g441 ( .A(n_442), .Y(n_441) );
INVx2_ASAP7_75t_SL g662 ( .A(n_442), .Y(n_662) );
BUFx6f_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
OAI22xp5_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_451), .B1(n_454), .B2(n_455), .Y(n_449) );
OAI22xp5_ASAP7_75t_L g490 ( .A1(n_451), .A2(n_455), .B1(n_491), .B2(n_492), .Y(n_490) );
INVx2_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx4_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
BUFx3_ASAP7_75t_L g632 ( .A(n_453), .Y(n_632) );
OAI22xp5_ASAP7_75t_L g660 ( .A1(n_453), .A2(n_661), .B1(n_662), .B2(n_663), .Y(n_660) );
INVx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx2_ASAP7_75t_L g496 ( .A(n_459), .Y(n_496) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g494 ( .A(n_461), .Y(n_494) );
AND2x2_ASAP7_75t_SL g461 ( .A(n_462), .B(n_477), .Y(n_461) );
NOR2xp33_ASAP7_75t_SL g462 ( .A(n_463), .B(n_470), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_464), .B(n_467), .Y(n_463) );
INVx1_ASAP7_75t_L g536 ( .A(n_468), .Y(n_536) );
BUFx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_471), .B(n_474), .Y(n_470) );
BUFx6f_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx2_ASAP7_75t_L g527 ( .A(n_476), .Y(n_527) );
NOR3xp33_ASAP7_75t_L g477 ( .A(n_478), .B(n_483), .C(n_490), .Y(n_477) );
INVx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx2_ASAP7_75t_L g622 ( .A(n_481), .Y(n_622) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
OAI22xp5_ASAP7_75t_SL g498 ( .A1(n_499), .A2(n_537), .B1(n_564), .B2(n_565), .Y(n_498) );
INVx1_ASAP7_75t_L g564 ( .A(n_499), .Y(n_564) );
XNOR2x1_ASAP7_75t_L g499 ( .A(n_500), .B(n_501), .Y(n_499) );
AND2x2_ASAP7_75t_L g501 ( .A(n_502), .B(n_521), .Y(n_501) );
INVx3_ASAP7_75t_L g543 ( .A(n_503), .Y(n_543) );
OAI211xp5_ASAP7_75t_L g504 ( .A1(n_505), .A2(n_506), .B(n_507), .C(n_510), .Y(n_504) );
BUFx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx1_ASAP7_75t_SL g512 ( .A(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx3_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
BUFx4f_ASAP7_75t_SL g612 ( .A(n_520), .Y(n_612) );
NOR3xp33_ASAP7_75t_L g521 ( .A(n_522), .B(n_528), .C(n_533), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_523), .B(n_525), .Y(n_522) );
INVx3_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
OAI22xp5_ASAP7_75t_L g528 ( .A1(n_529), .A2(n_530), .B1(n_531), .B2(n_532), .Y(n_528) );
INVx1_ASAP7_75t_L g565 ( .A(n_537), .Y(n_565) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx1_ASAP7_75t_L g563 ( .A(n_540), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_541), .B(n_553), .Y(n_540) );
NOR2xp67_ASAP7_75t_L g541 ( .A(n_542), .B(n_546), .Y(n_541) );
OAI21xp5_ASAP7_75t_SL g542 ( .A1(n_543), .A2(n_544), .B(n_545), .Y(n_542) );
OAI21xp33_ASAP7_75t_L g625 ( .A1(n_543), .A2(n_626), .B(n_627), .Y(n_625) );
OAI21xp5_ASAP7_75t_SL g703 ( .A1(n_543), .A2(n_704), .B(n_705), .Y(n_703) );
NAND3xp33_ASAP7_75t_L g546 ( .A(n_547), .B(n_549), .C(n_550), .Y(n_546) );
NOR2x1_ASAP7_75t_L g553 ( .A(n_554), .B(n_558), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_555), .B(n_556), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_559), .B(n_562), .Y(n_558) );
CKINVDCx16_ASAP7_75t_R g674 ( .A(n_566), .Y(n_674) );
AOI22xp5_ASAP7_75t_L g566 ( .A1(n_567), .A2(n_568), .B1(n_614), .B2(n_615), .Y(n_566) );
INVx2_ASAP7_75t_SL g567 ( .A(n_568), .Y(n_567) );
XNOR2x2_ASAP7_75t_L g568 ( .A(n_569), .B(n_593), .Y(n_568) );
XOR2x2_ASAP7_75t_L g569 ( .A(n_570), .B(n_592), .Y(n_569) );
NAND3x1_ASAP7_75t_L g570 ( .A(n_571), .B(n_581), .C(n_586), .Y(n_570) );
NOR2xp33_ASAP7_75t_L g571 ( .A(n_572), .B(n_576), .Y(n_571) );
OAI21xp5_ASAP7_75t_SL g572 ( .A1(n_573), .A2(n_574), .B(n_575), .Y(n_572) );
NAND3xp33_ASAP7_75t_L g576 ( .A(n_577), .B(n_579), .C(n_580), .Y(n_576) );
AND2x2_ASAP7_75t_L g581 ( .A(n_582), .B(n_584), .Y(n_581) );
AND2x2_ASAP7_75t_L g586 ( .A(n_587), .B(n_589), .Y(n_586) );
INVx1_ASAP7_75t_L g641 ( .A(n_590), .Y(n_641) );
XOR2x2_ASAP7_75t_L g593 ( .A(n_594), .B(n_613), .Y(n_593) );
NAND4xp75_ASAP7_75t_L g594 ( .A(n_595), .B(n_600), .C(n_605), .D(n_609), .Y(n_594) );
AND2x2_ASAP7_75t_L g595 ( .A(n_596), .B(n_598), .Y(n_595) );
CKINVDCx20_ASAP7_75t_R g630 ( .A(n_604), .Y(n_630) );
AND2x2_ASAP7_75t_L g605 ( .A(n_606), .B(n_608), .Y(n_605) );
INVx2_ASAP7_75t_L g646 ( .A(n_607), .Y(n_646) );
INVx4_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
OAI21xp5_ASAP7_75t_SL g657 ( .A1(n_611), .A2(n_658), .B(n_659), .Y(n_657) );
OAI21xp5_ASAP7_75t_L g723 ( .A1(n_611), .A2(n_724), .B(n_725), .Y(n_723) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
OAI22xp5_ASAP7_75t_SL g615 ( .A1(n_616), .A2(n_649), .B1(n_650), .B2(n_672), .Y(n_615) );
INVx2_ASAP7_75t_L g672 ( .A(n_616), .Y(n_672) );
INVx2_ASAP7_75t_SL g618 ( .A(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g619 ( .A(n_620), .B(n_633), .Y(n_619) );
NOR3xp33_ASAP7_75t_L g620 ( .A(n_621), .B(n_625), .C(n_628), .Y(n_620) );
OAI22xp33_ASAP7_75t_L g628 ( .A1(n_629), .A2(n_630), .B1(n_631), .B2(n_632), .Y(n_628) );
NOR3xp33_ASAP7_75t_L g633 ( .A(n_634), .B(n_639), .C(n_645), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_635), .B(n_637), .Y(n_634) );
OAI22xp5_ASAP7_75t_L g639 ( .A1(n_640), .A2(n_641), .B1(n_642), .B2(n_643), .Y(n_639) );
INVx1_ASAP7_75t_SL g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
XOR2x2_ASAP7_75t_L g650 ( .A(n_651), .B(n_671), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_652), .B(n_664), .Y(n_651) );
NOR3xp33_ASAP7_75t_L g652 ( .A(n_653), .B(n_657), .C(n_660), .Y(n_652) );
NOR2xp33_ASAP7_75t_L g664 ( .A(n_665), .B(n_668), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_666), .B(n_667), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_669), .B(n_670), .Y(n_668) );
INVx2_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
NOR2x1_ASAP7_75t_L g676 ( .A(n_677), .B(n_681), .Y(n_676) );
OR2x2_ASAP7_75t_SL g737 ( .A(n_677), .B(n_682), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_678), .B(n_680), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
HB1xp67_ASAP7_75t_L g706 ( .A(n_679), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_679), .B(n_709), .Y(n_712) );
CKINVDCx16_ASAP7_75t_R g709 ( .A(n_680), .Y(n_709) );
CKINVDCx20_ASAP7_75t_R g681 ( .A(n_682), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_683), .B(n_684), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_686), .B(n_687), .Y(n_685) );
OAI322xp33_ASAP7_75t_L g688 ( .A1(n_689), .A2(n_706), .A3(n_707), .B1(n_710), .B2(n_713), .C1(n_714), .C2(n_734), .Y(n_688) );
HB1xp67_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
NOR4xp75_ASAP7_75t_L g691 ( .A(n_692), .B(n_696), .C(n_699), .D(n_703), .Y(n_691) );
NAND2xp5_ASAP7_75t_SL g692 ( .A(n_693), .B(n_695), .Y(n_692) );
NAND2xp5_ASAP7_75t_SL g696 ( .A(n_697), .B(n_698), .Y(n_696) );
HB1xp67_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
CKINVDCx16_ASAP7_75t_R g710 ( .A(n_711), .Y(n_710) );
XOR2x2_ASAP7_75t_L g716 ( .A(n_713), .B(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx2_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
NAND3x1_ASAP7_75t_L g717 ( .A(n_718), .B(n_722), .C(n_730), .Y(n_717) );
AND2x2_ASAP7_75t_L g718 ( .A(n_719), .B(n_720), .Y(n_718) );
NOR2x1_ASAP7_75t_L g722 ( .A(n_723), .B(n_726), .Y(n_722) );
NAND3xp33_ASAP7_75t_L g726 ( .A(n_727), .B(n_728), .C(n_729), .Y(n_726) );
AND2x2_ASAP7_75t_L g730 ( .A(n_731), .B(n_733), .Y(n_730) );
HB1xp67_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
CKINVDCx20_ASAP7_75t_R g735 ( .A(n_736), .Y(n_735) );
CKINVDCx20_ASAP7_75t_R g736 ( .A(n_737), .Y(n_736) );
endmodule