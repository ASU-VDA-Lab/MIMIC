module fake_jpeg_6083_n_215 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_215);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_215;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_122;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx13_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_11),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_4),
.B(n_10),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_32),
.B(n_34),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_15),
.B(n_0),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_35),
.B(n_39),
.Y(n_54)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_37),
.B(n_40),
.Y(n_62)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

CKINVDCx6p67_ASAP7_75t_R g41 ( 
.A(n_28),
.Y(n_41)
);

BUFx6f_ASAP7_75t_SL g79 ( 
.A(n_41),
.Y(n_79)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_42),
.A2(n_48),
.B1(n_16),
.B2(n_30),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_43),
.Y(n_86)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_47),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_19),
.B(n_0),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_45),
.B(n_13),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_32),
.A2(n_26),
.B1(n_21),
.B2(n_29),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_50),
.A2(n_24),
.B1(n_2),
.B2(n_3),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_44),
.A2(n_26),
.B1(n_23),
.B2(n_29),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_52),
.A2(n_72),
.B1(n_17),
.B2(n_14),
.Y(n_104)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_56),
.B(n_59),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_43),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_57),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_58),
.Y(n_99)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_60),
.B(n_65),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_39),
.B(n_19),
.Y(n_64)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

BUFx16f_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_33),
.B(n_22),
.Y(n_66)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_41),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_67),
.B(n_70),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_48),
.A2(n_16),
.B1(n_30),
.B2(n_27),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_68),
.A2(n_78),
.B1(n_31),
.B2(n_25),
.Y(n_87)
);

BUFx4f_ASAP7_75t_SL g70 ( 
.A(n_42),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_40),
.B(n_16),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_71),
.B(n_83),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_47),
.A2(n_21),
.B1(n_23),
.B2(n_27),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_33),
.B(n_22),
.Y(n_73)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_73),
.Y(n_95)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_74),
.B(n_76),
.Y(n_97)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_35),
.Y(n_76)
);

BUFx16f_ASAP7_75t_L g77 ( 
.A(n_38),
.Y(n_77)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_77),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_49),
.A2(n_31),
.B1(n_30),
.B2(n_27),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_36),
.B(n_22),
.Y(n_80)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_46),
.B(n_14),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_82),
.Y(n_94)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_41),
.Y(n_83)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_41),
.Y(n_84)
);

NOR2x1_ASAP7_75t_L g105 ( 
.A(n_84),
.B(n_77),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_85),
.B(n_13),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_87),
.A2(n_107),
.B1(n_111),
.B2(n_53),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_62),
.B(n_25),
.C(n_31),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_90),
.B(n_70),
.Y(n_133)
);

AND2x6_ASAP7_75t_L g100 ( 
.A(n_65),
.B(n_20),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_100),
.B(n_101),
.Y(n_115)
);

AND2x6_ASAP7_75t_L g101 ( 
.A(n_65),
.B(n_24),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_72),
.B(n_24),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_102),
.B(n_5),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_103),
.B(n_104),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_105),
.B(n_84),
.Y(n_114)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_106),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_61),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_107)
);

A2O1A1Ixp33_ASAP7_75t_L g109 ( 
.A1(n_71),
.A2(n_1),
.B(n_5),
.C(n_6),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_109),
.B(n_110),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_62),
.B(n_1),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_56),
.A2(n_53),
.B1(n_60),
.B2(n_76),
.Y(n_111)
);

NOR3xp33_ASAP7_75t_L g155 ( 
.A(n_114),
.B(n_136),
.C(n_6),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_110),
.B(n_69),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_116),
.B(n_122),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_117),
.B(n_107),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_105),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_118),
.B(n_133),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_119),
.B(n_124),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_110),
.B(n_83),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_99),
.A2(n_70),
.B(n_77),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_123),
.A2(n_125),
.B(n_95),
.Y(n_148)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_97),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_101),
.A2(n_102),
.B(n_100),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_92),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_126),
.B(n_129),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_89),
.B(n_86),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_127),
.B(n_128),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_89),
.B(n_86),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_89),
.B(n_54),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_109),
.B(n_51),
.Y(n_130)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_130),
.Y(n_140)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_112),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_131),
.B(n_132),
.Y(n_142)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_88),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_96),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_134),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_91),
.B(n_90),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_135),
.Y(n_152)
);

OAI21xp33_ASAP7_75t_L g136 ( 
.A1(n_104),
.A2(n_59),
.B(n_7),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_94),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_137),
.B(n_108),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_127),
.A2(n_91),
.B(n_94),
.Y(n_143)
);

AOI221xp5_ASAP7_75t_L g170 ( 
.A1(n_143),
.A2(n_155),
.B1(n_121),
.B2(n_122),
.C(n_130),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_144),
.B(n_149),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_117),
.B(n_103),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_145),
.B(n_133),
.Y(n_162)
);

AO22x1_ASAP7_75t_L g146 ( 
.A1(n_136),
.A2(n_82),
.B1(n_75),
.B2(n_51),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_146),
.A2(n_128),
.B1(n_119),
.B2(n_129),
.Y(n_164)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_147),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_148),
.A2(n_123),
.B(n_114),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_125),
.B(n_95),
.C(n_93),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_125),
.A2(n_63),
.B1(n_93),
.B2(n_98),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_153),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_115),
.A2(n_63),
.B1(n_98),
.B2(n_55),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_154),
.B(n_118),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_137),
.B(n_112),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_156),
.B(n_157),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_115),
.B(n_79),
.C(n_75),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_147),
.B(n_120),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_160),
.B(n_163),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_161),
.A2(n_164),
.B1(n_146),
.B2(n_151),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_162),
.B(n_160),
.C(n_166),
.Y(n_175)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_156),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_140),
.B(n_116),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_165),
.B(n_168),
.Y(n_178)
);

FAx1_ASAP7_75t_SL g174 ( 
.A(n_167),
.B(n_158),
.CI(n_153),
.CON(n_174),
.SN(n_174)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_142),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_170),
.B(n_133),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_140),
.B(n_143),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_171),
.B(n_172),
.Y(n_182)
);

OAI32xp33_ASAP7_75t_L g172 ( 
.A1(n_151),
.A2(n_120),
.A3(n_148),
.B1(n_146),
.B2(n_138),
.Y(n_172)
);

AOI321xp33_ASAP7_75t_L g186 ( 
.A1(n_174),
.A2(n_179),
.A3(n_167),
.B1(n_166),
.B2(n_169),
.C(n_138),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_175),
.B(n_184),
.Y(n_187)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_177),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_168),
.B(n_131),
.Y(n_180)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_180),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_171),
.B(n_131),
.Y(n_181)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_181),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_163),
.B(n_132),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_183),
.B(n_185),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_162),
.B(n_157),
.C(n_149),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_169),
.Y(n_185)
);

AND2x2_ASAP7_75t_SL g195 ( 
.A(n_186),
.B(n_175),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_182),
.A2(n_173),
.B(n_159),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_188),
.A2(n_190),
.B(n_191),
.Y(n_196)
);

NOR3xp33_ASAP7_75t_SL g190 ( 
.A(n_174),
.B(n_172),
.C(n_173),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_176),
.A2(n_159),
.B(n_164),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_195),
.A2(n_133),
.B(n_186),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_187),
.B(n_184),
.C(n_145),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_197),
.A2(n_198),
.B(n_199),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_187),
.B(n_152),
.C(n_193),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_189),
.B(n_178),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_192),
.B(n_124),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_200),
.A2(n_165),
.B1(n_121),
.B2(n_185),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_201),
.B(n_141),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_196),
.A2(n_194),
.B(n_152),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_203),
.B(n_205),
.C(n_139),
.Y(n_206)
);

OAI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_196),
.A2(n_177),
.B1(n_190),
.B2(n_174),
.Y(n_204)
);

AOI322xp5_ASAP7_75t_L g209 ( 
.A1(n_204),
.A2(n_113),
.A3(n_123),
.B1(n_118),
.B2(n_150),
.C1(n_79),
.C2(n_9),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_206),
.B(n_209),
.C(n_113),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_207),
.B(n_118),
.Y(n_210)
);

OAI221xp5_ASAP7_75t_L g208 ( 
.A1(n_202),
.A2(n_135),
.B1(n_154),
.B2(n_144),
.C(n_150),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_208),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_210),
.A2(n_7),
.B(n_8),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_212),
.B(n_211),
.C(n_8),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_213),
.B(n_214),
.Y(n_215)
);


endmodule