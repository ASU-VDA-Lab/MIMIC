module real_jpeg_19444_n_17 (n_8, n_0, n_2, n_348, n_10, n_9, n_12, n_349, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_17);

input n_8;
input n_0;
input n_2;
input n_348;
input n_10;
input n_9;
input n_12;
input n_349;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx13_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_1),
.A2(n_24),
.B1(n_26),
.B2(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_1),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_1),
.A2(n_64),
.B1(n_71),
.B2(n_72),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g243 ( 
.A1(n_1),
.A2(n_54),
.B1(n_55),
.B2(n_64),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_1),
.A2(n_32),
.B1(n_33),
.B2(n_64),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_2),
.A2(n_54),
.B1(n_55),
.B2(n_95),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_2),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_2),
.A2(n_71),
.B1(n_72),
.B2(n_95),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_2),
.A2(n_32),
.B1(n_33),
.B2(n_95),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_2),
.A2(n_24),
.B1(n_26),
.B2(n_95),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_3),
.A2(n_54),
.B1(n_55),
.B2(n_107),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_3),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_3),
.A2(n_71),
.B1(n_72),
.B2(n_107),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_3),
.A2(n_32),
.B1(n_33),
.B2(n_107),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_3),
.A2(n_24),
.B1(n_26),
.B2(n_107),
.Y(n_223)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_5),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_5),
.B(n_116),
.Y(n_115)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_5),
.Y(n_125)
);

A2O1A1O1Ixp25_ASAP7_75t_L g91 ( 
.A1(n_6),
.A2(n_55),
.B(n_67),
.C(n_92),
.D(n_93),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_6),
.B(n_55),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_6),
.B(n_53),
.Y(n_103)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_6),
.Y(n_133)
);

OAI21xp33_ASAP7_75t_L g135 ( 
.A1(n_6),
.A2(n_113),
.B(n_115),
.Y(n_135)
);

A2O1A1O1Ixp25_ASAP7_75t_L g148 ( 
.A1(n_6),
.A2(n_32),
.B(n_48),
.C(n_149),
.D(n_150),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_6),
.B(n_32),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_6),
.B(n_36),
.Y(n_177)
);

AOI21xp33_ASAP7_75t_L g195 ( 
.A1(n_6),
.A2(n_33),
.B(n_196),
.Y(n_195)
);

OAI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_6),
.A2(n_24),
.B1(n_26),
.B2(n_133),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

BUFx12_ASAP7_75t_L g71 ( 
.A(n_8),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_9),
.A2(n_71),
.B1(n_72),
.B2(n_112),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_9),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_9),
.A2(n_54),
.B1(n_55),
.B2(n_112),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_9),
.A2(n_32),
.B1(n_33),
.B2(n_112),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_9),
.A2(n_24),
.B1(n_26),
.B2(n_112),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_10),
.A2(n_71),
.B1(n_72),
.B2(n_160),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_10),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_10),
.A2(n_54),
.B1(n_55),
.B2(n_160),
.Y(n_206)
);

OAI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_10),
.A2(n_32),
.B1(n_33),
.B2(n_160),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g296 ( 
.A1(n_10),
.A2(n_24),
.B1(n_26),
.B2(n_160),
.Y(n_296)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_12),
.A2(n_24),
.B1(n_26),
.B2(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_12),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_12),
.A2(n_62),
.B1(n_71),
.B2(n_72),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_12),
.A2(n_54),
.B1(n_55),
.B2(n_62),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_12),
.A2(n_32),
.B1(n_33),
.B2(n_62),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_13),
.A2(n_23),
.B1(n_24),
.B2(n_26),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_13),
.A2(n_23),
.B1(n_32),
.B2(n_33),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_13),
.A2(n_23),
.B1(n_71),
.B2(n_72),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_13),
.A2(n_23),
.B1(n_54),
.B2(n_55),
.Y(n_275)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_14),
.A2(n_29),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_15),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_16),
.A2(n_24),
.B1(n_26),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_16),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_16),
.A2(n_32),
.B1(n_33),
.B2(n_35),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_16),
.A2(n_35),
.B1(n_54),
.B2(n_55),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_16),
.A2(n_35),
.B1(n_71),
.B2(n_72),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_40),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_38),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_37),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_21),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_21),
.B(n_39),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_21),
.B(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_21),
.B(n_42),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_27),
.B1(n_34),
.B2(n_36),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_22),
.A2(n_27),
.B1(n_36),
.B2(n_77),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_24),
.Y(n_26)
);

A2O1A1Ixp33_ASAP7_75t_L g28 ( 
.A1(n_24),
.A2(n_29),
.B(n_30),
.C(n_31),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_29),
.Y(n_30)
);

A2O1A1Ixp33_ASAP7_75t_L g194 ( 
.A1(n_24),
.A2(n_29),
.B(n_133),
.C(n_195),
.Y(n_194)
);

BUFx2_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_SL g37 ( 
.A1(n_27),
.A2(n_34),
.B(n_36),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_27),
.A2(n_212),
.B(n_213),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_27),
.B(n_215),
.Y(n_224)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_28),
.A2(n_31),
.B1(n_61),
.B2(n_63),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_28),
.A2(n_31),
.B1(n_223),
.B2(n_252),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_28),
.A2(n_214),
.B(n_252),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_28),
.A2(n_31),
.B1(n_61),
.B2(n_296),
.Y(n_316)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_29),
.Y(n_196)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

OAI21xp33_ASAP7_75t_L g222 ( 
.A1(n_31),
.A2(n_223),
.B(n_224),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_31),
.A2(n_224),
.B(n_296),
.Y(n_295)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

O2A1O1Ixp33_ASAP7_75t_SL g48 ( 
.A1(n_33),
.A2(n_49),
.B(n_52),
.C(n_53),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_33),
.B(n_49),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_36),
.B(n_215),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_37),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_81),
.B(n_346),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_76),
.C(n_78),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_43),
.A2(n_44),
.B1(n_341),
.B2(n_343),
.Y(n_340)
);

CKINVDCx14_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_59),
.C(n_65),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_45),
.A2(n_46),
.B1(n_65),
.B2(n_321),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_47),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_47),
.A2(n_57),
.B1(n_171),
.B2(n_209),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_47),
.A2(n_209),
.B(n_227),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_47),
.A2(n_56),
.B1(n_57),
.B2(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_48),
.A2(n_53),
.B(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_48),
.B(n_173),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_48),
.A2(n_53),
.B1(n_249),
.B2(n_268),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_48),
.A2(n_53),
.B1(n_268),
.B2(n_287),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_49),
.A2(n_50),
.B1(n_54),
.B2(n_55),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_49),
.B(n_55),
.Y(n_157)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_52),
.A2(n_54),
.B1(n_156),
.B2(n_157),
.Y(n_155)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_53),
.Y(n_57)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_54),
.Y(n_55)
);

O2A1O1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_54),
.A2(n_68),
.B(n_69),
.C(n_70),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_68),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_57),
.B(n_151),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_57),
.A2(n_171),
.B(n_172),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_57),
.A2(n_172),
.B(n_248),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_58),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_59),
.A2(n_60),
.B1(n_329),
.B2(n_330),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_63),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_65),
.A2(n_319),
.B1(n_321),
.B2(n_322),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_65),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_SL g65 ( 
.A1(n_66),
.A2(n_74),
.B(n_75),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_66),
.A2(n_74),
.B1(n_106),
.B2(n_147),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_66),
.A2(n_147),
.B(n_184),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_66),
.A2(n_74),
.B1(n_206),
.B2(n_234),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_66),
.A2(n_74),
.B1(n_234),
.B2(n_243),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_66),
.A2(n_74),
.B1(n_243),
.B2(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_67),
.B(n_109),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_67),
.A2(n_70),
.B1(n_284),
.B2(n_285),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_68),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.Y(n_70)
);

CKINVDCx9p33_ASAP7_75t_R g73 ( 
.A(n_68),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_68),
.B(n_72),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_69),
.A2(n_71),
.B1(n_98),
.B2(n_99),
.Y(n_97)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_70),
.Y(n_74)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_71),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_71),
.B(n_114),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_72),
.B(n_137),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_74),
.B(n_94),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_74),
.A2(n_106),
.B(n_108),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_74),
.B(n_133),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_74),
.A2(n_108),
.B(n_206),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g285 ( 
.A(n_75),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_76),
.A2(n_78),
.B1(n_79),
.B2(n_342),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_76),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_339),
.B(n_345),
.Y(n_81)
);

OAI321xp33_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_312),
.A3(n_332),
.B1(n_337),
.B2(n_338),
.C(n_348),
.Y(n_82)
);

AOI321xp33_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_260),
.A3(n_300),
.B1(n_306),
.B2(n_311),
.C(n_349),
.Y(n_83)
);

NOR3xp33_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_217),
.C(n_256),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_188),
.B(n_216),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_87),
.A2(n_165),
.B(n_187),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_141),
.B(n_164),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_89),
.A2(n_117),
.B(n_140),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_100),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_90),
.B(n_100),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_91),
.B(n_96),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_91),
.A2(n_96),
.B1(n_97),
.B2(n_127),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_91),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_92),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_93),
.Y(n_184)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_94),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_110),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_103),
.B1(n_104),
.B2(n_105),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_102),
.B(n_105),
.C(n_110),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_111),
.A2(n_113),
.B(n_115),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_111),
.Y(n_123)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_113),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_113),
.A2(n_125),
.B1(n_159),
.B2(n_176),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_113),
.A2(n_114),
.B1(n_176),
.B2(n_199),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_113),
.A2(n_161),
.B1(n_199),
.B2(n_232),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_113),
.A2(n_161),
.B1(n_232),
.B2(n_241),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_113),
.A2(n_125),
.B(n_241),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_114),
.A2(n_121),
.B(n_131),
.Y(n_130)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_114),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_116),
.B(n_122),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_128),
.B(n_139),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_126),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_119),
.B(n_126),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_120),
.A2(n_122),
.B1(n_123),
.B2(n_124),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_125),
.B(n_133),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_129),
.A2(n_134),
.B(n_138),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_132),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_130),
.B(n_132),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_131),
.A2(n_159),
.B(n_161),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_135),
.B(n_136),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_143),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_142),
.B(n_143),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_144),
.A2(n_145),
.B1(n_154),
.B2(n_163),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_148),
.B1(n_152),
.B2(n_153),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_146),
.Y(n_153)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_148),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_148),
.B(n_153),
.C(n_163),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_149),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_150),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_151),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_154),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_158),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_155),
.B(n_158),
.Y(n_182)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_167),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_166),
.B(n_167),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_181),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_168),
.B(n_183),
.C(n_185),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_169),
.A2(n_170),
.B1(n_174),
.B2(n_180),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_169),
.B(n_177),
.C(n_178),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_174),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_177),
.B1(n_178),
.B2(n_179),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_175),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_177),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_182),
.A2(n_183),
.B1(n_185),
.B2(n_186),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_182),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_183),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_190),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_189),
.B(n_190),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_203),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_200),
.B1(n_201),
.B2(n_202),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_192),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_192),
.B(n_202),
.C(n_203),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_194),
.B1(n_197),
.B2(n_198),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_193),
.B(n_198),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_194),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_198),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_200),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_211),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_205),
.A2(n_207),
.B1(n_208),
.B2(n_210),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_205),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_207),
.B(n_210),
.C(n_211),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_208),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

AOI21xp33_ASAP7_75t_L g307 ( 
.A1(n_218),
.A2(n_308),
.B(n_309),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_236),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_219),
.B(n_236),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_230),
.C(n_235),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_220),
.B(n_259),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_229),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_225),
.B1(n_226),
.B2(n_228),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_222),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_225),
.B(n_228),
.C(n_229),
.Y(n_254)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_230),
.B(n_235),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_233),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_231),
.B(n_233),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_237),
.A2(n_238),
.B1(n_254),
.B2(n_255),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_244),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_239),
.B(n_244),
.C(n_255),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_242),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_240),
.B(n_242),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_245),
.B(n_250),
.C(n_253),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_247),
.A2(n_250),
.B1(n_251),
.B2(n_253),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_247),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_249),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_251),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_254),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_257),
.B(n_258),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_278),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_261),
.B(n_278),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_271),
.C(n_277),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_262),
.A2(n_263),
.B1(n_271),
.B2(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_265),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_264),
.B(n_267),
.C(n_269),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_266),
.A2(n_267),
.B1(n_269),
.B2(n_270),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_267),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_271),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_272),
.A2(n_273),
.B1(n_274),
.B2(n_276),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_272),
.A2(n_273),
.B1(n_294),
.B2(n_295),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_272),
.A2(n_291),
.B(n_295),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_273),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_273),
.B(n_274),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_274),
.Y(n_276)
);

CKINVDCx14_ASAP7_75t_R g284 ( 
.A(n_275),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_277),
.B(n_304),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_279),
.A2(n_280),
.B1(n_298),
.B2(n_299),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_282),
.B1(n_289),
.B2(n_290),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_281),
.B(n_290),
.C(n_299),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_282),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_283),
.A2(n_286),
.B(n_288),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_283),
.B(n_286),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_287),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_288),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_288),
.A2(n_314),
.B1(n_323),
.B2(n_336),
.Y(n_335)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_290),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_291),
.A2(n_292),
.B1(n_293),
.B2(n_297),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_293),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_295),
.Y(n_294)
);

CKINVDCx14_ASAP7_75t_R g299 ( 
.A(n_298),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_301),
.A2(n_307),
.B(n_310),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_303),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_302),
.B(n_303),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_325),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_313),
.B(n_325),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_323),
.C(n_324),
.Y(n_313)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_314),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_315),
.A2(n_316),
.B1(n_317),
.B2(n_318),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_315),
.A2(n_316),
.B1(n_327),
.B2(n_328),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_316),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_316),
.B(n_321),
.C(n_322),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_316),
.B(n_327),
.C(n_331),
.Y(n_344)
);

CKINVDCx16_ASAP7_75t_R g317 ( 
.A(n_318),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_319),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_324),
.B(n_335),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_331),
.Y(n_325)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_334),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_333),
.B(n_334),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_344),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_340),
.B(n_344),
.Y(n_345)
);

CKINVDCx14_ASAP7_75t_R g343 ( 
.A(n_341),
.Y(n_343)
);


endmodule