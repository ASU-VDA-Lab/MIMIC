module fake_jpeg_13399_n_601 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_601);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_601;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_15),
.B(n_6),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_5),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

BUFx8_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_2),
.B(n_7),
.Y(n_49)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_10),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

BUFx24_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_5),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_11),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_11),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_57),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_58),
.Y(n_123)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_59),
.Y(n_188)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_60),
.Y(n_144)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

INVx13_ASAP7_75t_L g130 ( 
.A(n_61),
.Y(n_130)
);

BUFx4f_ASAP7_75t_SL g62 ( 
.A(n_24),
.Y(n_62)
);

INVx13_ASAP7_75t_L g152 ( 
.A(n_62),
.Y(n_152)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_63),
.Y(n_153)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_64),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_40),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_65),
.B(n_66),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_40),
.Y(n_66)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_67),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_18),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_68),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_18),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_69),
.Y(n_141)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_70),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_49),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_71),
.B(n_75),
.Y(n_134)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_28),
.Y(n_72)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_72),
.Y(n_125)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_20),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_73),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_49),
.B(n_15),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_74),
.B(n_15),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_17),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_29),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_76),
.Y(n_159)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_77),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_24),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g135 ( 
.A(n_78),
.Y(n_135)
);

BUFx12_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g155 ( 
.A(n_79),
.Y(n_155)
);

BUFx8_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g167 ( 
.A(n_80),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_29),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_81),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_17),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_82),
.B(n_87),
.Y(n_142)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_30),
.Y(n_83)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_83),
.Y(n_189)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_38),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_84),
.B(n_97),
.Y(n_129)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_20),
.Y(n_85)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_85),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_29),
.Y(n_86)
);

INVx6_ASAP7_75t_L g165 ( 
.A(n_86),
.Y(n_165)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_41),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_17),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_88),
.B(n_100),
.Y(n_151)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_34),
.Y(n_89)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_89),
.Y(n_137)
);

INVx6_ASAP7_75t_SL g90 ( 
.A(n_53),
.Y(n_90)
);

CKINVDCx12_ASAP7_75t_R g148 ( 
.A(n_90),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

INVx6_ASAP7_75t_L g182 ( 
.A(n_91),
.Y(n_182)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_92),
.Y(n_187)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_93),
.Y(n_138)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_52),
.Y(n_94)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_94),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

INVx6_ASAP7_75t_L g192 ( 
.A(n_95),
.Y(n_192)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_48),
.Y(n_96)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_96),
.Y(n_145)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_38),
.Y(n_97)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_28),
.Y(n_98)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_98),
.Y(n_147)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_28),
.Y(n_99)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_99),
.Y(n_170)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_43),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_47),
.Y(n_101)
);

INVx8_ASAP7_75t_L g132 ( 
.A(n_101),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_51),
.Y(n_102)
);

INVx8_ASAP7_75t_L g157 ( 
.A(n_102),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_51),
.Y(n_103)
);

INVx8_ASAP7_75t_L g164 ( 
.A(n_103),
.Y(n_164)
);

BUFx12f_ASAP7_75t_L g104 ( 
.A(n_34),
.Y(n_104)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_104),
.Y(n_162)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_43),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_105),
.B(n_106),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_42),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_16),
.Y(n_107)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_107),
.Y(n_183)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_39),
.Y(n_108)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_108),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_42),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_109),
.B(n_110),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_42),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_51),
.Y(n_111)
);

INVx8_ASAP7_75t_L g172 ( 
.A(n_111),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_16),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_112),
.B(n_115),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_27),
.Y(n_113)
);

INVx8_ASAP7_75t_L g175 ( 
.A(n_113),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_27),
.Y(n_114)
);

INVx8_ASAP7_75t_L g178 ( 
.A(n_114),
.Y(n_178)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_19),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_32),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_116),
.B(n_52),
.Y(n_177)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_52),
.Y(n_117)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_117),
.Y(n_199)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_27),
.Y(n_118)
);

INVx3_ASAP7_75t_SL g126 ( 
.A(n_118),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_52),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g179 ( 
.A(n_119),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_36),
.Y(n_120)
);

INVx8_ASAP7_75t_L g194 ( 
.A(n_120),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_36),
.Y(n_121)
);

INVx8_ASAP7_75t_L g196 ( 
.A(n_121),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_94),
.B(n_56),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_122),
.B(n_150),
.Y(n_202)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_92),
.Y(n_127)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_127),
.Y(n_201)
);

OR2x2_ASAP7_75t_L g143 ( 
.A(n_117),
.B(n_32),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_143),
.B(n_174),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_146),
.B(n_193),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_61),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_149),
.B(n_168),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_72),
.B(n_56),
.Y(n_150)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_92),
.Y(n_160)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_160),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_67),
.A2(n_31),
.B1(n_37),
.B2(n_36),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_163),
.A2(n_197),
.B1(n_13),
.B2(n_11),
.Y(n_266)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_104),
.Y(n_166)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_166),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_61),
.Y(n_168)
);

BUFx10_ASAP7_75t_L g169 ( 
.A(n_80),
.Y(n_169)
);

CKINVDCx14_ASAP7_75t_R g226 ( 
.A(n_169),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_99),
.B(n_26),
.C(n_22),
.Y(n_174)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_119),
.Y(n_176)
);

INVx4_ASAP7_75t_L g241 ( 
.A(n_176),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_177),
.B(n_50),
.Y(n_254)
);

INVx5_ASAP7_75t_L g180 ( 
.A(n_104),
.Y(n_180)
);

INVx4_ASAP7_75t_L g261 ( 
.A(n_180),
.Y(n_261)
);

INVx11_ASAP7_75t_L g181 ( 
.A(n_80),
.Y(n_181)
);

INVx11_ASAP7_75t_L g203 ( 
.A(n_181),
.Y(n_203)
);

INVxp67_ASAP7_75t_SL g184 ( 
.A(n_79),
.Y(n_184)
);

INVx5_ASAP7_75t_SL g234 ( 
.A(n_184),
.Y(n_234)
);

INVx3_ASAP7_75t_SL g185 ( 
.A(n_89),
.Y(n_185)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_185),
.Y(n_207)
);

BUFx16f_ASAP7_75t_L g186 ( 
.A(n_79),
.Y(n_186)
);

INVx13_ASAP7_75t_L g246 ( 
.A(n_186),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_73),
.A2(n_31),
.B1(n_44),
.B2(n_37),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_190),
.A2(n_54),
.B1(n_45),
.B2(n_35),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_62),
.B(n_23),
.Y(n_193)
);

OAI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_113),
.A2(n_44),
.B1(n_37),
.B2(n_39),
.Y(n_197)
);

BUFx10_ASAP7_75t_L g198 ( 
.A(n_78),
.Y(n_198)
);

INVx4_ASAP7_75t_SL g267 ( 
.A(n_198),
.Y(n_267)
);

INVx8_ASAP7_75t_L g200 ( 
.A(n_58),
.Y(n_200)
);

INVx5_ASAP7_75t_L g210 ( 
.A(n_200),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_204),
.A2(n_244),
.B1(n_248),
.B2(n_255),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_131),
.B(n_55),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_206),
.B(n_208),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_134),
.B(n_55),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_123),
.Y(n_209)
);

INVx8_ASAP7_75t_L g274 ( 
.A(n_209),
.Y(n_274)
);

A2O1A1Ixp33_ASAP7_75t_L g211 ( 
.A1(n_143),
.A2(n_19),
.B(n_26),
.C(n_22),
.Y(n_211)
);

NOR2x1_ASAP7_75t_L g285 ( 
.A(n_211),
.B(n_155),
.Y(n_285)
);

OAI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_197),
.A2(n_86),
.B1(n_81),
.B2(n_76),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_212),
.A2(n_178),
.B1(n_179),
.B2(n_7),
.Y(n_314)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_125),
.Y(n_213)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_213),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_185),
.A2(n_50),
.B1(n_39),
.B2(n_108),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_214),
.A2(n_253),
.B1(n_258),
.B2(n_265),
.Y(n_273)
);

INVx5_ASAP7_75t_L g215 ( 
.A(n_167),
.Y(n_215)
);

BUFx2_ASAP7_75t_L g327 ( 
.A(n_215),
.Y(n_327)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_167),
.Y(n_216)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_216),
.Y(n_289)
);

INVx8_ASAP7_75t_L g218 ( 
.A(n_169),
.Y(n_218)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_218),
.Y(n_294)
);

BUFx12f_ASAP7_75t_L g219 ( 
.A(n_187),
.Y(n_219)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_219),
.Y(n_283)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_167),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g291 ( 
.A(n_220),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_169),
.A2(n_45),
.B(n_33),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_221),
.A2(n_228),
.B(n_162),
.Y(n_279)
);

INVx11_ASAP7_75t_L g222 ( 
.A(n_198),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g328 ( 
.A(n_222),
.Y(n_328)
);

CKINVDCx12_ASAP7_75t_R g223 ( 
.A(n_148),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_223),
.B(n_227),
.Y(n_323)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_133),
.Y(n_224)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_224),
.Y(n_286)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_186),
.Y(n_225)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_225),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_161),
.Y(n_227)
);

NAND2xp33_ASAP7_75t_SL g228 ( 
.A(n_198),
.B(n_187),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_129),
.B(n_52),
.Y(n_229)
);

XNOR2x1_ASAP7_75t_L g317 ( 
.A(n_229),
.B(n_236),
.Y(n_317)
);

AOI21xp33_ASAP7_75t_L g231 ( 
.A1(n_173),
.A2(n_23),
.B(n_54),
.Y(n_231)
);

OR2x2_ASAP7_75t_L g290 ( 
.A(n_231),
.B(n_235),
.Y(n_290)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_188),
.Y(n_232)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_232),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_158),
.B(n_21),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_129),
.B(n_154),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_123),
.Y(n_237)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_237),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_189),
.B(n_0),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_238),
.B(n_239),
.C(n_264),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_144),
.B(n_153),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_191),
.Y(n_240)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_240),
.Y(n_322)
);

INVx5_ASAP7_75t_L g242 ( 
.A(n_135),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g304 ( 
.A(n_242),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_139),
.Y(n_243)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_243),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_142),
.A2(n_118),
.B1(n_85),
.B2(n_121),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_155),
.Y(n_245)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_245),
.Y(n_298)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_140),
.Y(n_247)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_247),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_151),
.A2(n_120),
.B1(n_114),
.B2(n_111),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_183),
.Y(n_249)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_249),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_139),
.Y(n_250)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_250),
.Y(n_315)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_199),
.Y(n_252)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_252),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_184),
.A2(n_50),
.B1(n_31),
.B2(n_44),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_254),
.B(n_260),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_136),
.A2(n_103),
.B1(n_102),
.B2(n_101),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_136),
.A2(n_91),
.B1(n_69),
.B2(n_68),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_256),
.A2(n_270),
.B1(n_196),
.B2(n_194),
.Y(n_281)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_176),
.Y(n_257)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_257),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_141),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_L g259 ( 
.A1(n_132),
.A2(n_95),
.B1(n_35),
.B2(n_33),
.Y(n_259)
);

OAI22xp33_ASAP7_75t_L g277 ( 
.A1(n_259),
.A2(n_165),
.B1(n_182),
.B2(n_192),
.Y(n_277)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_179),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_124),
.B(n_21),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_262),
.B(n_155),
.Y(n_275)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_170),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_263),
.B(n_269),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_138),
.B(n_0),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_145),
.A2(n_137),
.B1(n_126),
.B2(n_147),
.Y(n_265)
);

OA22x2_ASAP7_75t_L g287 ( 
.A1(n_266),
.A2(n_171),
.B1(n_159),
.B2(n_194),
.Y(n_287)
);

INVx6_ASAP7_75t_L g268 ( 
.A(n_141),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_268),
.A2(n_200),
.B1(n_157),
.B2(n_132),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_195),
.B(n_13),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_126),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_270)
);

HAxp5_ASAP7_75t_SL g271 ( 
.A(n_130),
.B(n_13),
.CON(n_271),
.SN(n_271)
);

OR2x2_ASAP7_75t_L g307 ( 
.A(n_271),
.B(n_130),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g353 ( 
.A(n_275),
.B(n_302),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_277),
.A2(n_301),
.B1(n_325),
.B2(n_326),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_217),
.B(n_192),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_278),
.B(n_282),
.Y(n_332)
);

CKINVDCx16_ASAP7_75t_R g330 ( 
.A(n_279),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_281),
.B(n_287),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_238),
.B(n_165),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_238),
.B(n_182),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_284),
.B(n_302),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_285),
.B(n_271),
.Y(n_329)
);

OAI22x1_ASAP7_75t_L g352 ( 
.A1(n_292),
.A2(n_293),
.B1(n_218),
.B2(n_203),
.Y(n_352)
);

AOI22xp33_ASAP7_75t_SL g293 ( 
.A1(n_234),
.A2(n_135),
.B1(n_157),
.B2(n_164),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_236),
.B(n_135),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_299),
.B(n_307),
.Y(n_337)
);

AOI22xp33_ASAP7_75t_L g300 ( 
.A1(n_266),
.A2(n_172),
.B1(n_164),
.B2(n_175),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_300),
.A2(n_306),
.B1(n_308),
.B2(n_320),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_202),
.A2(n_128),
.B1(n_156),
.B2(n_171),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_211),
.B(n_172),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_236),
.A2(n_128),
.B1(n_156),
.B2(n_196),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_229),
.A2(n_264),
.B1(n_270),
.B2(n_239),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_264),
.B(n_175),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_309),
.B(n_311),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_228),
.A2(n_152),
.B(n_179),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g350 ( 
.A(n_310),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_230),
.B(n_178),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_229),
.B(n_152),
.C(n_159),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_313),
.B(n_267),
.Y(n_367)
);

OAI22xp33_ASAP7_75t_SL g365 ( 
.A1(n_314),
.A2(n_321),
.B1(n_203),
.B2(n_220),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_239),
.A2(n_13),
.B1(n_8),
.B2(n_7),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_213),
.A2(n_8),
.B1(n_1),
.B2(n_3),
.Y(n_321)
);

OAI22xp33_ASAP7_75t_SL g325 ( 
.A1(n_221),
.A2(n_8),
.B1(n_1),
.B2(n_4),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_268),
.A2(n_0),
.B1(n_4),
.B2(n_5),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g374 ( 
.A1(n_329),
.A2(n_366),
.B(n_367),
.Y(n_374)
);

AND2x6_ASAP7_75t_L g331 ( 
.A(n_278),
.B(n_234),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_331),
.B(n_336),
.Y(n_385)
);

BUFx2_ASAP7_75t_L g333 ( 
.A(n_274),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g386 ( 
.A(n_333),
.Y(n_386)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_286),
.Y(n_334)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_334),
.Y(n_372)
);

AND2x6_ASAP7_75t_L g336 ( 
.A(n_290),
.B(n_251),
.Y(n_336)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_286),
.Y(n_338)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_338),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_323),
.B(n_201),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g393 ( 
.A(n_339),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_311),
.B(n_233),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_340),
.Y(n_408)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_322),
.Y(n_342)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_342),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_303),
.B(n_226),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_344),
.B(n_347),
.Y(n_383)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_322),
.Y(n_345)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_345),
.Y(n_392)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_324),
.Y(n_346)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_346),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_275),
.B(n_225),
.Y(n_347)
);

INVx5_ASAP7_75t_L g348 ( 
.A(n_274),
.Y(n_348)
);

HB1xp67_ASAP7_75t_L g406 ( 
.A(n_348),
.Y(n_406)
);

CKINVDCx14_ASAP7_75t_R g349 ( 
.A(n_288),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_349),
.B(n_353),
.Y(n_399)
);

AOI22xp33_ASAP7_75t_SL g382 ( 
.A1(n_352),
.A2(n_357),
.B1(n_361),
.B2(n_215),
.Y(n_382)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_280),
.Y(n_354)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_354),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_319),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_355),
.B(n_356),
.Y(n_407)
);

BUFx3_ASAP7_75t_L g356 ( 
.A(n_327),
.Y(n_356)
);

AOI22xp33_ASAP7_75t_L g357 ( 
.A1(n_287),
.A2(n_207),
.B1(n_257),
.B2(n_243),
.Y(n_357)
);

INVx13_ASAP7_75t_L g359 ( 
.A(n_327),
.Y(n_359)
);

CKINVDCx16_ASAP7_75t_R g397 ( 
.A(n_359),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_282),
.B(n_241),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_360),
.B(n_364),
.Y(n_391)
);

AOI22xp33_ASAP7_75t_L g361 ( 
.A1(n_287),
.A2(n_207),
.B1(n_237),
.B2(n_209),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_280),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_362),
.B(n_363),
.Y(n_398)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_305),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_316),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_365),
.A2(n_299),
.B1(n_288),
.B2(n_297),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_296),
.B(n_241),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g368 ( 
.A(n_299),
.B(n_310),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_SL g384 ( 
.A1(n_368),
.A2(n_370),
.B(n_371),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_272),
.B(n_261),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_369),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_290),
.B(n_261),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_284),
.B(n_210),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_330),
.A2(n_341),
.B1(n_343),
.B2(n_350),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_373),
.A2(n_396),
.B1(n_402),
.B2(n_371),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_L g376 ( 
.A1(n_368),
.A2(n_279),
.B(n_307),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_376),
.A2(n_379),
.B(n_381),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_L g379 ( 
.A1(n_368),
.A2(n_285),
.B(n_273),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_380),
.B(n_404),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_330),
.A2(n_288),
.B(n_308),
.Y(n_381)
);

CKINVDCx16_ASAP7_75t_R g435 ( 
.A(n_382),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_335),
.A2(n_287),
.B1(n_301),
.B2(n_277),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_387),
.A2(n_388),
.B1(n_395),
.B2(n_400),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_335),
.A2(n_297),
.B1(n_309),
.B2(n_296),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g389 ( 
.A1(n_350),
.A2(n_313),
.B(n_314),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_L g433 ( 
.A1(n_389),
.A2(n_403),
.B(n_222),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_366),
.B(n_332),
.C(n_317),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_390),
.B(n_367),
.C(n_337),
.Y(n_422)
);

AOI22xp33_ASAP7_75t_SL g395 ( 
.A1(n_358),
.A2(n_294),
.B1(n_289),
.B2(n_291),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_341),
.A2(n_276),
.B1(n_281),
.B2(n_306),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_335),
.A2(n_297),
.B1(n_276),
.B2(n_326),
.Y(n_400)
);

AOI22xp33_ASAP7_75t_SL g401 ( 
.A1(n_358),
.A2(n_352),
.B1(n_333),
.B2(n_294),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_L g436 ( 
.A1(n_401),
.A2(n_328),
.B1(n_348),
.B2(n_333),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_L g402 ( 
.A1(n_343),
.A2(n_321),
.B1(n_317),
.B2(n_320),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_L g403 ( 
.A1(n_329),
.A2(n_289),
.B(n_283),
.Y(n_403)
);

OAI32xp33_ASAP7_75t_L g404 ( 
.A1(n_353),
.A2(n_312),
.A3(n_295),
.B1(n_315),
.B2(n_319),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_378),
.B(n_332),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_SL g464 ( 
.A(n_410),
.B(n_419),
.Y(n_464)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_398),
.Y(n_412)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_412),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_391),
.B(n_351),
.Y(n_413)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_413),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_391),
.B(n_351),
.Y(n_414)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_414),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_398),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_415),
.B(n_425),
.Y(n_470)
);

MAJx2_ASAP7_75t_L g416 ( 
.A(n_390),
.B(n_337),
.C(n_367),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_416),
.B(n_418),
.C(n_422),
.Y(n_459)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_394),
.Y(n_417)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_417),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_390),
.B(n_337),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_378),
.B(n_318),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_394),
.Y(n_420)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_420),
.Y(n_460)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_405),
.Y(n_421)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_421),
.Y(n_463)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_405),
.Y(n_423)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_423),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_406),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_426),
.A2(n_380),
.B1(n_387),
.B2(n_389),
.Y(n_455)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_372),
.Y(n_427)
);

INVx1_ASAP7_75t_SL g457 ( 
.A(n_427),
.Y(n_457)
);

XOR2x1_ASAP7_75t_L g428 ( 
.A(n_388),
.B(n_331),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_SL g458 ( 
.A(n_428),
.B(n_383),
.C(n_379),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_406),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_429),
.B(n_432),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_374),
.B(n_360),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_430),
.B(n_434),
.C(n_438),
.Y(n_471)
);

INVx4_ASAP7_75t_L g431 ( 
.A(n_397),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_431),
.B(n_441),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_408),
.B(n_364),
.Y(n_432)
);

INVxp67_ASAP7_75t_L g467 ( 
.A(n_433),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_374),
.B(n_346),
.C(n_363),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_436),
.A2(n_437),
.B1(n_396),
.B2(n_403),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_L g437 ( 
.A1(n_400),
.A2(n_336),
.B1(n_355),
.B2(n_258),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_381),
.B(n_304),
.C(n_298),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_376),
.B(n_362),
.C(n_354),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_439),
.B(n_376),
.Y(n_450)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_372),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_440),
.B(n_442),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_385),
.B(n_318),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_407),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_434),
.B(n_385),
.Y(n_445)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_445),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_432),
.B(n_383),
.Y(n_446)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_446),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_415),
.B(n_399),
.Y(n_447)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_447),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_L g448 ( 
.A1(n_426),
.A2(n_401),
.B1(n_395),
.B2(n_387),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_448),
.A2(n_455),
.B1(n_473),
.B2(n_436),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_SL g495 ( 
.A(n_450),
.B(n_375),
.Y(n_495)
);

OAI31xp33_ASAP7_75t_SL g454 ( 
.A1(n_424),
.A2(n_373),
.A3(n_399),
.B(n_379),
.Y(n_454)
);

AOI21xp5_ASAP7_75t_SL g480 ( 
.A1(n_454),
.A2(n_438),
.B(n_409),
.Y(n_480)
);

CKINVDCx16_ASAP7_75t_R g456 ( 
.A(n_411),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_456),
.B(n_411),
.Y(n_475)
);

AOI21xp5_ASAP7_75t_L g490 ( 
.A1(n_458),
.A2(n_461),
.B(n_454),
.Y(n_490)
);

AOI21xp5_ASAP7_75t_L g461 ( 
.A1(n_424),
.A2(n_403),
.B(n_384),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_418),
.B(n_384),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_462),
.B(n_422),
.C(n_416),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_L g478 ( 
.A1(n_466),
.A2(n_435),
.B1(n_433),
.B2(n_412),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_413),
.B(n_414),
.Y(n_469)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_469),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_442),
.B(n_393),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_472),
.B(n_430),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_L g473 ( 
.A1(n_435),
.A2(n_382),
.B1(n_402),
.B2(n_404),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g507 ( 
.A(n_474),
.B(n_495),
.Y(n_507)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_475),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_459),
.B(n_439),
.C(n_416),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_476),
.B(n_485),
.C(n_462),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_471),
.B(n_428),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_477),
.B(n_482),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g524 ( 
.A1(n_478),
.A2(n_460),
.B1(n_453),
.B2(n_345),
.Y(n_524)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_479),
.Y(n_503)
);

OAI21xp5_ASAP7_75t_SL g520 ( 
.A1(n_480),
.A2(n_490),
.B(n_500),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_447),
.B(n_425),
.Y(n_481)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_481),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_471),
.B(n_409),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_464),
.B(n_429),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_483),
.B(n_499),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_459),
.B(n_437),
.C(n_440),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_L g486 ( 
.A1(n_466),
.A2(n_427),
.B1(n_423),
.B2(n_421),
.Y(n_486)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_486),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_465),
.B(n_420),
.Y(n_487)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_487),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_L g505 ( 
.A1(n_488),
.A2(n_491),
.B1(n_493),
.B2(n_494),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_448),
.A2(n_455),
.B1(n_473),
.B2(n_456),
.Y(n_491)
);

OAI21xp5_ASAP7_75t_L g492 ( 
.A1(n_467),
.A2(n_417),
.B(n_407),
.Y(n_492)
);

OAI21xp5_ASAP7_75t_L g514 ( 
.A1(n_492),
.A2(n_452),
.B(n_470),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_467),
.A2(n_443),
.B1(n_452),
.B2(n_465),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_443),
.A2(n_431),
.B1(n_392),
.B2(n_377),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_469),
.B(n_375),
.Y(n_496)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_496),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_464),
.B(n_356),
.Y(n_499)
);

MAJx2_ASAP7_75t_R g500 ( 
.A(n_458),
.B(n_386),
.C(n_397),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_449),
.A2(n_392),
.B1(n_377),
.B2(n_355),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_L g506 ( 
.A1(n_501),
.A2(n_457),
.B1(n_468),
.B2(n_463),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_506),
.A2(n_492),
.B1(n_489),
.B2(n_498),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_481),
.B(n_470),
.Y(n_511)
);

INVxp67_ASAP7_75t_L g530 ( 
.A(n_511),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_514),
.B(n_517),
.Y(n_536)
);

XNOR2xp5_ASAP7_75t_L g537 ( 
.A(n_515),
.B(n_523),
.Y(n_537)
);

XOR2xp5_ASAP7_75t_L g516 ( 
.A(n_482),
.B(n_450),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g526 ( 
.A(n_516),
.B(n_518),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_476),
.B(n_461),
.C(n_449),
.Y(n_517)
);

XOR2xp5_ASAP7_75t_L g518 ( 
.A(n_474),
.B(n_444),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_485),
.B(n_451),
.C(n_457),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_519),
.B(n_521),
.Y(n_543)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_487),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_477),
.B(n_451),
.C(n_463),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_522),
.B(n_493),
.C(n_484),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_L g523 ( 
.A(n_495),
.B(n_468),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_SL g541 ( 
.A1(n_524),
.A2(n_216),
.B1(n_242),
.B2(n_359),
.Y(n_541)
);

AOI21x1_ASAP7_75t_L g525 ( 
.A1(n_520),
.A2(n_490),
.B(n_500),
.Y(n_525)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_525),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_527),
.B(n_533),
.Y(n_546)
);

XOR2xp5_ASAP7_75t_L g558 ( 
.A(n_528),
.B(n_507),
.Y(n_558)
);

AOI22xp5_ASAP7_75t_L g529 ( 
.A1(n_505),
.A2(n_475),
.B1(n_489),
.B2(n_496),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_529),
.B(n_535),
.Y(n_547)
);

INVxp33_ASAP7_75t_L g531 ( 
.A(n_512),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_531),
.B(n_540),
.Y(n_553)
);

AO221x1_ASAP7_75t_L g532 ( 
.A1(n_503),
.A2(n_497),
.B1(n_460),
.B2(n_453),
.C(n_480),
.Y(n_532)
);

AOI21xp5_ASAP7_75t_L g552 ( 
.A1(n_532),
.A2(n_534),
.B(n_513),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_519),
.B(n_494),
.Y(n_533)
);

OAI21xp5_ASAP7_75t_SL g534 ( 
.A1(n_517),
.A2(n_491),
.B(n_488),
.Y(n_534)
);

AOI22xp5_ASAP7_75t_L g535 ( 
.A1(n_509),
.A2(n_501),
.B1(n_334),
.B2(n_342),
.Y(n_535)
);

AOI22xp5_ASAP7_75t_L g538 ( 
.A1(n_502),
.A2(n_338),
.B1(n_250),
.B2(n_210),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_538),
.B(n_539),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_522),
.B(n_283),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_508),
.Y(n_540)
);

AOI22xp5_ASAP7_75t_L g549 ( 
.A1(n_541),
.A2(n_510),
.B1(n_513),
.B2(n_511),
.Y(n_549)
);

A2O1A1Ixp33_ASAP7_75t_SL g542 ( 
.A1(n_520),
.A2(n_359),
.B(n_267),
.C(n_219),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_542),
.B(n_523),
.C(n_260),
.Y(n_556)
);

XNOR2xp5_ASAP7_75t_L g544 ( 
.A(n_537),
.B(n_518),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_544),
.B(n_554),
.Y(n_562)
);

OAI21xp5_ASAP7_75t_L g545 ( 
.A1(n_530),
.A2(n_514),
.B(n_502),
.Y(n_545)
);

OAI21xp5_ASAP7_75t_L g561 ( 
.A1(n_545),
.A2(n_556),
.B(n_547),
.Y(n_561)
);

XOR2x2_ASAP7_75t_L g548 ( 
.A(n_536),
.B(n_511),
.Y(n_548)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_548),
.Y(n_564)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_549),
.Y(n_568)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_552),
.Y(n_571)
);

XNOR2xp5_ASAP7_75t_L g554 ( 
.A(n_537),
.B(n_504),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_531),
.B(n_524),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_555),
.B(n_557),
.Y(n_565)
);

XOR2xp5_ASAP7_75t_L g569 ( 
.A(n_556),
.B(n_558),
.Y(n_569)
);

AOI22xp5_ASAP7_75t_L g557 ( 
.A1(n_530),
.A2(n_516),
.B1(n_507),
.B2(n_515),
.Y(n_557)
);

XOR2xp5_ASAP7_75t_L g559 ( 
.A(n_543),
.B(n_504),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_559),
.B(n_541),
.Y(n_570)
);

HB1xp67_ASAP7_75t_L g560 ( 
.A(n_559),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_560),
.B(n_561),
.Y(n_580)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_544),
.B(n_526),
.C(n_527),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_563),
.B(n_566),
.Y(n_581)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_554),
.B(n_526),
.C(n_529),
.Y(n_566)
);

OAI21xp5_ASAP7_75t_SL g567 ( 
.A1(n_550),
.A2(n_528),
.B(n_535),
.Y(n_567)
);

OAI21xp5_ASAP7_75t_L g573 ( 
.A1(n_567),
.A2(n_545),
.B(n_553),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_570),
.B(n_205),
.Y(n_582)
);

OAI21xp33_ASAP7_75t_L g572 ( 
.A1(n_547),
.A2(n_542),
.B(n_538),
.Y(n_572)
);

AOI31xp67_ASAP7_75t_L g575 ( 
.A1(n_572),
.A2(n_551),
.A3(n_548),
.B(n_542),
.Y(n_575)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_573),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_562),
.B(n_546),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_574),
.B(n_576),
.Y(n_589)
);

XNOR2xp5_ASAP7_75t_L g584 ( 
.A(n_575),
.B(n_578),
.Y(n_584)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_565),
.B(n_558),
.C(n_542),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_571),
.B(n_219),
.Y(n_577)
);

OAI22xp5_ASAP7_75t_L g583 ( 
.A1(n_577),
.A2(n_568),
.B1(n_561),
.B2(n_563),
.Y(n_583)
);

OAI22xp5_ASAP7_75t_L g578 ( 
.A1(n_564),
.A2(n_245),
.B1(n_205),
.B2(n_246),
.Y(n_578)
);

XOR2xp5_ASAP7_75t_L g579 ( 
.A(n_569),
.B(n_246),
.Y(n_579)
);

MAJIxp5_ASAP7_75t_L g585 ( 
.A(n_579),
.B(n_582),
.C(n_567),
.Y(n_585)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_583),
.Y(n_590)
);

XNOR2xp5_ASAP7_75t_L g591 ( 
.A(n_585),
.B(n_576),
.Y(n_591)
);

MAJIxp5_ASAP7_75t_L g587 ( 
.A(n_581),
.B(n_566),
.C(n_569),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_587),
.B(n_589),
.Y(n_592)
);

INVx6_ASAP7_75t_L g588 ( 
.A(n_580),
.Y(n_588)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_588),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_591),
.B(n_592),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_593),
.B(n_587),
.Y(n_594)
);

AOI21xp5_ASAP7_75t_L g596 ( 
.A1(n_594),
.A2(n_586),
.B(n_590),
.Y(n_596)
);

OAI22xp33_ASAP7_75t_SL g598 ( 
.A1(n_596),
.A2(n_597),
.B1(n_588),
.B2(n_584),
.Y(n_598)
);

XOR2xp5_ASAP7_75t_L g597 ( 
.A(n_595),
.B(n_585),
.Y(n_597)
);

AO21x1_ASAP7_75t_L g599 ( 
.A1(n_598),
.A2(n_584),
.B(n_572),
.Y(n_599)
);

OAI22xp33_ASAP7_75t_L g600 ( 
.A1(n_599),
.A2(n_579),
.B1(n_4),
.B2(n_5),
.Y(n_600)
);

AOI21xp5_ASAP7_75t_L g601 ( 
.A1(n_600),
.A2(n_0),
.B(n_5),
.Y(n_601)
);


endmodule