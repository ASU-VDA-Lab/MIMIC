module real_aes_6275_n_98 (n_17, n_28, n_76, n_56, n_34, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_98);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_98;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_656;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_193;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g423 ( .A(n_0), .Y(n_423) );
INVx1_ASAP7_75t_L g479 ( .A(n_1), .Y(n_479) );
INVx1_ASAP7_75t_L g129 ( .A(n_2), .Y(n_129) );
AOI22xp33_ASAP7_75t_L g464 ( .A1(n_3), .A2(n_36), .B1(n_154), .B2(n_435), .Y(n_464) );
AOI21xp33_ASAP7_75t_L g173 ( .A1(n_4), .A2(n_145), .B(n_174), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_5), .B(n_143), .Y(n_490) );
AND2x6_ASAP7_75t_L g122 ( .A(n_6), .B(n_123), .Y(n_122) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_7), .A2(n_227), .B(n_228), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g424 ( .A(n_8), .B(n_37), .Y(n_424) );
INVx1_ASAP7_75t_L g179 ( .A(n_9), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_10), .B(n_208), .Y(n_207) );
INVx1_ASAP7_75t_L g114 ( .A(n_11), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_12), .B(n_135), .Y(n_443) );
INVx1_ASAP7_75t_L g233 ( .A(n_13), .Y(n_233) );
INVx1_ASAP7_75t_L g473 ( .A(n_14), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_15), .B(n_110), .Y(n_495) );
AO32x2_ASAP7_75t_L g462 ( .A1(n_16), .A2(n_109), .A3(n_143), .B1(n_437), .B2(n_463), .Y(n_462) );
NAND2xp5_ASAP7_75t_SL g446 ( .A(n_17), .B(n_154), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_18), .B(n_150), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_19), .B(n_110), .Y(n_481) );
AOI22xp33_ASAP7_75t_L g466 ( .A1(n_20), .A2(n_48), .B1(n_154), .B2(n_435), .Y(n_466) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_21), .B(n_145), .Y(n_190) );
AOI22xp33_ASAP7_75t_SL g436 ( .A1(n_22), .A2(n_74), .B1(n_135), .B2(n_154), .Y(n_436) );
NAND2xp5_ASAP7_75t_SL g458 ( .A(n_23), .B(n_154), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_24), .B(n_157), .Y(n_156) );
A2O1A1Ixp33_ASAP7_75t_L g230 ( .A1(n_25), .A2(n_231), .B(n_232), .C(n_234), .Y(n_230) );
BUFx6f_ASAP7_75t_L g121 ( .A(n_26), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_27), .B(n_140), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_28), .B(n_133), .Y(n_132) );
AOI222xp33_ASAP7_75t_L g98 ( .A1(n_29), .A2(n_99), .B1(n_710), .B2(n_719), .C1(n_727), .C2(n_733), .Y(n_98) );
OAI22xp5_ASAP7_75t_L g721 ( .A1(n_29), .A2(n_102), .B1(n_704), .B2(n_722), .Y(n_721) );
CKINVDCx20_ASAP7_75t_R g722 ( .A(n_29), .Y(n_722) );
INVx1_ASAP7_75t_L g168 ( .A(n_30), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_31), .B(n_140), .Y(n_460) );
INVx2_ASAP7_75t_L g120 ( .A(n_32), .Y(n_120) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_33), .B(n_154), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_34), .B(n_140), .Y(n_448) );
A2O1A1Ixp33_ASAP7_75t_L g191 ( .A1(n_35), .A2(n_122), .B(n_125), .C(n_192), .Y(n_191) );
INVx1_ASAP7_75t_L g166 ( .A(n_38), .Y(n_166) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_39), .B(n_133), .Y(n_220) );
NAND2xp5_ASAP7_75t_SL g485 ( .A(n_40), .B(n_154), .Y(n_485) );
CKINVDCx20_ASAP7_75t_R g725 ( .A(n_41), .Y(n_725) );
AOI22xp33_ASAP7_75t_L g434 ( .A1(n_42), .A2(n_84), .B1(n_197), .B2(n_435), .Y(n_434) );
NAND2xp5_ASAP7_75t_SL g488 ( .A(n_43), .B(n_154), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_44), .B(n_154), .Y(n_474) );
CKINVDCx16_ASAP7_75t_R g169 ( .A(n_45), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_46), .B(n_478), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_47), .B(n_145), .Y(n_210) );
AOI22xp33_ASAP7_75t_SL g499 ( .A1(n_49), .A2(n_58), .B1(n_135), .B2(n_154), .Y(n_499) );
AOI22xp5_ASAP7_75t_L g163 ( .A1(n_50), .A2(n_125), .B1(n_135), .B2(n_164), .Y(n_163) );
CKINVDCx20_ASAP7_75t_R g200 ( .A(n_51), .Y(n_200) );
NAND2xp5_ASAP7_75t_SL g442 ( .A(n_52), .B(n_154), .Y(n_442) );
CKINVDCx16_ASAP7_75t_R g116 ( .A(n_53), .Y(n_116) );
NAND2xp5_ASAP7_75t_SL g513 ( .A(n_54), .B(n_154), .Y(n_513) );
A2O1A1Ixp33_ASAP7_75t_L g176 ( .A1(n_55), .A2(n_153), .B(n_177), .C(n_178), .Y(n_176) );
CKINVDCx20_ASAP7_75t_R g224 ( .A(n_56), .Y(n_224) );
INVx1_ASAP7_75t_L g175 ( .A(n_57), .Y(n_175) );
INVx1_ASAP7_75t_L g123 ( .A(n_59), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_60), .B(n_154), .Y(n_480) );
INVx1_ASAP7_75t_L g113 ( .A(n_61), .Y(n_113) );
CKINVDCx20_ASAP7_75t_R g715 ( .A(n_62), .Y(n_715) );
AO32x2_ASAP7_75t_L g432 ( .A1(n_63), .A2(n_143), .A3(n_202), .B1(n_433), .B2(n_437), .Y(n_432) );
INVx1_ASAP7_75t_L g512 ( .A(n_64), .Y(n_512) );
INVx1_ASAP7_75t_L g455 ( .A(n_65), .Y(n_455) );
AOI222xp33_ASAP7_75t_L g100 ( .A1(n_66), .A2(n_67), .B1(n_101), .B2(n_703), .C1(n_707), .C2(n_708), .Y(n_100) );
INVx1_ASAP7_75t_L g707 ( .A(n_67), .Y(n_707) );
A2O1A1Ixp33_ASAP7_75t_SL g149 ( .A1(n_68), .A2(n_150), .B(n_151), .C(n_153), .Y(n_149) );
INVxp67_ASAP7_75t_L g152 ( .A(n_69), .Y(n_152) );
NAND2xp5_ASAP7_75t_SL g456 ( .A(n_70), .B(n_135), .Y(n_456) );
INVx1_ASAP7_75t_L g714 ( .A(n_71), .Y(n_714) );
CKINVDCx20_ASAP7_75t_R g171 ( .A(n_72), .Y(n_171) );
INVx1_ASAP7_75t_L g217 ( .A(n_73), .Y(n_217) );
A2O1A1Ixp33_ASAP7_75t_L g218 ( .A1(n_75), .A2(n_122), .B(n_125), .C(n_219), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_76), .B(n_435), .Y(n_447) );
NAND2xp5_ASAP7_75t_SL g459 ( .A(n_77), .B(n_135), .Y(n_459) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_78), .B(n_130), .Y(n_193) );
INVx2_ASAP7_75t_L g111 ( .A(n_79), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_80), .B(n_150), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_81), .B(n_135), .Y(n_486) );
A2O1A1Ixp33_ASAP7_75t_L g124 ( .A1(n_82), .A2(n_122), .B(n_125), .C(n_128), .Y(n_124) );
OR2x2_ASAP7_75t_L g421 ( .A(n_83), .B(n_422), .Y(n_421) );
INVx2_ASAP7_75t_L g702 ( .A(n_83), .Y(n_702) );
OR2x2_ASAP7_75t_L g718 ( .A(n_83), .B(n_709), .Y(n_718) );
AOI22xp33_ASAP7_75t_L g498 ( .A1(n_85), .A2(n_97), .B1(n_135), .B2(n_136), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_86), .B(n_140), .Y(n_180) );
CKINVDCx20_ASAP7_75t_R g138 ( .A(n_87), .Y(n_138) );
A2O1A1Ixp33_ASAP7_75t_L g204 ( .A1(n_88), .A2(n_122), .B(n_125), .C(n_205), .Y(n_204) );
CKINVDCx20_ASAP7_75t_R g212 ( .A(n_89), .Y(n_212) );
INVx1_ASAP7_75t_L g148 ( .A(n_90), .Y(n_148) );
CKINVDCx16_ASAP7_75t_R g229 ( .A(n_91), .Y(n_229) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_92), .B(n_130), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_93), .B(n_135), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_94), .B(n_143), .Y(n_235) );
AOI21xp5_ASAP7_75t_L g144 ( .A1(n_95), .A2(n_145), .B(n_146), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_96), .B(n_714), .Y(n_713) );
INVxp67_ASAP7_75t_L g99 ( .A(n_100), .Y(n_99) );
OAI22xp5_ASAP7_75t_SL g101 ( .A1(n_102), .A2(n_419), .B1(n_425), .B2(n_699), .Y(n_101) );
INVx2_ASAP7_75t_L g704 ( .A(n_102), .Y(n_704) );
OR4x1_ASAP7_75t_L g102 ( .A(n_103), .B(n_308), .C(n_368), .D(n_395), .Y(n_102) );
NAND4xp25_ASAP7_75t_SL g103 ( .A(n_104), .B(n_256), .C(n_287), .D(n_304), .Y(n_103) );
O2A1O1Ixp33_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_181), .B(n_183), .C(n_236), .Y(n_104) );
NOR2xp33_ASAP7_75t_L g105 ( .A(n_106), .B(n_159), .Y(n_105) );
INVx1_ASAP7_75t_L g298 ( .A(n_106), .Y(n_298) );
OAI22xp5_ASAP7_75t_L g416 ( .A1(n_106), .A2(n_339), .B1(n_387), .B2(n_417), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_107), .B(n_141), .Y(n_106) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_107), .B(n_243), .Y(n_242) );
OR2x2_ASAP7_75t_L g249 ( .A(n_107), .B(n_161), .Y(n_249) );
AND2x2_ASAP7_75t_L g291 ( .A(n_107), .B(n_292), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_107), .B(n_182), .Y(n_303) );
INVx1_ASAP7_75t_L g343 ( .A(n_107), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_107), .B(n_397), .Y(n_396) );
INVx3_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
AND2x2_ASAP7_75t_L g271 ( .A(n_108), .B(n_161), .Y(n_271) );
INVx3_ASAP7_75t_L g275 ( .A(n_108), .Y(n_275) );
NAND2xp5_ASAP7_75t_SL g332 ( .A(n_108), .B(n_333), .Y(n_332) );
AO21x2_ASAP7_75t_L g108 ( .A1(n_109), .A2(n_115), .B(n_137), .Y(n_108) );
AO21x2_ASAP7_75t_L g161 ( .A1(n_109), .A2(n_162), .B(n_170), .Y(n_161) );
NOR2xp33_ASAP7_75t_L g170 ( .A(n_109), .B(n_171), .Y(n_170) );
INVx2_ASAP7_75t_L g198 ( .A(n_109), .Y(n_198) );
INVx1_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_110), .Y(n_143) );
AND2x2_ASAP7_75t_L g110 ( .A(n_111), .B(n_112), .Y(n_110) );
AND2x2_ASAP7_75t_SL g140 ( .A(n_111), .B(n_112), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_113), .B(n_114), .Y(n_112) );
OAI21xp5_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_117), .B(n_124), .Y(n_115) );
OAI22xp33_ASAP7_75t_L g162 ( .A1(n_117), .A2(n_155), .B1(n_163), .B2(n_169), .Y(n_162) );
OAI21xp5_ASAP7_75t_L g216 ( .A1(n_117), .A2(n_217), .B(n_218), .Y(n_216) );
NAND2x1p5_ASAP7_75t_L g117 ( .A(n_118), .B(n_122), .Y(n_117) );
AND2x4_ASAP7_75t_L g145 ( .A(n_118), .B(n_122), .Y(n_145) );
AND2x2_ASAP7_75t_L g118 ( .A(n_119), .B(n_121), .Y(n_118) );
INVx1_ASAP7_75t_L g478 ( .A(n_119), .Y(n_478) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx2_ASAP7_75t_L g126 ( .A(n_120), .Y(n_126) );
INVx1_ASAP7_75t_L g136 ( .A(n_120), .Y(n_136) );
INVx1_ASAP7_75t_L g127 ( .A(n_121), .Y(n_127) );
INVx3_ASAP7_75t_L g131 ( .A(n_121), .Y(n_131) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_121), .Y(n_133) );
INVx1_ASAP7_75t_L g150 ( .A(n_121), .Y(n_150) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_121), .Y(n_165) );
INVx4_ASAP7_75t_SL g155 ( .A(n_122), .Y(n_155) );
BUFx3_ASAP7_75t_L g437 ( .A(n_122), .Y(n_437) );
OAI21xp5_ASAP7_75t_L g440 ( .A1(n_122), .A2(n_441), .B(n_445), .Y(n_440) );
OAI21xp5_ASAP7_75t_L g453 ( .A1(n_122), .A2(n_454), .B(n_457), .Y(n_453) );
OAI21xp5_ASAP7_75t_L g471 ( .A1(n_122), .A2(n_472), .B(n_476), .Y(n_471) );
OAI21xp5_ASAP7_75t_L g483 ( .A1(n_122), .A2(n_484), .B(n_487), .Y(n_483) );
INVx5_ASAP7_75t_L g147 ( .A(n_125), .Y(n_147) );
AND2x6_ASAP7_75t_L g125 ( .A(n_126), .B(n_127), .Y(n_125) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_126), .Y(n_154) );
BUFx3_ASAP7_75t_L g197 ( .A(n_126), .Y(n_197) );
INVx1_ASAP7_75t_L g435 ( .A(n_126), .Y(n_435) );
O2A1O1Ixp33_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_130), .B(n_132), .C(n_134), .Y(n_128) );
O2A1O1Ixp5_ASAP7_75t_SL g454 ( .A1(n_130), .A2(n_153), .B(n_455), .C(n_456), .Y(n_454) );
INVx2_ASAP7_75t_L g465 ( .A(n_130), .Y(n_465) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_130), .A2(n_485), .B(n_486), .Y(n_484) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_130), .A2(n_509), .B(n_510), .Y(n_508) );
INVx5_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
NOR2xp33_ASAP7_75t_L g151 ( .A(n_131), .B(n_152), .Y(n_151) );
NOR2xp33_ASAP7_75t_L g178 ( .A(n_131), .B(n_179), .Y(n_178) );
OAI22xp5_ASAP7_75t_SL g433 ( .A1(n_131), .A2(n_133), .B1(n_434), .B2(n_436), .Y(n_433) );
INVx2_ASAP7_75t_L g177 ( .A(n_133), .Y(n_177) );
INVx4_ASAP7_75t_L g208 ( .A(n_133), .Y(n_208) );
OAI22xp5_ASAP7_75t_L g463 ( .A1(n_133), .A2(n_464), .B1(n_465), .B2(n_466), .Y(n_463) );
OAI22xp5_ASAP7_75t_L g497 ( .A1(n_133), .A2(n_465), .B1(n_498), .B2(n_499), .Y(n_497) );
O2A1O1Ixp33_ASAP7_75t_L g472 ( .A1(n_134), .A2(n_473), .B(n_474), .C(n_475), .Y(n_472) );
INVx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx3_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
NOR2xp33_ASAP7_75t_L g137 ( .A(n_138), .B(n_139), .Y(n_137) );
NOR2xp33_ASAP7_75t_L g211 ( .A(n_139), .B(n_212), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_139), .B(n_224), .Y(n_223) );
INVx1_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx2_ASAP7_75t_L g202 ( .A(n_140), .Y(n_202) );
OA21x2_ASAP7_75t_L g225 ( .A1(n_140), .A2(n_226), .B(n_235), .Y(n_225) );
OA21x2_ASAP7_75t_L g439 ( .A1(n_140), .A2(n_440), .B(n_448), .Y(n_439) );
OA21x2_ASAP7_75t_L g452 ( .A1(n_140), .A2(n_453), .B(n_460), .Y(n_452) );
AND2x2_ASAP7_75t_L g362 ( .A(n_141), .B(n_172), .Y(n_362) );
NOR2xp33_ASAP7_75t_L g381 ( .A(n_141), .B(n_275), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_141), .B(n_390), .Y(n_389) );
INVx3_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
AND2x2_ASAP7_75t_L g182 ( .A(n_142), .B(n_161), .Y(n_182) );
INVx1_ASAP7_75t_L g244 ( .A(n_142), .Y(n_244) );
BUFx2_ASAP7_75t_L g248 ( .A(n_142), .Y(n_248) );
AND2x2_ASAP7_75t_L g292 ( .A(n_142), .B(n_160), .Y(n_292) );
OR2x2_ASAP7_75t_L g331 ( .A(n_142), .B(n_160), .Y(n_331) );
AND2x2_ASAP7_75t_L g356 ( .A(n_142), .B(n_172), .Y(n_356) );
AND2x2_ASAP7_75t_L g415 ( .A(n_142), .B(n_245), .Y(n_415) );
OA21x2_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_144), .B(n_156), .Y(n_142) );
INVx4_ASAP7_75t_L g158 ( .A(n_143), .Y(n_158) );
OA21x2_ASAP7_75t_L g482 ( .A1(n_143), .A2(n_483), .B(n_490), .Y(n_482) );
BUFx2_ASAP7_75t_L g227 ( .A(n_145), .Y(n_227) );
O2A1O1Ixp33_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_148), .B(n_149), .C(n_155), .Y(n_146) );
O2A1O1Ixp33_ASAP7_75t_L g174 ( .A1(n_147), .A2(n_155), .B(n_175), .C(n_176), .Y(n_174) );
O2A1O1Ixp33_ASAP7_75t_L g228 ( .A1(n_147), .A2(n_155), .B(n_229), .C(n_230), .Y(n_228) );
INVx1_ASAP7_75t_L g444 ( .A(n_150), .Y(n_444) );
INVx3_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
HB1xp67_ASAP7_75t_L g209 ( .A(n_154), .Y(n_209) );
OA21x2_ASAP7_75t_L g172 ( .A1(n_157), .A2(n_173), .B(n_180), .Y(n_172) );
INVx3_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
NOR2xp33_ASAP7_75t_SL g199 ( .A(n_158), .B(n_200), .Y(n_199) );
NAND3xp33_ASAP7_75t_L g496 ( .A(n_158), .B(n_437), .C(n_497), .Y(n_496) );
AO21x1_ASAP7_75t_L g543 ( .A1(n_158), .A2(n_497), .B(n_544), .Y(n_543) );
INVx1_ASAP7_75t_L g390 ( .A(n_159), .Y(n_390) );
OR2x2_ASAP7_75t_L g159 ( .A(n_160), .B(n_172), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_160), .B(n_172), .Y(n_276) );
AND2x2_ASAP7_75t_L g286 ( .A(n_160), .B(n_275), .Y(n_286) );
BUFx2_ASAP7_75t_L g297 ( .A(n_160), .Y(n_297) );
INVx3_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
AND2x2_ASAP7_75t_L g319 ( .A(n_161), .B(n_172), .Y(n_319) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_161), .Y(n_374) );
OAI22xp5_ASAP7_75t_SL g164 ( .A1(n_165), .A2(n_166), .B1(n_167), .B2(n_168), .Y(n_164) );
INVx2_ASAP7_75t_L g167 ( .A(n_165), .Y(n_167) );
INVx4_ASAP7_75t_L g231 ( .A(n_165), .Y(n_231) );
AND2x2_ASAP7_75t_SL g181 ( .A(n_172), .B(n_182), .Y(n_181) );
INVx1_ASAP7_75t_SL g245 ( .A(n_172), .Y(n_245) );
BUFx2_ASAP7_75t_L g270 ( .A(n_172), .Y(n_270) );
INVx2_ASAP7_75t_L g289 ( .A(n_172), .Y(n_289) );
AND2x2_ASAP7_75t_L g351 ( .A(n_172), .B(n_275), .Y(n_351) );
AOI21xp5_ASAP7_75t_L g445 ( .A1(n_177), .A2(n_446), .B(n_447), .Y(n_445) );
O2A1O1Ixp5_ASAP7_75t_L g511 ( .A1(n_177), .A2(n_477), .B(n_512), .C(n_513), .Y(n_511) );
AOI321xp33_ASAP7_75t_L g370 ( .A1(n_181), .A2(n_371), .A3(n_372), .B1(n_373), .B2(n_375), .C(n_376), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_182), .B(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_182), .B(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g364 ( .A(n_182), .B(n_343), .Y(n_364) );
AND2x2_ASAP7_75t_L g397 ( .A(n_182), .B(n_289), .Y(n_397) );
INVx1_ASAP7_75t_SL g183 ( .A(n_184), .Y(n_183) );
OR2x2_ASAP7_75t_L g184 ( .A(n_185), .B(n_213), .Y(n_184) );
OR2x2_ASAP7_75t_L g299 ( .A(n_185), .B(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
AND2x2_ASAP7_75t_L g186 ( .A(n_187), .B(n_201), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx3_ASAP7_75t_L g251 ( .A(n_188), .Y(n_251) );
AND2x2_ASAP7_75t_L g261 ( .A(n_188), .B(n_215), .Y(n_261) );
AND2x2_ASAP7_75t_L g266 ( .A(n_188), .B(n_241), .Y(n_266) );
INVx1_ASAP7_75t_L g283 ( .A(n_188), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_188), .B(n_264), .Y(n_302) );
AND2x2_ASAP7_75t_L g307 ( .A(n_188), .B(n_240), .Y(n_307) );
OR2x2_ASAP7_75t_L g339 ( .A(n_188), .B(n_328), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_188), .B(n_252), .Y(n_378) );
AND2x2_ASAP7_75t_L g412 ( .A(n_188), .B(n_238), .Y(n_412) );
OR2x6_ASAP7_75t_L g188 ( .A(n_189), .B(n_199), .Y(n_188) );
AOI21xp5_ASAP7_75t_SL g189 ( .A1(n_190), .A2(n_191), .B(n_198), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g192 ( .A1(n_193), .A2(n_194), .B(n_195), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_195), .A2(n_220), .B(n_221), .Y(n_219) );
INVx2_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
INVx1_ASAP7_75t_L g234 ( .A(n_197), .Y(n_234) );
INVx1_ASAP7_75t_L g222 ( .A(n_198), .Y(n_222) );
OA21x2_ASAP7_75t_L g470 ( .A1(n_198), .A2(n_471), .B(n_481), .Y(n_470) );
OA21x2_ASAP7_75t_L g506 ( .A1(n_198), .A2(n_507), .B(n_514), .Y(n_506) );
INVx1_ASAP7_75t_L g239 ( .A(n_201), .Y(n_239) );
INVx2_ASAP7_75t_L g254 ( .A(n_201), .Y(n_254) );
AND2x2_ASAP7_75t_L g294 ( .A(n_201), .B(n_265), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_201), .B(n_241), .Y(n_316) );
AO21x2_ASAP7_75t_L g201 ( .A1(n_202), .A2(n_203), .B(n_211), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_204), .B(n_210), .Y(n_203) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_206), .A2(n_207), .B(n_209), .Y(n_205) );
INVx1_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
AND2x2_ASAP7_75t_L g400 ( .A(n_214), .B(n_251), .Y(n_400) );
AND2x2_ASAP7_75t_L g214 ( .A(n_215), .B(n_225), .Y(n_214) );
INVx2_ASAP7_75t_L g241 ( .A(n_215), .Y(n_241) );
AND2x2_ASAP7_75t_L g394 ( .A(n_215), .B(n_254), .Y(n_394) );
AO21x2_ASAP7_75t_L g215 ( .A1(n_216), .A2(n_222), .B(n_223), .Y(n_215) );
AND2x2_ASAP7_75t_L g240 ( .A(n_225), .B(n_241), .Y(n_240) );
INVx2_ASAP7_75t_L g255 ( .A(n_225), .Y(n_255) );
INVx1_ASAP7_75t_L g265 ( .A(n_225), .Y(n_265) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_231), .B(n_233), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g457 ( .A1(n_231), .A2(n_458), .B(n_459), .Y(n_457) );
INVx1_ASAP7_75t_L g475 ( .A(n_231), .Y(n_475) );
OAI22xp33_ASAP7_75t_L g236 ( .A1(n_237), .A2(n_242), .B1(n_246), .B2(n_250), .Y(n_236) );
OAI22xp33_ASAP7_75t_L g391 ( .A1(n_237), .A2(n_355), .B1(n_392), .B2(n_393), .Y(n_391) );
INVx1_ASAP7_75t_SL g237 ( .A(n_238), .Y(n_237) );
AND2x2_ASAP7_75t_L g238 ( .A(n_239), .B(n_240), .Y(n_238) );
INVx1_ASAP7_75t_L g306 ( .A(n_239), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_240), .B(n_283), .Y(n_282) );
INVx2_ASAP7_75t_L g301 ( .A(n_241), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_241), .B(n_254), .Y(n_328) );
INVx1_ASAP7_75t_L g344 ( .A(n_241), .Y(n_344) );
AND2x2_ASAP7_75t_L g285 ( .A(n_243), .B(n_286), .Y(n_285) );
INVx3_ASAP7_75t_SL g324 ( .A(n_243), .Y(n_324) );
NOR2xp33_ASAP7_75t_L g401 ( .A(n_243), .B(n_249), .Y(n_401) );
AND2x4_ASAP7_75t_L g243 ( .A(n_244), .B(n_245), .Y(n_243) );
INVx1_ASAP7_75t_L g410 ( .A(n_246), .Y(n_410) );
OR2x2_ASAP7_75t_L g246 ( .A(n_247), .B(n_249), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_247), .B(n_343), .Y(n_385) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
INVx3_ASAP7_75t_SL g290 ( .A(n_249), .Y(n_290) );
NAND2x1_ASAP7_75t_SL g250 ( .A(n_251), .B(n_252), .Y(n_250) );
AND2x2_ASAP7_75t_L g311 ( .A(n_251), .B(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g318 ( .A(n_251), .B(n_255), .Y(n_318) );
AND2x2_ASAP7_75t_L g323 ( .A(n_251), .B(n_264), .Y(n_323) );
HB1xp67_ASAP7_75t_L g372 ( .A(n_251), .Y(n_372) );
OAI311xp33_ASAP7_75t_L g395 ( .A1(n_252), .A2(n_396), .A3(n_398), .B1(n_399), .C1(n_409), .Y(n_395) );
INVx2_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
OR2x2_ASAP7_75t_L g408 ( .A(n_253), .B(n_281), .Y(n_408) );
OR2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
AND2x2_ASAP7_75t_L g264 ( .A(n_254), .B(n_265), .Y(n_264) );
AND2x2_ASAP7_75t_L g312 ( .A(n_254), .B(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g367 ( .A(n_254), .Y(n_367) );
INVx1_ASAP7_75t_L g260 ( .A(n_255), .Y(n_260) );
INVx1_ASAP7_75t_L g280 ( .A(n_255), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_255), .B(n_301), .Y(n_300) );
INVx2_ASAP7_75t_L g313 ( .A(n_255), .Y(n_313) );
AOI221xp5_ASAP7_75t_SL g256 ( .A1(n_257), .A2(n_259), .B1(n_267), .B2(n_272), .C(n_277), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_258), .B(n_262), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g259 ( .A(n_260), .B(n_261), .Y(n_259) );
INVx4_ASAP7_75t_L g281 ( .A(n_261), .Y(n_281) );
AND2x2_ASAP7_75t_L g375 ( .A(n_261), .B(n_294), .Y(n_375) );
AND2x2_ASAP7_75t_L g382 ( .A(n_261), .B(n_264), .Y(n_382) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g263 ( .A(n_264), .B(n_266), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_264), .B(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g293 ( .A(n_266), .B(n_294), .Y(n_293) );
INVx1_ASAP7_75t_SL g267 ( .A(n_268), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_269), .B(n_271), .Y(n_268) );
NOR2xp33_ASAP7_75t_L g341 ( .A(n_269), .B(n_342), .Y(n_341) );
INVx1_ASAP7_75t_SL g269 ( .A(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g418 ( .A(n_271), .B(n_362), .Y(n_418) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
OR2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_276), .Y(n_273) );
INVx1_ASAP7_75t_SL g274 ( .A(n_275), .Y(n_274) );
OR2x2_ASAP7_75t_L g403 ( .A(n_275), .B(n_331), .Y(n_403) );
OAI211xp5_ASAP7_75t_L g368 ( .A1(n_276), .A2(n_369), .B(n_370), .C(n_383), .Y(n_368) );
AOI21xp33_ASAP7_75t_SL g277 ( .A1(n_278), .A2(n_282), .B(n_284), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
NOR2xp67_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
INVx1_ASAP7_75t_L g347 ( .A(n_281), .Y(n_347) );
OAI221xp5_ASAP7_75t_L g376 ( .A1(n_282), .A2(n_377), .B1(n_378), .B2(n_379), .C(n_380), .Y(n_376) );
AND2x2_ASAP7_75t_L g353 ( .A(n_283), .B(n_294), .Y(n_353) );
AND2x2_ASAP7_75t_L g406 ( .A(n_283), .B(n_301), .Y(n_406) );
INVx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
NOR2xp33_ASAP7_75t_L g348 ( .A(n_286), .B(n_324), .Y(n_348) );
O2A1O1Ixp33_ASAP7_75t_L g287 ( .A1(n_288), .A2(n_291), .B(n_293), .C(n_295), .Y(n_287) );
AND2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_290), .Y(n_288) );
AND2x2_ASAP7_75t_L g334 ( .A(n_289), .B(n_292), .Y(n_334) );
OR2x2_ASAP7_75t_L g377 ( .A(n_289), .B(n_331), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_290), .B(n_356), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_290), .B(n_362), .Y(n_361) );
INVx1_ASAP7_75t_SL g321 ( .A(n_291), .Y(n_321) );
INVx1_ASAP7_75t_L g387 ( .A(n_294), .Y(n_387) );
OAI22xp5_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_299), .B1(n_302), .B2(n_303), .Y(n_295) );
INVx1_ASAP7_75t_L g310 ( .A(n_296), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_297), .B(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g373 ( .A(n_298), .B(n_374), .Y(n_373) );
INVxp67_ASAP7_75t_L g359 ( .A(n_300), .Y(n_359) );
NOR2xp33_ASAP7_75t_L g386 ( .A(n_301), .B(n_387), .Y(n_386) );
OAI22xp33_ASAP7_75t_L g360 ( .A1(n_302), .A2(n_361), .B1(n_363), .B2(n_365), .Y(n_360) );
INVx1_ASAP7_75t_L g369 ( .A(n_305), .Y(n_369) );
AND2x2_ASAP7_75t_L g305 ( .A(n_306), .B(n_307), .Y(n_305) );
AND2x2_ASAP7_75t_L g411 ( .A(n_306), .B(n_406), .Y(n_411) );
AOI222xp33_ASAP7_75t_L g340 ( .A1(n_307), .A2(n_341), .B1(n_344), .B2(n_345), .C1(n_348), .C2(n_349), .Y(n_340) );
NAND4xp25_ASAP7_75t_SL g308 ( .A(n_309), .B(n_329), .C(n_340), .D(n_352), .Y(n_308) );
AOI221xp5_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_311), .B1(n_314), .B2(n_319), .C(n_320), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_312), .B(n_347), .Y(n_346) );
INVxp67_ASAP7_75t_L g338 ( .A(n_313), .Y(n_338) );
AOI221xp5_ASAP7_75t_L g383 ( .A1(n_314), .A2(n_384), .B1(n_386), .B2(n_388), .C(n_391), .Y(n_383) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
OR2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g326 ( .A(n_318), .B(n_327), .Y(n_326) );
OAI21xp33_ASAP7_75t_L g380 ( .A1(n_319), .A2(n_381), .B(n_382), .Y(n_380) );
OAI22xp5_ASAP7_75t_L g320 ( .A1(n_321), .A2(n_322), .B1(n_324), .B2(n_325), .Y(n_320) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx2_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
OAI21xp5_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_332), .B(n_335), .Y(n_329) );
INVxp67_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
OR2x2_ASAP7_75t_L g336 ( .A(n_337), .B(n_339), .Y(n_336) );
HB1xp67_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g371 ( .A(n_342), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_343), .B(n_362), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_343), .B(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_347), .B(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_SL g379 ( .A(n_351), .Y(n_379) );
AOI221xp5_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_354), .B1(n_357), .B2(n_359), .C(n_360), .Y(n_352) );
INVxp67_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
AOI222xp33_ASAP7_75t_L g399 ( .A1(n_362), .A2(n_400), .B1(n_401), .B2(n_402), .C1(n_404), .C2(n_407), .Y(n_399) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_366), .B(n_406), .Y(n_405) );
INVxp67_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g398 ( .A(n_372), .Y(n_398) );
INVxp67_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVxp33_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
AOI221xp5_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_411), .B1(n_412), .B2(n_413), .C(n_416), .Y(n_409) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVxp67_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
OAI22xp5_ASAP7_75t_L g703 ( .A1(n_419), .A2(n_704), .B1(n_705), .B2(n_706), .Y(n_703) );
INVx2_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
OR2x2_ASAP7_75t_L g701 ( .A(n_422), .B(n_702), .Y(n_701) );
INVx2_ASAP7_75t_L g709 ( .A(n_422), .Y(n_709) );
AND2x2_ASAP7_75t_L g422 ( .A(n_423), .B(n_424), .Y(n_422) );
INVx2_ASAP7_75t_L g706 ( .A(n_425), .Y(n_706) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
AND3x1_ASAP7_75t_L g426 ( .A(n_427), .B(n_619), .C(n_667), .Y(n_426) );
NOR4xp25_ASAP7_75t_L g427 ( .A(n_428), .B(n_547), .C(n_592), .D(n_606), .Y(n_427) );
OAI311xp33_ASAP7_75t_L g428 ( .A1(n_429), .A2(n_467), .A3(n_491), .B1(n_500), .C1(n_515), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_430), .B(n_438), .Y(n_429) );
OAI21xp33_ASAP7_75t_L g500 ( .A1(n_430), .A2(n_501), .B(n_503), .Y(n_500) );
AND2x2_ASAP7_75t_L g608 ( .A(n_430), .B(n_535), .Y(n_608) );
AND2x2_ASAP7_75t_L g665 ( .A(n_430), .B(n_551), .Y(n_665) );
BUFx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
AND2x2_ASAP7_75t_L g558 ( .A(n_431), .B(n_461), .Y(n_558) );
AND2x2_ASAP7_75t_L g615 ( .A(n_431), .B(n_563), .Y(n_615) );
INVx1_ASAP7_75t_L g656 ( .A(n_431), .Y(n_656) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
BUFx6f_ASAP7_75t_L g524 ( .A(n_432), .Y(n_524) );
AND2x2_ASAP7_75t_L g565 ( .A(n_432), .B(n_461), .Y(n_565) );
AND2x2_ASAP7_75t_L g569 ( .A(n_432), .B(n_462), .Y(n_569) );
INVx1_ASAP7_75t_L g581 ( .A(n_432), .Y(n_581) );
OAI21xp5_ASAP7_75t_L g507 ( .A1(n_437), .A2(n_508), .B(n_511), .Y(n_507) );
AND2x2_ASAP7_75t_L g438 ( .A(n_439), .B(n_449), .Y(n_438) );
AND2x2_ASAP7_75t_L g502 ( .A(n_439), .B(n_461), .Y(n_502) );
INVx2_ASAP7_75t_L g536 ( .A(n_439), .Y(n_536) );
AND2x2_ASAP7_75t_L g551 ( .A(n_439), .B(n_462), .Y(n_551) );
HB1xp67_ASAP7_75t_L g557 ( .A(n_439), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_439), .B(n_563), .Y(n_562) );
OR2x2_ASAP7_75t_L g571 ( .A(n_439), .B(n_534), .Y(n_571) );
INVx1_ASAP7_75t_L g583 ( .A(n_439), .Y(n_583) );
INVx1_ASAP7_75t_L g624 ( .A(n_439), .Y(n_624) );
NOR2xp33_ASAP7_75t_L g677 ( .A(n_439), .B(n_524), .Y(n_677) );
AOI21xp5_ASAP7_75t_L g441 ( .A1(n_442), .A2(n_443), .B(n_444), .Y(n_441) );
NOR2xp67_ASAP7_75t_L g449 ( .A(n_450), .B(n_461), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
AND2x2_ASAP7_75t_L g501 ( .A(n_451), .B(n_502), .Y(n_501) );
HB1xp67_ASAP7_75t_L g529 ( .A(n_451), .Y(n_529) );
AND2x2_ASAP7_75t_SL g582 ( .A(n_451), .B(n_583), .Y(n_582) );
OR2x2_ASAP7_75t_L g586 ( .A(n_451), .B(n_461), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_451), .B(n_581), .Y(n_644) );
INVx2_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx2_ASAP7_75t_L g534 ( .A(n_452), .Y(n_534) );
HB1xp67_ASAP7_75t_L g550 ( .A(n_452), .Y(n_550) );
OR2x2_ASAP7_75t_L g623 ( .A(n_452), .B(n_624), .Y(n_623) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
BUFx2_ASAP7_75t_L g530 ( .A(n_462), .Y(n_530) );
AND2x2_ASAP7_75t_L g535 ( .A(n_462), .B(n_536), .Y(n_535) );
O2A1O1Ixp33_ASAP7_75t_L g476 ( .A1(n_465), .A2(n_477), .B(n_479), .C(n_480), .Y(n_476) );
AOI21xp5_ASAP7_75t_L g487 ( .A1(n_465), .A2(n_488), .B(n_489), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_467), .B(n_518), .Y(n_681) );
INVx1_ASAP7_75t_SL g467 ( .A(n_468), .Y(n_467) );
OR2x2_ASAP7_75t_L g651 ( .A(n_468), .B(n_493), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_469), .B(n_482), .Y(n_468) );
AND2x2_ASAP7_75t_L g527 ( .A(n_469), .B(n_518), .Y(n_527) );
INVx2_ASAP7_75t_L g539 ( .A(n_469), .Y(n_539) );
AND2x2_ASAP7_75t_L g573 ( .A(n_469), .B(n_521), .Y(n_573) );
AND2x2_ASAP7_75t_L g640 ( .A(n_469), .B(n_641), .Y(n_640) );
INVx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_470), .B(n_506), .Y(n_505) );
AND2x2_ASAP7_75t_L g520 ( .A(n_470), .B(n_521), .Y(n_520) );
AND2x2_ASAP7_75t_L g560 ( .A(n_470), .B(n_482), .Y(n_560) );
AND2x2_ASAP7_75t_L g577 ( .A(n_470), .B(n_578), .Y(n_577) );
INVx2_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
AND2x2_ASAP7_75t_L g503 ( .A(n_482), .B(n_504), .Y(n_503) );
INVx3_ASAP7_75t_L g521 ( .A(n_482), .Y(n_521) );
AND2x2_ASAP7_75t_L g526 ( .A(n_482), .B(n_506), .Y(n_526) );
AND2x2_ASAP7_75t_L g599 ( .A(n_482), .B(n_578), .Y(n_599) );
AND2x2_ASAP7_75t_L g664 ( .A(n_482), .B(n_654), .Y(n_664) );
OAI311xp33_ASAP7_75t_L g547 ( .A1(n_491), .A2(n_548), .A3(n_552), .B1(n_554), .C1(n_574), .Y(n_547) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
AND2x2_ASAP7_75t_L g559 ( .A(n_492), .B(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g618 ( .A(n_492), .B(n_526), .Y(n_618) );
AND2x2_ASAP7_75t_L g692 ( .A(n_492), .B(n_573), .Y(n_692) );
INVx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_493), .B(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g627 ( .A(n_493), .Y(n_627) );
INVx2_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx3_ASAP7_75t_L g518 ( .A(n_494), .Y(n_518) );
NOR2x1_ASAP7_75t_L g590 ( .A(n_494), .B(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g647 ( .A(n_494), .B(n_521), .Y(n_647) );
AND2x4_ASAP7_75t_L g494 ( .A(n_495), .B(n_496), .Y(n_494) );
INVx1_ASAP7_75t_L g544 ( .A(n_495), .Y(n_544) );
AND2x2_ASAP7_75t_L g522 ( .A(n_502), .B(n_523), .Y(n_522) );
AND2x2_ASAP7_75t_L g575 ( .A(n_502), .B(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g655 ( .A(n_502), .B(n_656), .Y(n_655) );
AOI221xp5_ASAP7_75t_L g554 ( .A1(n_503), .A2(n_535), .B1(n_555), .B2(n_559), .C(n_561), .Y(n_554) );
INVx1_ASAP7_75t_L g679 ( .A(n_504), .Y(n_679) );
OR2x2_ASAP7_75t_L g645 ( .A(n_505), .B(n_646), .Y(n_645) );
AND2x2_ASAP7_75t_L g540 ( .A(n_506), .B(n_521), .Y(n_540) );
OR2x2_ASAP7_75t_L g542 ( .A(n_506), .B(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g567 ( .A(n_506), .Y(n_567) );
INVx2_ASAP7_75t_L g578 ( .A(n_506), .Y(n_578) );
AND2x2_ASAP7_75t_L g605 ( .A(n_506), .B(n_543), .Y(n_605) );
HB1xp67_ASAP7_75t_L g634 ( .A(n_506), .Y(n_634) );
AOI221xp5_ASAP7_75t_L g515 ( .A1(n_516), .A2(n_522), .B1(n_525), .B2(n_528), .C(n_531), .Y(n_515) );
INVx1_ASAP7_75t_SL g516 ( .A(n_517), .Y(n_516) );
OR2x2_ASAP7_75t_L g517 ( .A(n_518), .B(n_519), .Y(n_517) );
AND2x2_ASAP7_75t_L g616 ( .A(n_518), .B(n_526), .Y(n_616) );
AND2x2_ASAP7_75t_L g666 ( .A(n_518), .B(n_520), .Y(n_666) );
INVx2_ASAP7_75t_SL g519 ( .A(n_520), .Y(n_519) );
AND2x2_ASAP7_75t_L g553 ( .A(n_520), .B(n_524), .Y(n_553) );
AND2x2_ASAP7_75t_L g632 ( .A(n_520), .B(n_605), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_521), .B(n_567), .Y(n_566) );
INVx2_ASAP7_75t_L g591 ( .A(n_521), .Y(n_591) );
OAI21xp33_ASAP7_75t_L g601 ( .A1(n_522), .A2(n_602), .B(n_604), .Y(n_601) );
OR2x2_ASAP7_75t_L g545 ( .A(n_523), .B(n_546), .Y(n_545) );
OR2x2_ASAP7_75t_L g611 ( .A(n_523), .B(n_571), .Y(n_611) );
NOR2xp33_ASAP7_75t_L g622 ( .A(n_523), .B(n_623), .Y(n_622) );
INVx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
AND2x2_ASAP7_75t_L g588 ( .A(n_524), .B(n_557), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_524), .B(n_671), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_525), .B(n_551), .Y(n_661) );
AND2x2_ASAP7_75t_L g525 ( .A(n_526), .B(n_527), .Y(n_525) );
AND2x2_ASAP7_75t_L g584 ( .A(n_526), .B(n_539), .Y(n_584) );
INVx1_ASAP7_75t_L g600 ( .A(n_527), .Y(n_600) );
NOR2xp33_ASAP7_75t_L g528 ( .A(n_529), .B(n_530), .Y(n_528) );
OAI22xp5_ASAP7_75t_L g531 ( .A1(n_532), .A2(n_537), .B1(n_541), .B2(n_545), .Y(n_531) );
INVx2_ASAP7_75t_SL g532 ( .A(n_533), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_534), .B(n_535), .Y(n_533) );
INVx2_ASAP7_75t_L g563 ( .A(n_534), .Y(n_563) );
INVx1_ASAP7_75t_L g576 ( .A(n_534), .Y(n_576) );
INVx1_ASAP7_75t_L g546 ( .A(n_535), .Y(n_546) );
AND2x2_ASAP7_75t_L g617 ( .A(n_535), .B(n_563), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_535), .B(n_643), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_538), .B(n_540), .Y(n_537) );
OR2x2_ASAP7_75t_L g541 ( .A(n_538), .B(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_538), .B(n_654), .Y(n_653) );
NOR2xp67_ASAP7_75t_L g685 ( .A(n_538), .B(n_686), .Y(n_685) );
INVx3_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
AND2x2_ASAP7_75t_L g688 ( .A(n_540), .B(n_640), .Y(n_688) );
INVx1_ASAP7_75t_SL g654 ( .A(n_542), .Y(n_654) );
AND2x2_ASAP7_75t_L g594 ( .A(n_543), .B(n_578), .Y(n_594) );
INVx1_ASAP7_75t_L g641 ( .A(n_543), .Y(n_641) );
OAI222xp33_ASAP7_75t_L g682 ( .A1(n_548), .A2(n_638), .B1(n_683), .B2(n_684), .C1(n_687), .C2(n_689), .Y(n_682) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_550), .B(n_551), .Y(n_549) );
INVx1_ASAP7_75t_L g603 ( .A(n_550), .Y(n_603) );
AND2x2_ASAP7_75t_L g614 ( .A(n_551), .B(n_615), .Y(n_614) );
NAND2xp5_ASAP7_75t_SL g683 ( .A(n_551), .B(n_656), .Y(n_683) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_553), .B(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g658 ( .A(n_555), .Y(n_658) );
AND2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_558), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx1_ASAP7_75t_SL g596 ( .A(n_558), .Y(n_596) );
AND2x2_ASAP7_75t_L g675 ( .A(n_558), .B(n_636), .Y(n_675) );
AND2x2_ASAP7_75t_L g698 ( .A(n_558), .B(n_582), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_560), .B(n_594), .Y(n_593) );
OAI32xp33_ASAP7_75t_L g561 ( .A1(n_562), .A2(n_564), .A3(n_566), .B1(n_568), .B2(n_572), .Y(n_561) );
BUFx2_ASAP7_75t_L g636 ( .A(n_563), .Y(n_636) );
NOR2xp33_ASAP7_75t_L g663 ( .A(n_564), .B(n_582), .Y(n_663) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g602 ( .A(n_565), .B(n_603), .Y(n_602) );
AND2x4_ASAP7_75t_L g670 ( .A(n_565), .B(n_671), .Y(n_670) );
OR2x2_ASAP7_75t_L g659 ( .A(n_566), .B(n_660), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_569), .B(n_570), .Y(n_568) );
AND2x2_ASAP7_75t_L g630 ( .A(n_569), .B(n_603), .Y(n_630) );
INVx2_ASAP7_75t_SL g570 ( .A(n_571), .Y(n_570) );
OAI221xp5_ASAP7_75t_SL g592 ( .A1(n_571), .A2(n_593), .B1(n_595), .B2(n_597), .C(n_601), .Y(n_592) );
INVx2_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g604 ( .A(n_573), .B(n_605), .Y(n_604) );
AND2x2_ASAP7_75t_L g610 ( .A(n_573), .B(n_594), .Y(n_610) );
AOI221xp5_ASAP7_75t_L g574 ( .A1(n_575), .A2(n_577), .B1(n_579), .B2(n_584), .C(n_585), .Y(n_574) );
INVx1_ASAP7_75t_L g693 ( .A(n_575), .Y(n_693) );
NAND2xp5_ASAP7_75t_SL g669 ( .A(n_576), .B(n_670), .Y(n_669) );
NAND2x1p5_ASAP7_75t_L g589 ( .A(n_577), .B(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g579 ( .A(n_580), .B(n_582), .Y(n_579) );
HB1xp67_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_582), .B(n_596), .Y(n_595) );
INVx2_ASAP7_75t_L g648 ( .A(n_582), .Y(n_648) );
BUFx3_ASAP7_75t_L g671 ( .A(n_583), .Y(n_671) );
INVx1_ASAP7_75t_SL g612 ( .A(n_584), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_584), .B(n_626), .Y(n_625) );
AOI21xp33_ASAP7_75t_SL g585 ( .A1(n_586), .A2(n_587), .B(n_589), .Y(n_585) );
OAI221xp5_ASAP7_75t_L g690 ( .A1(n_586), .A2(n_687), .B1(n_691), .B2(n_693), .C(n_694), .Y(n_690) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g633 ( .A(n_591), .B(n_594), .Y(n_633) );
INVx1_ASAP7_75t_L g697 ( .A(n_591), .Y(n_697) );
INVx2_ASAP7_75t_L g686 ( .A(n_594), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_594), .B(n_697), .Y(n_696) );
OR2x2_ASAP7_75t_L g597 ( .A(n_598), .B(n_600), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g639 ( .A(n_599), .B(n_640), .Y(n_639) );
OAI221xp5_ASAP7_75t_SL g606 ( .A1(n_607), .A2(n_609), .B1(n_611), .B2(n_612), .C(n_613), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx1_ASAP7_75t_SL g609 ( .A(n_610), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g613 ( .A1(n_614), .A2(n_616), .B1(n_617), .B2(n_618), .Y(n_613) );
AOI22xp5_ASAP7_75t_L g676 ( .A1(n_615), .A2(n_677), .B1(n_678), .B2(n_680), .Y(n_676) );
OAI21xp5_ASAP7_75t_L g694 ( .A1(n_618), .A2(n_695), .B(n_698), .Y(n_694) );
NOR4xp25_ASAP7_75t_SL g619 ( .A(n_620), .B(n_628), .C(n_637), .D(n_657), .Y(n_619) );
NOR2xp33_ASAP7_75t_L g620 ( .A(n_621), .B(n_625), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
OAI22xp5_ASAP7_75t_L g628 ( .A1(n_629), .A2(n_631), .B1(n_634), .B2(n_635), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
NOR2xp33_ASAP7_75t_L g631 ( .A(n_632), .B(n_633), .Y(n_631) );
INVx1_ASAP7_75t_L g673 ( .A(n_633), .Y(n_673) );
OAI221xp5_ASAP7_75t_L g637 ( .A1(n_638), .A2(n_642), .B1(n_645), .B2(n_648), .C(n_649), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g660 ( .A(n_640), .Y(n_660) );
INVx1_ASAP7_75t_SL g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
OAI21xp5_ASAP7_75t_SL g649 ( .A1(n_650), .A2(n_652), .B(n_655), .Y(n_649) );
INVx1_ASAP7_75t_SL g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
OAI211xp5_ASAP7_75t_L g657 ( .A1(n_658), .A2(n_659), .B(n_661), .C(n_662), .Y(n_657) );
AOI22xp5_ASAP7_75t_L g662 ( .A1(n_663), .A2(n_664), .B1(n_665), .B2(n_666), .Y(n_662) );
CKINVDCx14_ASAP7_75t_R g672 ( .A(n_666), .Y(n_672) );
NOR3xp33_ASAP7_75t_L g667 ( .A(n_668), .B(n_682), .C(n_690), .Y(n_667) );
OAI221xp5_ASAP7_75t_L g668 ( .A1(n_669), .A2(n_672), .B1(n_673), .B2(n_674), .C(n_676), .Y(n_668) );
INVxp67_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_SL g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
CKINVDCx16_ASAP7_75t_R g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx2_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx2_ASAP7_75t_L g705 ( .A(n_700), .Y(n_705) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
NOR2x2_ASAP7_75t_L g708 ( .A(n_702), .B(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
NAND2xp33_ASAP7_75t_L g711 ( .A(n_712), .B(n_716), .Y(n_711) );
NOR2xp33_ASAP7_75t_SL g712 ( .A(n_713), .B(n_715), .Y(n_712) );
INVx1_ASAP7_75t_SL g732 ( .A(n_713), .Y(n_732) );
INVx1_ASAP7_75t_L g731 ( .A(n_715), .Y(n_731) );
OA21x2_ASAP7_75t_L g734 ( .A1(n_715), .A2(n_732), .B(n_735), .Y(n_734) );
INVx1_ASAP7_75t_SL g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_SL g717 ( .A(n_718), .Y(n_717) );
HB1xp67_ASAP7_75t_L g723 ( .A(n_718), .Y(n_723) );
HB1xp67_ASAP7_75t_L g726 ( .A(n_718), .Y(n_726) );
BUFx2_ASAP7_75t_L g735 ( .A(n_718), .Y(n_735) );
INVxp67_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
AOI21xp5_ASAP7_75t_L g720 ( .A1(n_721), .A2(n_723), .B(n_724), .Y(n_720) );
NOR2xp33_ASAP7_75t_L g724 ( .A(n_725), .B(n_726), .Y(n_724) );
CKINVDCx20_ASAP7_75t_R g727 ( .A(n_728), .Y(n_727) );
CKINVDCx20_ASAP7_75t_R g728 ( .A(n_729), .Y(n_728) );
AND2x2_ASAP7_75t_L g729 ( .A(n_730), .B(n_732), .Y(n_729) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_SL g733 ( .A(n_734), .Y(n_733) );
endmodule