module real_aes_6344_n_286 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_285, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_283, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_281, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_284, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_282, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_286);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_285;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_283;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_281;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_284;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_282;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_286;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_624;
wire n_800;
wire n_778;
wire n_618;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_287;
wire n_503;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_878;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_766;
wire n_852;
wire n_329;
wire n_857;
wire n_461;
wire n_571;
wire n_549;
wire n_376;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_884;
wire n_560;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_767;
wire n_696;
wire n_889;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_415;
wire n_572;
wire n_815;
wire n_519;
wire n_638;
wire n_564;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_462;
wire n_289;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_356;
wire n_478;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_352;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_693;
wire n_496;
wire n_468;
wire n_746;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_874;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_671;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_867;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_807;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_361;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_296;
wire n_702;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_848;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_723;
wire n_662;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_692;
wire n_544;
wire n_789;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_472;
wire n_866;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_741;
wire n_314;
wire n_753;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_456;
wire n_359;
wire n_717;
wire n_712;
wire n_312;
wire n_433;
wire n_516;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_639;
wire n_546;
wire n_587;
wire n_811;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_836;
wire n_888;
wire n_793;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_652;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_842;
wire n_849;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
INVx1_ASAP7_75t_L g670 ( .A(n_0), .Y(n_670) );
AOI22xp5_ASAP7_75t_SL g750 ( .A1(n_1), .A2(n_239), .B1(n_547), .B2(n_658), .Y(n_750) );
AOI22xp33_ASAP7_75t_SL g802 ( .A1(n_2), .A2(n_17), .B1(n_402), .B2(n_523), .Y(n_802) );
AOI22xp5_ASAP7_75t_L g799 ( .A1(n_3), .A2(n_120), .B1(n_377), .B2(n_800), .Y(n_799) );
AOI22xp33_ASAP7_75t_L g497 ( .A1(n_4), .A2(n_19), .B1(n_498), .B2(n_499), .Y(n_497) );
CKINVDCx20_ASAP7_75t_R g549 ( .A(n_5), .Y(n_549) );
AOI22xp5_ASAP7_75t_L g690 ( .A1(n_6), .A2(n_61), .B1(n_346), .B2(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g654 ( .A(n_7), .Y(n_654) );
INVx1_ASAP7_75t_L g561 ( .A(n_8), .Y(n_561) );
CKINVDCx20_ASAP7_75t_R g553 ( .A(n_9), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g303 ( .A1(n_10), .A2(n_131), .B1(n_304), .B2(n_319), .Y(n_303) );
CKINVDCx20_ASAP7_75t_R g581 ( .A(n_11), .Y(n_581) );
CKINVDCx20_ASAP7_75t_R g715 ( .A(n_12), .Y(n_715) );
AOI22xp33_ASAP7_75t_SL g790 ( .A1(n_13), .A2(n_139), .B1(n_512), .B2(n_791), .Y(n_790) );
AOI22xp5_ASAP7_75t_L g702 ( .A1(n_14), .A2(n_150), .B1(n_356), .B2(n_513), .Y(n_702) );
AOI222xp33_ASAP7_75t_L g404 ( .A1(n_15), .A2(n_129), .B1(n_217), .B2(n_377), .C1(n_405), .C2(n_406), .Y(n_404) );
AOI22xp33_ASAP7_75t_SL g785 ( .A1(n_16), .A2(n_220), .B1(n_786), .B2(n_788), .Y(n_785) );
AOI22xp33_ASAP7_75t_L g882 ( .A1(n_18), .A2(n_36), .B1(n_394), .B2(n_482), .Y(n_882) );
AOI221xp5_ASAP7_75t_L g572 ( .A1(n_20), .A2(n_115), .B1(n_498), .B2(n_573), .C(n_574), .Y(n_572) );
CKINVDCx20_ASAP7_75t_R g754 ( .A(n_21), .Y(n_754) );
CKINVDCx20_ASAP7_75t_R g545 ( .A(n_22), .Y(n_545) );
AOI22xp33_ASAP7_75t_SL g480 ( .A1(n_23), .A2(n_169), .B1(n_481), .B2(n_482), .Y(n_480) );
AOI222xp33_ASAP7_75t_L g521 ( .A1(n_24), .A2(n_90), .B1(n_144), .B2(n_522), .C1(n_523), .C2(n_524), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g874 ( .A1(n_25), .A2(n_143), .B1(n_377), .B2(n_695), .Y(n_874) );
AOI22xp33_ASAP7_75t_L g455 ( .A1(n_26), .A2(n_106), .B1(n_456), .B2(n_458), .Y(n_455) );
INVx1_ASAP7_75t_L g663 ( .A(n_27), .Y(n_663) );
CKINVDCx20_ASAP7_75t_R g537 ( .A(n_28), .Y(n_537) );
NAND2xp5_ASAP7_75t_SL g474 ( .A(n_29), .B(n_475), .Y(n_474) );
AO22x2_ASAP7_75t_L g316 ( .A1(n_30), .A2(n_94), .B1(n_308), .B2(n_313), .Y(n_316) );
INVx1_ASAP7_75t_L g826 ( .A(n_30), .Y(n_826) );
AOI22xp33_ASAP7_75t_L g391 ( .A1(n_31), .A2(n_193), .B1(n_304), .B2(n_392), .Y(n_391) );
AOI211xp5_ASAP7_75t_L g286 ( .A1(n_32), .A2(n_287), .B(n_296), .C(n_828), .Y(n_286) );
AOI22xp33_ASAP7_75t_SL g758 ( .A1(n_33), .A2(n_208), .B1(n_371), .B2(n_402), .Y(n_758) );
AOI22xp5_ASAP7_75t_L g633 ( .A1(n_34), .A2(n_158), .B1(n_487), .B2(n_501), .Y(n_633) );
AOI22xp5_ASAP7_75t_L g697 ( .A1(n_35), .A2(n_260), .B1(n_332), .B2(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g660 ( .A(n_37), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_38), .B(n_400), .Y(n_399) );
CKINVDCx20_ASAP7_75t_R g839 ( .A(n_39), .Y(n_839) );
INVx1_ASAP7_75t_L g693 ( .A(n_40), .Y(n_693) );
AOI22xp5_ASAP7_75t_L g829 ( .A1(n_41), .A2(n_830), .B1(n_852), .B2(n_853), .Y(n_829) );
CKINVDCx20_ASAP7_75t_R g852 ( .A(n_41), .Y(n_852) );
AOI22xp33_ASAP7_75t_SL g476 ( .A1(n_42), .A2(n_177), .B1(n_346), .B2(n_350), .Y(n_476) );
AO22x2_ASAP7_75t_L g318 ( .A1(n_43), .A2(n_97), .B1(n_308), .B2(n_309), .Y(n_318) );
INVx1_ASAP7_75t_L g827 ( .A(n_43), .Y(n_827) );
AOI22xp5_ASAP7_75t_L g534 ( .A1(n_44), .A2(n_135), .B1(n_351), .B2(n_378), .Y(n_534) );
CKINVDCx20_ASAP7_75t_R g850 ( .A(n_45), .Y(n_850) );
AOI22xp33_ASAP7_75t_L g657 ( .A1(n_46), .A2(n_162), .B1(n_512), .B2(n_658), .Y(n_657) );
AOI22xp33_ASAP7_75t_L g803 ( .A1(n_47), .A2(n_269), .B1(n_342), .B2(n_517), .Y(n_803) );
AOI22xp33_ASAP7_75t_L g751 ( .A1(n_48), .A2(n_166), .B1(n_359), .B2(n_501), .Y(n_751) );
AOI22xp33_ASAP7_75t_L g507 ( .A1(n_49), .A2(n_91), .B1(n_456), .B2(n_508), .Y(n_507) );
CKINVDCx20_ASAP7_75t_R g893 ( .A(n_50), .Y(n_893) );
CKINVDCx20_ASAP7_75t_R g728 ( .A(n_51), .Y(n_728) );
AOI22xp33_ASAP7_75t_SL g609 ( .A1(n_52), .A2(n_114), .B1(n_461), .B2(n_503), .Y(n_609) );
CKINVDCx20_ASAP7_75t_R g470 ( .A(n_53), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_54), .B(n_430), .Y(n_429) );
AOI22xp33_ASAP7_75t_SL g607 ( .A1(n_55), .A2(n_75), .B1(n_499), .B2(n_608), .Y(n_607) );
CKINVDCx20_ASAP7_75t_R g870 ( .A(n_56), .Y(n_870) );
AOI22xp33_ASAP7_75t_SL g603 ( .A1(n_57), .A2(n_161), .B1(n_520), .B2(n_604), .Y(n_603) );
CKINVDCx20_ASAP7_75t_R g722 ( .A(n_58), .Y(n_722) );
AOI222xp33_ASAP7_75t_L g367 ( .A1(n_59), .A2(n_187), .B1(n_261), .B2(n_368), .C1(n_371), .C2(n_375), .Y(n_367) );
AOI22xp33_ASAP7_75t_L g459 ( .A1(n_60), .A2(n_121), .B1(n_460), .B2(n_461), .Y(n_459) );
AOI22xp33_ASAP7_75t_SL g612 ( .A1(n_62), .A2(n_64), .B1(n_394), .B2(n_449), .Y(n_612) );
CKINVDCx20_ASAP7_75t_R g876 ( .A(n_63), .Y(n_876) );
AOI22xp5_ASAP7_75t_SL g747 ( .A1(n_65), .A2(n_164), .B1(n_487), .B2(n_748), .Y(n_747) );
OAI22xp5_ASAP7_75t_L g765 ( .A1(n_66), .A2(n_766), .B1(n_767), .B2(n_768), .Y(n_765) );
INVx1_ASAP7_75t_L g766 ( .A(n_66), .Y(n_766) );
CKINVDCx20_ASAP7_75t_R g618 ( .A(n_67), .Y(n_618) );
AOI22xp5_ASAP7_75t_L g564 ( .A1(n_68), .A2(n_565), .B1(n_566), .B2(n_586), .Y(n_564) );
INVx1_ASAP7_75t_L g586 ( .A(n_68), .Y(n_586) );
AOI221xp5_ASAP7_75t_L g579 ( .A1(n_69), .A2(n_103), .B1(n_342), .B2(n_516), .C(n_580), .Y(n_579) );
CKINVDCx20_ASAP7_75t_R g629 ( .A(n_70), .Y(n_629) );
AOI22xp33_ASAP7_75t_L g635 ( .A1(n_71), .A2(n_277), .B1(n_385), .B2(n_479), .Y(n_635) );
CKINVDCx20_ASAP7_75t_R g846 ( .A(n_72), .Y(n_846) );
AOI22xp33_ASAP7_75t_L g401 ( .A1(n_73), .A2(n_152), .B1(n_402), .B2(n_403), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g844 ( .A1(n_74), .A2(n_191), .B1(n_481), .B2(n_667), .Y(n_844) );
AOI22xp33_ASAP7_75t_L g355 ( .A1(n_76), .A2(n_180), .B1(n_356), .B2(n_359), .Y(n_355) );
AOI22xp33_ASAP7_75t_SL g478 ( .A1(n_77), .A2(n_195), .B1(n_356), .B2(n_479), .Y(n_478) );
NAND2xp5_ASAP7_75t_SL g602 ( .A(n_78), .B(n_517), .Y(n_602) );
AOI22xp33_ASAP7_75t_L g793 ( .A1(n_79), .A2(n_170), .B1(n_392), .B2(n_569), .Y(n_793) );
AOI22xp5_ASAP7_75t_SL g746 ( .A1(n_80), .A2(n_145), .B1(n_324), .B2(n_698), .Y(n_746) );
CKINVDCx20_ASAP7_75t_R g624 ( .A(n_81), .Y(n_624) );
INVx1_ASAP7_75t_L g424 ( .A(n_82), .Y(n_424) );
AO22x2_ASAP7_75t_L g614 ( .A1(n_83), .A2(n_615), .B1(n_638), .B2(n_639), .Y(n_614) );
CKINVDCx20_ASAP7_75t_R g639 ( .A(n_83), .Y(n_639) );
AOI22xp33_ASAP7_75t_L g634 ( .A1(n_84), .A2(n_236), .B1(n_362), .B2(n_482), .Y(n_634) );
AOI22xp33_ASAP7_75t_L g759 ( .A1(n_85), .A2(n_224), .B1(n_343), .B2(n_517), .Y(n_759) );
CKINVDCx20_ASAP7_75t_R g833 ( .A(n_86), .Y(n_833) );
AOI211xp5_ASAP7_75t_L g831 ( .A1(n_87), .A2(n_522), .B(n_832), .C(n_836), .Y(n_831) );
CKINVDCx20_ASAP7_75t_R g886 ( .A(n_88), .Y(n_886) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_89), .A2(n_225), .B1(n_516), .B2(n_518), .Y(n_515) );
AOI22xp33_ASAP7_75t_L g806 ( .A1(n_92), .A2(n_151), .B1(n_304), .B2(n_485), .Y(n_806) );
INVx1_ASAP7_75t_L g703 ( .A(n_93), .Y(n_703) );
CKINVDCx20_ASAP7_75t_R g541 ( .A(n_95), .Y(n_541) );
AOI222xp33_ASAP7_75t_L g585 ( .A1(n_96), .A2(n_117), .B1(n_137), .B2(n_405), .C1(n_426), .C2(n_430), .Y(n_585) );
INVx1_ASAP7_75t_L g419 ( .A(n_98), .Y(n_419) );
AOI22xp33_ASAP7_75t_L g810 ( .A1(n_99), .A2(n_200), .B1(n_360), .B2(n_365), .Y(n_810) );
CKINVDCx20_ASAP7_75t_R g380 ( .A(n_100), .Y(n_380) );
INVx1_ASAP7_75t_L g294 ( .A(n_101), .Y(n_294) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_102), .A2(n_140), .B1(n_510), .B2(n_513), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g731 ( .A1(n_104), .A2(n_154), .B1(n_446), .B2(n_485), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_105), .B(n_678), .Y(n_677) );
AOI22xp5_ASAP7_75t_L g807 ( .A1(n_107), .A2(n_199), .B1(n_356), .B2(n_386), .Y(n_807) );
AOI22xp33_ASAP7_75t_SL g445 ( .A1(n_108), .A2(n_141), .B1(n_446), .B2(n_449), .Y(n_445) );
INVx1_ASAP7_75t_L g292 ( .A(n_109), .Y(n_292) );
AOI22xp33_ASAP7_75t_SL g471 ( .A1(n_110), .A2(n_149), .B1(n_371), .B2(n_378), .Y(n_471) );
AOI22xp33_ASAP7_75t_SL g809 ( .A1(n_111), .A2(n_171), .B1(n_389), .B2(n_392), .Y(n_809) );
AOI22xp33_ASAP7_75t_L g843 ( .A1(n_112), .A2(n_201), .B1(n_510), .B2(n_513), .Y(n_843) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_113), .B(n_342), .Y(n_689) );
INVx1_ASAP7_75t_L g536 ( .A(n_116), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g344 ( .A1(n_118), .A2(n_157), .B1(n_345), .B2(n_350), .Y(n_344) );
AOI22xp33_ASAP7_75t_L g393 ( .A1(n_119), .A2(n_244), .B1(n_319), .B2(n_394), .Y(n_393) );
CKINVDCx20_ASAP7_75t_R g760 ( .A(n_122), .Y(n_760) );
INVx1_ASAP7_75t_L g672 ( .A(n_123), .Y(n_672) );
INVx1_ASAP7_75t_L g681 ( .A(n_124), .Y(n_681) );
AOI22xp33_ASAP7_75t_L g736 ( .A1(n_125), .A2(n_206), .B1(n_394), .B2(n_737), .Y(n_736) );
XNOR2xp5_ASAP7_75t_L g590 ( .A(n_126), .B(n_591), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_127), .B(n_600), .Y(n_599) );
AOI22xp5_ASAP7_75t_L g649 ( .A1(n_128), .A2(n_650), .B1(n_682), .B2(n_683), .Y(n_649) );
CKINVDCx16_ASAP7_75t_R g682 ( .A(n_128), .Y(n_682) );
INVx1_ASAP7_75t_L g577 ( .A(n_130), .Y(n_577) );
INVx1_ASAP7_75t_L g562 ( .A(n_132), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g388 ( .A1(n_133), .A2(n_237), .B1(n_365), .B2(n_389), .Y(n_388) );
AOI22xp5_ASAP7_75t_SL g411 ( .A1(n_134), .A2(n_412), .B1(n_462), .B2(n_463), .Y(n_411) );
INVx1_ASAP7_75t_L g463 ( .A(n_134), .Y(n_463) );
AOI221xp5_ASAP7_75t_L g568 ( .A1(n_136), .A2(n_194), .B1(n_324), .B2(n_569), .C(n_570), .Y(n_568) );
AOI22xp5_ASAP7_75t_L g756 ( .A1(n_138), .A2(n_185), .B1(n_351), .B2(n_377), .Y(n_756) );
AOI22xp33_ASAP7_75t_L g835 ( .A1(n_142), .A2(n_211), .B1(n_520), .B2(n_604), .Y(n_835) );
CKINVDCx20_ASAP7_75t_R g407 ( .A(n_146), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g834 ( .A(n_147), .B(n_338), .Y(n_834) );
INVx2_ASAP7_75t_L g295 ( .A(n_148), .Y(n_295) );
AOI22xp33_ASAP7_75t_SL g596 ( .A1(n_153), .A2(n_222), .B1(n_426), .B2(n_597), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g519 ( .A1(n_155), .A2(n_234), .B1(n_351), .B2(n_520), .Y(n_519) );
CKINVDCx20_ASAP7_75t_R g837 ( .A(n_156), .Y(n_837) );
AND2x6_ASAP7_75t_L g291 ( .A(n_159), .B(n_292), .Y(n_291) );
HB1xp67_ASAP7_75t_L g820 ( .A(n_159), .Y(n_820) );
AO22x2_ASAP7_75t_L g307 ( .A1(n_160), .A2(n_233), .B1(n_308), .B2(n_309), .Y(n_307) );
AOI22xp33_ASAP7_75t_L g664 ( .A1(n_163), .A2(n_247), .B1(n_665), .B2(n_667), .Y(n_664) );
AOI22xp33_ASAP7_75t_L g384 ( .A1(n_165), .A2(n_257), .B1(n_385), .B2(n_386), .Y(n_384) );
AOI22xp33_ASAP7_75t_L g323 ( .A1(n_167), .A2(n_198), .B1(n_324), .B2(n_332), .Y(n_323) );
INVx1_ASAP7_75t_L g415 ( .A(n_168), .Y(n_415) );
CKINVDCx20_ASAP7_75t_R g539 ( .A(n_172), .Y(n_539) );
CKINVDCx20_ASAP7_75t_R g550 ( .A(n_173), .Y(n_550) );
CKINVDCx20_ASAP7_75t_R g396 ( .A(n_174), .Y(n_396) );
AOI22xp33_ASAP7_75t_SL g701 ( .A1(n_175), .A2(n_263), .B1(n_386), .B2(n_501), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_176), .B(n_524), .Y(n_724) );
CKINVDCx20_ASAP7_75t_R g811 ( .A(n_178), .Y(n_811) );
INVx1_ASAP7_75t_L g438 ( .A(n_179), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g452 ( .A1(n_181), .A2(n_204), .B1(n_392), .B2(n_453), .Y(n_452) );
AOI22xp33_ASAP7_75t_L g636 ( .A1(n_182), .A2(n_262), .B1(n_319), .B2(n_637), .Y(n_636) );
AOI22xp33_ASAP7_75t_SL g484 ( .A1(n_183), .A2(n_254), .B1(n_304), .B2(n_485), .Y(n_484) );
AO22x1_ASAP7_75t_L g570 ( .A1(n_184), .A2(n_227), .B1(n_458), .B2(n_571), .Y(n_570) );
AOI22xp5_ASAP7_75t_L g881 ( .A1(n_186), .A2(n_212), .B1(n_334), .B2(n_481), .Y(n_881) );
CKINVDCx20_ASAP7_75t_R g488 ( .A(n_188), .Y(n_488) );
AO22x2_ASAP7_75t_L g312 ( .A1(n_189), .A2(n_250), .B1(n_308), .B2(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g428 ( .A(n_190), .Y(n_428) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_192), .A2(n_256), .B1(n_375), .B2(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g533 ( .A(n_196), .Y(n_533) );
INVx1_ASAP7_75t_L g851 ( .A(n_197), .Y(n_851) );
CKINVDCx20_ASAP7_75t_R g873 ( .A(n_202), .Y(n_873) );
AOI22xp5_ASAP7_75t_L g694 ( .A1(n_203), .A2(n_279), .B1(n_431), .B2(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g558 ( .A(n_205), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_207), .B(n_400), .Y(n_688) );
AOI22xp33_ASAP7_75t_SL g486 ( .A1(n_209), .A2(n_255), .B1(n_324), .B2(n_487), .Y(n_486) );
AOI22xp33_ASAP7_75t_SL g610 ( .A1(n_210), .A2(n_232), .B1(n_456), .B2(n_611), .Y(n_610) );
AOI22xp33_ASAP7_75t_L g502 ( .A1(n_213), .A2(n_284), .B1(n_503), .B2(n_505), .Y(n_502) );
CKINVDCx20_ASAP7_75t_R g723 ( .A(n_214), .Y(n_723) );
NAND2xp5_ASAP7_75t_SL g546 ( .A(n_215), .B(n_547), .Y(n_546) );
INVx1_ASAP7_75t_L g779 ( .A(n_216), .Y(n_779) );
AOI22xp33_ASAP7_75t_L g361 ( .A1(n_218), .A2(n_251), .B1(n_362), .B2(n_365), .Y(n_361) );
INVx1_ASAP7_75t_L g676 ( .A(n_219), .Y(n_676) );
CKINVDCx20_ASAP7_75t_R g871 ( .A(n_221), .Y(n_871) );
CKINVDCx20_ASAP7_75t_R g631 ( .A(n_223), .Y(n_631) );
CKINVDCx20_ASAP7_75t_R g892 ( .A(n_226), .Y(n_892) );
CKINVDCx20_ASAP7_75t_R g848 ( .A(n_228), .Y(n_848) );
AOI22xp33_ASAP7_75t_SL g699 ( .A1(n_229), .A2(n_238), .B1(n_394), .B2(n_700), .Y(n_699) );
CKINVDCx20_ASAP7_75t_R g726 ( .A(n_230), .Y(n_726) );
INVx1_ASAP7_75t_L g775 ( .A(n_231), .Y(n_775) );
NOR2xp33_ASAP7_75t_L g824 ( .A(n_233), .B(n_825), .Y(n_824) );
NAND2xp5_ASAP7_75t_SL g473 ( .A(n_235), .B(n_342), .Y(n_473) );
AOI22xp33_ASAP7_75t_L g732 ( .A1(n_240), .A2(n_281), .B1(n_569), .B2(n_733), .Y(n_732) );
CKINVDCx20_ASAP7_75t_R g555 ( .A(n_241), .Y(n_555) );
AOI22xp33_ASAP7_75t_L g337 ( .A1(n_242), .A2(n_259), .B1(n_338), .B2(n_342), .Y(n_337) );
CKINVDCx20_ASAP7_75t_R g621 ( .A(n_243), .Y(n_621) );
INVx1_ASAP7_75t_L g433 ( .A(n_245), .Y(n_433) );
INVx1_ASAP7_75t_L g680 ( .A(n_246), .Y(n_680) );
INVx1_ASAP7_75t_L g575 ( .A(n_248), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g739 ( .A1(n_249), .A2(n_265), .B1(n_740), .B2(n_741), .Y(n_739) );
INVx1_ASAP7_75t_L g823 ( .A(n_250), .Y(n_823) );
AOI22xp33_ASAP7_75t_SL g782 ( .A1(n_252), .A2(n_253), .B1(n_783), .B2(n_784), .Y(n_782) );
INVx1_ASAP7_75t_L g656 ( .A(n_258), .Y(n_656) );
OA22x2_ASAP7_75t_L g710 ( .A1(n_264), .A2(n_711), .B1(n_712), .B2(n_742), .Y(n_710) );
INVx1_ASAP7_75t_L g711 ( .A(n_264), .Y(n_711) );
CKINVDCx20_ASAP7_75t_R g884 ( .A(n_266), .Y(n_884) );
CKINVDCx20_ASAP7_75t_R g582 ( .A(n_267), .Y(n_582) );
INVx1_ASAP7_75t_L g308 ( .A(n_268), .Y(n_308) );
INVx1_ASAP7_75t_L g310 ( .A(n_268), .Y(n_310) );
CKINVDCx20_ASAP7_75t_R g595 ( .A(n_270), .Y(n_595) );
INVx1_ASAP7_75t_L g772 ( .A(n_271), .Y(n_772) );
CKINVDCx20_ASAP7_75t_R g878 ( .A(n_272), .Y(n_878) );
INVx1_ASAP7_75t_L g674 ( .A(n_273), .Y(n_674) );
INVx1_ASAP7_75t_L g771 ( .A(n_274), .Y(n_771) );
AOI22xp33_ASAP7_75t_L g776 ( .A1(n_275), .A2(n_285), .B1(n_371), .B2(n_597), .Y(n_776) );
INVx1_ASAP7_75t_L g862 ( .A(n_276), .Y(n_862) );
OA22x2_ASAP7_75t_L g865 ( .A1(n_276), .A2(n_862), .B1(n_866), .B2(n_867), .Y(n_865) );
OA22x2_ASAP7_75t_L g493 ( .A1(n_278), .A2(n_494), .B1(n_495), .B2(n_525), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_278), .Y(n_494) );
INVx1_ASAP7_75t_L g778 ( .A(n_280), .Y(n_778) );
CKINVDCx20_ASAP7_75t_R g798 ( .A(n_282), .Y(n_798) );
CKINVDCx20_ASAP7_75t_R g717 ( .A(n_283), .Y(n_717) );
CKINVDCx20_ASAP7_75t_R g287 ( .A(n_288), .Y(n_287) );
CKINVDCx20_ASAP7_75t_R g288 ( .A(n_289), .Y(n_288) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AND2x4_ASAP7_75t_L g290 ( .A(n_291), .B(n_293), .Y(n_290) );
HB1xp67_ASAP7_75t_L g819 ( .A(n_292), .Y(n_819) );
OAI21xp5_ASAP7_75t_L g860 ( .A1(n_293), .A2(n_818), .B(n_861), .Y(n_860) );
AND2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_295), .Y(n_293) );
AOI221xp5_ASAP7_75t_L g296 ( .A1(n_297), .A2(n_491), .B1(n_813), .B2(n_814), .C(n_815), .Y(n_296) );
INVxp67_ASAP7_75t_L g814 ( .A(n_297), .Y(n_814) );
AOI22xp5_ASAP7_75t_SL g297 ( .A1(n_298), .A2(n_299), .B1(n_410), .B2(n_490), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
AO22x1_ASAP7_75t_SL g299 ( .A1(n_300), .A2(n_381), .B1(n_408), .B2(n_409), .Y(n_299) );
INVx2_ASAP7_75t_SL g408 ( .A(n_300), .Y(n_408) );
XOR2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_380), .Y(n_300) );
NAND4xp75_ASAP7_75t_L g301 ( .A(n_302), .B(n_336), .C(n_354), .D(n_367), .Y(n_301) );
AND2x2_ASAP7_75t_L g302 ( .A(n_303), .B(n_323), .Y(n_302) );
BUFx3_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
BUFx3_ASAP7_75t_L g448 ( .A(n_305), .Y(n_448) );
BUFx3_ASAP7_75t_L g501 ( .A(n_305), .Y(n_501) );
AND2x2_ASAP7_75t_L g305 ( .A(n_306), .B(n_314), .Y(n_305) );
AND2x2_ASAP7_75t_L g364 ( .A(n_306), .B(n_335), .Y(n_364) );
NAND2xp5_ASAP7_75t_SL g556 ( .A(n_306), .B(n_335), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_306), .B(n_314), .Y(n_559) );
AND2x2_ASAP7_75t_L g306 ( .A(n_307), .B(n_311), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_307), .B(n_312), .Y(n_322) );
INVx2_ASAP7_75t_L g330 ( .A(n_307), .Y(n_330) );
AND2x2_ASAP7_75t_L g349 ( .A(n_307), .B(n_316), .Y(n_349) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g313 ( .A(n_310), .Y(n_313) );
INVx1_ASAP7_75t_L g352 ( .A(n_311), .Y(n_352) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g331 ( .A(n_312), .Y(n_331) );
AND2x2_ASAP7_75t_L g341 ( .A(n_312), .B(n_330), .Y(n_341) );
INVx1_ASAP7_75t_L g374 ( .A(n_312), .Y(n_374) );
AND2x4_ASAP7_75t_L g320 ( .A(n_314), .B(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g358 ( .A(n_314), .B(n_329), .Y(n_358) );
AND2x4_ASAP7_75t_L g360 ( .A(n_314), .B(n_341), .Y(n_360) );
AND2x2_ASAP7_75t_L g314 ( .A(n_315), .B(n_317), .Y(n_314) );
OR2x2_ASAP7_75t_L g328 ( .A(n_315), .B(n_318), .Y(n_328) );
AND2x2_ASAP7_75t_L g335 ( .A(n_315), .B(n_318), .Y(n_335) );
INVx2_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g353 ( .A(n_316), .B(n_318), .Y(n_353) );
AND2x2_ASAP7_75t_L g373 ( .A(n_317), .B(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g437 ( .A(n_317), .Y(n_437) );
INVx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g348 ( .A(n_318), .Y(n_348) );
BUFx3_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
BUFx3_ASAP7_75t_L g451 ( .A(n_320), .Y(n_451) );
BUFx3_ASAP7_75t_L g485 ( .A(n_320), .Y(n_485) );
BUFx2_ASAP7_75t_L g513 ( .A(n_320), .Y(n_513) );
INVx1_ASAP7_75t_L g554 ( .A(n_320), .Y(n_554) );
BUFx3_ASAP7_75t_L g658 ( .A(n_320), .Y(n_658) );
BUFx2_ASAP7_75t_SL g784 ( .A(n_320), .Y(n_784) );
BUFx2_ASAP7_75t_SL g888 ( .A(n_320), .Y(n_888) );
AND2x2_ASAP7_75t_L g547 ( .A(n_321), .B(n_437), .Y(n_547) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
OR2x6_ASAP7_75t_L g366 ( .A(n_322), .B(n_348), .Y(n_366) );
INVx1_ASAP7_75t_L g847 ( .A(n_324), .Y(n_847) );
INVx3_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx2_ASAP7_75t_SL g508 ( .A(n_325), .Y(n_508) );
INVx11_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx11_ASAP7_75t_L g387 ( .A(n_326), .Y(n_387) );
AND2x6_ASAP7_75t_L g326 ( .A(n_327), .B(n_329), .Y(n_326) );
AND2x4_ASAP7_75t_L g340 ( .A(n_327), .B(n_341), .Y(n_340) );
INVx2_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
OR2x2_ASAP7_75t_L g417 ( .A(n_328), .B(n_418), .Y(n_417) );
AND2x4_ASAP7_75t_L g334 ( .A(n_329), .B(n_335), .Y(n_334) );
AND2x6_ASAP7_75t_L g370 ( .A(n_329), .B(n_353), .Y(n_370) );
AND2x2_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
INVx2_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx3_ASAP7_75t_L g392 ( .A(n_333), .Y(n_392) );
INVx2_ASAP7_75t_L g498 ( .A(n_333), .Y(n_498) );
OAI22xp5_ASAP7_75t_SL g548 ( .A1(n_333), .A2(n_357), .B1(n_549), .B2(n_550), .Y(n_548) );
OAI221xp5_ASAP7_75t_SL g659 ( .A1(n_333), .A2(n_660), .B1(n_661), .B2(n_663), .C(n_664), .Y(n_659) );
OAI22xp5_ASAP7_75t_L g845 ( .A1(n_333), .A2(n_846), .B1(n_847), .B2(n_848), .Y(n_845) );
INVx6_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
BUFx3_ASAP7_75t_L g487 ( .A(n_334), .Y(n_487) );
BUFx3_ASAP7_75t_L g608 ( .A(n_334), .Y(n_608) );
AND2x6_ASAP7_75t_L g343 ( .A(n_335), .B(n_341), .Y(n_343) );
NAND2x1p5_ASAP7_75t_L g398 ( .A(n_335), .B(n_341), .Y(n_398) );
AND2x2_ASAP7_75t_SL g336 ( .A(n_337), .B(n_344), .Y(n_336) );
INVx2_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx2_ASAP7_75t_L g400 ( .A(n_339), .Y(n_400) );
INVx2_ASAP7_75t_L g475 ( .A(n_339), .Y(n_475) );
INVx5_ASAP7_75t_L g517 ( .A(n_339), .Y(n_517) );
INVx4_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g418 ( .A(n_341), .Y(n_418) );
INVx1_ASAP7_75t_L g601 ( .A(n_342), .Y(n_601) );
BUFx4f_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
BUFx2_ASAP7_75t_L g518 ( .A(n_343), .Y(n_518) );
BUFx2_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
BUFx3_ASAP7_75t_L g402 ( .A(n_346), .Y(n_402) );
BUFx2_ASAP7_75t_L g520 ( .A(n_346), .Y(n_520) );
AND2x4_ASAP7_75t_L g346 ( .A(n_347), .B(n_349), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
AND2x4_ASAP7_75t_L g372 ( .A(n_349), .B(n_373), .Y(n_372) );
AND2x4_ASAP7_75t_L g378 ( .A(n_349), .B(n_379), .Y(n_378) );
NAND2x1p5_ASAP7_75t_L g436 ( .A(n_349), .B(n_437), .Y(n_436) );
BUFx3_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
BUFx6f_ASAP7_75t_L g403 ( .A(n_351), .Y(n_403) );
BUFx2_ASAP7_75t_SL g695 ( .A(n_351), .Y(n_695) );
BUFx2_ASAP7_75t_SL g800 ( .A(n_351), .Y(n_800) );
AND2x4_ASAP7_75t_L g351 ( .A(n_352), .B(n_353), .Y(n_351) );
INVx1_ASAP7_75t_L g442 ( .A(n_352), .Y(n_442) );
INVx1_ASAP7_75t_L g441 ( .A(n_353), .Y(n_441) );
AND2x2_ASAP7_75t_L g354 ( .A(n_355), .B(n_361), .Y(n_354) );
INVx3_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx3_ASAP7_75t_L g385 ( .A(n_357), .Y(n_385) );
INVx2_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
BUFx6f_ASAP7_75t_L g457 ( .A(n_358), .Y(n_457) );
BUFx2_ASAP7_75t_SL g748 ( .A(n_358), .Y(n_748) );
BUFx3_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
BUFx3_ASAP7_75t_L g394 ( .A(n_360), .Y(n_394) );
BUFx3_ASAP7_75t_L g479 ( .A(n_360), .Y(n_479) );
BUFx6f_ASAP7_75t_L g512 ( .A(n_360), .Y(n_512) );
INVx2_ASAP7_75t_L g544 ( .A(n_360), .Y(n_544) );
INVx2_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx5_ASAP7_75t_L g389 ( .A(n_363), .Y(n_389) );
INVx1_ASAP7_75t_L g481 ( .A(n_363), .Y(n_481) );
INVx4_ASAP7_75t_L g504 ( .A(n_363), .Y(n_504) );
BUFx3_ASAP7_75t_L g666 ( .A(n_363), .Y(n_666) );
INVx3_ASAP7_75t_L g698 ( .A(n_363), .Y(n_698) );
INVx8_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
BUFx4f_ASAP7_75t_SL g461 ( .A(n_365), .Y(n_461) );
BUFx2_ASAP7_75t_L g482 ( .A(n_365), .Y(n_482) );
BUFx2_ASAP7_75t_L g505 ( .A(n_365), .Y(n_505) );
BUFx2_ASAP7_75t_L g788 ( .A(n_365), .Y(n_788) );
INVx6_ASAP7_75t_SL g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_SL g667 ( .A(n_366), .Y(n_667) );
INVx1_ASAP7_75t_SL g700 ( .A(n_366), .Y(n_700) );
INVx1_ASAP7_75t_L g741 ( .A(n_366), .Y(n_741) );
INVx4_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
BUFx2_ASAP7_75t_L g721 ( .A(n_369), .Y(n_721) );
INVx4_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
BUFx6f_ASAP7_75t_L g405 ( .A(n_370), .Y(n_405) );
INVx2_ASAP7_75t_L g469 ( .A(n_370), .Y(n_469) );
BUFx3_ASAP7_75t_L g522 ( .A(n_370), .Y(n_522) );
INVx2_ASAP7_75t_SL g540 ( .A(n_370), .Y(n_540) );
INVx2_ASAP7_75t_L g755 ( .A(n_370), .Y(n_755) );
INVx4_ASAP7_75t_L g427 ( .A(n_371), .Y(n_427) );
BUFx6f_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
BUFx6f_ASAP7_75t_L g406 ( .A(n_372), .Y(n_406) );
BUFx4f_ASAP7_75t_SL g523 ( .A(n_372), .Y(n_523) );
BUFx2_ASAP7_75t_L g627 ( .A(n_372), .Y(n_627) );
BUFx6f_ASAP7_75t_L g691 ( .A(n_372), .Y(n_691) );
INVx1_ASAP7_75t_L g379 ( .A(n_374), .Y(n_379) );
INVx1_ASAP7_75t_L g840 ( .A(n_375), .Y(n_840) );
INVx3_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
BUFx4f_ASAP7_75t_SL g524 ( .A(n_377), .Y(n_524) );
BUFx12f_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
BUFx6f_ASAP7_75t_L g431 ( .A(n_378), .Y(n_431) );
BUFx6f_ASAP7_75t_L g597 ( .A(n_378), .Y(n_597) );
INVx2_ASAP7_75t_SL g409 ( .A(n_381), .Y(n_409) );
XOR2x2_ASAP7_75t_L g381 ( .A(n_382), .B(n_407), .Y(n_381) );
NAND4xp75_ASAP7_75t_L g382 ( .A(n_383), .B(n_390), .C(n_395), .D(n_404), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_384), .B(n_388), .Y(n_383) );
INVx1_ASAP7_75t_L g792 ( .A(n_386), .Y(n_792) );
INVx5_ASAP7_75t_SL g386 ( .A(n_387), .Y(n_386) );
INVx2_ASAP7_75t_L g453 ( .A(n_387), .Y(n_453) );
NOR2xp33_ASAP7_75t_L g560 ( .A(n_387), .B(n_561), .Y(n_560) );
INVx4_ASAP7_75t_L g611 ( .A(n_387), .Y(n_611) );
INVx2_ASAP7_75t_SL g637 ( .A(n_387), .Y(n_637) );
INVx1_ASAP7_75t_L g891 ( .A(n_387), .Y(n_891) );
BUFx6f_ASAP7_75t_L g460 ( .A(n_389), .Y(n_460) );
BUFx2_ASAP7_75t_L g740 ( .A(n_389), .Y(n_740) );
AND2x2_ASAP7_75t_L g390 ( .A(n_391), .B(n_393), .Y(n_390) );
BUFx2_ASAP7_75t_L g458 ( .A(n_394), .Y(n_458) );
OA211x2_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_397), .B(n_399), .C(n_401), .Y(n_395) );
OAI22xp5_ASAP7_75t_L g535 ( .A1(n_397), .A2(n_436), .B1(n_536), .B2(n_537), .Y(n_535) );
OAI22xp5_ASAP7_75t_L g669 ( .A1(n_397), .A2(n_670), .B1(n_671), .B2(n_672), .Y(n_669) );
INVx2_ASAP7_75t_L g719 ( .A(n_397), .Y(n_719) );
BUFx3_ASAP7_75t_L g773 ( .A(n_397), .Y(n_773) );
BUFx3_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g421 ( .A(n_398), .Y(n_421) );
INVx1_ASAP7_75t_SL g605 ( .A(n_403), .Y(n_605) );
INVx2_ASAP7_75t_SL g423 ( .A(n_405), .Y(n_423) );
INVx2_ASAP7_75t_L g594 ( .A(n_405), .Y(n_594) );
CKINVDCx20_ASAP7_75t_R g877 ( .A(n_406), .Y(n_877) );
INVx2_ASAP7_75t_SL g490 ( .A(n_410), .Y(n_490) );
OA22x2_ASAP7_75t_L g410 ( .A1(n_411), .A2(n_464), .B1(n_465), .B2(n_489), .Y(n_410) );
INVx1_ASAP7_75t_L g489 ( .A(n_411), .Y(n_489) );
INVx2_ASAP7_75t_SL g462 ( .A(n_412), .Y(n_462) );
AND2x2_ASAP7_75t_L g412 ( .A(n_413), .B(n_443), .Y(n_412) );
NOR3xp33_ASAP7_75t_L g413 ( .A(n_414), .B(n_422), .C(n_432), .Y(n_413) );
OAI22xp5_ASAP7_75t_L g414 ( .A1(n_415), .A2(n_416), .B1(n_419), .B2(n_420), .Y(n_414) );
BUFx6f_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
OAI21xp5_ASAP7_75t_L g532 ( .A1(n_417), .A2(n_533), .B(n_534), .Y(n_532) );
INVx2_ASAP7_75t_L g620 ( .A(n_417), .Y(n_620) );
INVx1_ASAP7_75t_SL g420 ( .A(n_421), .Y(n_420) );
INVx2_ASAP7_75t_L g622 ( .A(n_421), .Y(n_622) );
OAI221xp5_ASAP7_75t_L g422 ( .A1(n_423), .A2(n_424), .B1(n_425), .B2(n_428), .C(n_429), .Y(n_422) );
OAI221xp5_ASAP7_75t_SL g673 ( .A1(n_423), .A2(n_674), .B1(n_675), .B2(n_676), .C(n_677), .Y(n_673) );
OAI21xp33_ASAP7_75t_SL g774 ( .A1(n_423), .A2(n_775), .B(n_776), .Y(n_774) );
OAI221xp5_ASAP7_75t_L g720 ( .A1(n_425), .A2(n_721), .B1(n_722), .B2(n_723), .C(n_724), .Y(n_720) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx3_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
OAI22xp5_ASAP7_75t_L g538 ( .A1(n_427), .A2(n_539), .B1(n_540), .B2(n_541), .Y(n_538) );
BUFx3_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
OAI22xp5_ASAP7_75t_L g432 ( .A1(n_433), .A2(n_434), .B1(n_438), .B2(n_439), .Y(n_432) );
INVx3_ASAP7_75t_SL g434 ( .A(n_435), .Y(n_434) );
INVx2_ASAP7_75t_L g630 ( .A(n_435), .Y(n_630) );
INVx4_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
OAI22xp5_ASAP7_75t_L g580 ( .A1(n_436), .A2(n_581), .B1(n_582), .B2(n_583), .Y(n_580) );
BUFx3_ASAP7_75t_L g727 ( .A(n_436), .Y(n_727) );
OAI22xp5_ASAP7_75t_L g777 ( .A1(n_436), .A2(n_439), .B1(n_778), .B2(n_779), .Y(n_777) );
OAI22xp5_ASAP7_75t_L g725 ( .A1(n_439), .A2(n_726), .B1(n_727), .B2(n_728), .Y(n_725) );
BUFx2_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
CKINVDCx16_ASAP7_75t_R g584 ( .A(n_440), .Y(n_584) );
OAI22xp5_ASAP7_75t_L g628 ( .A1(n_440), .A2(n_629), .B1(n_630), .B2(n_631), .Y(n_628) );
OR2x6_ASAP7_75t_L g440 ( .A(n_441), .B(n_442), .Y(n_440) );
NOR2xp33_ASAP7_75t_L g443 ( .A(n_444), .B(n_454), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_445), .B(n_452), .Y(n_444) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
BUFx4f_ASAP7_75t_SL g783 ( .A(n_448), .Y(n_783) );
INVx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
HB1xp67_ASAP7_75t_L g571 ( .A(n_451), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_455), .B(n_459), .Y(n_454) );
BUFx3_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
BUFx6f_ASAP7_75t_L g569 ( .A(n_457), .Y(n_569) );
CKINVDCx20_ASAP7_75t_R g578 ( .A(n_461), .Y(n_578) );
INVx4_ASAP7_75t_SL g464 ( .A(n_465), .Y(n_464) );
XOR2x2_ASAP7_75t_L g465 ( .A(n_466), .B(n_488), .Y(n_465) );
NAND3x1_ASAP7_75t_L g466 ( .A(n_467), .B(n_477), .C(n_483), .Y(n_466) );
NOR2xp33_ASAP7_75t_L g467 ( .A(n_468), .B(n_472), .Y(n_467) );
OAI21xp5_ASAP7_75t_SL g468 ( .A1(n_469), .A2(n_470), .B(n_471), .Y(n_468) );
OAI21xp5_ASAP7_75t_L g692 ( .A1(n_469), .A2(n_693), .B(n_694), .Y(n_692) );
OAI21xp5_ASAP7_75t_L g797 ( .A1(n_469), .A2(n_798), .B(n_799), .Y(n_797) );
NAND3xp33_ASAP7_75t_L g472 ( .A(n_473), .B(n_474), .C(n_476), .Y(n_472) );
AND2x2_ASAP7_75t_L g477 ( .A(n_478), .B(n_480), .Y(n_477) );
AND2x2_ASAP7_75t_L g483 ( .A(n_484), .B(n_486), .Y(n_483) );
INVx1_ASAP7_75t_L g813 ( .A(n_491), .Y(n_813) );
XOR2xp5_ASAP7_75t_L g491 ( .A(n_492), .B(n_644), .Y(n_491) );
AOI22xp5_ASAP7_75t_L g492 ( .A1(n_493), .A2(n_526), .B1(n_642), .B2(n_643), .Y(n_492) );
INVx1_ASAP7_75t_L g642 ( .A(n_493), .Y(n_642) );
INVx1_ASAP7_75t_SL g525 ( .A(n_495), .Y(n_525) );
NAND4xp75_ASAP7_75t_L g495 ( .A(n_496), .B(n_506), .C(n_514), .D(n_521), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_497), .B(n_502), .Y(n_496) );
INVx2_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
BUFx2_ASAP7_75t_L g573 ( .A(n_501), .Y(n_573) );
BUFx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx2_ASAP7_75t_L g787 ( .A(n_504), .Y(n_787) );
AND2x2_ASAP7_75t_L g506 ( .A(n_507), .B(n_509), .Y(n_506) );
INVx1_ASAP7_75t_L g655 ( .A(n_508), .Y(n_655) );
INVx3_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx4_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
AND2x2_ASAP7_75t_SL g514 ( .A(n_515), .B(n_519), .Y(n_514) );
BUFx6f_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx3_ASAP7_75t_L g625 ( .A(n_522), .Y(n_625) );
INVx1_ASAP7_75t_L g643 ( .A(n_526), .Y(n_643) );
AOI22xp5_ASAP7_75t_L g526 ( .A1(n_527), .A2(n_528), .B1(n_563), .B2(n_641), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
BUFx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
XNOR2x1_ASAP7_75t_L g529 ( .A(n_530), .B(n_562), .Y(n_529) );
AND3x2_ASAP7_75t_L g530 ( .A(n_531), .B(n_542), .C(n_551), .Y(n_530) );
NOR3xp33_ASAP7_75t_L g531 ( .A(n_532), .B(n_535), .C(n_538), .Y(n_531) );
NOR2xp33_ASAP7_75t_L g542 ( .A(n_543), .B(n_548), .Y(n_542) );
OAI21xp5_ASAP7_75t_SL g543 ( .A1(n_544), .A2(n_545), .B(n_546), .Y(n_543) );
NOR3xp33_ASAP7_75t_L g551 ( .A(n_552), .B(n_557), .C(n_560), .Y(n_551) );
OAI22xp5_ASAP7_75t_L g552 ( .A1(n_553), .A2(n_554), .B1(n_555), .B2(n_556), .Y(n_552) );
BUFx2_ASAP7_75t_R g576 ( .A(n_556), .Y(n_576) );
NOR2xp33_ASAP7_75t_L g557 ( .A(n_558), .B(n_559), .Y(n_557) );
INVx1_ASAP7_75t_L g662 ( .A(n_559), .Y(n_662) );
INVx1_ASAP7_75t_L g641 ( .A(n_563), .Y(n_641) );
AOI22xp5_ASAP7_75t_L g563 ( .A1(n_564), .A2(n_587), .B1(n_588), .B2(n_640), .Y(n_563) );
INVx1_ASAP7_75t_L g640 ( .A(n_564), .Y(n_640) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
AND4x1_ASAP7_75t_L g567 ( .A(n_568), .B(n_572), .C(n_579), .D(n_585), .Y(n_567) );
INVx1_ASAP7_75t_SL g653 ( .A(n_569), .Y(n_653) );
OAI22xp5_ASAP7_75t_L g574 ( .A1(n_575), .A2(n_576), .B1(n_577), .B2(n_578), .Y(n_574) );
OAI22xp5_ASAP7_75t_L g679 ( .A1(n_583), .A2(n_630), .B1(n_680), .B2(n_681), .Y(n_679) );
INVx2_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx2_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
AO22x1_ASAP7_75t_L g588 ( .A1(n_589), .A2(n_590), .B1(n_613), .B2(n_614), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
NAND4xp75_ASAP7_75t_SL g591 ( .A(n_592), .B(n_606), .C(n_610), .D(n_612), .Y(n_591) );
NOR2xp67_ASAP7_75t_L g592 ( .A(n_593), .B(n_598), .Y(n_592) );
OAI21xp5_ASAP7_75t_SL g593 ( .A1(n_594), .A2(n_595), .B(n_596), .Y(n_593) );
BUFx4f_ASAP7_75t_L g678 ( .A(n_597), .Y(n_678) );
NAND3xp33_ASAP7_75t_L g598 ( .A(n_599), .B(n_602), .C(n_603), .Y(n_598) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
AND2x2_ASAP7_75t_L g606 ( .A(n_607), .B(n_609), .Y(n_606) );
INVx1_ASAP7_75t_L g734 ( .A(n_608), .Y(n_734) );
INVx2_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx1_ASAP7_75t_SL g638 ( .A(n_615), .Y(n_638) );
AND2x2_ASAP7_75t_SL g615 ( .A(n_616), .B(n_632), .Y(n_615) );
NOR3xp33_ASAP7_75t_L g616 ( .A(n_617), .B(n_623), .C(n_628), .Y(n_616) );
OAI22xp5_ASAP7_75t_L g617 ( .A1(n_618), .A2(n_619), .B1(n_621), .B2(n_622), .Y(n_617) );
OAI22xp5_ASAP7_75t_SL g869 ( .A1(n_619), .A2(n_718), .B1(n_870), .B2(n_871), .Y(n_869) );
INVx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx1_ASAP7_75t_SL g671 ( .A(n_620), .Y(n_671) );
INVx2_ASAP7_75t_L g716 ( .A(n_620), .Y(n_716) );
OAI21xp33_ASAP7_75t_L g623 ( .A1(n_624), .A2(n_625), .B(n_626), .Y(n_623) );
OAI21xp33_ASAP7_75t_L g872 ( .A1(n_625), .A2(n_873), .B(n_874), .Y(n_872) );
INVx1_ASAP7_75t_L g675 ( .A(n_627), .Y(n_675) );
AND4x1_ASAP7_75t_L g632 ( .A(n_633), .B(n_634), .C(n_635), .D(n_636), .Y(n_632) );
INVx1_ASAP7_75t_L g738 ( .A(n_637), .Y(n_738) );
OAI22xp5_ASAP7_75t_L g644 ( .A1(n_645), .A2(n_646), .B1(n_706), .B2(n_707), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
OAI22xp5_ASAP7_75t_SL g646 ( .A1(n_647), .A2(n_684), .B1(n_704), .B2(n_705), .Y(n_646) );
INVx1_ASAP7_75t_SL g704 ( .A(n_647), .Y(n_704) );
BUFx2_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g683 ( .A(n_650), .Y(n_683) );
AND2x2_ASAP7_75t_SL g650 ( .A(n_651), .B(n_668), .Y(n_650) );
NOR2xp33_ASAP7_75t_L g651 ( .A(n_652), .B(n_659), .Y(n_651) );
OAI221xp5_ASAP7_75t_SL g652 ( .A1(n_653), .A2(n_654), .B1(n_655), .B2(n_656), .C(n_657), .Y(n_652) );
OAI22xp5_ASAP7_75t_L g849 ( .A1(n_653), .A2(n_661), .B1(n_850), .B2(n_851), .Y(n_849) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g894 ( .A(n_662), .Y(n_894) );
INVx3_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
NOR3xp33_ASAP7_75t_L g668 ( .A(n_669), .B(n_673), .C(n_679), .Y(n_668) );
INVx1_ASAP7_75t_L g705 ( .A(n_684), .Y(n_705) );
XOR2x2_ASAP7_75t_L g684 ( .A(n_685), .B(n_703), .Y(n_684) );
NAND4xp75_ASAP7_75t_SL g685 ( .A(n_686), .B(n_696), .C(n_701), .D(n_702), .Y(n_685) );
NOR2xp67_ASAP7_75t_SL g686 ( .A(n_687), .B(n_692), .Y(n_686) );
NAND3xp33_ASAP7_75t_L g687 ( .A(n_688), .B(n_689), .C(n_690), .Y(n_687) );
INVx1_ASAP7_75t_L g838 ( .A(n_691), .Y(n_838) );
AND2x2_ASAP7_75t_L g696 ( .A(n_697), .B(n_699), .Y(n_696) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
AOI22xp5_ASAP7_75t_L g707 ( .A1(n_708), .A2(n_709), .B1(n_762), .B2(n_763), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
OAI22xp5_ASAP7_75t_L g709 ( .A1(n_710), .A2(n_743), .B1(n_744), .B2(n_761), .Y(n_709) );
INVx1_ASAP7_75t_L g761 ( .A(n_710), .Y(n_761) );
INVx1_ASAP7_75t_L g742 ( .A(n_712), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_713), .B(n_729), .Y(n_712) );
NOR3xp33_ASAP7_75t_L g713 ( .A(n_714), .B(n_720), .C(n_725), .Y(n_713) );
OAI22xp5_ASAP7_75t_L g714 ( .A1(n_715), .A2(n_716), .B1(n_717), .B2(n_718), .Y(n_714) );
OAI22xp5_ASAP7_75t_L g770 ( .A1(n_716), .A2(n_771), .B1(n_772), .B2(n_773), .Y(n_770) );
OAI211xp5_ASAP7_75t_L g832 ( .A1(n_718), .A2(n_833), .B(n_834), .C(n_835), .Y(n_832) );
INVx2_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
OAI22xp33_ASAP7_75t_L g875 ( .A1(n_727), .A2(n_876), .B1(n_877), .B2(n_878), .Y(n_875) );
NOR2xp67_ASAP7_75t_L g729 ( .A(n_730), .B(n_735), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_731), .B(n_732), .Y(n_730) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_736), .B(n_739), .Y(n_735) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx2_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
XOR2x2_ASAP7_75t_L g744 ( .A(n_745), .B(n_760), .Y(n_744) );
NAND4xp75_ASAP7_75t_SL g745 ( .A(n_746), .B(n_747), .C(n_749), .D(n_752), .Y(n_745) );
INVx1_ASAP7_75t_L g885 ( .A(n_748), .Y(n_885) );
AND2x2_ASAP7_75t_L g749 ( .A(n_750), .B(n_751), .Y(n_749) );
NOR2xp33_ASAP7_75t_L g752 ( .A(n_753), .B(n_757), .Y(n_752) );
OAI21xp5_ASAP7_75t_L g753 ( .A1(n_754), .A2(n_755), .B(n_756), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_758), .B(n_759), .Y(n_757) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
AO22x1_ASAP7_75t_L g763 ( .A1(n_764), .A2(n_765), .B1(n_794), .B2(n_812), .Y(n_763) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
INVx1_ASAP7_75t_SL g767 ( .A(n_768), .Y(n_767) );
AND2x2_ASAP7_75t_L g768 ( .A(n_769), .B(n_780), .Y(n_768) );
NOR3xp33_ASAP7_75t_L g769 ( .A(n_770), .B(n_774), .C(n_777), .Y(n_769) );
NOR2xp33_ASAP7_75t_L g780 ( .A(n_781), .B(n_789), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_782), .B(n_785), .Y(n_781) );
INVx3_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_790), .B(n_793), .Y(n_789) );
INVx2_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
INVx3_ASAP7_75t_SL g812 ( .A(n_794), .Y(n_812) );
XOR2x2_ASAP7_75t_L g794 ( .A(n_795), .B(n_811), .Y(n_794) );
NAND2xp5_ASAP7_75t_SL g795 ( .A(n_796), .B(n_804), .Y(n_795) );
NOR2xp33_ASAP7_75t_L g796 ( .A(n_797), .B(n_801), .Y(n_796) );
NAND2xp5_ASAP7_75t_L g801 ( .A(n_802), .B(n_803), .Y(n_801) );
NOR2xp33_ASAP7_75t_L g804 ( .A(n_805), .B(n_808), .Y(n_804) );
NAND2xp5_ASAP7_75t_L g805 ( .A(n_806), .B(n_807), .Y(n_805) );
NAND2xp5_ASAP7_75t_L g808 ( .A(n_809), .B(n_810), .Y(n_808) );
INVx1_ASAP7_75t_SL g815 ( .A(n_816), .Y(n_815) );
NOR2x1_ASAP7_75t_L g816 ( .A(n_817), .B(n_821), .Y(n_816) );
OR2x2_ASAP7_75t_SL g897 ( .A(n_817), .B(n_822), .Y(n_897) );
NAND2xp5_ASAP7_75t_L g817 ( .A(n_818), .B(n_820), .Y(n_817) );
CKINVDCx20_ASAP7_75t_R g856 ( .A(n_818), .Y(n_856) );
INVx1_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g861 ( .A(n_819), .B(n_858), .Y(n_861) );
CKINVDCx16_ASAP7_75t_R g858 ( .A(n_820), .Y(n_858) );
CKINVDCx20_ASAP7_75t_R g821 ( .A(n_822), .Y(n_821) );
NAND2xp5_ASAP7_75t_L g822 ( .A(n_823), .B(n_824), .Y(n_822) );
NAND2xp5_ASAP7_75t_L g825 ( .A(n_826), .B(n_827), .Y(n_825) );
OAI322xp33_ASAP7_75t_L g828 ( .A1(n_829), .A2(n_854), .A3(n_857), .B1(n_859), .B2(n_862), .C1(n_863), .C2(n_895), .Y(n_828) );
INVx1_ASAP7_75t_L g853 ( .A(n_830), .Y(n_853) );
AND2x2_ASAP7_75t_L g830 ( .A(n_831), .B(n_841), .Y(n_830) );
OAI22xp5_ASAP7_75t_L g836 ( .A1(n_837), .A2(n_838), .B1(n_839), .B2(n_840), .Y(n_836) );
NOR3xp33_ASAP7_75t_L g841 ( .A(n_842), .B(n_845), .C(n_849), .Y(n_841) );
NAND2xp5_ASAP7_75t_L g842 ( .A(n_843), .B(n_844), .Y(n_842) );
HB1xp67_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
HB1xp67_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
INVx1_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
CKINVDCx16_ASAP7_75t_R g859 ( .A(n_860), .Y(n_859) );
INVx1_ASAP7_75t_SL g863 ( .A(n_864), .Y(n_863) );
INVx2_ASAP7_75t_L g864 ( .A(n_865), .Y(n_864) );
INVx2_ASAP7_75t_SL g866 ( .A(n_867), .Y(n_866) );
AND2x2_ASAP7_75t_L g867 ( .A(n_868), .B(n_879), .Y(n_867) );
NOR3xp33_ASAP7_75t_L g868 ( .A(n_869), .B(n_872), .C(n_875), .Y(n_868) );
NOR3xp33_ASAP7_75t_L g879 ( .A(n_880), .B(n_883), .C(n_889), .Y(n_879) );
NAND2xp5_ASAP7_75t_L g880 ( .A(n_881), .B(n_882), .Y(n_880) );
OAI22xp5_ASAP7_75t_L g883 ( .A1(n_884), .A2(n_885), .B1(n_886), .B2(n_887), .Y(n_883) );
INVx1_ASAP7_75t_SL g887 ( .A(n_888), .Y(n_887) );
OAI22xp5_ASAP7_75t_L g889 ( .A1(n_890), .A2(n_892), .B1(n_893), .B2(n_894), .Y(n_889) );
INVx2_ASAP7_75t_L g890 ( .A(n_891), .Y(n_890) );
CKINVDCx20_ASAP7_75t_R g895 ( .A(n_896), .Y(n_895) );
CKINVDCx20_ASAP7_75t_R g896 ( .A(n_897), .Y(n_896) );
endmodule