module fake_netlist_6_4426_n_800 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_157, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_800);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_157;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_800;

wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_208;
wire n_161;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_783;
wire n_725;
wire n_358;
wire n_160;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_255;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_222;
wire n_300;
wire n_248;
wire n_179;
wire n_517;
wire n_718;
wire n_747;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_658;
wire n_616;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_693;
wire n_167;
wire n_758;
wire n_174;
wire n_516;
wire n_720;
wire n_525;
wire n_631;
wire n_611;
wire n_491;
wire n_656;
wire n_772;
wire n_797;
wire n_666;
wire n_371;
wire n_795;
wire n_770;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_779;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_777;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_163;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_594;
wire n_565;
wire n_719;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_599;
wire n_513;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_792;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_788;
wire n_325;
wire n_767;
wire n_329;
wire n_464;
wire n_600;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_159;
wire n_162;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_775;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_728;
wire n_681;
wire n_729;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_697;
wire n_687;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_736;
wire n_613;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_663;
wire n_379;
wire n_170;
wire n_778;
wire n_332;
wire n_336;
wire n_410;
wire n_398;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_171;
wire n_678;
wire n_192;
wire n_169;
wire n_649;
wire n_283;

INVx1_ASAP7_75t_L g159 ( 
.A(n_11),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_45),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_124),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_12),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_79),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_75),
.Y(n_164)
);

BUFx2_ASAP7_75t_L g165 ( 
.A(n_135),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_104),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_145),
.Y(n_167)
);

CKINVDCx14_ASAP7_75t_R g168 ( 
.A(n_15),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_33),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_133),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_122),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_62),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_41),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_71),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_89),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_139),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_102),
.Y(n_177)
);

INVx2_ASAP7_75t_SL g178 ( 
.A(n_96),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_40),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_39),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_24),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_66),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_153),
.Y(n_183)
);

INVx2_ASAP7_75t_SL g184 ( 
.A(n_87),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_110),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_6),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_113),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_97),
.Y(n_188)
);

BUFx2_ASAP7_75t_L g189 ( 
.A(n_155),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_65),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_128),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_37),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_29),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_109),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_130),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_134),
.Y(n_196)
);

BUFx2_ASAP7_75t_SL g197 ( 
.A(n_157),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_23),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_114),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_63),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_106),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_9),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_99),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_100),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_112),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_6),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_150),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_9),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_4),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_72),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_151),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_25),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_126),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_59),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_108),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_83),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_162),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_159),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_208),
.Y(n_219)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_173),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_212),
.B(n_186),
.Y(n_221)
);

AND2x6_ASAP7_75t_L g222 ( 
.A(n_173),
.B(n_19),
.Y(n_222)
);

AND2x4_ASAP7_75t_L g223 ( 
.A(n_169),
.B(n_20),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_173),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_168),
.B(n_0),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_164),
.Y(n_226)
);

AND2x4_ASAP7_75t_L g227 ( 
.A(n_169),
.B(n_21),
.Y(n_227)
);

AND2x4_ASAP7_75t_L g228 ( 
.A(n_181),
.B(n_22),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_166),
.Y(n_229)
);

OA21x2_ASAP7_75t_L g230 ( 
.A1(n_181),
.A2(n_0),
.B(n_1),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g231 ( 
.A(n_202),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_173),
.Y(n_232)
);

BUFx2_ASAP7_75t_L g233 ( 
.A(n_168),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_170),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_206),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_174),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_165),
.B(n_189),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_176),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_200),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g240 ( 
.A(n_209),
.Y(n_240)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_187),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_214),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_200),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_200),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_200),
.Y(n_245)
);

AND2x4_ASAP7_75t_L g246 ( 
.A(n_187),
.B(n_26),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_195),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_195),
.Y(n_248)
);

AND2x4_ASAP7_75t_L g249 ( 
.A(n_178),
.B(n_184),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_177),
.Y(n_250)
);

BUFx12f_ASAP7_75t_L g251 ( 
.A(n_214),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_180),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_182),
.B(n_2),
.Y(n_253)
);

NOR2x1_ASAP7_75t_L g254 ( 
.A(n_198),
.B(n_203),
.Y(n_254)
);

BUFx2_ASAP7_75t_L g255 ( 
.A(n_193),
.Y(n_255)
);

BUFx2_ASAP7_75t_L g256 ( 
.A(n_193),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_188),
.B(n_3),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_210),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_205),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_233),
.B(n_210),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_243),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_233),
.B(n_160),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_243),
.Y(n_263)
);

INVx5_ASAP7_75t_L g264 ( 
.A(n_222),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_244),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_244),
.Y(n_266)
);

OAI22xp33_ASAP7_75t_L g267 ( 
.A1(n_235),
.A2(n_207),
.B1(n_211),
.B2(n_213),
.Y(n_267)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_224),
.Y(n_268)
);

OR2x2_ASAP7_75t_L g269 ( 
.A(n_217),
.B(n_4),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_237),
.B(n_216),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_245),
.Y(n_271)
);

BUFx3_ASAP7_75t_L g272 ( 
.A(n_223),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_245),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_248),
.Y(n_274)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_224),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_224),
.Y(n_276)
);

INVx4_ASAP7_75t_L g277 ( 
.A(n_222),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_248),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_248),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_248),
.Y(n_280)
);

NAND3xp33_ASAP7_75t_L g281 ( 
.A(n_225),
.B(n_215),
.C(n_204),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_249),
.B(n_161),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_224),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_221),
.B(n_163),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_232),
.Y(n_285)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_232),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_232),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_232),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_239),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_225),
.B(n_167),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_239),
.Y(n_291)
);

BUFx6f_ASAP7_75t_SL g292 ( 
.A(n_249),
.Y(n_292)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_239),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_239),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_218),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_247),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_218),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_249),
.B(n_242),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_247),
.Y(n_299)
);

OR2x2_ASAP7_75t_L g300 ( 
.A(n_231),
.B(n_5),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_241),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_251),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_241),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_241),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_257),
.B(n_171),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_219),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_250),
.Y(n_307)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_223),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_274),
.Y(n_309)
);

AOI221xp5_ASAP7_75t_L g310 ( 
.A1(n_267),
.A2(n_257),
.B1(n_221),
.B2(n_253),
.C(n_256),
.Y(n_310)
);

BUFx3_ASAP7_75t_L g311 ( 
.A(n_306),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_272),
.B(n_223),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_272),
.B(n_227),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_306),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_274),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_308),
.B(n_227),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_278),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_284),
.B(n_251),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_279),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_278),
.Y(n_320)
);

NAND2xp33_ASAP7_75t_SL g321 ( 
.A(n_269),
.B(n_240),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_308),
.A2(n_254),
.B(n_228),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_270),
.B(n_258),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_282),
.B(n_252),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_298),
.B(n_258),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_283),
.Y(n_326)
);

BUFx3_ASAP7_75t_L g327 ( 
.A(n_301),
.Y(n_327)
);

INVx4_ASAP7_75t_L g328 ( 
.A(n_268),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_282),
.B(n_226),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_305),
.B(n_227),
.Y(n_330)
);

INVx3_ASAP7_75t_L g331 ( 
.A(n_276),
.Y(n_331)
);

AND2x4_ASAP7_75t_L g332 ( 
.A(n_269),
.B(n_228),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_281),
.B(n_228),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_290),
.B(n_246),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g335 ( 
.A(n_276),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_283),
.Y(n_336)
);

BUFx5_ASAP7_75t_L g337 ( 
.A(n_265),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_291),
.Y(n_338)
);

NOR3xp33_ASAP7_75t_L g339 ( 
.A(n_260),
.B(n_255),
.C(n_256),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_279),
.B(n_246),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_280),
.B(n_246),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_280),
.B(n_220),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_291),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_268),
.B(n_220),
.Y(n_344)
);

AND2x4_ASAP7_75t_L g345 ( 
.A(n_300),
.B(n_229),
.Y(n_345)
);

NAND2x1_ASAP7_75t_L g346 ( 
.A(n_277),
.B(n_222),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_268),
.B(n_220),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_262),
.B(n_234),
.Y(n_348)
);

NAND3xp33_ASAP7_75t_L g349 ( 
.A(n_300),
.B(n_238),
.C(n_236),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_302),
.B(n_172),
.Y(n_350)
);

BUFx5_ASAP7_75t_L g351 ( 
.A(n_265),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_302),
.B(n_175),
.Y(n_352)
);

NOR2xp67_ASAP7_75t_L g353 ( 
.A(n_264),
.B(n_179),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_275),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_275),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_275),
.B(n_250),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_286),
.B(n_250),
.Y(n_357)
);

O2A1O1Ixp33_ASAP7_75t_L g358 ( 
.A1(n_295),
.A2(n_230),
.B(n_255),
.C(n_197),
.Y(n_358)
);

BUFx5_ASAP7_75t_L g359 ( 
.A(n_266),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_286),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_286),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_264),
.B(n_183),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_293),
.B(n_250),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_293),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_293),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_285),
.B(n_250),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_264),
.B(n_185),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_285),
.B(n_259),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_292),
.B(n_259),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_287),
.B(n_259),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_287),
.B(n_259),
.Y(n_371)
);

AND2x4_ASAP7_75t_L g372 ( 
.A(n_301),
.B(n_190),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_292),
.Y(n_373)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_276),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_312),
.B(n_307),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g376 ( 
.A1(n_313),
.A2(n_277),
.B(n_264),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_316),
.B(n_307),
.Y(n_377)
);

HB1xp67_ASAP7_75t_L g378 ( 
.A(n_332),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_L g379 ( 
.A1(n_340),
.A2(n_277),
.B(n_264),
.Y(n_379)
);

O2A1O1Ixp33_ASAP7_75t_L g380 ( 
.A1(n_358),
.A2(n_297),
.B(n_295),
.C(n_299),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_334),
.B(n_296),
.Y(n_381)
);

O2A1O1Ixp33_ASAP7_75t_L g382 ( 
.A1(n_333),
.A2(n_297),
.B(n_296),
.C(n_299),
.Y(n_382)
);

NOR3xp33_ASAP7_75t_L g383 ( 
.A(n_310),
.B(n_191),
.C(n_192),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_327),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_332),
.B(n_288),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g386 ( 
.A1(n_341),
.A2(n_289),
.B(n_288),
.Y(n_386)
);

O2A1O1Ixp33_ASAP7_75t_L g387 ( 
.A1(n_330),
.A2(n_230),
.B(n_303),
.C(n_304),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_L g388 ( 
.A1(n_322),
.A2(n_289),
.B(n_294),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_311),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_L g390 ( 
.A1(n_342),
.A2(n_294),
.B(n_276),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_309),
.Y(n_391)
);

NAND2xp33_ASAP7_75t_L g392 ( 
.A(n_348),
.B(n_222),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_318),
.B(n_194),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_344),
.A2(n_294),
.B(n_276),
.Y(n_394)
);

O2A1O1Ixp33_ASAP7_75t_L g395 ( 
.A1(n_314),
.A2(n_230),
.B(n_303),
.C(n_304),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_315),
.Y(n_396)
);

AOI21x1_ASAP7_75t_L g397 ( 
.A1(n_347),
.A2(n_273),
.B(n_266),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_319),
.Y(n_398)
);

AOI21xp5_ASAP7_75t_L g399 ( 
.A1(n_346),
.A2(n_294),
.B(n_261),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_317),
.Y(n_400)
);

INVx3_ASAP7_75t_L g401 ( 
.A(n_328),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_L g402 ( 
.A1(n_329),
.A2(n_261),
.B(n_271),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_356),
.A2(n_294),
.B(n_263),
.Y(n_403)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_357),
.A2(n_271),
.B(n_263),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_320),
.B(n_259),
.Y(n_405)
);

AOI21x1_ASAP7_75t_L g406 ( 
.A1(n_354),
.A2(n_273),
.B(n_292),
.Y(n_406)
);

HB1xp67_ASAP7_75t_L g407 ( 
.A(n_345),
.Y(n_407)
);

BUFx2_ASAP7_75t_L g408 ( 
.A(n_321),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_323),
.B(n_196),
.Y(n_409)
);

O2A1O1Ixp33_ASAP7_75t_L g410 ( 
.A1(n_324),
.A2(n_325),
.B(n_345),
.C(n_367),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_326),
.B(n_336),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_363),
.A2(n_201),
.B(n_199),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_372),
.B(n_5),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_372),
.A2(n_222),
.B1(n_80),
.B2(n_81),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_349),
.B(n_222),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_339),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_338),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_337),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g419 ( 
.A1(n_366),
.A2(n_78),
.B(n_156),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_335),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_343),
.B(n_27),
.Y(n_421)
);

BUFx2_ASAP7_75t_L g422 ( 
.A(n_373),
.Y(n_422)
);

AOI21xp5_ASAP7_75t_L g423 ( 
.A1(n_368),
.A2(n_77),
.B(n_154),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_L g424 ( 
.A1(n_369),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_370),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_328),
.B(n_28),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_371),
.A2(n_362),
.B(n_353),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_350),
.B(n_11),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_337),
.B(n_30),
.Y(n_429)
);

AOI21x1_ASAP7_75t_L g430 ( 
.A1(n_355),
.A2(n_85),
.B(n_152),
.Y(n_430)
);

NAND3xp33_ASAP7_75t_L g431 ( 
.A(n_352),
.B(n_365),
.C(n_360),
.Y(n_431)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_361),
.A2(n_84),
.B(n_149),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_364),
.A2(n_82),
.B(n_148),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_337),
.B(n_31),
.Y(n_434)
);

INVx1_ASAP7_75t_SL g435 ( 
.A(n_337),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_337),
.B(n_32),
.Y(n_436)
);

O2A1O1Ixp33_ASAP7_75t_L g437 ( 
.A1(n_331),
.A2(n_12),
.B(n_13),
.C(n_14),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_L g438 ( 
.A1(n_331),
.A2(n_88),
.B(n_147),
.Y(n_438)
);

AO22x1_ASAP7_75t_L g439 ( 
.A1(n_335),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_439)
);

BUFx8_ASAP7_75t_L g440 ( 
.A(n_351),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_335),
.B(n_16),
.Y(n_441)
);

AOI21xp5_ASAP7_75t_L g442 ( 
.A1(n_374),
.A2(n_90),
.B(n_146),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_351),
.B(n_34),
.Y(n_443)
);

AND3x1_ASAP7_75t_SL g444 ( 
.A(n_417),
.B(n_416),
.C(n_424),
.Y(n_444)
);

OAI21x1_ASAP7_75t_L g445 ( 
.A1(n_427),
.A2(n_359),
.B(n_351),
.Y(n_445)
);

INVx2_ASAP7_75t_SL g446 ( 
.A(n_384),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g447 ( 
.A1(n_401),
.A2(n_374),
.B(n_359),
.Y(n_447)
);

OAI21x1_ASAP7_75t_L g448 ( 
.A1(n_397),
.A2(n_376),
.B(n_386),
.Y(n_448)
);

AOI21x1_ASAP7_75t_SL g449 ( 
.A1(n_443),
.A2(n_359),
.B(n_351),
.Y(n_449)
);

AOI21x1_ASAP7_75t_L g450 ( 
.A1(n_399),
.A2(n_359),
.B(n_351),
.Y(n_450)
);

INVx4_ASAP7_75t_L g451 ( 
.A(n_389),
.Y(n_451)
);

OAI22x1_ASAP7_75t_L g452 ( 
.A1(n_408),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_385),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_389),
.B(n_374),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_407),
.B(n_359),
.Y(n_455)
);

OAI21x1_ASAP7_75t_L g456 ( 
.A1(n_379),
.A2(n_158),
.B(n_91),
.Y(n_456)
);

OAI21x1_ASAP7_75t_L g457 ( 
.A1(n_388),
.A2(n_144),
.B(n_86),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_L g458 ( 
.A1(n_387),
.A2(n_76),
.B(n_142),
.Y(n_458)
);

AOI21xp5_ASAP7_75t_L g459 ( 
.A1(n_401),
.A2(n_74),
.B(n_141),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_378),
.Y(n_460)
);

INVx1_ASAP7_75t_SL g461 ( 
.A(n_413),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_409),
.B(n_17),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_389),
.B(n_92),
.Y(n_463)
);

NOR2xp67_ASAP7_75t_L g464 ( 
.A(n_431),
.B(n_73),
.Y(n_464)
);

OAI21x1_ASAP7_75t_L g465 ( 
.A1(n_418),
.A2(n_93),
.B(n_35),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_435),
.B(n_94),
.Y(n_466)
);

OAI21x1_ASAP7_75t_L g467 ( 
.A1(n_406),
.A2(n_143),
.B(n_36),
.Y(n_467)
);

NOR2x1_ASAP7_75t_SL g468 ( 
.A(n_420),
.B(n_70),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_411),
.Y(n_469)
);

OAI21x1_ASAP7_75t_L g470 ( 
.A1(n_394),
.A2(n_95),
.B(n_38),
.Y(n_470)
);

AOI21xp5_ASAP7_75t_L g471 ( 
.A1(n_435),
.A2(n_98),
.B(n_42),
.Y(n_471)
);

OR2x2_ASAP7_75t_L g472 ( 
.A(n_422),
.B(n_18),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_410),
.B(n_43),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_400),
.Y(n_474)
);

OAI21x1_ASAP7_75t_L g475 ( 
.A1(n_402),
.A2(n_44),
.B(n_46),
.Y(n_475)
);

AOI21xp5_ASAP7_75t_L g476 ( 
.A1(n_375),
.A2(n_47),
.B(n_48),
.Y(n_476)
);

NAND2x1p5_ASAP7_75t_L g477 ( 
.A(n_420),
.B(n_49),
.Y(n_477)
);

NAND2x1p5_ASAP7_75t_L g478 ( 
.A(n_420),
.B(n_50),
.Y(n_478)
);

A2O1A1Ixp33_ASAP7_75t_L g479 ( 
.A1(n_383),
.A2(n_51),
.B(n_52),
.C(n_53),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_425),
.B(n_54),
.Y(n_480)
);

INVx4_ASAP7_75t_L g481 ( 
.A(n_391),
.Y(n_481)
);

INVx1_ASAP7_75t_SL g482 ( 
.A(n_428),
.Y(n_482)
);

OAI21x1_ASAP7_75t_SL g483 ( 
.A1(n_421),
.A2(n_55),
.B(n_56),
.Y(n_483)
);

AOI21xp5_ASAP7_75t_L g484 ( 
.A1(n_377),
.A2(n_57),
.B(n_58),
.Y(n_484)
);

OAI21xp5_ASAP7_75t_L g485 ( 
.A1(n_395),
.A2(n_60),
.B(n_61),
.Y(n_485)
);

AOI21xp5_ASAP7_75t_L g486 ( 
.A1(n_381),
.A2(n_64),
.B(n_67),
.Y(n_486)
);

BUFx3_ASAP7_75t_L g487 ( 
.A(n_441),
.Y(n_487)
);

INVx3_ASAP7_75t_L g488 ( 
.A(n_396),
.Y(n_488)
);

OAI22x1_ASAP7_75t_L g489 ( 
.A1(n_393),
.A2(n_68),
.B1(n_69),
.B2(n_101),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_416),
.B(n_103),
.Y(n_490)
);

NOR2x1_ASAP7_75t_L g491 ( 
.A(n_443),
.B(n_105),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_402),
.B(n_107),
.Y(n_492)
);

OAI21x1_ASAP7_75t_L g493 ( 
.A1(n_390),
.A2(n_111),
.B(n_115),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_398),
.B(n_116),
.Y(n_494)
);

BUFx2_ASAP7_75t_L g495 ( 
.A(n_439),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_429),
.B(n_117),
.Y(n_496)
);

AOI21xp5_ASAP7_75t_L g497 ( 
.A1(n_392),
.A2(n_118),
.B(n_119),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_380),
.B(n_120),
.Y(n_498)
);

O2A1O1Ixp5_ASAP7_75t_L g499 ( 
.A1(n_415),
.A2(n_121),
.B(n_123),
.C(n_125),
.Y(n_499)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_440),
.Y(n_500)
);

BUFx3_ASAP7_75t_L g501 ( 
.A(n_500),
.Y(n_501)
);

AND2x4_ASAP7_75t_L g502 ( 
.A(n_451),
.B(n_414),
.Y(n_502)
);

OAI21x1_ASAP7_75t_L g503 ( 
.A1(n_449),
.A2(n_430),
.B(n_436),
.Y(n_503)
);

INVx4_ASAP7_75t_L g504 ( 
.A(n_451),
.Y(n_504)
);

INVx1_ASAP7_75t_SL g505 ( 
.A(n_472),
.Y(n_505)
);

OAI21x1_ASAP7_75t_L g506 ( 
.A1(n_445),
.A2(n_434),
.B(n_426),
.Y(n_506)
);

OAI21x1_ASAP7_75t_L g507 ( 
.A1(n_448),
.A2(n_382),
.B(n_403),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_453),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_488),
.Y(n_509)
);

AO21x2_ASAP7_75t_L g510 ( 
.A1(n_458),
.A2(n_485),
.B(n_473),
.Y(n_510)
);

INVx1_ASAP7_75t_SL g511 ( 
.A(n_461),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_488),
.Y(n_512)
);

BUFx3_ASAP7_75t_L g513 ( 
.A(n_500),
.Y(n_513)
);

OR2x6_ASAP7_75t_L g514 ( 
.A(n_455),
.B(n_437),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_L g515 ( 
.A1(n_469),
.A2(n_466),
.B1(n_461),
.B2(n_487),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_474),
.B(n_440),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_482),
.B(n_412),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_482),
.B(n_405),
.Y(n_518)
);

AOI22xp33_ASAP7_75t_L g519 ( 
.A1(n_490),
.A2(n_424),
.B1(n_404),
.B2(n_423),
.Y(n_519)
);

AOI22xp33_ASAP7_75t_L g520 ( 
.A1(n_462),
.A2(n_495),
.B1(n_485),
.B2(n_458),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_480),
.Y(n_521)
);

AOI22xp33_ASAP7_75t_L g522 ( 
.A1(n_489),
.A2(n_419),
.B1(n_442),
.B2(n_438),
.Y(n_522)
);

OAI21x1_ASAP7_75t_SL g523 ( 
.A1(n_468),
.A2(n_433),
.B(n_432),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_481),
.Y(n_524)
);

BUFx2_ASAP7_75t_R g525 ( 
.A(n_463),
.Y(n_525)
);

OAI21x1_ASAP7_75t_L g526 ( 
.A1(n_450),
.A2(n_127),
.B(n_129),
.Y(n_526)
);

OAI21x1_ASAP7_75t_L g527 ( 
.A1(n_457),
.A2(n_131),
.B(n_132),
.Y(n_527)
);

OAI21x1_ASAP7_75t_L g528 ( 
.A1(n_475),
.A2(n_136),
.B(n_137),
.Y(n_528)
);

BUFx2_ASAP7_75t_L g529 ( 
.A(n_460),
.Y(n_529)
);

OAI21xp5_ASAP7_75t_L g530 ( 
.A1(n_492),
.A2(n_138),
.B(n_140),
.Y(n_530)
);

OAI21x1_ASAP7_75t_L g531 ( 
.A1(n_470),
.A2(n_493),
.B(n_456),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_480),
.Y(n_532)
);

OAI21x1_ASAP7_75t_L g533 ( 
.A1(n_465),
.A2(n_467),
.B(n_496),
.Y(n_533)
);

OAI21x1_ASAP7_75t_L g534 ( 
.A1(n_496),
.A2(n_447),
.B(n_466),
.Y(n_534)
);

OAI21x1_ASAP7_75t_L g535 ( 
.A1(n_494),
.A2(n_497),
.B(n_491),
.Y(n_535)
);

HB1xp67_ASAP7_75t_L g536 ( 
.A(n_446),
.Y(n_536)
);

OA21x2_ASAP7_75t_L g537 ( 
.A1(n_498),
.A2(n_499),
.B(n_479),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_481),
.B(n_478),
.Y(n_538)
);

OAI21x1_ASAP7_75t_L g539 ( 
.A1(n_483),
.A2(n_459),
.B(n_484),
.Y(n_539)
);

AND2x4_ASAP7_75t_L g540 ( 
.A(n_454),
.B(n_464),
.Y(n_540)
);

NAND2x1p5_ASAP7_75t_L g541 ( 
.A(n_471),
.B(n_476),
.Y(n_541)
);

OA21x2_ASAP7_75t_L g542 ( 
.A1(n_486),
.A2(n_444),
.B(n_477),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_477),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_478),
.Y(n_544)
);

NOR2x1_ASAP7_75t_R g545 ( 
.A(n_452),
.B(n_258),
.Y(n_545)
);

OAI21x1_ASAP7_75t_L g546 ( 
.A1(n_449),
.A2(n_445),
.B(n_448),
.Y(n_546)
);

AOI21xp5_ASAP7_75t_L g547 ( 
.A1(n_466),
.A2(n_435),
.B(n_401),
.Y(n_547)
);

AO21x2_ASAP7_75t_L g548 ( 
.A1(n_458),
.A2(n_485),
.B(n_473),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_500),
.Y(n_549)
);

NOR2x1_ASAP7_75t_R g550 ( 
.A(n_500),
.B(n_258),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_508),
.Y(n_551)
);

BUFx3_ASAP7_75t_L g552 ( 
.A(n_501),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_508),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_546),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_515),
.B(n_520),
.Y(n_555)
);

CKINVDCx11_ASAP7_75t_R g556 ( 
.A(n_505),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_509),
.Y(n_557)
);

BUFx3_ASAP7_75t_L g558 ( 
.A(n_501),
.Y(n_558)
);

AOI21x1_ASAP7_75t_L g559 ( 
.A1(n_546),
.A2(n_503),
.B(n_533),
.Y(n_559)
);

OAI22xp33_ASAP7_75t_L g560 ( 
.A1(n_511),
.A2(n_516),
.B1(n_549),
.B2(n_529),
.Y(n_560)
);

AOI22xp33_ASAP7_75t_SL g561 ( 
.A1(n_510),
.A2(n_548),
.B1(n_549),
.B2(n_529),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_507),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_509),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_521),
.B(n_532),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_536),
.B(n_545),
.Y(n_565)
);

INVx2_ASAP7_75t_SL g566 ( 
.A(n_538),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_507),
.Y(n_567)
);

INVx2_ASAP7_75t_SL g568 ( 
.A(n_538),
.Y(n_568)
);

HB1xp67_ASAP7_75t_L g569 ( 
.A(n_512),
.Y(n_569)
);

AO21x2_ASAP7_75t_L g570 ( 
.A1(n_510),
.A2(n_548),
.B(n_531),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_512),
.Y(n_571)
);

AOI22xp33_ASAP7_75t_L g572 ( 
.A1(n_502),
.A2(n_510),
.B1(n_548),
.B2(n_514),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_526),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_524),
.Y(n_574)
);

AO21x1_ASAP7_75t_SL g575 ( 
.A1(n_530),
.A2(n_532),
.B(n_521),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_524),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_526),
.Y(n_577)
);

AND2x2_ASAP7_75t_L g578 ( 
.A(n_514),
.B(n_518),
.Y(n_578)
);

INVxp67_ASAP7_75t_SL g579 ( 
.A(n_543),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_531),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_543),
.Y(n_581)
);

HB1xp67_ASAP7_75t_L g582 ( 
.A(n_513),
.Y(n_582)
);

AND2x2_ASAP7_75t_L g583 ( 
.A(n_514),
.B(n_502),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_544),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_513),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_527),
.Y(n_586)
);

AOI22xp33_ASAP7_75t_L g587 ( 
.A1(n_502),
.A2(n_514),
.B1(n_519),
.B2(n_517),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_544),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_542),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_542),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_527),
.Y(n_591)
);

INVx3_ASAP7_75t_L g592 ( 
.A(n_504),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_542),
.B(n_540),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_542),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_528),
.Y(n_595)
);

BUFx3_ASAP7_75t_L g596 ( 
.A(n_552),
.Y(n_596)
);

HB1xp67_ASAP7_75t_L g597 ( 
.A(n_582),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_564),
.B(n_540),
.Y(n_598)
);

HB1xp67_ASAP7_75t_L g599 ( 
.A(n_552),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_551),
.Y(n_600)
);

AND2x4_ASAP7_75t_SL g601 ( 
.A(n_592),
.B(n_504),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_551),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_578),
.B(n_540),
.Y(n_603)
);

OR2x2_ASAP7_75t_L g604 ( 
.A(n_555),
.B(n_537),
.Y(n_604)
);

INVx2_ASAP7_75t_SL g605 ( 
.A(n_552),
.Y(n_605)
);

INVx2_ASAP7_75t_SL g606 ( 
.A(n_558),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_578),
.B(n_528),
.Y(n_607)
);

OR2x2_ASAP7_75t_L g608 ( 
.A(n_572),
.B(n_537),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_553),
.B(n_537),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_553),
.B(n_537),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_553),
.Y(n_611)
);

AOI22xp33_ASAP7_75t_L g612 ( 
.A1(n_583),
.A2(n_541),
.B1(n_522),
.B2(n_504),
.Y(n_612)
);

BUFx3_ASAP7_75t_L g613 ( 
.A(n_558),
.Y(n_613)
);

OR2x2_ASAP7_75t_L g614 ( 
.A(n_587),
.B(n_534),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_583),
.B(n_525),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g616 ( 
.A(n_571),
.B(n_541),
.Y(n_616)
);

OR2x2_ASAP7_75t_L g617 ( 
.A(n_593),
.B(n_534),
.Y(n_617)
);

HB1xp67_ASAP7_75t_L g618 ( 
.A(n_558),
.Y(n_618)
);

AO31x2_ASAP7_75t_L g619 ( 
.A1(n_589),
.A2(n_547),
.A3(n_503),
.B(n_506),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_557),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_557),
.B(n_541),
.Y(n_621)
);

OAI22xp5_ASAP7_75t_L g622 ( 
.A1(n_560),
.A2(n_550),
.B1(n_523),
.B2(n_539),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_566),
.B(n_550),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_563),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_563),
.Y(n_625)
);

OR2x2_ASAP7_75t_L g626 ( 
.A(n_593),
.B(n_533),
.Y(n_626)
);

INVxp67_ASAP7_75t_SL g627 ( 
.A(n_579),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_566),
.B(n_539),
.Y(n_628)
);

INVx2_ASAP7_75t_SL g629 ( 
.A(n_585),
.Y(n_629)
);

BUFx6f_ASAP7_75t_L g630 ( 
.A(n_568),
.Y(n_630)
);

NOR2x1p5_ASAP7_75t_L g631 ( 
.A(n_592),
.B(n_523),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_568),
.B(n_535),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_556),
.Y(n_633)
);

OR2x2_ASAP7_75t_L g634 ( 
.A(n_561),
.B(n_594),
.Y(n_634)
);

INVx1_ASAP7_75t_SL g635 ( 
.A(n_565),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_569),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_574),
.B(n_535),
.Y(n_637)
);

OR2x6_ASAP7_75t_L g638 ( 
.A(n_586),
.B(n_506),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_574),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_576),
.Y(n_640)
);

INVx4_ASAP7_75t_L g641 ( 
.A(n_592),
.Y(n_641)
);

BUFx3_ASAP7_75t_L g642 ( 
.A(n_592),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_581),
.B(n_584),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_581),
.B(n_584),
.Y(n_644)
);

OR2x2_ASAP7_75t_L g645 ( 
.A(n_589),
.B(n_594),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_598),
.B(n_588),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_643),
.B(n_590),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_603),
.B(n_588),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_620),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_636),
.B(n_576),
.Y(n_650)
);

AND2x4_ASAP7_75t_L g651 ( 
.A(n_643),
.B(n_554),
.Y(n_651)
);

INVx1_ASAP7_75t_SL g652 ( 
.A(n_635),
.Y(n_652)
);

BUFx2_ASAP7_75t_L g653 ( 
.A(n_626),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_639),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_629),
.B(n_590),
.Y(n_655)
);

OAI22xp5_ASAP7_75t_L g656 ( 
.A1(n_623),
.A2(n_595),
.B1(n_591),
.B2(n_586),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_644),
.B(n_607),
.Y(n_657)
);

INVxp67_ASAP7_75t_SL g658 ( 
.A(n_627),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_645),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_644),
.B(n_607),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_597),
.B(n_570),
.Y(n_661)
);

AOI22xp33_ASAP7_75t_L g662 ( 
.A1(n_622),
.A2(n_575),
.B1(n_595),
.B2(n_570),
.Y(n_662)
);

HB1xp67_ASAP7_75t_L g663 ( 
.A(n_599),
.Y(n_663)
);

AOI22xp33_ASAP7_75t_L g664 ( 
.A1(n_615),
.A2(n_575),
.B1(n_570),
.B2(n_591),
.Y(n_664)
);

INVxp67_ASAP7_75t_SL g665 ( 
.A(n_639),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_645),
.Y(n_666)
);

INVx4_ASAP7_75t_L g667 ( 
.A(n_601),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_615),
.B(n_567),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_604),
.B(n_554),
.Y(n_669)
);

BUFx2_ASAP7_75t_L g670 ( 
.A(n_626),
.Y(n_670)
);

BUFx2_ASAP7_75t_L g671 ( 
.A(n_617),
.Y(n_671)
);

AOI222xp33_ASAP7_75t_L g672 ( 
.A1(n_629),
.A2(n_562),
.B1(n_567),
.B2(n_591),
.C1(n_586),
.C2(n_554),
.Y(n_672)
);

HB1xp67_ASAP7_75t_L g673 ( 
.A(n_618),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_617),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_600),
.Y(n_675)
);

AOI22xp33_ASAP7_75t_L g676 ( 
.A1(n_614),
.A2(n_573),
.B1(n_577),
.B2(n_567),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_637),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_624),
.Y(n_678)
);

NOR2x1_ASAP7_75t_L g679 ( 
.A(n_596),
.B(n_573),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_625),
.Y(n_680)
);

INVx2_ASAP7_75t_SL g681 ( 
.A(n_596),
.Y(n_681)
);

AND2x4_ASAP7_75t_L g682 ( 
.A(n_630),
.B(n_580),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_609),
.Y(n_683)
);

HB1xp67_ASAP7_75t_L g684 ( 
.A(n_605),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_640),
.B(n_562),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_609),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_657),
.B(n_634),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_657),
.B(n_634),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_649),
.Y(n_689)
);

AND2x4_ASAP7_75t_L g690 ( 
.A(n_674),
.B(n_628),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_660),
.B(n_671),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_654),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_678),
.Y(n_693)
);

O2A1O1Ixp5_ASAP7_75t_L g694 ( 
.A1(n_656),
.A2(n_632),
.B(n_614),
.C(n_604),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_680),
.Y(n_695)
);

AND2x4_ASAP7_75t_SL g696 ( 
.A(n_667),
.B(n_630),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_648),
.B(n_621),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_659),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_660),
.B(n_608),
.Y(n_699)
);

BUFx2_ASAP7_75t_SL g700 ( 
.A(n_681),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_646),
.B(n_621),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_658),
.B(n_612),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_659),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_666),
.Y(n_704)
);

AND2x2_ASAP7_75t_L g705 ( 
.A(n_671),
.B(n_670),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_666),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_655),
.B(n_663),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_674),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_673),
.B(n_616),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_653),
.B(n_608),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_668),
.B(n_616),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_653),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_670),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_650),
.B(n_610),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_677),
.B(n_610),
.Y(n_715)
);

AOI22xp5_ASAP7_75t_L g716 ( 
.A1(n_702),
.A2(n_664),
.B1(n_652),
.B2(n_662),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_689),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_699),
.B(n_669),
.Y(n_718)
);

HB1xp67_ASAP7_75t_L g719 ( 
.A(n_705),
.Y(n_719)
);

NAND4xp25_ASAP7_75t_L g720 ( 
.A(n_707),
.B(n_661),
.C(n_672),
.D(n_676),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_692),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_693),
.Y(n_722)
);

AOI33xp33_ASAP7_75t_L g723 ( 
.A1(n_695),
.A2(n_677),
.A3(n_681),
.B1(n_647),
.B2(n_654),
.B3(n_686),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_691),
.B(n_686),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_708),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_698),
.Y(n_726)
);

NOR2xp67_ASAP7_75t_L g727 ( 
.A(n_703),
.B(n_684),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_692),
.Y(n_728)
);

NOR3xp33_ASAP7_75t_L g729 ( 
.A(n_702),
.B(n_605),
.C(n_606),
.Y(n_729)
);

AND2x2_ASAP7_75t_L g730 ( 
.A(n_699),
.B(n_691),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_701),
.B(n_665),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_704),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_706),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_690),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_697),
.B(n_688),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_687),
.B(n_683),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_717),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_722),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_725),
.Y(n_739)
);

INVxp67_ASAP7_75t_L g740 ( 
.A(n_719),
.Y(n_740)
);

AOI22xp33_ASAP7_75t_L g741 ( 
.A1(n_716),
.A2(n_710),
.B1(n_688),
.B2(n_687),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_735),
.B(n_709),
.Y(n_742)
);

OR2x2_ASAP7_75t_L g743 ( 
.A(n_719),
.B(n_710),
.Y(n_743)
);

AOI22xp5_ASAP7_75t_L g744 ( 
.A1(n_729),
.A2(n_690),
.B1(n_705),
.B2(n_711),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_718),
.B(n_713),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_726),
.Y(n_746)
);

A2O1A1Ixp33_ASAP7_75t_L g747 ( 
.A1(n_723),
.A2(n_694),
.B(n_633),
.C(n_696),
.Y(n_747)
);

INVxp67_ASAP7_75t_L g748 ( 
.A(n_732),
.Y(n_748)
);

XOR2x2_ASAP7_75t_L g749 ( 
.A(n_730),
.B(n_633),
.Y(n_749)
);

XOR2x2_ASAP7_75t_L g750 ( 
.A(n_730),
.B(n_714),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_748),
.B(n_718),
.Y(n_751)
);

OAI211xp5_ASAP7_75t_L g752 ( 
.A1(n_747),
.A2(n_720),
.B(n_727),
.C(n_731),
.Y(n_752)
);

A2O1A1Ixp33_ASAP7_75t_L g753 ( 
.A1(n_744),
.A2(n_723),
.B(n_734),
.C(n_733),
.Y(n_753)
);

OAI21xp33_ASAP7_75t_L g754 ( 
.A1(n_741),
.A2(n_712),
.B(n_736),
.Y(n_754)
);

AOI21xp5_ASAP7_75t_L g755 ( 
.A1(n_742),
.A2(n_679),
.B(n_696),
.Y(n_755)
);

OAI21xp33_ASAP7_75t_L g756 ( 
.A1(n_750),
.A2(n_690),
.B(n_734),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_751),
.Y(n_757)
);

XOR2x2_ASAP7_75t_L g758 ( 
.A(n_755),
.B(n_749),
.Y(n_758)
);

AOI21xp5_ASAP7_75t_L g759 ( 
.A1(n_752),
.A2(n_737),
.B(n_738),
.Y(n_759)
);

OAI21xp5_ASAP7_75t_SL g760 ( 
.A1(n_753),
.A2(n_740),
.B(n_745),
.Y(n_760)
);

AOI22xp5_ASAP7_75t_L g761 ( 
.A1(n_754),
.A2(n_745),
.B1(n_746),
.B2(n_739),
.Y(n_761)
);

NAND4xp25_ASAP7_75t_SL g762 ( 
.A(n_756),
.B(n_743),
.C(n_724),
.D(n_728),
.Y(n_762)
);

AND2x2_ASAP7_75t_L g763 ( 
.A(n_757),
.B(n_728),
.Y(n_763)
);

NAND4xp25_ASAP7_75t_L g764 ( 
.A(n_760),
.B(n_613),
.C(n_715),
.D(n_721),
.Y(n_764)
);

AO21x1_ASAP7_75t_L g765 ( 
.A1(n_759),
.A2(n_721),
.B(n_667),
.Y(n_765)
);

AOI221xp5_ASAP7_75t_L g766 ( 
.A1(n_762),
.A2(n_700),
.B1(n_630),
.B2(n_683),
.C(n_682),
.Y(n_766)
);

OAI21xp33_ASAP7_75t_L g767 ( 
.A1(n_761),
.A2(n_613),
.B(n_606),
.Y(n_767)
);

NOR2x1_ASAP7_75t_L g768 ( 
.A(n_764),
.B(n_758),
.Y(n_768)
);

NAND3xp33_ASAP7_75t_L g769 ( 
.A(n_767),
.B(n_630),
.C(n_628),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_769),
.Y(n_770)
);

NOR4xp75_ASAP7_75t_L g771 ( 
.A(n_768),
.B(n_765),
.C(n_763),
.D(n_766),
.Y(n_771)
);

NOR4xp25_ASAP7_75t_L g772 ( 
.A(n_769),
.B(n_602),
.C(n_685),
.D(n_573),
.Y(n_772)
);

NOR2x1_ASAP7_75t_L g773 ( 
.A(n_770),
.B(n_700),
.Y(n_773)
);

NOR2x1_ASAP7_75t_L g774 ( 
.A(n_771),
.B(n_667),
.Y(n_774)
);

AND2x4_ASAP7_75t_L g775 ( 
.A(n_772),
.B(n_682),
.Y(n_775)
);

NOR2xp67_ASAP7_75t_L g776 ( 
.A(n_770),
.B(n_682),
.Y(n_776)
);

NAND4xp75_ASAP7_75t_L g777 ( 
.A(n_770),
.B(n_647),
.C(n_669),
.D(n_577),
.Y(n_777)
);

AOI22xp5_ASAP7_75t_L g778 ( 
.A1(n_770),
.A2(n_651),
.B1(n_631),
.B2(n_675),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_773),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_776),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_774),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_778),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_775),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_777),
.Y(n_784)
);

INVxp67_ASAP7_75t_L g785 ( 
.A(n_781),
.Y(n_785)
);

NOR4xp75_ASAP7_75t_SL g786 ( 
.A(n_780),
.B(n_601),
.C(n_642),
.D(n_619),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_783),
.Y(n_787)
);

AO22x2_ASAP7_75t_L g788 ( 
.A1(n_779),
.A2(n_641),
.B1(n_675),
.B2(n_611),
.Y(n_788)
);

AOI21xp5_ASAP7_75t_L g789 ( 
.A1(n_787),
.A2(n_780),
.B(n_782),
.Y(n_789)
);

AOI21xp5_ASAP7_75t_L g790 ( 
.A1(n_785),
.A2(n_784),
.B(n_638),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_788),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_789),
.Y(n_792)
);

AOI21xp33_ASAP7_75t_L g793 ( 
.A1(n_791),
.A2(n_786),
.B(n_638),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_790),
.B(n_651),
.Y(n_794)
);

OAI22xp5_ASAP7_75t_SL g795 ( 
.A1(n_792),
.A2(n_642),
.B1(n_641),
.B2(n_600),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_794),
.B(n_651),
.Y(n_796)
);

AOI21xp5_ASAP7_75t_L g797 ( 
.A1(n_795),
.A2(n_793),
.B(n_577),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_797),
.Y(n_798)
);

OR2x6_ASAP7_75t_L g799 ( 
.A(n_798),
.B(n_796),
.Y(n_799)
);

OAI21xp5_ASAP7_75t_L g800 ( 
.A1(n_799),
.A2(n_559),
.B(n_638),
.Y(n_800)
);


endmodule