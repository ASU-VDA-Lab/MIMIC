module fake_jpeg_23117_n_288 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_288);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_288;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

INVx4_ASAP7_75t_SL g29 ( 
.A(n_20),
.Y(n_29)
);

OR2x2_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_16),
.Y(n_41)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx3_ASAP7_75t_SL g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

NAND2xp33_ASAP7_75t_SL g74 ( 
.A(n_41),
.B(n_52),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_31),
.A2(n_25),
.B1(n_13),
.B2(n_17),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_42),
.A2(n_29),
.B1(n_13),
.B2(n_17),
.Y(n_72)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_30),
.B(n_27),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_44),
.B(n_51),
.Y(n_60)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_50),
.B(n_29),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_33),
.B(n_27),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_32),
.B(n_12),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_46),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_55),
.Y(n_83)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_53),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g76 ( 
.A(n_57),
.Y(n_76)
);

BUFx4f_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_44),
.B(n_24),
.Y(n_61)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_63),
.Y(n_93)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_66),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_49),
.B(n_24),
.Y(n_67)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_69),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_48),
.B(n_37),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_41),
.Y(n_84)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_72),
.A2(n_29),
.B1(n_54),
.B2(n_21),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_73),
.B(n_75),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_60),
.B(n_51),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_77),
.B(n_84),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_80),
.A2(n_68),
.B1(n_65),
.B2(n_58),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_74),
.B(n_41),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_90),
.B(n_96),
.C(n_52),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_62),
.A2(n_74),
.B1(n_31),
.B2(n_70),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_91),
.A2(n_94),
.B1(n_58),
.B2(n_64),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_60),
.A2(n_31),
.B1(n_29),
.B2(n_36),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_55),
.A2(n_38),
.B(n_50),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_95),
.A2(n_49),
.B(n_28),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_72),
.B(n_52),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_98),
.B(n_34),
.Y(n_140)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_76),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_99),
.B(n_100),
.Y(n_130)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_76),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_95),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_101),
.B(n_102),
.Y(n_132)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_87),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_103),
.Y(n_138)
);

OAI21xp33_ASAP7_75t_SL g134 ( 
.A1(n_104),
.A2(n_115),
.B(n_117),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_87),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_105),
.B(n_106),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_94),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_89),
.A2(n_96),
.B1(n_90),
.B2(n_84),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_107),
.A2(n_114),
.B1(n_115),
.B2(n_117),
.Y(n_121)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_85),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_108),
.B(n_110),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_81),
.B(n_48),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_109),
.B(n_79),
.Y(n_127)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_111),
.A2(n_101),
.B(n_106),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_81),
.A2(n_32),
.B1(n_30),
.B2(n_35),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_113),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_86),
.A2(n_36),
.B1(n_40),
.B2(n_38),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_86),
.A2(n_32),
.B1(n_37),
.B2(n_30),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_78),
.B(n_56),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_116),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_83),
.A2(n_32),
.B1(n_35),
.B2(n_37),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_118),
.A2(n_56),
.B1(n_71),
.B2(n_78),
.Y(n_142)
);

MAJx2_ASAP7_75t_L g119 ( 
.A(n_82),
.B(n_35),
.C(n_46),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_28),
.C(n_64),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_120),
.B(n_126),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_107),
.B(n_98),
.C(n_102),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_122),
.B(n_135),
.C(n_136),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_123),
.A2(n_23),
.B(n_22),
.Y(n_167)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_109),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_125),
.B(n_129),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g126 ( 
.A(n_118),
.B(n_82),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_127),
.B(n_131),
.Y(n_149)
);

XOR2x1_ASAP7_75t_L g128 ( 
.A(n_111),
.B(n_46),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g163 ( 
.A(n_128),
.B(n_26),
.Y(n_163)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_114),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_99),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_103),
.A2(n_43),
.B(n_93),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_133),
.A2(n_100),
.B(n_88),
.Y(n_150)
);

OAI21xp33_ASAP7_75t_SL g162 ( 
.A1(n_134),
.A2(n_142),
.B(n_66),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_112),
.B(n_105),
.C(n_119),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_108),
.B(n_85),
.C(n_97),
.Y(n_136)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_113),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_139),
.A2(n_92),
.B1(n_63),
.B2(n_19),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_140),
.B(n_69),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_132),
.A2(n_104),
.B1(n_88),
.B2(n_59),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_144),
.A2(n_155),
.B1(n_156),
.B2(n_164),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_143),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_146),
.Y(n_172)
);

XNOR2x1_ASAP7_75t_SL g147 ( 
.A(n_128),
.B(n_135),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_147),
.A2(n_20),
.B1(n_18),
.B2(n_14),
.Y(n_182)
);

CKINVDCx14_ASAP7_75t_R g183 ( 
.A(n_150),
.Y(n_183)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_127),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_151),
.B(n_159),
.Y(n_173)
);

INVx2_ASAP7_75t_SL g152 ( 
.A(n_131),
.Y(n_152)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_152),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_122),
.B(n_110),
.C(n_57),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_153),
.B(n_154),
.C(n_157),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_124),
.A2(n_19),
.B(n_26),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_120),
.B(n_66),
.C(n_26),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_130),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_123),
.A2(n_0),
.B(n_1),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_160),
.B(n_161),
.Y(n_184)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_136),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_162),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_163),
.B(n_167),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_133),
.A2(n_139),
.B(n_124),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_137),
.A2(n_23),
.B(n_22),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_165),
.A2(n_121),
.B1(n_129),
.B2(n_125),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_140),
.B(n_23),
.C(n_22),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_166),
.B(n_121),
.C(n_141),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_142),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_168),
.B(n_18),
.Y(n_185)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_149),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_171),
.B(n_174),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_176),
.B(n_178),
.C(n_188),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_148),
.B(n_126),
.C(n_138),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_149),
.Y(n_179)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_179),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_158),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_180),
.Y(n_194)
);

AO22x1_ASAP7_75t_SL g181 ( 
.A1(n_147),
.A2(n_138),
.B1(n_18),
.B2(n_14),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_181),
.A2(n_185),
.B(n_169),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_182),
.B(n_167),
.Y(n_193)
);

CKINVDCx14_ASAP7_75t_R g186 ( 
.A(n_165),
.Y(n_186)
);

CKINVDCx14_ASAP7_75t_R g210 ( 
.A(n_186),
.Y(n_210)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_152),
.Y(n_187)
);

INVx11_ASAP7_75t_L g204 ( 
.A(n_187),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_148),
.B(n_20),
.C(n_1),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_152),
.Y(n_189)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_189),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_190),
.A2(n_144),
.B1(n_168),
.B2(n_160),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_150),
.Y(n_191)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_191),
.Y(n_197)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_193),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_196),
.A2(n_202),
.B1(n_207),
.B2(n_170),
.Y(n_225)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_187),
.Y(n_199)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_199),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_178),
.B(n_145),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_200),
.B(n_209),
.C(n_211),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_183),
.A2(n_164),
.B1(n_156),
.B2(n_157),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_181),
.B(n_145),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_203),
.B(n_177),
.Y(n_222)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_205),
.Y(n_214)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_173),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_206),
.B(n_208),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_190),
.A2(n_153),
.B1(n_163),
.B2(n_166),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_185),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_175),
.B(n_154),
.C(n_3),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_175),
.B(n_0),
.C(n_4),
.Y(n_211)
);

A2O1A1Ixp33_ASAP7_75t_L g216 ( 
.A1(n_205),
.A2(n_181),
.B(n_184),
.C(n_182),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_216),
.A2(n_210),
.B(n_197),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_199),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_217),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_201),
.B(n_209),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_219),
.B(n_224),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_204),
.B(n_172),
.Y(n_220)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_220),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_204),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_221),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_SL g231 ( 
.A(n_222),
.B(n_203),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_195),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_223),
.A2(n_213),
.B1(n_217),
.B2(n_222),
.Y(n_242)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_198),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_225),
.A2(n_228),
.B1(n_229),
.B2(n_218),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_194),
.B(n_174),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_226),
.B(n_227),
.Y(n_233)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_195),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_194),
.B(n_176),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_197),
.A2(n_170),
.B1(n_188),
.B2(n_177),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_218),
.B(n_201),
.C(n_200),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_230),
.B(n_244),
.C(n_4),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_231),
.B(n_11),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_232),
.A2(n_239),
.B1(n_242),
.B2(n_5),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_214),
.A2(n_215),
.B(n_212),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_235),
.B(n_10),
.C(n_11),
.Y(n_252)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_237),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_223),
.A2(n_192),
.B1(n_208),
.B2(n_206),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_216),
.A2(n_192),
.B1(n_193),
.B2(n_211),
.Y(n_240)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_240),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_221),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_241),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_218),
.B(n_4),
.C(n_5),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_245),
.B(n_250),
.C(n_255),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_236),
.B(n_12),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_246),
.B(n_252),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_230),
.B(n_12),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_247),
.B(n_254),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_239),
.B(n_4),
.C(n_5),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_251),
.B(n_244),
.Y(n_261)
);

XNOR2x1_ASAP7_75t_L g266 ( 
.A(n_253),
.B(n_7),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_234),
.B(n_10),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_231),
.B(n_5),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_235),
.B(n_6),
.C(n_7),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_256),
.B(n_233),
.C(n_232),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_257),
.B(n_243),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_260),
.B(n_262),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_261),
.B(n_264),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_250),
.B(n_238),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_263),
.B(n_7),
.C(n_8),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_245),
.B(n_233),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_256),
.B(n_240),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_265),
.B(n_268),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_266),
.A2(n_255),
.B1(n_251),
.B2(n_9),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_248),
.B(n_9),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_258),
.B(n_249),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_269),
.A2(n_275),
.B(n_267),
.Y(n_278)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_270),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_273),
.B(n_276),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_263),
.B(n_7),
.C(n_8),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_259),
.B(n_8),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_271),
.B(n_259),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_277),
.B(n_278),
.C(n_274),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_274),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_280),
.A2(n_266),
.B(n_272),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_282),
.B(n_283),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_284),
.Y(n_285)
);

BUFx24_ASAP7_75t_SL g286 ( 
.A(n_285),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_286),
.B(n_279),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_287),
.B(n_281),
.Y(n_288)
);


endmodule