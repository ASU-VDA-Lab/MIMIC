module real_jpeg_15819_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_288;
wire n_78;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_470;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_155;
wire n_120;
wire n_405;
wire n_319;
wire n_493;
wire n_93;
wire n_242;
wire n_487;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_0),
.A2(n_19),
.B(n_495),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_0),
.B(n_496),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_1),
.A2(n_14),
.B1(n_44),
.B2(n_45),
.Y(n_43)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_1),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_1),
.B(n_142),
.Y(n_141)
);

AND2x2_ASAP7_75t_SL g158 ( 
.A(n_1),
.B(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_1),
.B(n_370),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_1),
.B(n_389),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_1),
.B(n_414),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_2),
.Y(n_62)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_2),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_2),
.Y(n_160)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_2),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_3),
.B(n_39),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_3),
.B(n_83),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_3),
.B(n_113),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_3),
.B(n_123),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_3),
.B(n_138),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_3),
.B(n_197),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_3),
.B(n_318),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_3),
.B(n_453),
.Y(n_452)
);

AND2x2_ASAP7_75t_SL g58 ( 
.A(n_4),
.B(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_4),
.B(n_72),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_4),
.B(n_109),
.Y(n_108)
);

AND2x2_ASAP7_75t_SL g161 ( 
.A(n_4),
.B(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_4),
.B(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_4),
.B(n_343),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_4),
.B(n_349),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_4),
.B(n_156),
.Y(n_386)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_5),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_5),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_5),
.Y(n_168)
);

BUFx5_ASAP7_75t_L g346 ( 
.A(n_5),
.Y(n_346)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_5),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_6),
.B(n_76),
.Y(n_75)
);

NAND2x1p5_ASAP7_75t_L g96 ( 
.A(n_6),
.B(n_72),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_6),
.B(n_127),
.Y(n_126)
);

AND2x2_ASAP7_75t_SL g131 ( 
.A(n_6),
.B(n_132),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_6),
.B(n_166),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_6),
.B(n_204),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_6),
.B(n_209),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_6),
.B(n_303),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_7),
.B(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_7),
.B(n_238),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_7),
.B(n_272),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_7),
.B(n_367),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_7),
.B(n_401),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_7),
.B(n_422),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_7),
.B(n_428),
.Y(n_427)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g127 ( 
.A(n_8),
.Y(n_127)
);

BUFx5_ASAP7_75t_L g156 ( 
.A(n_8),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_9),
.B(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_9),
.B(n_70),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_9),
.B(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_9),
.B(n_155),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_9),
.B(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_9),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_10),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_10),
.Y(n_106)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_10),
.Y(n_140)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_10),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_10),
.Y(n_270)
);

INVxp33_ASAP7_75t_L g496 ( 
.A(n_11),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_12),
.Y(n_66)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_12),
.Y(n_111)
);

BUFx5_ASAP7_75t_L g144 ( 
.A(n_12),
.Y(n_144)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_12),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_13),
.B(n_31),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_13),
.B(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_13),
.B(n_232),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_13),
.B(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_13),
.B(n_362),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_13),
.B(n_166),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_13),
.B(n_412),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_13),
.B(n_414),
.Y(n_430)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_14),
.B(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_14),
.B(n_95),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_14),
.B(n_162),
.Y(n_220)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_14),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_14),
.B(n_322),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_14),
.B(n_451),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_14),
.B(n_493),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_15),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_16),
.Y(n_125)
);

BUFx4f_ASAP7_75t_L g211 ( 
.A(n_16),
.Y(n_211)
);

BUFx8_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_17),
.Y(n_81)
);

BUFx5_ASAP7_75t_L g303 ( 
.A(n_17),
.Y(n_303)
);

BUFx5_ASAP7_75t_L g455 ( 
.A(n_17),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_470),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_437),
.B(n_469),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2x1_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_328),
.Y(n_22)
);

A2O1A1O1Ixp25_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_224),
.B(n_287),
.C(n_288),
.D(n_327),
.Y(n_23)
);

NAND4xp25_ASAP7_75t_L g328 ( 
.A(n_24),
.B(n_288),
.C(n_329),
.D(n_331),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_177),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_25),
.B(n_177),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_101),
.C(n_147),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_26),
.A2(n_27),
.B1(n_102),
.B2(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_27),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_67),
.Y(n_27)
);

INVxp33_ASAP7_75t_SL g179 ( 
.A(n_28),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_42),
.C(n_50),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_29),
.B(n_279),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_32),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_30),
.B(n_34),
.C(n_38),
.Y(n_90)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_31),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g485 ( 
.A(n_31),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_34),
.B1(n_38),
.B2(n_41),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_37),
.Y(n_350)
);

INVx1_ASAP7_75t_SL g41 ( 
.A(n_38),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_38),
.B(n_208),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_39),
.Y(n_249)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_41),
.B(n_208),
.Y(n_340)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_42),
.A2(n_43),
.B1(n_50),
.B2(n_51),
.Y(n_279)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_43),
.A2(n_241),
.B(n_246),
.Y(n_240)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_48),
.Y(n_273)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g197 ( 
.A(n_49),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_49),
.Y(n_245)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_58),
.C(n_63),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_52),
.B(n_63),
.Y(n_150)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx4_ASAP7_75t_L g390 ( 
.A(n_57),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_57),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_58),
.B(n_150),
.Y(n_149)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_62),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_62),
.Y(n_219)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_66),
.Y(n_319)
);

INVx4_ASAP7_75t_L g464 ( 
.A(n_66),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_68),
.A2(n_89),
.B1(n_99),
.B2(n_100),
.Y(n_67)
);

INVxp67_ASAP7_75t_SL g99 ( 
.A(n_68),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_68),
.Y(n_180)
);

A2O1A1Ixp33_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_71),
.B(n_74),
.C(n_86),
.Y(n_68)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_69),
.A2(n_71),
.B1(n_87),
.B2(n_88),
.Y(n_176)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

INVx6_ASAP7_75t_L g313 ( 
.A(n_72),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_73),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_74),
.B(n_176),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_78),
.C(n_82),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_75),
.A2(n_82),
.B1(n_252),
.B2(n_253),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_75),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_75),
.A2(n_165),
.B1(n_252),
.B2(n_262),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_75),
.B(n_262),
.C(n_462),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_75),
.A2(n_130),
.B1(n_131),
.B2(n_252),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_78),
.B(n_251),
.Y(n_250)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_81),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_82),
.B(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_82),
.Y(n_253)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_88),
.Y(n_86)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_89),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_90),
.A2(n_91),
.B1(n_92),
.B2(n_98),
.Y(n_89)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_90),
.Y(n_98)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_94),
.B1(n_96),
.B2(n_97),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_93),
.B(n_97),
.C(n_98),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_96),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_100),
.Y(n_181)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_102),
.Y(n_285)
);

XNOR2x1_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_115),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_103),
.B(n_129),
.C(n_145),
.Y(n_185)
);

XNOR2x2_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_107),
.Y(n_103)
);

MAJx2_ASAP7_75t_L g198 ( 
.A(n_104),
.B(n_108),
.C(n_112),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_SL g107 ( 
.A(n_108),
.B(n_112),
.Y(n_107)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_110),
.Y(n_493)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_111),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_112),
.A2(n_448),
.B1(n_449),
.B2(n_450),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_112),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_112),
.B(n_449),
.C(n_452),
.Y(n_489)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_114),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_129),
.B1(n_145),
.B2(n_146),
.Y(n_115)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_116),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_120),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_117),
.B(n_121),
.C(n_128),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_119),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_118),
.B(n_242),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_118),
.B(n_269),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_122),
.B1(n_126),
.B2(n_128),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_121),
.A2(n_122),
.B1(n_153),
.B2(n_154),
.Y(n_263)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_122),
.B(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_126),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_126),
.A2(n_128),
.B1(n_208),
.B2(n_212),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_126),
.B(n_348),
.Y(n_392)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_127),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_128),
.B(n_203),
.C(n_208),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_128),
.B(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_129),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_136),
.C(n_141),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_130),
.A2(n_131),
.B1(n_141),
.B2(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_136),
.A2(n_137),
.B1(n_171),
.B2(n_172),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_136),
.A2(n_137),
.B1(n_321),
.B2(n_326),
.Y(n_320)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_137),
.B(n_317),
.C(n_326),
.Y(n_466)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_140),
.Y(n_402)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_141),
.Y(n_173)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_147),
.B(n_284),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_169),
.C(n_174),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_148),
.B(n_276),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_151),
.C(n_157),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_149),
.B(n_256),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_151),
.A2(n_152),
.B1(n_157),
.B2(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

BUFx12f_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_157),
.Y(n_257)
);

MAJx2_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_161),
.C(n_165),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_158),
.A2(n_165),
.B1(n_261),
.B2(n_262),
.Y(n_260)
);

CKINVDCx14_ASAP7_75t_R g261 ( 
.A(n_158),
.Y(n_261)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_161),
.B(n_260),
.Y(n_259)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_SL g262 ( 
.A(n_165),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_165),
.A2(n_208),
.B1(n_212),
.B2(n_262),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_165),
.B(n_212),
.C(n_311),
.Y(n_467)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx8_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_170),
.B(n_175),
.Y(n_276)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_182),
.Y(n_177)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_178),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_180),
.C(n_181),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_183),
.A2(n_201),
.B1(n_222),
.B2(n_223),
.Y(n_182)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_183),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_185),
.B1(n_186),
.B2(n_200),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_184),
.B(n_187),
.C(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_186),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_188),
.B1(n_189),
.B2(n_199),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_189),
.Y(n_199)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_189),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_198),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_192),
.B1(n_195),
.B2(n_196),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

MAJx2_ASAP7_75t_L g299 ( 
.A(n_192),
.B(n_195),
.C(n_198),
.Y(n_299)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g490 ( 
.A1(n_195),
.A2(n_196),
.B1(n_491),
.B2(n_492),
.Y(n_490)
);

INVx2_ASAP7_75t_SL g195 ( 
.A(n_196),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_196),
.B(n_302),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_196),
.B(n_306),
.C(n_458),
.Y(n_457)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_201),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_201),
.B(n_222),
.C(n_290),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_213),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_202),
.B(n_214),
.C(n_215),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_207),
.Y(n_202)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_208),
.Y(n_212)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_218),
.B1(n_220),
.B2(n_221),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_217),
.B(n_221),
.C(n_253),
.Y(n_315)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_218),
.Y(n_217)
);

INVx5_ASAP7_75t_L g368 ( 
.A(n_219),
.Y(n_368)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_220),
.Y(n_221)
);

OAI21x1_ASAP7_75t_SL g224 ( 
.A1(n_225),
.A2(n_281),
.B(n_286),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_274),
.Y(n_225)
);

NOR2x1_ASAP7_75t_L g330 ( 
.A(n_226),
.B(n_274),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_254),
.C(n_258),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_227),
.B(n_352),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_228),
.B(n_239),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_228),
.B(n_240),
.C(n_250),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.C(n_236),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_229),
.B(n_338),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_230),
.A2(n_231),
.B1(n_236),
.B2(n_237),
.Y(n_338)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_250),
.Y(n_239)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_254),
.A2(n_255),
.B1(n_258),
.B2(n_353),
.Y(n_352)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_258),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_263),
.C(n_264),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_SL g335 ( 
.A(n_259),
.B(n_336),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_263),
.B(n_264),
.Y(n_336)
);

MAJx2_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_268),
.C(n_271),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_265),
.B(n_271),
.Y(n_374)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_268),
.B(n_374),
.Y(n_373)
);

INVx4_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx4_ASAP7_75t_L g365 ( 
.A(n_270),
.Y(n_365)
);

INVx4_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx8_ASAP7_75t_L g451 ( 
.A(n_273),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_277),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_275),
.B(n_278),
.C(n_280),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_280),
.Y(n_277)
);

NOR2x1_ASAP7_75t_L g329 ( 
.A(n_281),
.B(n_330),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

OR2x2_ASAP7_75t_L g286 ( 
.A(n_282),
.B(n_283),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_291),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_289),
.B(n_291),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_294),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_292),
.B(n_295),
.C(n_308),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_308),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_296),
.A2(n_297),
.B1(n_298),
.B2(n_307),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_296),
.B(n_299),
.C(n_300),
.Y(n_440)
);

INVx1_ASAP7_75t_SL g296 ( 
.A(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_298),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_SL g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

AO22x1_ASAP7_75t_SL g300 ( 
.A1(n_301),
.A2(n_304),
.B1(n_305),
.B2(n_306),
.Y(n_300)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_301),
.Y(n_305)
);

CKINVDCx14_ASAP7_75t_R g458 ( 
.A(n_302),
.Y(n_458)
);

INVx1_ASAP7_75t_SL g306 ( 
.A(n_304),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_314),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_309),
.B(n_315),
.C(n_316),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_SL g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_313),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_312),
.B(n_463),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_312),
.B(n_484),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_320),
.Y(n_316)
);

INVx1_ASAP7_75t_SL g318 ( 
.A(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_SL g326 ( 
.A(n_321),
.Y(n_326)
);

BUFx2_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_332),
.A2(n_354),
.B(n_436),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_351),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_333),
.B(n_351),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_337),
.C(n_339),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_334),
.A2(n_335),
.B1(n_376),
.B2(n_377),
.Y(n_375)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_SL g377 ( 
.A(n_337),
.B(n_339),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_341),
.C(n_347),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_340),
.A2(n_341),
.B1(n_342),
.B2(n_359),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_340),
.Y(n_359)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

BUFx2_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_345),
.Y(n_424)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_SL g357 ( 
.A(n_347),
.B(n_358),
.Y(n_357)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_349),
.Y(n_429)
);

INVx5_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

AOI21x1_ASAP7_75t_SL g354 ( 
.A1(n_355),
.A2(n_378),
.B(n_435),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_375),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_SL g435 ( 
.A(n_356),
.B(n_375),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_360),
.C(n_373),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_357),
.B(n_394),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_360),
.B(n_373),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_366),
.C(n_369),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_361),
.B(n_383),
.Y(n_382)
);

INVx1_ASAP7_75t_SL g362 ( 
.A(n_363),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_366),
.B(n_369),
.Y(n_383)
);

INVx5_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx4_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

BUFx3_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

OAI21x1_ASAP7_75t_L g378 ( 
.A1(n_379),
.A2(n_395),
.B(n_434),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_393),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_380),
.B(n_393),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_384),
.C(n_391),
.Y(n_380)
);

AOI22xp33_ASAP7_75t_SL g404 ( 
.A1(n_381),
.A2(n_382),
.B1(n_405),
.B2(n_407),
.Y(n_404)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_384),
.A2(n_391),
.B1(n_392),
.B2(n_406),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_384),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_387),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_385),
.A2(n_386),
.B1(n_387),
.B2(n_388),
.Y(n_398)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_L g395 ( 
.A1(n_396),
.A2(n_408),
.B(n_433),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_404),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_SL g433 ( 
.A(n_397),
.B(n_404),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_399),
.C(n_403),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_398),
.B(n_417),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_399),
.A2(n_400),
.B1(n_403),
.B2(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

HB1xp67_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

CKINVDCx16_ASAP7_75t_R g418 ( 
.A(n_403),
.Y(n_418)
);

INVxp67_ASAP7_75t_SL g407 ( 
.A(n_405),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_SL g408 ( 
.A1(n_409),
.A2(n_419),
.B(n_432),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_416),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_410),
.B(n_416),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_413),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_411),
.B(n_413),
.Y(n_425)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

AOI21xp5_ASAP7_75t_L g419 ( 
.A1(n_420),
.A2(n_426),
.B(n_431),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_421),
.B(n_425),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_SL g431 ( 
.A(n_421),
.B(n_425),
.Y(n_431)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_430),
.Y(n_426)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

CKINVDCx14_ASAP7_75t_R g437 ( 
.A(n_438),
.Y(n_437)
);

OR2x6_ASAP7_75t_SL g438 ( 
.A(n_439),
.B(n_468),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_439),
.B(n_468),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_440),
.B(n_441),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_440),
.B(n_442),
.C(n_459),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_459),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_443),
.B(n_444),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_443),
.B(n_445),
.C(n_457),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_457),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_446),
.A2(n_447),
.B1(n_452),
.B2(n_456),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_452),
.Y(n_456)
);

INVx1_ASAP7_75t_SL g453 ( 
.A(n_454),
.Y(n_453)
);

INVx8_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_460),
.B(n_465),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_460),
.B(n_466),
.C(n_467),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_462),
.Y(n_460)
);

HB1xp67_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_466),
.B(n_467),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_471),
.B(n_494),
.Y(n_470)
);

INVxp33_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_473),
.B(n_474),
.Y(n_472)
);

NOR2xp67_ASAP7_75t_SL g494 ( 
.A(n_473),
.B(n_474),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_475),
.B(n_476),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_477),
.B(n_478),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_479),
.A2(n_480),
.B1(n_487),
.B2(n_488),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_SL g480 ( 
.A(n_481),
.B(n_482),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_483),
.B(n_486),
.Y(n_482)
);

INVx4_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_SL g488 ( 
.A(n_489),
.B(n_490),
.Y(n_488)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);


endmodule