module fake_jpeg_26434_n_164 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_164);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_164;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx4f_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_4),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_5),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_8),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g53 ( 
.A(n_30),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

BUFx4f_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

BUFx24_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_11),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_6),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_11),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_13),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_8),
.Y(n_63)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_14),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_1),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_51),
.B(n_0),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_70),
.B(n_66),
.Y(n_76)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_73),
.Y(n_74)
);

INVx6_ASAP7_75t_SL g75 ( 
.A(n_72),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_76),
.B(n_0),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_49),
.Y(n_77)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_77),
.Y(n_92)
);

INVx2_ASAP7_75t_R g82 ( 
.A(n_69),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_82),
.B(n_67),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_73),
.A2(n_46),
.B1(n_64),
.B2(n_61),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_84),
.A2(n_52),
.B1(n_2),
.B2(n_3),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_71),
.A2(n_63),
.B1(n_55),
.B2(n_45),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_85),
.A2(n_63),
.B1(n_68),
.B2(n_51),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_60),
.Y(n_86)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_86),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_67),
.B(n_59),
.Y(n_87)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_90),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_89),
.A2(n_94),
.B1(n_6),
.B2(n_7),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_82),
.B(n_66),
.Y(n_90)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_84),
.B(n_68),
.Y(n_93)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_93),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_85),
.A2(n_53),
.B1(n_65),
.B2(n_48),
.Y(n_94)
);

AO22x1_ASAP7_75t_L g95 ( 
.A1(n_74),
.A2(n_50),
.B1(n_56),
.B2(n_58),
.Y(n_95)
);

OA22x2_ASAP7_75t_L g107 ( 
.A1(n_95),
.A2(n_96),
.B1(n_99),
.B2(n_81),
.Y(n_107)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_75),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_L g97 ( 
.A1(n_80),
.A2(n_62),
.B1(n_54),
.B2(n_28),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_97),
.A2(n_80),
.B1(n_78),
.B2(n_83),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_98),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_79),
.B(n_1),
.Y(n_99)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_101),
.Y(n_110)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_74),
.Y(n_104)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_104),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_105),
.B(n_107),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_111),
.B(n_113),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_88),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_114),
.A2(n_100),
.B1(n_97),
.B2(n_103),
.Y(n_117)
);

BUFx24_ASAP7_75t_L g116 ( 
.A(n_112),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_116),
.B(n_102),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_117),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_106),
.B(n_109),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_119),
.B(n_120),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_108),
.B(n_93),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_105),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_121),
.B(n_123),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_110),
.B(n_92),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_122),
.B(n_124),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_114),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_107),
.B(n_96),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_120),
.B(n_107),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_125),
.A2(n_131),
.B(n_139),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_115),
.A2(n_99),
.B(n_102),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_126),
.A2(n_125),
.B(n_138),
.Y(n_145)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_128),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_118),
.B(n_95),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_129),
.Y(n_149)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_116),
.Y(n_130)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_130),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_116),
.Y(n_131)
);

OAI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_117),
.A2(n_31),
.B1(n_44),
.B2(n_43),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_132),
.A2(n_136),
.B1(n_22),
.B2(n_23),
.Y(n_144)
);

OAI32xp33_ASAP7_75t_L g133 ( 
.A1(n_115),
.A2(n_7),
.A3(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_133)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_133),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_120),
.B(n_26),
.C(n_42),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_135),
.B(n_19),
.C(n_20),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_122),
.B(n_33),
.Y(n_137)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_137),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_119),
.B(n_13),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_127),
.A2(n_15),
.B1(n_16),
.B2(n_18),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_142),
.Y(n_152)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_143),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_144),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_151),
.B(n_145),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_153),
.A2(n_154),
.B1(n_149),
.B2(n_126),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_150),
.A2(n_148),
.B1(n_145),
.B2(n_144),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_153),
.C(n_147),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_140),
.C(n_134),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_157),
.A2(n_146),
.B1(n_152),
.B2(n_132),
.Y(n_158)
);

AOI31xp67_ASAP7_75t_L g159 ( 
.A1(n_158),
.A2(n_141),
.A3(n_135),
.B(n_36),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_159),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_160),
.B(n_143),
.Y(n_161)
);

NOR3x1_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_32),
.C(n_34),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_37),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_38),
.Y(n_164)
);


endmodule