module fake_jpeg_2892_n_119 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_119);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_119;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_4),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_1),
.B(n_2),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx10_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_5),
.B(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx4_ASAP7_75t_SL g54 ( 
.A(n_29),
.Y(n_54)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_12),
.B(n_19),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_31),
.B(n_3),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_11),
.B(n_8),
.Y(n_32)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_34),
.Y(n_47)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_11),
.B(n_9),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_38),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_17),
.B(n_0),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_40),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_17),
.B(n_0),
.Y(n_40)
);

OA22x2_ASAP7_75t_L g44 ( 
.A1(n_30),
.A2(n_35),
.B1(n_26),
.B2(n_36),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_44),
.A2(n_53),
.B1(n_58),
.B2(n_29),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_28),
.A2(n_25),
.B1(n_13),
.B2(n_22),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_46),
.A2(n_56),
.B1(n_58),
.B2(n_44),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_32),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_49),
.B(n_5),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_31),
.B(n_25),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_59),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_27),
.A2(n_24),
.B1(n_15),
.B2(n_20),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_28),
.A2(n_23),
.B1(n_20),
.B2(n_24),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_55),
.A2(n_33),
.B1(n_39),
.B2(n_29),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_36),
.A2(n_13),
.B1(n_22),
.B2(n_18),
.Y(n_56)
);

OA22x2_ASAP7_75t_L g58 ( 
.A1(n_37),
.A2(n_15),
.B1(n_16),
.B2(n_23),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_34),
.B(n_0),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_61),
.B(n_3),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_62),
.B(n_64),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_61),
.B(n_29),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_63),
.B(n_75),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_49),
.B(n_3),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_39),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_66),
.B(n_67),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_39),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_68),
.A2(n_77),
.B1(n_56),
.B2(n_54),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_70),
.B(n_44),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_72),
.B(n_76),
.Y(n_81)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_73),
.Y(n_80)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_50),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_6),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_58),
.A2(n_6),
.B1(n_16),
.B2(n_45),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_78),
.A2(n_79),
.B1(n_87),
.B2(n_54),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_58),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_83),
.B(n_70),
.C(n_75),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_77),
.A2(n_44),
.B1(n_57),
.B2(n_48),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_65),
.B(n_48),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_88),
.B(n_64),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_91),
.B(n_93),
.Y(n_103)
);

NOR3xp33_ASAP7_75t_L g100 ( 
.A(n_92),
.B(n_94),
.C(n_95),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_90),
.B(n_73),
.C(n_74),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_90),
.B(n_62),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_86),
.A2(n_69),
.B(n_68),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_96),
.B(n_98),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_85),
.B(n_69),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_97),
.B(n_99),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_52),
.C(n_43),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_78),
.A2(n_83),
.B1(n_88),
.B2(n_80),
.Y(n_99)
);

A2O1A1O1Ixp25_ASAP7_75t_L g102 ( 
.A1(n_91),
.A2(n_83),
.B(n_78),
.C(n_81),
.D(n_84),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_102),
.B(n_101),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_81),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_98),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_106),
.B(n_109),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_103),
.B(n_80),
.C(n_89),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_107),
.B(n_108),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_101),
.A2(n_89),
.B1(n_82),
.B2(n_57),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_100),
.Y(n_110)
);

AOI322xp5_ASAP7_75t_L g111 ( 
.A1(n_110),
.A2(n_104),
.A3(n_102),
.B1(n_103),
.B2(n_82),
.C1(n_41),
.C2(n_50),
.Y(n_111)
);

AOI31xp67_ASAP7_75t_L g114 ( 
.A1(n_111),
.A2(n_107),
.A3(n_108),
.B(n_43),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_114),
.B(n_115),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_113),
.B(n_6),
.Y(n_115)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_116),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_112),
.C(n_41),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_112),
.Y(n_119)
);


endmodule