module fake_netlist_1_3968_n_584 (n_44, n_81, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_584);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_584;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_461;
wire n_305;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_540;
wire n_563;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_554;
wire n_447;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_583;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_493;
wire n_418;
wire n_555;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx2_ASAP7_75t_L g82 ( .A(n_62), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_18), .Y(n_83) );
CKINVDCx5p33_ASAP7_75t_R g84 ( .A(n_54), .Y(n_84) );
BUFx6f_ASAP7_75t_L g85 ( .A(n_10), .Y(n_85) );
NOR2xp67_ASAP7_75t_L g86 ( .A(n_68), .B(n_64), .Y(n_86) );
CKINVDCx5p33_ASAP7_75t_R g87 ( .A(n_1), .Y(n_87) );
CKINVDCx5p33_ASAP7_75t_R g88 ( .A(n_59), .Y(n_88) );
BUFx3_ASAP7_75t_L g89 ( .A(n_19), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_16), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_5), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_75), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_2), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_30), .Y(n_94) );
INVx2_ASAP7_75t_L g95 ( .A(n_76), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_44), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_8), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_7), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_36), .Y(n_99) );
BUFx2_ASAP7_75t_SL g100 ( .A(n_53), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_65), .Y(n_101) );
INVx2_ASAP7_75t_SL g102 ( .A(n_15), .Y(n_102) );
CKINVDCx14_ASAP7_75t_R g103 ( .A(n_24), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_58), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_73), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_12), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_80), .Y(n_107) );
CKINVDCx16_ASAP7_75t_R g108 ( .A(n_56), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_39), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_14), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_69), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_60), .Y(n_112) );
BUFx2_ASAP7_75t_L g113 ( .A(n_37), .Y(n_113) );
INVxp67_ASAP7_75t_SL g114 ( .A(n_78), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_5), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_50), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_51), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_63), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_26), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_6), .Y(n_120) );
NAND2xp33_ASAP7_75t_L g121 ( .A(n_84), .B(n_32), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_92), .Y(n_122) );
AOI22xp5_ASAP7_75t_L g123 ( .A1(n_87), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_92), .Y(n_124) );
BUFx6f_ASAP7_75t_L g125 ( .A(n_89), .Y(n_125) );
INVx4_ASAP7_75t_L g126 ( .A(n_113), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_82), .Y(n_127) );
INVx2_ASAP7_75t_L g128 ( .A(n_82), .Y(n_128) );
OAI22xp5_ASAP7_75t_L g129 ( .A1(n_83), .A2(n_0), .B1(n_3), .B2(n_4), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_94), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_113), .B(n_102), .Y(n_131) );
NOR2xp33_ASAP7_75t_SL g132 ( .A(n_108), .B(n_34), .Y(n_132) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_89), .Y(n_133) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_85), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_95), .Y(n_135) );
OA21x2_ASAP7_75t_L g136 ( .A1(n_94), .A2(n_33), .B(n_79), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_95), .Y(n_137) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_85), .Y(n_138) );
NAND2x1_ASAP7_75t_L g139 ( .A(n_102), .B(n_3), .Y(n_139) );
OA21x2_ASAP7_75t_L g140 ( .A1(n_96), .A2(n_35), .B(n_77), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_96), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_99), .Y(n_142) );
HB1xp67_ASAP7_75t_L g143 ( .A(n_87), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_101), .Y(n_144) );
AND2x6_ASAP7_75t_L g145 ( .A(n_122), .B(n_83), .Y(n_145) );
OAI22xp5_ASAP7_75t_SL g146 ( .A1(n_123), .A2(n_120), .B1(n_90), .B2(n_93), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_134), .Y(n_147) );
INVx3_ASAP7_75t_L g148 ( .A(n_127), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_127), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_126), .B(n_105), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_126), .B(n_107), .Y(n_151) );
NAND2xp5_ASAP7_75t_SL g152 ( .A(n_122), .B(n_109), .Y(n_152) );
NAND2xp5_ASAP7_75t_SL g153 ( .A(n_126), .B(n_84), .Y(n_153) );
AND2x4_ASAP7_75t_L g154 ( .A(n_126), .B(n_124), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_124), .B(n_111), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_134), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_128), .Y(n_157) );
INVx2_ASAP7_75t_SL g158 ( .A(n_130), .Y(n_158) );
NOR2xp33_ASAP7_75t_L g159 ( .A(n_131), .B(n_112), .Y(n_159) );
NOR3xp33_ASAP7_75t_L g160 ( .A(n_129), .B(n_106), .C(n_91), .Y(n_160) );
INVx2_ASAP7_75t_SL g161 ( .A(n_130), .Y(n_161) );
BUFx3_ASAP7_75t_L g162 ( .A(n_125), .Y(n_162) );
INVx4_ASAP7_75t_L g163 ( .A(n_125), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_134), .Y(n_164) );
AND2x2_ASAP7_75t_L g165 ( .A(n_141), .B(n_103), .Y(n_165) );
INVx5_ASAP7_75t_L g166 ( .A(n_125), .Y(n_166) );
AOI22xp33_ASAP7_75t_L g167 ( .A1(n_141), .A2(n_93), .B1(n_97), .B2(n_98), .Y(n_167) );
INVx5_ASAP7_75t_L g168 ( .A(n_125), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_134), .Y(n_169) );
AND2x4_ASAP7_75t_L g170 ( .A(n_142), .B(n_97), .Y(n_170) );
INVx2_ASAP7_75t_SL g171 ( .A(n_142), .Y(n_171) );
BUFx3_ASAP7_75t_L g172 ( .A(n_125), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_158), .Y(n_173) );
AOI22xp5_ASAP7_75t_L g174 ( .A1(n_146), .A2(n_132), .B1(n_123), .B2(n_144), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_154), .B(n_143), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_162), .Y(n_176) );
NOR3xp33_ASAP7_75t_L g177 ( .A(n_146), .B(n_139), .C(n_120), .Y(n_177) );
AOI21xp5_ASAP7_75t_L g178 ( .A1(n_158), .A2(n_121), .B(n_140), .Y(n_178) );
AND2x6_ASAP7_75t_SL g179 ( .A(n_159), .B(n_98), .Y(n_179) );
CKINVDCx20_ASAP7_75t_R g180 ( .A(n_165), .Y(n_180) );
OR2x2_ASAP7_75t_L g181 ( .A(n_165), .B(n_90), .Y(n_181) );
BUFx3_ASAP7_75t_L g182 ( .A(n_154), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_154), .B(n_144), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_162), .Y(n_184) );
NOR2xp33_ASAP7_75t_SL g185 ( .A(n_165), .B(n_88), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_154), .B(n_88), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_162), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_154), .B(n_104), .Y(n_188) );
AND2x4_ASAP7_75t_L g189 ( .A(n_170), .B(n_139), .Y(n_189) );
INVx2_ASAP7_75t_SL g190 ( .A(n_170), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_158), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_161), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_172), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_153), .B(n_119), .Y(n_194) );
AOI22xp5_ASAP7_75t_L g195 ( .A1(n_160), .A2(n_115), .B1(n_110), .B2(n_137), .Y(n_195) );
INVx2_ASAP7_75t_SL g196 ( .A(n_170), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_159), .B(n_119), .Y(n_197) );
INVx8_ASAP7_75t_L g198 ( .A(n_145), .Y(n_198) );
AND2x2_ASAP7_75t_L g199 ( .A(n_170), .B(n_137), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_161), .Y(n_200) );
OAI21xp5_ASAP7_75t_L g201 ( .A1(n_161), .A2(n_140), .B(n_136), .Y(n_201) );
AOI22xp33_ASAP7_75t_L g202 ( .A1(n_160), .A2(n_85), .B1(n_133), .B2(n_135), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_150), .B(n_104), .Y(n_203) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_171), .A2(n_140), .B(n_136), .Y(n_204) );
BUFx6f_ASAP7_75t_L g205 ( .A(n_145), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_171), .B(n_118), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_150), .B(n_118), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_172), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_151), .B(n_128), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g210 ( .A(n_181), .B(n_151), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_173), .A2(n_171), .B(n_152), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_173), .A2(n_152), .B(n_155), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_191), .A2(n_155), .B(n_136), .Y(n_213) );
INVxp67_ASAP7_75t_L g214 ( .A(n_185), .Y(n_214) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_205), .B(n_170), .Y(n_215) );
OR2x6_ASAP7_75t_SL g216 ( .A(n_181), .B(n_149), .Y(n_216) );
INVxp67_ASAP7_75t_L g217 ( .A(n_197), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_203), .B(n_167), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_205), .B(n_167), .Y(n_219) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_191), .A2(n_140), .B(n_136), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_182), .Y(n_221) );
BUFx3_ASAP7_75t_L g222 ( .A(n_180), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_182), .Y(n_223) );
AOI22xp5_ASAP7_75t_L g224 ( .A1(n_180), .A2(n_145), .B1(n_149), .B2(n_157), .Y(n_224) );
OAI22xp5_ASAP7_75t_L g225 ( .A1(n_190), .A2(n_157), .B1(n_148), .B2(n_135), .Y(n_225) );
NOR2xp67_ASAP7_75t_L g226 ( .A(n_174), .B(n_148), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_192), .A2(n_163), .B(n_172), .Y(n_227) );
CKINVDCx5p33_ASAP7_75t_R g228 ( .A(n_179), .Y(n_228) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_205), .B(n_148), .Y(n_229) );
AOI22xp33_ASAP7_75t_L g230 ( .A1(n_190), .A2(n_145), .B1(n_148), .B2(n_85), .Y(n_230) );
INVx1_ASAP7_75t_SL g231 ( .A(n_199), .Y(n_231) );
BUFx2_ASAP7_75t_L g232 ( .A(n_189), .Y(n_232) );
AND2x4_ASAP7_75t_L g233 ( .A(n_189), .B(n_148), .Y(n_233) );
NOR2xp33_ASAP7_75t_L g234 ( .A(n_175), .B(n_145), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_189), .B(n_145), .Y(n_235) );
OAI22xp5_ASAP7_75t_L g236 ( .A1(n_196), .A2(n_114), .B1(n_85), .B2(n_116), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_192), .A2(n_163), .B(n_117), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_179), .B(n_145), .Y(n_238) );
AND2x4_ASAP7_75t_L g239 ( .A(n_189), .B(n_145), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_196), .B(n_145), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_200), .A2(n_178), .B(n_204), .Y(n_241) );
NAND2xp5_ASAP7_75t_SL g242 ( .A(n_205), .B(n_163), .Y(n_242) );
NAND2xp5_ASAP7_75t_SL g243 ( .A(n_205), .B(n_163), .Y(n_243) );
AOI21xp5_ASAP7_75t_L g244 ( .A1(n_200), .A2(n_163), .B(n_147), .Y(n_244) );
O2A1O1Ixp5_ASAP7_75t_L g245 ( .A1(n_201), .A2(n_169), .B(n_147), .C(n_156), .Y(n_245) );
HB1xp67_ASAP7_75t_L g246 ( .A(n_222), .Y(n_246) );
OR2x6_ASAP7_75t_L g247 ( .A(n_239), .B(n_198), .Y(n_247) );
OAI21x1_ASAP7_75t_L g248 ( .A1(n_241), .A2(n_220), .B(n_213), .Y(n_248) );
INVx2_ASAP7_75t_L g249 ( .A(n_245), .Y(n_249) );
OAI21xp5_ASAP7_75t_L g250 ( .A1(n_212), .A2(n_183), .B(n_186), .Y(n_250) );
OAI21xp5_ASAP7_75t_L g251 ( .A1(n_218), .A2(n_188), .B(n_207), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_210), .B(n_174), .Y(n_252) );
INVx3_ASAP7_75t_L g253 ( .A(n_239), .Y(n_253) );
O2A1O1Ixp33_ASAP7_75t_L g254 ( .A1(n_217), .A2(n_177), .B(n_209), .C(n_206), .Y(n_254) );
INVxp67_ASAP7_75t_SL g255 ( .A(n_232), .Y(n_255) );
AND2x2_ASAP7_75t_L g256 ( .A(n_210), .B(n_199), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_233), .Y(n_257) );
OAI22xp5_ASAP7_75t_L g258 ( .A1(n_224), .A2(n_195), .B1(n_198), .B2(n_202), .Y(n_258) );
AND2x4_ASAP7_75t_L g259 ( .A(n_226), .B(n_195), .Y(n_259) );
OR2x2_ASAP7_75t_L g260 ( .A(n_231), .B(n_194), .Y(n_260) );
NOR2x1_ASAP7_75t_SL g261 ( .A(n_215), .B(n_198), .Y(n_261) );
AO22x2_ASAP7_75t_L g262 ( .A1(n_214), .A2(n_100), .B1(n_193), .B2(n_187), .Y(n_262) );
AOI21xp5_ASAP7_75t_L g263 ( .A1(n_211), .A2(n_208), .B(n_193), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_216), .B(n_198), .Y(n_264) );
NAND3xp33_ASAP7_75t_L g265 ( .A(n_230), .B(n_133), .C(n_168), .Y(n_265) );
INVx4_ASAP7_75t_L g266 ( .A(n_233), .Y(n_266) );
OAI22xp5_ASAP7_75t_L g267 ( .A1(n_235), .A2(n_208), .B1(n_187), .B2(n_184), .Y(n_267) );
INVx1_ASAP7_75t_SL g268 ( .A(n_228), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_221), .Y(n_269) );
AOI31xp67_ASAP7_75t_L g270 ( .A1(n_219), .A2(n_147), .A3(n_156), .B(n_169), .Y(n_270) );
AOI22xp5_ASAP7_75t_L g271 ( .A1(n_238), .A2(n_145), .B1(n_176), .B2(n_184), .Y(n_271) );
A2O1A1Ixp33_ASAP7_75t_L g272 ( .A1(n_237), .A2(n_86), .B(n_100), .C(n_176), .Y(n_272) );
AOI21xp5_ASAP7_75t_L g273 ( .A1(n_244), .A2(n_169), .B(n_156), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_235), .B(n_133), .Y(n_274) );
OAI21xp5_ASAP7_75t_L g275 ( .A1(n_227), .A2(n_240), .B(n_225), .Y(n_275) );
BUFx6f_ASAP7_75t_L g276 ( .A(n_248), .Y(n_276) );
NAND2x1p5_ASAP7_75t_L g277 ( .A(n_266), .B(n_223), .Y(n_277) );
INVx6_ASAP7_75t_L g278 ( .A(n_266), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_252), .B(n_234), .Y(n_279) );
AOI21xp5_ASAP7_75t_L g280 ( .A1(n_249), .A2(n_229), .B(n_242), .Y(n_280) );
NAND2x1p5_ASAP7_75t_L g281 ( .A(n_266), .B(n_243), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_269), .Y(n_282) );
OA21x2_ASAP7_75t_L g283 ( .A1(n_248), .A2(n_230), .B(n_164), .Y(n_283) );
OAI21xp5_ASAP7_75t_L g284 ( .A1(n_251), .A2(n_236), .B(n_234), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_269), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_249), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_270), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_250), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_274), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_256), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_262), .Y(n_291) );
OAI21x1_ASAP7_75t_L g292 ( .A1(n_263), .A2(n_164), .B(n_133), .Y(n_292) );
AO31x2_ASAP7_75t_L g293 ( .A1(n_272), .A2(n_164), .A3(n_138), .B(n_134), .Y(n_293) );
NAND2x1p5_ASAP7_75t_L g294 ( .A(n_253), .B(n_168), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_262), .Y(n_295) );
AOI21x1_ASAP7_75t_L g296 ( .A1(n_262), .A2(n_133), .B(n_138), .Y(n_296) );
OAI21x1_ASAP7_75t_L g297 ( .A1(n_275), .A2(n_168), .B(n_166), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_257), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_256), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_259), .B(n_4), .Y(n_300) );
OA21x2_ASAP7_75t_L g301 ( .A1(n_287), .A2(n_272), .B(n_273), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_286), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_282), .Y(n_303) );
AND2x4_ASAP7_75t_L g304 ( .A(n_282), .B(n_259), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_286), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_286), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_285), .Y(n_307) );
HB1xp67_ASAP7_75t_L g308 ( .A(n_291), .Y(n_308) );
AND2x2_ASAP7_75t_L g309 ( .A(n_285), .B(n_259), .Y(n_309) );
AND2x2_ASAP7_75t_L g310 ( .A(n_290), .B(n_253), .Y(n_310) );
BUFx2_ASAP7_75t_L g311 ( .A(n_291), .Y(n_311) );
OR2x2_ASAP7_75t_L g312 ( .A(n_290), .B(n_264), .Y(n_312) );
AO21x2_ASAP7_75t_L g313 ( .A1(n_296), .A2(n_265), .B(n_267), .Y(n_313) );
AND2x2_ASAP7_75t_L g314 ( .A(n_299), .B(n_253), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_276), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_288), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_288), .Y(n_317) );
HB1xp67_ASAP7_75t_L g318 ( .A(n_291), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_298), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_299), .B(n_255), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_298), .Y(n_321) );
HB1xp67_ASAP7_75t_L g322 ( .A(n_300), .Y(n_322) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_300), .Y(n_323) );
AND2x2_ASAP7_75t_L g324 ( .A(n_298), .B(n_260), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_316), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_309), .B(n_276), .Y(n_326) );
AND2x2_ASAP7_75t_L g327 ( .A(n_309), .B(n_276), .Y(n_327) );
AOI22xp5_ASAP7_75t_L g328 ( .A1(n_322), .A2(n_279), .B1(n_258), .B2(n_284), .Y(n_328) );
AND2x2_ASAP7_75t_L g329 ( .A(n_319), .B(n_276), .Y(n_329) );
OAI22xp5_ASAP7_75t_L g330 ( .A1(n_323), .A2(n_295), .B1(n_289), .B2(n_277), .Y(n_330) );
AND2x2_ASAP7_75t_L g331 ( .A(n_319), .B(n_276), .Y(n_331) );
OR2x2_ASAP7_75t_L g332 ( .A(n_321), .B(n_276), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_316), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_321), .B(n_295), .Y(n_334) );
INVx3_ASAP7_75t_L g335 ( .A(n_315), .Y(n_335) );
AND2x2_ASAP7_75t_L g336 ( .A(n_303), .B(n_295), .Y(n_336) );
AND2x2_ASAP7_75t_L g337 ( .A(n_303), .B(n_293), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_302), .Y(n_338) );
HB1xp67_ASAP7_75t_L g339 ( .A(n_302), .Y(n_339) );
HB1xp67_ASAP7_75t_L g340 ( .A(n_302), .Y(n_340) );
OR2x2_ASAP7_75t_L g341 ( .A(n_317), .B(n_293), .Y(n_341) );
AND2x2_ASAP7_75t_L g342 ( .A(n_307), .B(n_293), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_307), .B(n_293), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_317), .Y(n_344) );
OR2x2_ASAP7_75t_L g345 ( .A(n_305), .B(n_293), .Y(n_345) );
NAND2x1p5_ASAP7_75t_L g346 ( .A(n_312), .B(n_304), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_305), .Y(n_347) );
BUFx3_ASAP7_75t_L g348 ( .A(n_305), .Y(n_348) );
INVx2_ASAP7_75t_SL g349 ( .A(n_306), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_306), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_306), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_304), .B(n_293), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_315), .Y(n_353) );
AND2x2_ASAP7_75t_L g354 ( .A(n_304), .B(n_287), .Y(n_354) );
INVx1_ASAP7_75t_SL g355 ( .A(n_324), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_325), .Y(n_356) );
OR2x2_ASAP7_75t_SL g357 ( .A(n_341), .B(n_308), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_325), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_338), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_338), .Y(n_360) );
NOR2xp33_ASAP7_75t_SL g361 ( .A(n_355), .B(n_312), .Y(n_361) );
BUFx2_ASAP7_75t_L g362 ( .A(n_339), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_355), .B(n_324), .Y(n_363) );
BUFx3_ASAP7_75t_L g364 ( .A(n_348), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_326), .B(n_311), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_326), .B(n_311), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_327), .B(n_308), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_327), .B(n_318), .Y(n_368) );
AND2x2_ASAP7_75t_L g369 ( .A(n_352), .B(n_318), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_333), .Y(n_370) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_339), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_352), .B(n_315), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_333), .B(n_304), .Y(n_373) );
NAND4xp25_ASAP7_75t_L g374 ( .A(n_328), .B(n_254), .C(n_320), .D(n_268), .Y(n_374) );
AND2x2_ASAP7_75t_L g375 ( .A(n_337), .B(n_301), .Y(n_375) );
NOR2xp33_ASAP7_75t_L g376 ( .A(n_346), .B(n_246), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_344), .B(n_310), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_337), .B(n_301), .Y(n_378) );
OR2x2_ASAP7_75t_L g379 ( .A(n_340), .B(n_320), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_342), .B(n_301), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_344), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_342), .B(n_301), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_343), .B(n_310), .Y(n_383) );
INVx2_ASAP7_75t_SL g384 ( .A(n_348), .Y(n_384) );
OR2x2_ASAP7_75t_L g385 ( .A(n_340), .B(n_314), .Y(n_385) );
INVx1_ASAP7_75t_SL g386 ( .A(n_348), .Y(n_386) );
OR2x2_ASAP7_75t_L g387 ( .A(n_349), .B(n_314), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_328), .B(n_289), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_343), .Y(n_389) );
AND2x4_ASAP7_75t_L g390 ( .A(n_354), .B(n_287), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_329), .B(n_283), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_329), .B(n_283), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_331), .B(n_283), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_347), .Y(n_394) );
OR2x2_ASAP7_75t_L g395 ( .A(n_349), .B(n_313), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_347), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_350), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_338), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_350), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_346), .B(n_284), .Y(n_400) );
OR2x2_ASAP7_75t_L g401 ( .A(n_349), .B(n_313), .Y(n_401) );
OR2x2_ASAP7_75t_L g402 ( .A(n_389), .B(n_341), .Y(n_402) );
OR2x2_ASAP7_75t_L g403 ( .A(n_363), .B(n_332), .Y(n_403) );
NOR2x1_ASAP7_75t_L g404 ( .A(n_374), .B(n_330), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_356), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_372), .B(n_354), .Y(n_406) );
OR2x2_ASAP7_75t_L g407 ( .A(n_379), .B(n_332), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_389), .B(n_336), .Y(n_408) );
OR2x2_ASAP7_75t_L g409 ( .A(n_379), .B(n_351), .Y(n_409) );
NOR2x1_ASAP7_75t_L g410 ( .A(n_374), .B(n_330), .Y(n_410) );
OAI21xp33_ASAP7_75t_SL g411 ( .A1(n_384), .A2(n_351), .B(n_345), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_359), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_359), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_361), .B(n_336), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_372), .B(n_331), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_359), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_383), .B(n_334), .Y(n_417) );
OR2x2_ASAP7_75t_L g418 ( .A(n_385), .B(n_346), .Y(n_418) );
OR2x2_ASAP7_75t_L g419 ( .A(n_357), .B(n_345), .Y(n_419) );
NOR2xp33_ASAP7_75t_L g420 ( .A(n_388), .B(n_6), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_383), .B(n_334), .Y(n_421) );
INVx2_ASAP7_75t_SL g422 ( .A(n_371), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_377), .B(n_353), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_356), .B(n_353), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_375), .B(n_353), .Y(n_425) );
INVx2_ASAP7_75t_SL g426 ( .A(n_362), .Y(n_426) );
NOR2xp33_ASAP7_75t_L g427 ( .A(n_376), .B(n_7), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_358), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_358), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_370), .B(n_335), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_370), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_375), .B(n_335), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_378), .B(n_335), .Y(n_433) );
AND2x4_ASAP7_75t_SL g434 ( .A(n_367), .B(n_335), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_381), .Y(n_435) );
AND2x4_ASAP7_75t_SL g436 ( .A(n_367), .B(n_247), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_360), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_381), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_394), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_378), .B(n_296), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_394), .Y(n_441) );
OR2x2_ASAP7_75t_L g442 ( .A(n_357), .B(n_313), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_380), .B(n_313), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_396), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_360), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_380), .B(n_297), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_396), .Y(n_447) );
INVx3_ASAP7_75t_L g448 ( .A(n_364), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_397), .Y(n_449) );
OR2x2_ASAP7_75t_L g450 ( .A(n_385), .B(n_138), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_382), .B(n_297), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_397), .Y(n_452) );
BUFx2_ASAP7_75t_L g453 ( .A(n_362), .Y(n_453) );
BUFx2_ASAP7_75t_L g454 ( .A(n_364), .Y(n_454) );
INVx3_ASAP7_75t_SL g455 ( .A(n_384), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_382), .B(n_283), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_453), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_421), .B(n_369), .Y(n_458) );
OAI22xp33_ASAP7_75t_L g459 ( .A1(n_419), .A2(n_387), .B1(n_364), .B2(n_386), .Y(n_459) );
HB1xp67_ASAP7_75t_L g460 ( .A(n_422), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_450), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_450), .Y(n_462) );
INVx1_ASAP7_75t_SL g463 ( .A(n_455), .Y(n_463) );
AND2x4_ASAP7_75t_L g464 ( .A(n_434), .B(n_369), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_412), .Y(n_465) );
HB1xp67_ASAP7_75t_L g466 ( .A(n_422), .Y(n_466) );
NOR2xp33_ASAP7_75t_L g467 ( .A(n_411), .B(n_373), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_405), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_421), .B(n_365), .Y(n_469) );
AOI32xp33_ASAP7_75t_L g470 ( .A1(n_404), .A2(n_366), .A3(n_365), .B1(n_368), .B2(n_391), .Y(n_470) );
NOR2xp33_ASAP7_75t_L g471 ( .A(n_420), .B(n_387), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_428), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_417), .B(n_368), .Y(n_473) );
OR2x2_ASAP7_75t_L g474 ( .A(n_403), .B(n_366), .Y(n_474) );
OR2x2_ASAP7_75t_L g475 ( .A(n_407), .B(n_399), .Y(n_475) );
AND2x2_ASAP7_75t_SL g476 ( .A(n_434), .B(n_399), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_429), .Y(n_477) );
INVxp67_ASAP7_75t_SL g478 ( .A(n_440), .Y(n_478) );
AOI321xp33_ASAP7_75t_L g479 ( .A1(n_410), .A2(n_400), .A3(n_390), .B1(n_392), .B2(n_391), .C(n_393), .Y(n_479) );
INVxp67_ASAP7_75t_L g480 ( .A(n_426), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_431), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_425), .B(n_392), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_415), .B(n_390), .Y(n_483) );
INVxp67_ASAP7_75t_L g484 ( .A(n_426), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_435), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_438), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_439), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_441), .Y(n_488) );
NAND2x1_ASAP7_75t_L g489 ( .A(n_448), .B(n_398), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_425), .B(n_393), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_402), .B(n_390), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_444), .Y(n_492) );
OAI322xp33_ASAP7_75t_L g493 ( .A1(n_420), .A2(n_395), .A3(n_401), .B1(n_398), .B2(n_360), .C1(n_138), .C2(n_277), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_447), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_402), .B(n_390), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_449), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_415), .B(n_398), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_406), .B(n_401), .Y(n_498) );
OR2x2_ASAP7_75t_L g499 ( .A(n_409), .B(n_395), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_452), .Y(n_500) );
OR2x2_ASAP7_75t_L g501 ( .A(n_406), .B(n_138), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_408), .B(n_8), .Y(n_502) );
INVx1_ASAP7_75t_SL g503 ( .A(n_455), .Y(n_503) );
AOI211xp5_ASAP7_75t_SL g504 ( .A1(n_493), .A2(n_427), .B(n_419), .C(n_448), .Y(n_504) );
OAI211xp5_ASAP7_75t_SL g505 ( .A1(n_470), .A2(n_427), .B(n_442), .C(n_448), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_501), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_468), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_472), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_477), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_467), .B(n_443), .Y(n_510) );
AOI321xp33_ASAP7_75t_SL g511 ( .A1(n_463), .A2(n_9), .A3(n_10), .B1(n_11), .B2(n_12), .C(n_13), .Y(n_511) );
NAND3x2_ASAP7_75t_L g512 ( .A(n_464), .B(n_454), .C(n_442), .Y(n_512) );
OAI33xp33_ASAP7_75t_L g513 ( .A1(n_459), .A2(n_414), .A3(n_423), .B1(n_430), .B2(n_418), .B3(n_424), .Y(n_513) );
BUFx2_ASAP7_75t_L g514 ( .A(n_476), .Y(n_514) );
OR2x2_ASAP7_75t_L g515 ( .A(n_478), .B(n_432), .Y(n_515) );
A2O1A1Ixp33_ASAP7_75t_SL g516 ( .A1(n_502), .A2(n_443), .B(n_416), .C(n_412), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_471), .A2(n_436), .B1(n_451), .B2(n_446), .Y(n_517) );
OAI21xp33_ASAP7_75t_L g518 ( .A1(n_467), .A2(n_432), .B(n_433), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_465), .Y(n_519) );
OAI21xp5_ASAP7_75t_L g520 ( .A1(n_503), .A2(n_440), .B(n_433), .Y(n_520) );
O2A1O1Ixp33_ASAP7_75t_L g521 ( .A1(n_460), .A2(n_413), .B(n_445), .C(n_437), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_461), .B(n_451), .Y(n_522) );
NOR3xp33_ASAP7_75t_L g523 ( .A(n_459), .B(n_260), .C(n_445), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_481), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_462), .B(n_446), .Y(n_525) );
OAI22xp5_ASAP7_75t_L g526 ( .A1(n_476), .A2(n_436), .B1(n_456), .B2(n_437), .Y(n_526) );
AOI21xp33_ASAP7_75t_SL g527 ( .A1(n_460), .A2(n_456), .B(n_11), .Y(n_527) );
OAI31xp33_ASAP7_75t_L g528 ( .A1(n_466), .A2(n_416), .A3(n_413), .B(n_277), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_483), .B(n_292), .Y(n_529) );
INVx2_ASAP7_75t_L g530 ( .A(n_466), .Y(n_530) );
OAI22xp33_ASAP7_75t_SL g531 ( .A1(n_489), .A2(n_278), .B1(n_281), .B2(n_294), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_498), .B(n_292), .Y(n_532) );
INVxp67_ASAP7_75t_L g533 ( .A(n_457), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_485), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_486), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_505), .A2(n_471), .B1(n_464), .B2(n_478), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_507), .Y(n_537) );
AOI22xp5_ASAP7_75t_L g538 ( .A1(n_518), .A2(n_480), .B1(n_484), .B2(n_491), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_508), .Y(n_539) );
OAI22xp5_ASAP7_75t_L g540 ( .A1(n_512), .A2(n_480), .B1(n_484), .B2(n_473), .Y(n_540) );
AOI222xp33_ASAP7_75t_L g541 ( .A1(n_513), .A2(n_495), .B1(n_487), .B2(n_492), .C1(n_496), .C2(n_500), .Y(n_541) );
OAI211xp5_ASAP7_75t_L g542 ( .A1(n_527), .A2(n_479), .B(n_499), .C(n_494), .Y(n_542) );
AOI211xp5_ASAP7_75t_L g543 ( .A1(n_523), .A2(n_475), .B(n_488), .C(n_458), .Y(n_543) );
OAI221xp5_ASAP7_75t_L g544 ( .A1(n_514), .A2(n_474), .B1(n_490), .B2(n_482), .C(n_465), .Y(n_544) );
AOI22xp5_ASAP7_75t_L g545 ( .A1(n_517), .A2(n_497), .B1(n_469), .B2(n_278), .Y(n_545) );
NOR4xp25_ASAP7_75t_L g546 ( .A(n_533), .B(n_9), .C(n_13), .D(n_14), .Y(n_546) );
OAI31xp33_ASAP7_75t_SL g547 ( .A1(n_526), .A2(n_15), .A3(n_16), .B(n_17), .Y(n_547) );
OAI211xp5_ASAP7_75t_SL g548 ( .A1(n_504), .A2(n_17), .B(n_18), .C(n_271), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g549 ( .A1(n_523), .A2(n_278), .B1(n_281), .B2(n_294), .Y(n_549) );
OAI221xp5_ASAP7_75t_L g550 ( .A1(n_517), .A2(n_278), .B1(n_281), .B2(n_294), .C(n_280), .Y(n_550) );
AO221x1_ASAP7_75t_L g551 ( .A1(n_513), .A2(n_278), .B1(n_21), .B2(n_22), .C(n_23), .Y(n_551) );
AOI22xp5_ASAP7_75t_L g552 ( .A1(n_506), .A2(n_247), .B1(n_168), .B2(n_166), .Y(n_552) );
CKINVDCx14_ASAP7_75t_R g553 ( .A(n_515), .Y(n_553) );
OAI222xp33_ASAP7_75t_L g554 ( .A1(n_510), .A2(n_247), .B1(n_168), .B2(n_166), .C1(n_261), .C2(n_29), .Y(n_554) );
AOI221x1_ASAP7_75t_L g555 ( .A1(n_531), .A2(n_20), .B1(n_25), .B2(n_27), .C(n_28), .Y(n_555) );
AOI22xp33_ASAP7_75t_L g556 ( .A1(n_520), .A2(n_168), .B1(n_166), .B2(n_247), .Y(n_556) );
OAI32xp33_ASAP7_75t_L g557 ( .A1(n_533), .A2(n_31), .A3(n_38), .B1(n_40), .B2(n_41), .Y(n_557) );
OAI222xp33_ASAP7_75t_L g558 ( .A1(n_521), .A2(n_168), .B1(n_166), .B2(n_45), .C1(n_46), .C2(n_47), .Y(n_558) );
NAND4xp25_ASAP7_75t_L g559 ( .A(n_516), .B(n_42), .C(n_43), .D(n_48), .Y(n_559) );
OAI221xp5_ASAP7_75t_L g560 ( .A1(n_528), .A2(n_168), .B1(n_166), .B2(n_55), .C(n_57), .Y(n_560) );
AOI22xp5_ASAP7_75t_L g561 ( .A1(n_522), .A2(n_166), .B1(n_52), .B2(n_61), .Y(n_561) );
OAI211xp5_ASAP7_75t_SL g562 ( .A1(n_516), .A2(n_49), .B(n_66), .C(n_67), .Y(n_562) );
AOI21xp5_ASAP7_75t_L g563 ( .A1(n_530), .A2(n_166), .B(n_71), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_509), .Y(n_564) );
AOI322xp5_ASAP7_75t_L g565 ( .A1(n_525), .A2(n_70), .A3(n_72), .B1(n_74), .B2(n_81), .C1(n_511), .C2(n_535), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_541), .B(n_543), .Y(n_566) );
NOR2x1_ASAP7_75t_L g567 ( .A(n_559), .B(n_548), .Y(n_567) );
NAND3xp33_ASAP7_75t_SL g568 ( .A(n_546), .B(n_565), .C(n_536), .Y(n_568) );
NAND4xp25_ASAP7_75t_L g569 ( .A(n_547), .B(n_548), .C(n_556), .D(n_549), .Y(n_569) );
NAND4xp25_ASAP7_75t_L g570 ( .A(n_555), .B(n_562), .C(n_545), .D(n_542), .Y(n_570) );
NAND3xp33_ASAP7_75t_SL g571 ( .A(n_560), .B(n_540), .C(n_551), .Y(n_571) );
NOR4xp25_ASAP7_75t_L g572 ( .A(n_568), .B(n_544), .C(n_558), .D(n_564), .Y(n_572) );
NAND3xp33_ASAP7_75t_SL g573 ( .A(n_566), .B(n_538), .C(n_552), .Y(n_573) );
INVx2_ASAP7_75t_L g574 ( .A(n_567), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_574), .B(n_553), .Y(n_575) );
NOR2x1_ASAP7_75t_L g576 ( .A(n_573), .B(n_571), .Y(n_576) );
OR2x6_ASAP7_75t_L g577 ( .A(n_575), .B(n_572), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_576), .Y(n_578) );
XNOR2xp5_ASAP7_75t_L g579 ( .A(n_577), .B(n_569), .Y(n_579) );
AOI22xp5_ASAP7_75t_L g580 ( .A1(n_579), .A2(n_578), .B1(n_570), .B2(n_539), .Y(n_580) );
OAI22x1_ASAP7_75t_L g581 ( .A1(n_580), .A2(n_561), .B1(n_537), .B2(n_524), .Y(n_581) );
OAI21xp5_ASAP7_75t_L g582 ( .A1(n_581), .A2(n_563), .B(n_557), .Y(n_582) );
AO21x2_ASAP7_75t_L g583 ( .A1(n_582), .A2(n_554), .B(n_534), .Y(n_583) );
AOI222xp33_ASAP7_75t_L g584 ( .A1(n_583), .A2(n_519), .B1(n_529), .B2(n_532), .C1(n_550), .C2(n_578), .Y(n_584) );
endmodule