module fake_jpeg_32138_n_506 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_506);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_506;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVxp67_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_16),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_16),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

CKINVDCx14_ASAP7_75t_R g32 ( 
.A(n_17),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_7),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_3),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

BUFx6f_ASAP7_75t_SL g50 ( 
.A(n_6),
.Y(n_50)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_51),
.Y(n_143)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_27),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_53),
.B(n_55),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_19),
.B(n_29),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_54),
.B(n_70),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_19),
.B(n_17),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_27),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_56),
.B(n_58),
.Y(n_119)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_57),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_29),
.B(n_15),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_32),
.B(n_15),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_59),
.B(n_68),
.Y(n_126)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_60),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_61),
.Y(n_107)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

INVx11_ASAP7_75t_L g158 ( 
.A(n_62),
.Y(n_158)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_63),
.Y(n_161)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_64),
.Y(n_104)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_65),
.Y(n_125)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_66),
.Y(n_108)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_67),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_27),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_32),
.B(n_14),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_69),
.B(n_73),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_23),
.B(n_14),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_28),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_71),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_72),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_18),
.B(n_14),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_21),
.Y(n_74)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_74),
.Y(n_134)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_75),
.Y(n_132)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_31),
.Y(n_76)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_76),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_50),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_77),
.B(n_78),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_38),
.B(n_0),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_79),
.Y(n_157)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_31),
.Y(n_80)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_80),
.Y(n_136)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_21),
.Y(n_81)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_81),
.Y(n_152)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_31),
.Y(n_82)
);

INVx8_ASAP7_75t_L g156 ( 
.A(n_82),
.Y(n_156)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_28),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_83),
.Y(n_138)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_84),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_30),
.Y(n_85)
);

BUFx8_ASAP7_75t_L g114 ( 
.A(n_85),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_28),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_86),
.Y(n_150)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_50),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_88),
.B(n_100),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_23),
.B(n_39),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_89),
.B(n_98),
.Y(n_133)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_35),
.Y(n_90)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_90),
.Y(n_140)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_91),
.Y(n_117)
);

INVx2_ASAP7_75t_SL g92 ( 
.A(n_30),
.Y(n_92)
);

CKINVDCx6p67_ASAP7_75t_R g149 ( 
.A(n_92),
.Y(n_149)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_44),
.Y(n_93)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_93),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_35),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_94),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_35),
.Y(n_95)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_95),
.Y(n_135)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_37),
.Y(n_96)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_96),
.Y(n_142)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_43),
.Y(n_97)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_97),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_24),
.B(n_0),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_30),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_99),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_45),
.B(n_0),
.Y(n_100)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_43),
.Y(n_101)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_101),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_37),
.Y(n_102)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_102),
.Y(n_159)
);

NOR2x1_ASAP7_75t_L g106 ( 
.A(n_63),
.B(n_24),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_106),
.B(n_153),
.Y(n_213)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_85),
.B(n_25),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_115),
.B(n_118),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_72),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_79),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_120),
.B(n_123),
.Y(n_174)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_85),
.B(n_25),
.Y(n_123)
);

BUFx10_ASAP7_75t_L g128 ( 
.A(n_99),
.Y(n_128)
);

INVx3_ASAP7_75t_SL g180 ( 
.A(n_128),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_102),
.A2(n_49),
.B1(n_48),
.B2(n_37),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_129),
.A2(n_95),
.B1(n_86),
.B2(n_61),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_92),
.B(n_34),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_137),
.B(n_147),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_99),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_141),
.B(n_145),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_94),
.A2(n_43),
.B1(n_41),
.B2(n_39),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_144),
.A2(n_145),
.B1(n_22),
.B2(n_36),
.Y(n_197)
);

OR2x2_ASAP7_75t_L g145 ( 
.A(n_80),
.B(n_41),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_75),
.B(n_34),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_90),
.Y(n_148)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_148),
.Y(n_184)
);

A2O1A1Ixp33_ASAP7_75t_L g153 ( 
.A1(n_57),
.A2(n_40),
.B(n_36),
.C(n_26),
.Y(n_153)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_96),
.Y(n_155)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_155),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_103),
.B(n_84),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_162),
.B(n_200),
.Y(n_222)
);

AO22x1_ASAP7_75t_L g163 ( 
.A1(n_106),
.A2(n_83),
.B1(n_52),
.B2(n_91),
.Y(n_163)
);

A2O1A1Ixp33_ASAP7_75t_L g229 ( 
.A1(n_163),
.A2(n_205),
.B(n_212),
.C(n_178),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_160),
.Y(n_164)
);

BUFx2_ASAP7_75t_L g252 ( 
.A(n_164),
.Y(n_252)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_112),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g261 ( 
.A(n_165),
.Y(n_261)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_121),
.Y(n_166)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_166),
.Y(n_245)
);

INVx8_ASAP7_75t_L g168 ( 
.A(n_114),
.Y(n_168)
);

INVx6_ASAP7_75t_L g236 ( 
.A(n_168),
.Y(n_236)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_121),
.Y(n_169)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_169),
.Y(n_220)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_110),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_171),
.Y(n_223)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_134),
.Y(n_172)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_172),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_160),
.Y(n_173)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_173),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_149),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_175),
.B(n_186),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_176),
.A2(n_181),
.B1(n_197),
.B2(n_204),
.Y(n_231)
);

BUFx12f_ASAP7_75t_L g177 ( 
.A(n_149),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g258 ( 
.A(n_177),
.Y(n_258)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_152),
.Y(n_179)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_179),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_135),
.A2(n_71),
.B1(n_82),
.B2(n_76),
.Y(n_181)
);

CKINVDCx14_ASAP7_75t_R g182 ( 
.A(n_149),
.Y(n_182)
);

NAND3xp33_ASAP7_75t_L g248 ( 
.A(n_182),
.B(n_210),
.C(n_215),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_107),
.Y(n_183)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_183),
.Y(n_254)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_132),
.Y(n_185)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_185),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_115),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_161),
.Y(n_187)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_187),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_107),
.Y(n_188)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_188),
.Y(n_251)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_124),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_190),
.Y(n_239)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_136),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_191),
.B(n_193),
.Y(n_250)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_131),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_192),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_105),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_122),
.Y(n_194)
);

BUFx24_ASAP7_75t_L g230 ( 
.A(n_194),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_133),
.B(n_26),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_195),
.B(n_196),
.Y(n_221)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_125),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_113),
.B(n_93),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_198),
.B(n_203),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_112),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_199),
.A2(n_208),
.B1(n_209),
.B2(n_216),
.Y(n_218)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_140),
.Y(n_200)
);

INVx13_ASAP7_75t_L g201 ( 
.A(n_114),
.Y(n_201)
);

OR2x2_ASAP7_75t_L g228 ( 
.A(n_201),
.B(n_205),
.Y(n_228)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_142),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_202),
.B(n_211),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_139),
.B(n_20),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_104),
.A2(n_97),
.B1(n_87),
.B2(n_67),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_153),
.A2(n_20),
.B1(n_22),
.B2(n_40),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_119),
.B(n_101),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_206),
.B(n_207),
.Y(n_238)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_109),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_109),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_130),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_126),
.B(n_66),
.Y(n_210)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_131),
.Y(n_211)
);

OA22x2_ASAP7_75t_L g212 ( 
.A1(n_123),
.A2(n_62),
.B1(n_51),
.B2(n_49),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_212),
.B(n_214),
.Y(n_243)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_117),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_146),
.B(n_151),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_130),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_162),
.B(n_154),
.C(n_127),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_217),
.B(n_226),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_L g219 ( 
.A1(n_163),
.A2(n_213),
.B1(n_159),
.B2(n_135),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_219),
.A2(n_237),
.B1(n_240),
.B2(n_183),
.Y(n_279)
);

MAJx2_ASAP7_75t_L g226 ( 
.A(n_170),
.B(n_128),
.C(n_114),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_229),
.A2(n_247),
.B(n_181),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_197),
.B(n_159),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_234),
.B(n_242),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_167),
.A2(n_122),
.B1(n_150),
.B2(n_138),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_174),
.A2(n_150),
.B1(n_138),
.B2(n_156),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_212),
.B(n_154),
.C(n_156),
.Y(n_241)
);

MAJx2_ASAP7_75t_L g274 ( 
.A(n_241),
.B(n_249),
.C(n_111),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_187),
.B(n_128),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_200),
.B(n_116),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_244),
.B(n_259),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_204),
.A2(n_157),
.B(n_143),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_202),
.B(n_116),
.C(n_108),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_192),
.A2(n_108),
.B1(n_117),
.B2(n_158),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_255),
.B(n_256),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_177),
.A2(n_158),
.B(n_157),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_177),
.A2(n_111),
.B1(n_49),
.B2(n_48),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_257),
.A2(n_180),
.B1(n_168),
.B2(n_165),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_184),
.B(n_48),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_243),
.A2(n_211),
.B1(n_190),
.B2(n_166),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_263),
.A2(n_300),
.B(n_261),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_242),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_264),
.B(n_265),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_227),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_228),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_266),
.B(n_272),
.Y(n_313)
);

CKINVDCx14_ASAP7_75t_R g311 ( 
.A(n_267),
.Y(n_311)
);

INVx4_ASAP7_75t_L g268 ( 
.A(n_236),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_268),
.Y(n_330)
);

INVx13_ASAP7_75t_L g270 ( 
.A(n_245),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_270),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_241),
.A2(n_176),
.B1(n_164),
.B2(n_173),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_271),
.A2(n_299),
.B1(n_247),
.B2(n_251),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_228),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_224),
.B(n_189),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_273),
.B(n_281),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_SL g314 ( 
.A(n_274),
.B(n_249),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_225),
.Y(n_275)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_275),
.Y(n_302)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_244),
.Y(n_276)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_276),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g278 ( 
.A(n_220),
.Y(n_278)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_278),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_279),
.A2(n_239),
.B1(n_252),
.B2(n_254),
.Y(n_327)
);

AND2x6_ASAP7_75t_L g280 ( 
.A(n_248),
.B(n_201),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_280),
.B(n_283),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_235),
.B(n_169),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_246),
.Y(n_282)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_282),
.Y(n_315)
);

CKINVDCx14_ASAP7_75t_R g283 ( 
.A(n_243),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_SL g333 ( 
.A1(n_285),
.A2(n_298),
.B1(n_252),
.B2(n_254),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_227),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_286),
.B(n_291),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_221),
.B(n_214),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_287),
.B(n_288),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_222),
.B(n_194),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_246),
.Y(n_289)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_289),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_229),
.B(n_0),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_290),
.B(n_293),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_223),
.B(n_199),
.Y(n_291)
);

INVx13_ASAP7_75t_L g292 ( 
.A(n_245),
.Y(n_292)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_292),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_227),
.Y(n_293)
);

INVx13_ASAP7_75t_L g294 ( 
.A(n_258),
.Y(n_294)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_294),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_238),
.B(n_180),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_295),
.B(n_297),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_243),
.A2(n_47),
.B(n_2),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_296),
.A2(n_218),
.B(n_259),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_222),
.B(n_188),
.Y(n_297)
);

INVx5_ASAP7_75t_L g298 ( 
.A(n_236),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_231),
.A2(n_13),
.B1(n_2),
.B2(n_3),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_232),
.B(n_1),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_301),
.A2(n_307),
.B1(n_322),
.B2(n_268),
.Y(n_358)
);

NOR2x1_ASAP7_75t_R g305 ( 
.A(n_266),
.B(n_272),
.Y(n_305)
);

OR2x2_ASAP7_75t_SL g361 ( 
.A(n_305),
.B(n_294),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_271),
.A2(n_299),
.B1(n_277),
.B2(n_276),
.Y(n_307)
);

OAI22xp33_ASAP7_75t_SL g308 ( 
.A1(n_290),
.A2(n_234),
.B1(n_231),
.B2(n_226),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_308),
.A2(n_321),
.B1(n_325),
.B2(n_327),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_277),
.A2(n_222),
.B1(n_217),
.B2(n_253),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g340 ( 
.A(n_310),
.B(n_334),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_312),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_314),
.B(n_331),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_262),
.B(n_232),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_316),
.B(n_326),
.C(n_274),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_269),
.A2(n_255),
.B1(n_256),
.B2(n_251),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_277),
.A2(n_233),
.B1(n_250),
.B2(n_239),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_269),
.A2(n_264),
.B1(n_284),
.B2(n_279),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_262),
.B(n_253),
.C(n_233),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_SL g331 ( 
.A(n_274),
.B(n_261),
.Y(n_331)
);

INVx13_ASAP7_75t_L g365 ( 
.A(n_333),
.Y(n_365)
);

OAI22xp33_ASAP7_75t_SL g335 ( 
.A1(n_267),
.A2(n_225),
.B1(n_220),
.B2(n_260),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_335),
.B(n_263),
.Y(n_337)
);

INVx8_ASAP7_75t_L g336 ( 
.A(n_330),
.Y(n_336)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_336),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_337),
.A2(n_302),
.B1(n_330),
.B2(n_275),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_306),
.B(n_284),
.Y(n_338)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_338),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_329),
.Y(n_339)
);

OR2x2_ASAP7_75t_L g395 ( 
.A(n_339),
.B(n_346),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_306),
.B(n_287),
.Y(n_341)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_341),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_325),
.B(n_300),
.Y(n_342)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_342),
.Y(n_377)
);

AND2x6_ASAP7_75t_L g344 ( 
.A(n_311),
.B(n_280),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_SL g373 ( 
.A1(n_344),
.A2(n_350),
.B(n_356),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_304),
.B(n_273),
.Y(n_345)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_345),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_304),
.B(n_281),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_348),
.B(n_230),
.Y(n_396)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_315),
.Y(n_349)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_349),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g350 ( 
.A1(n_334),
.A2(n_293),
.B(n_286),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_332),
.B(n_265),
.Y(n_351)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_351),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_332),
.B(n_297),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_352),
.Y(n_382)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_321),
.B(n_288),
.Y(n_353)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_353),
.B(n_319),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_303),
.B(n_296),
.Y(n_354)
);

CKINVDCx16_ASAP7_75t_R g369 ( 
.A(n_354),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_303),
.B(n_323),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_355),
.B(n_318),
.Y(n_368)
);

OR2x2_ASAP7_75t_L g356 ( 
.A(n_305),
.B(n_282),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_322),
.A2(n_313),
.B(n_310),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g384 ( 
.A(n_357),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_358),
.A2(n_359),
.B1(n_362),
.B2(n_327),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_307),
.A2(n_289),
.B1(n_298),
.B2(n_275),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_361),
.A2(n_328),
.B1(n_312),
.B2(n_324),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_301),
.A2(n_317),
.B1(n_323),
.B2(n_320),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_324),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_363),
.B(n_292),
.Y(n_389)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_315),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_364),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_328),
.B(n_294),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_SL g378 ( 
.A(n_366),
.B(n_367),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_SL g367 ( 
.A(n_318),
.B(n_260),
.Y(n_367)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_368),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_343),
.B(n_314),
.C(n_331),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_371),
.B(n_372),
.C(n_381),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_343),
.B(n_326),
.C(n_316),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_376),
.A2(n_393),
.B1(n_394),
.B2(n_361),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_SL g399 ( 
.A(n_380),
.B(n_340),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_348),
.B(n_309),
.C(n_319),
.Y(n_381)
);

NOR2x1_ASAP7_75t_L g383 ( 
.A(n_340),
.B(n_309),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_383),
.B(n_350),
.Y(n_401)
);

INVx1_ASAP7_75t_SL g402 ( 
.A(n_385),
.Y(n_402)
);

CKINVDCx14_ASAP7_75t_R g421 ( 
.A(n_386),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_339),
.A2(n_330),
.B1(n_302),
.B2(n_230),
.Y(n_387)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_387),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_389),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_355),
.B(n_292),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_390),
.B(n_363),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_340),
.A2(n_230),
.B1(n_270),
.B2(n_5),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_358),
.A2(n_230),
.B1(n_270),
.B2(n_5),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_396),
.B(n_353),
.C(n_357),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_397),
.A2(n_384),
.B1(n_375),
.B2(n_383),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_SL g398 ( 
.A(n_369),
.B(n_362),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_398),
.B(n_406),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_399),
.B(n_414),
.Y(n_437)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_378),
.Y(n_400)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_400),
.Y(n_426)
);

CKINVDCx14_ASAP7_75t_R g440 ( 
.A(n_401),
.Y(n_440)
);

BUFx24_ASAP7_75t_SL g404 ( 
.A(n_395),
.Y(n_404)
);

BUFx24_ASAP7_75t_SL g422 ( 
.A(n_404),
.Y(n_422)
);

XNOR2x1_ASAP7_75t_L g405 ( 
.A(n_371),
.B(n_342),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_405),
.B(n_411),
.Y(n_427)
);

AOI21xp5_ASAP7_75t_L g406 ( 
.A1(n_373),
.A2(n_347),
.B(n_353),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_378),
.Y(n_407)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_407),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_SL g409 ( 
.A(n_374),
.B(n_346),
.Y(n_409)
);

CKINVDCx16_ASAP7_75t_R g424 ( 
.A(n_409),
.Y(n_424)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_388),
.Y(n_410)
);

HB1xp67_ASAP7_75t_L g431 ( 
.A(n_410),
.Y(n_431)
);

AOI21xp33_ASAP7_75t_L g412 ( 
.A1(n_373),
.A2(n_344),
.B(n_354),
.Y(n_412)
);

NOR2xp67_ASAP7_75t_SL g429 ( 
.A(n_412),
.B(n_399),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_396),
.B(n_360),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_415),
.A2(n_400),
.B1(n_407),
.B2(n_395),
.Y(n_433)
);

AOI21xp5_ASAP7_75t_L g416 ( 
.A1(n_380),
.A2(n_356),
.B(n_360),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g432 ( 
.A1(n_416),
.A2(n_418),
.B1(n_394),
.B2(n_337),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_376),
.A2(n_377),
.B1(n_392),
.B2(n_382),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_417),
.A2(n_377),
.B1(n_359),
.B2(n_385),
.Y(n_423)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_388),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_381),
.B(n_338),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_420),
.B(n_408),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_423),
.B(n_429),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_425),
.B(n_434),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_420),
.B(n_372),
.C(n_384),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_428),
.B(n_408),
.C(n_411),
.Y(n_442)
);

A2O1A1Ixp33_ASAP7_75t_SL g430 ( 
.A1(n_401),
.A2(n_385),
.B(n_344),
.C(n_392),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_430),
.B(n_439),
.Y(n_446)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_432),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_433),
.B(n_436),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_405),
.B(n_374),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_421),
.A2(n_375),
.B1(n_382),
.B2(n_379),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_413),
.A2(n_379),
.B1(n_365),
.B2(n_391),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_441),
.B(n_416),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_442),
.B(n_451),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_441),
.B(n_414),
.C(n_406),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_444),
.B(n_449),
.C(n_454),
.Y(n_461)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_426),
.Y(n_445)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_445),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_428),
.B(n_417),
.C(n_402),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_438),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_450),
.B(n_452),
.Y(n_469)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_435),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_427),
.B(n_402),
.C(n_419),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_424),
.B(n_403),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_455),
.B(n_456),
.Y(n_468)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_431),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_427),
.B(n_391),
.C(n_397),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_457),
.B(n_437),
.C(n_434),
.Y(n_462)
);

INVxp67_ASAP7_75t_L g458 ( 
.A(n_446),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_458),
.B(n_463),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_442),
.B(n_437),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_459),
.B(n_462),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_451),
.B(n_423),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_453),
.B(n_393),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_464),
.B(n_453),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_457),
.B(n_430),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_465),
.B(n_341),
.Y(n_483)
);

OR2x2_ASAP7_75t_L g466 ( 
.A(n_448),
.B(n_351),
.Y(n_466)
);

CKINVDCx16_ASAP7_75t_R g476 ( 
.A(n_466),
.Y(n_476)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_447),
.A2(n_430),
.B(n_418),
.Y(n_470)
);

AOI21xp5_ASAP7_75t_L g474 ( 
.A1(n_470),
.A2(n_471),
.B(n_444),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_449),
.B(n_440),
.C(n_352),
.Y(n_471)
);

AOI211xp5_ASAP7_75t_SL g472 ( 
.A1(n_458),
.A2(n_430),
.B(n_466),
.C(n_467),
.Y(n_472)
);

AOI21xp5_ASAP7_75t_SL g489 ( 
.A1(n_472),
.A2(n_479),
.B(n_356),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_474),
.B(n_477),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_475),
.B(n_480),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_468),
.A2(n_443),
.B1(n_460),
.B2(n_465),
.Y(n_477)
);

NOR2xp67_ASAP7_75t_SL g478 ( 
.A(n_461),
.B(n_454),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_SL g491 ( 
.A(n_478),
.B(n_481),
.Y(n_491)
);

AOI21xp5_ASAP7_75t_SL g479 ( 
.A1(n_469),
.A2(n_471),
.B(n_410),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_461),
.A2(n_349),
.B1(n_364),
.B2(n_370),
.Y(n_480)
);

NOR2xp67_ASAP7_75t_SL g481 ( 
.A(n_462),
.B(n_422),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_483),
.B(n_345),
.Y(n_487)
);

FAx1_ASAP7_75t_SL g484 ( 
.A(n_472),
.B(n_483),
.CI(n_473),
.CON(n_484),
.SN(n_484)
);

NOR2xp33_ASAP7_75t_SL g495 ( 
.A(n_484),
.B(n_485),
.Y(n_495)
);

NOR2xp67_ASAP7_75t_SL g485 ( 
.A(n_482),
.B(n_370),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_487),
.B(n_489),
.Y(n_494)
);

AOI21xp5_ASAP7_75t_L g490 ( 
.A1(n_479),
.A2(n_366),
.B(n_367),
.Y(n_490)
);

AOI322xp5_ASAP7_75t_L g496 ( 
.A1(n_490),
.A2(n_336),
.A3(n_4),
.B1(n_5),
.B2(n_7),
.C1(n_8),
.C2(n_3),
.Y(n_496)
);

OAI21xp33_ASAP7_75t_L g492 ( 
.A1(n_491),
.A2(n_476),
.B(n_365),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_492),
.B(n_493),
.Y(n_499)
);

AOI322xp5_ASAP7_75t_L g493 ( 
.A1(n_484),
.A2(n_486),
.A3(n_489),
.B1(n_488),
.B2(n_365),
.C1(n_336),
.C2(n_9),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_496),
.B(n_4),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_497),
.B(n_498),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_495),
.B(n_4),
.C(n_5),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_499),
.B(n_494),
.C(n_9),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_500),
.B(n_8),
.Y(n_502)
);

AOI21xp5_ASAP7_75t_L g503 ( 
.A1(n_502),
.A2(n_501),
.B(n_10),
.Y(n_503)
);

OAI21xp5_ASAP7_75t_SL g504 ( 
.A1(n_503),
.A2(n_8),
.B(n_10),
.Y(n_504)
);

AOI21xp5_ASAP7_75t_L g505 ( 
.A1(n_504),
.A2(n_12),
.B(n_13),
.Y(n_505)
);

AOI21xp5_ASAP7_75t_SL g506 ( 
.A1(n_505),
.A2(n_13),
.B(n_503),
.Y(n_506)
);


endmodule