module fake_jpeg_6998_n_317 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_317);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_317;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_7),
.B(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_38),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_36),
.B(n_37),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_16),
.B(n_15),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_16),
.B(n_15),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_41),
.Y(n_51)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_40),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_25),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_43),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_33),
.A2(n_28),
.B1(n_19),
.B2(n_30),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_44),
.A2(n_54),
.B1(n_27),
.B2(n_32),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_36),
.B(n_16),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_45),
.B(n_48),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_L g46 ( 
.A1(n_40),
.A2(n_28),
.B1(n_24),
.B2(n_26),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_46),
.A2(n_50),
.B1(n_23),
.B2(n_29),
.Y(n_80)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_39),
.A2(n_30),
.B1(n_19),
.B2(n_28),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_33),
.A2(n_40),
.B1(n_39),
.B2(n_19),
.Y(n_54)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_57),
.B(n_63),
.Y(n_76)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_34),
.A2(n_30),
.B1(n_24),
.B2(n_22),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_59),
.A2(n_62),
.B(n_23),
.Y(n_82)
);

AND2x2_ASAP7_75t_SL g60 ( 
.A(n_43),
.B(n_20),
.Y(n_60)
);

AOI21xp33_ASAP7_75t_L g78 ( 
.A1(n_60),
.A2(n_20),
.B(n_29),
.Y(n_78)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_35),
.A2(n_22),
.B1(n_31),
.B2(n_27),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_35),
.B(n_22),
.Y(n_63)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_66),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_43),
.B(n_31),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_68),
.B(n_26),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_69),
.B(n_83),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_60),
.A2(n_31),
.B1(n_27),
.B2(n_21),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_70),
.A2(n_75),
.B1(n_93),
.B2(n_58),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_72),
.A2(n_73),
.B1(n_59),
.B2(n_52),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_60),
.A2(n_32),
.B1(n_21),
.B2(n_29),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_63),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_91),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_60),
.A2(n_10),
.B1(n_13),
.B2(n_14),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_78),
.A2(n_82),
.B(n_53),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_80),
.A2(n_54),
.B1(n_64),
.B2(n_49),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_47),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_60),
.B(n_43),
.C(n_20),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_94),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_45),
.B(n_43),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_85),
.B(n_53),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_47),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_86),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_44),
.B(n_20),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_SL g104 ( 
.A(n_87),
.B(n_54),
.Y(n_104)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_51),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_92),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_58),
.A2(n_14),
.B1(n_13),
.B2(n_11),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_50),
.B(n_20),
.C(n_25),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_96),
.Y(n_123)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_88),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_97),
.B(n_98),
.Y(n_127)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_76),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_76),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_99),
.B(n_101),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_64),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_100),
.B(n_112),
.Y(n_121)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_103),
.A2(n_94),
.B1(n_71),
.B2(n_75),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_104),
.B(n_116),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_80),
.A2(n_55),
.B1(n_52),
.B2(n_51),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_105),
.A2(n_74),
.B1(n_70),
.B2(n_89),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_86),
.B(n_53),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_106),
.B(n_118),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_82),
.Y(n_108)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_108),
.Y(n_134)
);

AOI21xp33_ASAP7_75t_L g109 ( 
.A1(n_85),
.A2(n_68),
.B(n_29),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_109),
.A2(n_100),
.B(n_114),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_71),
.B(n_48),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_111),
.B(n_120),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_79),
.B(n_62),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_79),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_113),
.B(n_117),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_69),
.B(n_50),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_115),
.B(n_87),
.Y(n_140)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_72),
.Y(n_117)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_85),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_119),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_SL g122 ( 
.A(n_112),
.B(n_78),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_122),
.B(n_142),
.C(n_120),
.Y(n_167)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_95),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_124),
.B(n_128),
.Y(n_159)
);

OR2x2_ASAP7_75t_SL g128 ( 
.A(n_110),
.B(n_69),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_95),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_129),
.B(n_136),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_131),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_133),
.A2(n_120),
.B(n_107),
.Y(n_165)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_135),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_98),
.B(n_69),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_99),
.B(n_89),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_137),
.B(n_143),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_117),
.A2(n_87),
.B1(n_73),
.B2(n_94),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_138),
.Y(n_150)
);

OAI22x1_ASAP7_75t_SL g139 ( 
.A1(n_116),
.A2(n_87),
.B1(n_84),
.B2(n_93),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_139),
.A2(n_119),
.B1(n_114),
.B2(n_115),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_140),
.B(n_145),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_102),
.B(n_84),
.C(n_67),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_111),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_103),
.A2(n_105),
.B1(n_104),
.B2(n_118),
.Y(n_144)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_144),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_110),
.B(n_90),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_106),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_146),
.B(n_77),
.Y(n_171)
);

OA22x2_ASAP7_75t_L g151 ( 
.A1(n_139),
.A2(n_104),
.B1(n_106),
.B2(n_120),
.Y(n_151)
);

A2O1A1Ixp33_ASAP7_75t_SL g178 ( 
.A1(n_151),
.A2(n_171),
.B(n_138),
.C(n_141),
.Y(n_178)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_145),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_152),
.B(n_153),
.Y(n_195)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_132),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_154),
.B(n_135),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_127),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_155),
.B(n_156),
.Y(n_197)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_132),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_121),
.B(n_102),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_157),
.B(n_161),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_121),
.A2(n_109),
.B(n_113),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_158),
.A2(n_140),
.B(n_130),
.Y(n_174)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_127),
.Y(n_161)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_141),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_164),
.B(n_168),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_165),
.A2(n_173),
.B(n_130),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_167),
.B(n_122),
.C(n_129),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_126),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_133),
.B(n_90),
.Y(n_169)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_169),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_126),
.Y(n_170)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_170),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_143),
.B(n_101),
.Y(n_172)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_172),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_125),
.B(n_77),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_174),
.B(n_179),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_172),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_175),
.B(n_168),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_162),
.A2(n_147),
.B1(n_131),
.B2(n_144),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_176),
.A2(n_177),
.B1(n_178),
.B2(n_184),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_162),
.A2(n_147),
.B1(n_154),
.B2(n_148),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_149),
.A2(n_123),
.B1(n_134),
.B2(n_146),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_180),
.A2(n_190),
.B1(n_159),
.B2(n_160),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_167),
.B(n_125),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_181),
.B(n_185),
.C(n_189),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_182),
.B(n_194),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_151),
.A2(n_134),
.B(n_142),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_183),
.A2(n_191),
.B1(n_193),
.B2(n_151),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_151),
.A2(n_147),
.B1(n_128),
.B2(n_124),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_163),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_188),
.B(n_164),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_167),
.B(n_122),
.C(n_67),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_151),
.B(n_136),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_151),
.A2(n_137),
.B(n_17),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_148),
.A2(n_52),
.B1(n_101),
.B2(n_81),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_173),
.B(n_97),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_157),
.B(n_66),
.C(n_57),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_196),
.B(n_173),
.C(n_169),
.Y(n_204)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_200),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_198),
.B(n_155),
.Y(n_202)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_202),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_177),
.A2(n_193),
.B1(n_178),
.B2(n_176),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_203),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_204),
.B(n_205),
.C(n_201),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_181),
.B(n_157),
.C(n_158),
.Y(n_205)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_206),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_187),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_207),
.B(n_214),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_178),
.A2(n_191),
.B1(n_183),
.B2(n_149),
.Y(n_208)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_208),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_197),
.B(n_163),
.Y(n_209)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_209),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_186),
.B(n_166),
.Y(n_211)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_211),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_186),
.B(n_166),
.Y(n_212)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_212),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_199),
.B(n_156),
.Y(n_213)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_213),
.Y(n_241)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_187),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_192),
.B(n_152),
.Y(n_215)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_215),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_216),
.A2(n_165),
.B(n_174),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_218),
.B(n_190),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_194),
.B(n_153),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_219),
.B(n_223),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_190),
.A2(n_150),
.B1(n_158),
.B2(n_159),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_220),
.A2(n_184),
.B1(n_189),
.B2(n_179),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_178),
.A2(n_165),
.B1(n_170),
.B2(n_161),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_222),
.A2(n_195),
.B1(n_160),
.B2(n_175),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_196),
.B(n_81),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_205),
.B(n_185),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_229),
.B(n_239),
.C(n_201),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_230),
.A2(n_210),
.B1(n_182),
.B2(n_211),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_214),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_232),
.B(n_242),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_233),
.A2(n_217),
.B(n_212),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_235),
.A2(n_240),
.B1(n_217),
.B2(n_204),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_207),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_230),
.B(n_221),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_245),
.B(n_249),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_236),
.B(n_215),
.Y(n_246)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_246),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_237),
.A2(n_220),
.B1(n_216),
.B2(n_218),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_247),
.B(n_257),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_248),
.B(n_256),
.C(n_234),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_239),
.B(n_221),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_250),
.A2(n_255),
.B1(n_261),
.B2(n_0),
.Y(n_276)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_226),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_251),
.B(n_253),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_252),
.B(n_259),
.Y(n_267)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_231),
.Y(n_253)
);

XNOR2x1_ASAP7_75t_L g254 ( 
.A(n_233),
.B(n_210),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_254),
.A2(n_241),
.B1(n_1),
.B2(n_2),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_229),
.B(n_171),
.C(n_56),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_225),
.A2(n_81),
.B1(n_91),
.B2(n_14),
.Y(n_257)
);

INVxp67_ASAP7_75t_SL g258 ( 
.A(n_224),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_258),
.B(n_243),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_240),
.B(n_17),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_241),
.B(n_11),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_260),
.B(n_244),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_243),
.A2(n_228),
.B1(n_227),
.B2(n_224),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_262),
.B(n_271),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_250),
.A2(n_228),
.B1(n_227),
.B2(n_238),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_263),
.A2(n_276),
.B1(n_245),
.B2(n_249),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_265),
.A2(n_272),
.B(n_274),
.Y(n_289)
);

NOR2xp67_ASAP7_75t_SL g278 ( 
.A(n_266),
.B(n_0),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_248),
.B(n_65),
.C(n_1),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_254),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_273),
.B(n_3),
.Y(n_288)
);

NAND4xp25_ASAP7_75t_L g274 ( 
.A(n_261),
.B(n_65),
.C(n_11),
.D(n_2),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_256),
.B(n_65),
.C(n_1),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_275),
.B(n_3),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_263),
.A2(n_247),
.B(n_259),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_277),
.A2(n_285),
.B(n_4),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_278),
.A2(n_287),
.B(n_4),
.Y(n_299)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_279),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_264),
.B(n_0),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_280),
.B(n_281),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_269),
.B(n_1),
.Y(n_281)
);

INVx6_ASAP7_75t_L g282 ( 
.A(n_272),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_282),
.B(n_286),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_284),
.B(n_275),
.C(n_268),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_267),
.A2(n_3),
.B(n_4),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_270),
.B(n_265),
.Y(n_286)
);

OAI21x1_ASAP7_75t_L g287 ( 
.A1(n_266),
.A2(n_3),
.B(n_4),
.Y(n_287)
);

CKINVDCx14_ASAP7_75t_R g295 ( 
.A(n_288),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_290),
.B(n_292),
.Y(n_300)
);

FAx1_ASAP7_75t_L g292 ( 
.A(n_277),
.B(n_267),
.CI(n_268),
.CON(n_292),
.SN(n_292)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_282),
.B(n_283),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_293),
.A2(n_296),
.B(n_5),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_279),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_297),
.B(n_285),
.Y(n_301)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_299),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_301),
.A2(n_305),
.B(n_306),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_298),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_302),
.B(n_303),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_294),
.A2(n_289),
.B1(n_65),
.B2(n_7),
.Y(n_303)
);

NOR2x1_ASAP7_75t_L g305 ( 
.A(n_292),
.B(n_5),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_298),
.A2(n_5),
.B(n_6),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_307),
.A2(n_291),
.B(n_295),
.Y(n_308)
);

OAI21xp33_ASAP7_75t_L g313 ( 
.A1(n_308),
.A2(n_304),
.B(n_8),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_300),
.B(n_6),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_309),
.A2(n_310),
.B(n_8),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_305),
.A2(n_7),
.B(n_8),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_313),
.B(n_314),
.C(n_312),
.Y(n_315)
);

AO21x2_ASAP7_75t_L g316 ( 
.A1(n_315),
.A2(n_311),
.B(n_9),
.Y(n_316)
);

BUFx24_ASAP7_75t_SL g317 ( 
.A(n_316),
.Y(n_317)
);


endmodule