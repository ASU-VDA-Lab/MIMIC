module fake_jpeg_11378_n_187 (n_13, n_21, n_53, n_33, n_54, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_187);

input n_13;
input n_21;
input n_53;
input n_33;
input n_54;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_187;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx4_ASAP7_75t_L g55 ( 
.A(n_52),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

BUFx16f_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_10),
.Y(n_58)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_11),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_2),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_9),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_5),
.Y(n_64)
);

BUFx4f_ASAP7_75t_L g65 ( 
.A(n_12),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_30),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_27),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_18),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_20),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_28),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_53),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_22),
.Y(n_79)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_15),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_2),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_0),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_13),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_63),
.B(n_0),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_84),
.B(n_88),
.Y(n_95)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

INVxp67_ASAP7_75t_SL g94 ( 
.A(n_86),
.Y(n_94)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_61),
.Y(n_89)
);

AOI21xp33_ASAP7_75t_L g106 ( 
.A1(n_89),
.A2(n_73),
.B(n_77),
.Y(n_106)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_67),
.Y(n_90)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_90),
.Y(n_100)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_59),
.Y(n_91)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_91),
.Y(n_105)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_92),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_85),
.A2(n_60),
.B1(n_82),
.B2(n_83),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_93),
.A2(n_99),
.B1(n_71),
.B2(n_67),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_92),
.B(n_81),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_96),
.B(n_103),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_69),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_97),
.B(n_78),
.C(n_76),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_90),
.A2(n_80),
.B1(n_62),
.B2(n_64),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_85),
.A2(n_60),
.B1(n_62),
.B2(n_55),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_84),
.B(n_79),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_57),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_107),
.B(n_109),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_101),
.A2(n_80),
.B1(n_70),
.B2(n_72),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_108),
.A2(n_13),
.B(n_14),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_75),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_110),
.B(n_122),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_111),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_136)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_100),
.Y(n_112)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_112),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_97),
.A2(n_74),
.B1(n_68),
.B2(n_66),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_113),
.A2(n_121),
.B1(n_10),
.B2(n_11),
.Y(n_140)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_104),
.Y(n_114)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_114),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_98),
.A2(n_71),
.B1(n_65),
.B2(n_25),
.Y(n_115)
);

BUFx4f_ASAP7_75t_SL g116 ( 
.A(n_100),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_116),
.B(n_117),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_102),
.C(n_94),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_101),
.Y(n_118)
);

HB1xp67_ASAP7_75t_L g132 ( 
.A(n_118),
.Y(n_132)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_105),
.Y(n_119)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_119),
.Y(n_142)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_104),
.Y(n_120)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_120),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_105),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_103),
.B(n_3),
.Y(n_122)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_104),
.Y(n_124)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_124),
.Y(n_146)
);

OAI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_98),
.A2(n_23),
.B1(n_48),
.B2(n_47),
.Y(n_125)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_100),
.Y(n_126)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_126),
.Y(n_128)
);

NOR2x1_ASAP7_75t_L g129 ( 
.A(n_123),
.B(n_4),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_129),
.B(n_134),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_125),
.B(n_5),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_111),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_135),
.B(n_29),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_126),
.B(n_6),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_137),
.A2(n_116),
.B(n_17),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_115),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_140),
.A2(n_143),
.B1(n_137),
.B2(n_133),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_121),
.B(n_12),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_141),
.B(n_144),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_118),
.B(n_14),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_147),
.B(n_157),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_139),
.A2(n_16),
.B1(n_19),
.B2(n_26),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_148),
.B(n_150),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_127),
.B(n_31),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_151),
.B(n_149),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_152),
.B(n_155),
.Y(n_169)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_130),
.Y(n_154)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_154),
.Y(n_166)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_131),
.Y(n_155)
);

OR2x2_ASAP7_75t_SL g156 ( 
.A(n_145),
.B(n_34),
.Y(n_156)
);

A2O1A1O1Ixp25_ASAP7_75t_L g161 ( 
.A1(n_156),
.A2(n_39),
.B(n_40),
.C(n_41),
.D(n_43),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_129),
.A2(n_35),
.B(n_37),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_133),
.B(n_38),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_158),
.B(n_159),
.C(n_132),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_142),
.A2(n_146),
.B1(n_138),
.B2(n_136),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_160),
.B(n_161),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_158),
.B(n_132),
.C(n_46),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_163),
.B(n_164),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_153),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_156),
.B(n_45),
.C(n_128),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_165),
.B(n_162),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_168),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_166),
.Y(n_171)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_171),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_172),
.B(n_167),
.C(n_169),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_169),
.Y(n_173)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_173),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_175),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_179),
.B(n_170),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_180),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_181),
.B(n_174),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_182),
.B(n_176),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_183),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_184),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_185),
.B(n_177),
.Y(n_186)
);

BUFx24_ASAP7_75t_SL g187 ( 
.A(n_186),
.Y(n_187)
);


endmodule