module real_jpeg_32467_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_712, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_712;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_661;
wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_630;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_663;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_648;
wire n_95;
wire n_541;
wire n_441;
wire n_696;
wire n_657;
wire n_656;
wire n_643;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_669;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_679;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_640;
wire n_666;
wire n_160;
wire n_211;
wire n_574;
wire n_627;
wire n_595;
wire n_490;
wire n_39;
wire n_685;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_680;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_678;
wire n_30;
wire n_328;
wire n_578;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_620;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_668;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_605;
wire n_483;
wire n_367;
wire n_639;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_682;
wire n_317;
wire n_658;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_674;
wire n_252;
wire n_601;
wire n_655;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_525;
wire n_393;
wire n_221;
wire n_489;
wire n_611;
wire n_104;
wire n_153;
wire n_634;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_684;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_646;
wire n_214;
wire n_671;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_704;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_631;
wire n_673;
wire n_175;
wire n_338;
wire n_653;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_650;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_652;
wire n_334;
wire n_647;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_707;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_710;
wire n_703;
wire n_110;
wire n_195;
wire n_533;
wire n_592;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_651;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_689;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_615;
wire n_212;
wire n_697;
wire n_579;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_672;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_670;
wire n_524;
wire n_589;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_644;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_693;
wire n_419;
wire n_632;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_692;
wire n_49;
wire n_514;
wire n_68;
wire n_633;
wire n_497;
wire n_638;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_596;
wire n_312;
wire n_617;
wire n_325;
wire n_316;
wire n_307;
wire n_594;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_604;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_688;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_572;
wire n_586;
wire n_548;
wire n_319;
wire n_664;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_637;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_698;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_613;
wire n_231;
wire n_44;
wire n_635;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_642;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_654;
wire n_616;
wire n_377;
wire n_686;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_699;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_667;
wire n_708;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_683;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_691;
wire n_458;
wire n_677;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_701;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_628;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_675;
wire n_695;
wire n_138;
wire n_662;
wire n_217;
wire n_709;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_649;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_343;
wire n_292;
wire n_702;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_681;
wire n_287;
wire n_400;
wire n_388;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_636;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_706;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_597;
wire n_618;
wire n_609;
wire n_700;
wire n_94;
wire n_645;
wire n_687;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_705;
wire n_530;
wire n_694;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_641;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_690;
wire n_24;
wire n_92;
wire n_676;
wire n_187;
wire n_436;
wire n_629;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_659;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_660;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_625;
wire n_96;
wire n_665;
wire n_308;
wire n_433;
wire n_364;

BUFx12f_ASAP7_75t_L g144 ( 
.A(n_0),
.Y(n_144)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_0),
.Y(n_155)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_0),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_0),
.Y(n_355)
);

BUFx3_ASAP7_75t_L g577 ( 
.A(n_0),
.Y(n_577)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_1),
.A2(n_126),
.B1(n_129),
.B2(n_130),
.Y(n_125)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_1),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_1),
.A2(n_129),
.B1(n_228),
.B2(n_232),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_1),
.A2(n_129),
.B1(n_286),
.B2(n_288),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_L g653 ( 
.A1(n_1),
.A2(n_60),
.B1(n_129),
.B2(n_654),
.Y(n_653)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_2),
.A2(n_246),
.B1(n_247),
.B2(n_248),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_2),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_2),
.A2(n_246),
.B1(n_400),
.B2(n_402),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_2),
.A2(n_246),
.B1(n_501),
.B2(n_502),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_L g580 ( 
.A1(n_2),
.A2(n_246),
.B1(n_581),
.B2(n_585),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_4),
.A2(n_50),
.B1(n_51),
.B2(n_58),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_4),
.A2(n_50),
.B1(n_135),
.B2(n_138),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_4),
.A2(n_50),
.B1(n_108),
.B2(n_126),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g626 ( 
.A1(n_4),
.A2(n_50),
.B1(n_627),
.B2(n_628),
.Y(n_626)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_5),
.A2(n_207),
.B1(n_208),
.B2(n_209),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_5),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_5),
.A2(n_208),
.B1(n_235),
.B2(n_238),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_5),
.A2(n_208),
.B1(n_305),
.B2(n_309),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_5),
.A2(n_208),
.B1(n_418),
.B2(n_420),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_6),
.A2(n_63),
.B1(n_64),
.B2(n_67),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_6),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_6),
.A2(n_63),
.B1(n_148),
.B2(n_150),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_6),
.A2(n_63),
.B1(n_116),
.B2(n_275),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g647 ( 
.A1(n_6),
.A2(n_63),
.B1(n_337),
.B2(n_648),
.Y(n_647)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_7),
.A2(n_162),
.B1(n_169),
.B2(n_170),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_7),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_7),
.A2(n_170),
.B1(n_256),
.B2(n_258),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_7),
.A2(n_170),
.B1(n_384),
.B2(n_388),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_7),
.A2(n_170),
.B1(n_480),
.B2(n_483),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_8),
.Y(n_710)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_9),
.A2(n_160),
.B1(n_161),
.B2(n_164),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_9),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_9),
.A2(n_160),
.B1(n_317),
.B2(n_320),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_SL g446 ( 
.A1(n_9),
.A2(n_160),
.B1(n_447),
.B2(n_451),
.Y(n_446)
);

AOI22xp33_ASAP7_75t_SL g557 ( 
.A1(n_9),
.A2(n_160),
.B1(n_544),
.B2(n_558),
.Y(n_557)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_10),
.A2(n_115),
.B1(n_118),
.B2(n_119),
.Y(n_114)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_10),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_10),
.A2(n_118),
.B1(n_186),
.B2(n_191),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g357 ( 
.A1(n_10),
.A2(n_118),
.B1(n_358),
.B2(n_360),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g636 ( 
.A1(n_10),
.A2(n_118),
.B1(n_637),
.B2(n_639),
.Y(n_636)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_11),
.Y(n_57)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_12),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_12),
.Y(n_184)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_13),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_13),
.Y(n_140)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_13),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_13),
.Y(n_152)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_14),
.Y(n_91)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_14),
.Y(n_99)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_14),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_15),
.B(n_704),
.Y(n_703)
);

CKINVDCx11_ASAP7_75t_R g709 ( 
.A(n_15),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_16),
.B(n_343),
.Y(n_342)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_16),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_16),
.B(n_71),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_16),
.B(n_472),
.Y(n_471)
);

AOI22xp33_ASAP7_75t_L g508 ( 
.A1(n_16),
.A2(n_395),
.B1(n_509),
.B2(n_514),
.Y(n_508)
);

OAI21xp33_ASAP7_75t_L g598 ( 
.A1(n_16),
.A2(n_141),
.B(n_561),
.Y(n_598)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_17),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_17),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_17),
.Y(n_122)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_17),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_18),
.Y(n_190)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_18),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_705),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_74),
.B(n_703),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_72),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g693 ( 
.A(n_22),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_22),
.B(n_692),
.Y(n_700)
);

AOI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_49),
.B1(n_62),
.B2(n_70),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_L g73 ( 
.A1(n_23),
.A2(n_62),
.B(n_70),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g635 ( 
.A1(n_23),
.A2(n_70),
.B1(n_304),
.B2(n_636),
.Y(n_635)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_23),
.Y(n_652)
);

AOI22xp5_ASAP7_75t_L g685 ( 
.A1(n_23),
.A2(n_49),
.B1(n_70),
.B2(n_686),
.Y(n_685)
);

HB1xp67_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_24),
.B(n_159),
.Y(n_158)
);

AO22x1_ASAP7_75t_SL g244 ( 
.A1(n_24),
.A2(n_71),
.B1(n_159),
.B2(n_245),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_24),
.B(n_168),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_24),
.B(n_394),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_38),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_29),
.B1(n_32),
.B2(n_34),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g638 ( 
.A(n_26),
.Y(n_638)
);

INVx4_ASAP7_75t_SL g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g654 ( 
.A(n_27),
.Y(n_654)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g336 ( 
.A(n_31),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_31),
.Y(n_351)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_42),
.B1(n_45),
.B2(n_47),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_43),
.Y(n_209)
);

INVx4_ASAP7_75t_L g648 ( 
.A(n_43),
.Y(n_648)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_44),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_44),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_44),
.Y(n_341)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_44),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_44),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx8_ASAP7_75t_L g322 ( 
.A(n_46),
.Y(n_322)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_SL g394 ( 
.A1(n_51),
.A2(n_395),
.B(n_396),
.Y(n_394)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_56),
.Y(n_169)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_56),
.Y(n_332)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_57),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_57),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_57),
.Y(n_250)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_57),
.Y(n_308)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVxp67_ASAP7_75t_SL g309 ( 
.A(n_69),
.Y(n_309)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_70),
.Y(n_655)
);

HB1xp67_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_71),
.B(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_71),
.B(n_304),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_71),
.B(n_245),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_73),
.B(n_693),
.Y(n_704)
);

AO21x1_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_619),
.B(n_694),
.Y(n_74)
);

NAND2x1_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_434),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_371),
.B(n_430),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_78),
.B(n_616),
.Y(n_615)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_265),
.B(n_310),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_79),
.B(n_265),
.Y(n_433)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g432 ( 
.A(n_80),
.B(n_266),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_210),
.C(n_220),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_82),
.A2(n_83),
.B1(n_211),
.B2(n_370),
.Y(n_369)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_156),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_84),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_133),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_85),
.B(n_133),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_114),
.B1(n_123),
.B2(n_125),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_86),
.A2(n_123),
.B1(n_125),
.B2(n_218),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_86),
.A2(n_114),
.B1(n_123),
.B2(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_86),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g499 ( 
.A1(n_86),
.A2(n_123),
.B1(n_446),
.B2(n_500),
.Y(n_499)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_100),
.Y(n_86)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_87),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_92),
.B1(n_95),
.B2(n_97),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_88),
.A2(n_92),
.B1(n_95),
.B2(n_97),
.Y(n_124)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx6_ASAP7_75t_L g532 ( 
.A(n_90),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_93),
.Y(n_137)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_93),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_94),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_94),
.Y(n_146)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_94),
.Y(n_359)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_94),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_94),
.Y(n_487)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_96),
.Y(n_232)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx3_ASAP7_75t_L g551 ( 
.A(n_98),
.Y(n_551)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVxp67_ASAP7_75t_SL g282 ( 
.A(n_100),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_105),
.B1(n_108),
.B2(n_111),
.Y(n_100)
);

AOI22x1_ASAP7_75t_SL g173 ( 
.A1(n_101),
.A2(n_174),
.B1(n_177),
.B2(n_181),
.Y(n_173)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_103),
.Y(n_237)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_104),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_104),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_104),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_107),
.Y(n_113)
);

BUFx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_110),
.Y(n_117)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_110),
.Y(n_505)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx5_ASAP7_75t_L g390 ( 
.A(n_117),
.Y(n_390)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_117),
.Y(n_453)
);

BUFx4f_ASAP7_75t_SL g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_122),
.Y(n_128)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_124),
.B(n_283),
.Y(n_298)
);

INVxp67_ASAP7_75t_SL g296 ( 
.A(n_125),
.Y(n_296)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx3_ASAP7_75t_SL g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_SL g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

OAI22x1_ASAP7_75t_SL g133 ( 
.A1(n_134),
.A2(n_141),
.B1(n_147),
.B2(n_153),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_134),
.A2(n_224),
.B(n_226),
.Y(n_223)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx2_ASAP7_75t_SL g138 ( 
.A(n_139),
.Y(n_138)
);

BUFx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_140),
.Y(n_482)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_140),
.Y(n_549)
);

AOI21x1_ASAP7_75t_SL g212 ( 
.A1(n_141),
.A2(n_147),
.B(n_213),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_141),
.A2(n_357),
.B1(n_417),
.B2(n_423),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_L g556 ( 
.A1(n_141),
.A2(n_557),
.B(n_561),
.Y(n_556)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_142),
.B(n_227),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_142),
.A2(n_227),
.B1(n_353),
.B2(n_356),
.Y(n_352)
);

AO22x1_ASAP7_75t_SL g478 ( 
.A1(n_142),
.A2(n_479),
.B1(n_488),
.B2(n_489),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g575 ( 
.A1(n_142),
.A2(n_576),
.B1(n_578),
.B2(n_579),
.Y(n_575)
);

NAND2xp33_ASAP7_75t_R g596 ( 
.A(n_142),
.B(n_479),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_145),
.Y(n_142)
);

INVx8_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx8_ASAP7_75t_L g225 ( 
.A(n_144),
.Y(n_225)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_150),
.Y(n_560)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx6_ASAP7_75t_L g231 ( 
.A(n_152),
.Y(n_231)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_152),
.Y(n_419)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_152),
.Y(n_537)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_152),
.Y(n_607)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_153),
.Y(n_489)
);

INVx2_ASAP7_75t_SL g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_155),
.Y(n_595)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_171),
.Y(n_156)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_157),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_167),
.Y(n_157)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx11_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

BUFx12f_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_167),
.B(n_393),
.Y(n_392)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_169),
.Y(n_247)
);

INVxp33_ASAP7_75t_SL g269 ( 
.A(n_171),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_185),
.B1(n_194),
.B2(n_206),
.Y(n_171)
);

INVx2_ASAP7_75t_SL g263 ( 
.A(n_172),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_172),
.A2(n_185),
.B1(n_285),
.B2(n_292),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_172),
.B(n_255),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_172),
.A2(n_194),
.B1(n_398),
.B2(n_399),
.Y(n_397)
);

AO22x1_ASAP7_75t_L g625 ( 
.A1(n_172),
.A2(n_194),
.B1(n_285),
.B2(n_626),
.Y(n_625)
);

AOI22xp5_ASAP7_75t_L g646 ( 
.A1(n_172),
.A2(n_194),
.B1(n_626),
.B2(n_647),
.Y(n_646)
);

OAI21xp33_ASAP7_75t_SL g684 ( 
.A1(n_172),
.A2(n_194),
.B(n_647),
.Y(n_684)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

AND2x4_ASAP7_75t_L g194 ( 
.A(n_173),
.B(n_195),
.Y(n_194)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_175),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_179),
.Y(n_477)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_180),
.Y(n_241)
);

BUFx5_ASAP7_75t_L g278 ( 
.A(n_180),
.Y(n_278)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_184),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g469 ( 
.A(n_184),
.Y(n_469)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_189),
.Y(n_207)
);

INVx8_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx4_ASAP7_75t_L g633 ( 
.A(n_192),
.Y(n_633)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_193),
.Y(n_197)
);

BUFx5_ASAP7_75t_L g202 ( 
.A(n_193),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g513 ( 
.A(n_193),
.Y(n_513)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_194),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g292 ( 
.A(n_194),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_194),
.B(n_255),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_198),
.B1(n_200),
.B2(n_203),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_197),
.Y(n_465)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_202),
.Y(n_287)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_206),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVxp67_ASAP7_75t_SL g370 ( 
.A(n_211),
.Y(n_370)
);

OAI21xp33_ASAP7_75t_SL g211 ( 
.A1(n_212),
.A2(n_216),
.B(n_219),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_212),
.B(n_216),
.Y(n_219)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_212),
.Y(n_299)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

BUFx4f_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVxp67_ASAP7_75t_SL g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_218),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_219),
.B(n_301),
.Y(n_663)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_221),
.B(n_369),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_242),
.B(n_264),
.Y(n_221)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_222),
.Y(n_365)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_233),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_223),
.B(n_233),
.Y(n_405)
);

BUFx3_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx5_ASAP7_75t_L g562 ( 
.A(n_225),
.Y(n_562)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

BUFx2_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_231),
.Y(n_361)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_234),
.Y(n_391)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_236),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx2_ASAP7_75t_SL g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx5_ASAP7_75t_L g461 ( 
.A(n_241),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_251),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_243),
.B(n_251),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_243),
.A2(n_244),
.B1(n_252),
.B2(n_367),
.Y(n_366)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVxp33_ASAP7_75t_SL g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_252),
.Y(n_367)
);

OAI22x1_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_254),
.B1(n_262),
.B2(n_263),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_253),
.A2(n_316),
.B(n_323),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g507 ( 
.A1(n_253),
.A2(n_323),
.B(n_508),
.Y(n_507)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_257),
.Y(n_291)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx2_ASAP7_75t_SL g319 ( 
.A(n_261),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_261),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_L g413 ( 
.A1(n_263),
.A2(n_414),
.B(n_415),
.Y(n_413)
);

NOR2x1_ASAP7_75t_R g564 ( 
.A(n_263),
.B(n_395),
.Y(n_564)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_271),
.Y(n_266)
);

INVxp67_ASAP7_75t_SL g669 ( 
.A(n_267),
.Y(n_669)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.C(n_270),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_293),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g668 ( 
.A(n_272),
.Y(n_668)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_284),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_273),
.B(n_284),
.Y(n_664)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_279),
.B1(n_281),
.B2(n_283),
.Y(n_273)
);

OA21x2_ASAP7_75t_L g641 ( 
.A1(n_274),
.A2(n_279),
.B(n_281),
.Y(n_641)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

HB1xp67_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_278),
.Y(n_387)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_278),
.Y(n_542)
);

AOI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_279),
.A2(n_281),
.B1(n_383),
.B2(n_391),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_279),
.B(n_383),
.Y(n_454)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_280),
.B(n_282),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g568 ( 
.A(n_280),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_281),
.B(n_554),
.Y(n_553)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_281),
.Y(n_566)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

BUFx3_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g667 ( 
.A(n_293),
.Y(n_667)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_300),
.Y(n_293)
);

AO21x1_ASAP7_75t_L g294 ( 
.A1(n_295),
.A2(n_298),
.B(n_299),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_297),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_301),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_303),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_302),
.B(n_326),
.Y(n_325)
);

INVx3_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx4_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_308),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_368),
.Y(n_310)
);

OR2x2_ASAP7_75t_L g431 ( 
.A(n_311),
.B(n_368),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_362),
.C(n_363),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_312),
.B(n_374),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_324),
.C(n_327),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_314),
.A2(n_315),
.B1(n_324),
.B2(n_325),
.Y(n_380)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_316),
.Y(n_398)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

BUFx2_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx4_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_328),
.B(n_380),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_352),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_329),
.B(n_352),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_330),
.A2(n_333),
.B1(n_342),
.B2(n_345),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_337),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_341),
.Y(n_401)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_342),
.Y(n_396)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_343),
.Y(n_640)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

NAND2xp33_ASAP7_75t_SL g345 ( 
.A(n_346),
.B(n_349),
.Y(n_345)
);

BUFx2_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

HB1xp67_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

BUFx3_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

HB1xp67_ASAP7_75t_L g424 ( 
.A(n_355),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_355),
.Y(n_604)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx3_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_362),
.A2(n_364),
.B1(n_375),
.B2(n_376),
.Y(n_374)
);

INVxp67_ASAP7_75t_SL g376 ( 
.A(n_362),
.Y(n_376)
);

INVxp67_ASAP7_75t_SL g363 ( 
.A(n_364),
.Y(n_363)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_364),
.Y(n_375)
);

XNOR2x1_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_366),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_377),
.C(n_406),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_L g616 ( 
.A1(n_373),
.A2(n_617),
.B(n_618),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_377),
.Y(n_617)
);

MAJx2_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_381),
.C(n_404),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_378),
.A2(n_379),
.B1(n_428),
.B2(n_429),
.Y(n_427)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

XNOR2x1_ASAP7_75t_L g428 ( 
.A(n_381),
.B(n_405),
.Y(n_428)
);

MAJx2_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_392),
.C(n_397),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_382),
.B(n_397),
.Y(n_409)
);

INVxp67_ASAP7_75t_SL g567 ( 
.A(n_383),
.Y(n_567)
);

INVx4_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx3_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

BUFx2_ASAP7_75t_L g501 ( 
.A(n_387),
.Y(n_501)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_392),
.B(n_409),
.Y(n_408)
);

OAI211xp5_ASAP7_75t_L g457 ( 
.A1(n_395),
.A2(n_458),
.B(n_462),
.C(n_466),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_395),
.B(n_540),
.Y(n_539)
);

OAI21xp33_ASAP7_75t_SL g554 ( 
.A1(n_395),
.A2(n_448),
.B(n_539),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_395),
.B(n_568),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_395),
.B(n_601),
.Y(n_600)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_399),
.Y(n_414)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_402),
.Y(n_627)
);

INVx4_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_403),
.Y(n_472)
);

HB1xp67_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

OR2x2_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_427),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_407),
.B(n_427),
.Y(n_618)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_410),
.C(n_411),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_SL g490 ( 
.A(n_408),
.B(n_491),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_410),
.A2(n_411),
.B1(n_412),
.B2(n_492),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_410),
.Y(n_492)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_413),
.B(n_416),
.C(n_425),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_413),
.B(n_441),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_416),
.A2(n_425),
.B1(n_426),
.B2(n_442),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_416),
.Y(n_442)
);

INVxp33_ASAP7_75t_SL g488 ( 
.A(n_417),
.Y(n_488)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

BUFx2_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g587 ( 
.A(n_422),
.Y(n_587)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_428),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_L g430 ( 
.A1(n_431),
.A2(n_432),
.B(n_433),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_435),
.B(n_615),
.Y(n_434)
);

OAI21x1_ASAP7_75t_L g435 ( 
.A1(n_436),
.A2(n_493),
.B(n_613),
.Y(n_435)
);

AND2x4_ASAP7_75t_L g436 ( 
.A(n_437),
.B(n_490),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_438),
.B(n_614),
.Y(n_613)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_439),
.B(n_443),
.C(n_455),
.Y(n_438)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_440),
.B(n_496),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_L g496 ( 
.A1(n_443),
.A2(n_444),
.B1(n_455),
.B2(n_497),
.Y(n_496)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

OAI21xp5_ASAP7_75t_SL g444 ( 
.A1(n_445),
.A2(n_446),
.B(n_454),
.Y(n_444)
);

INVx1_ASAP7_75t_SL g447 ( 
.A(n_448),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

INVx4_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

INVx1_ASAP7_75t_SL g451 ( 
.A(n_452),
.Y(n_451)
);

BUFx2_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g552 ( 
.A(n_454),
.B(n_553),
.Y(n_552)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_455),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_456),
.B(n_478),
.Y(n_455)
);

XOR2x1_ASAP7_75t_L g518 ( 
.A(n_456),
.B(n_478),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_457),
.B(n_470),
.Y(n_456)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

HB1xp67_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

INVx3_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_471),
.B(n_473),
.Y(n_470)
);

INVxp67_ASAP7_75t_SL g473 ( 
.A(n_474),
.Y(n_473)
);

BUFx2_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

NAND2xp33_ASAP7_75t_SL g561 ( 
.A(n_479),
.B(n_562),
.Y(n_561)
);

INVx1_ASAP7_75t_SL g480 ( 
.A(n_481),
.Y(n_480)
);

BUFx2_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

INVx4_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

INVxp67_ASAP7_75t_SL g614 ( 
.A(n_490),
.Y(n_614)
);

AOI21x1_ASAP7_75t_L g493 ( 
.A1(n_494),
.A2(n_519),
.B(n_612),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_495),
.B(n_498),
.Y(n_494)
);

NOR2x1_ASAP7_75t_L g612 ( 
.A(n_495),
.B(n_498),
.Y(n_612)
);

MAJIxp5_ASAP7_75t_SL g498 ( 
.A(n_499),
.B(n_506),
.C(n_518),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_L g572 ( 
.A(n_499),
.B(n_507),
.Y(n_572)
);

OAI22xp5_ASAP7_75t_L g565 ( 
.A1(n_500),
.A2(n_566),
.B1(n_567),
.B2(n_568),
.Y(n_565)
);

BUFx4f_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

INVx4_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

INVx4_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

HB1xp67_ASAP7_75t_L g506 ( 
.A(n_507),
.Y(n_506)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

BUFx2_ASAP7_75t_SL g510 ( 
.A(n_511),
.Y(n_510)
);

HB1xp67_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

BUFx3_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

INVx3_ASAP7_75t_L g515 ( 
.A(n_516),
.Y(n_515)
);

INVx4_ASAP7_75t_L g516 ( 
.A(n_517),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g571 ( 
.A(n_518),
.B(n_572),
.Y(n_571)
);

OAI321xp33_ASAP7_75t_L g519 ( 
.A1(n_520),
.A2(n_569),
.A3(n_573),
.B1(n_610),
.B2(n_611),
.C(n_712),
.Y(n_519)
);

NOR2xp67_ASAP7_75t_L g520 ( 
.A(n_521),
.B(n_555),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_521),
.B(n_555),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_522),
.B(n_552),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g588 ( 
.A(n_522),
.B(n_552),
.Y(n_588)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_523),
.A2(n_533),
.B1(n_538),
.B2(n_543),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_524),
.B(n_528),
.Y(n_523)
);

HB1xp67_ASAP7_75t_L g524 ( 
.A(n_525),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_526),
.Y(n_525)
);

HB1xp67_ASAP7_75t_L g526 ( 
.A(n_527),
.Y(n_526)
);

BUFx2_ASAP7_75t_L g528 ( 
.A(n_529),
.Y(n_528)
);

HB1xp67_ASAP7_75t_L g529 ( 
.A(n_530),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_531),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_532),
.Y(n_531)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_534),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_535),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_536),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_537),
.Y(n_536)
);

INVxp67_ASAP7_75t_L g538 ( 
.A(n_539),
.Y(n_538)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_541),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_542),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_544),
.B(n_550),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_545),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_546),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_547),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_548),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_549),
.Y(n_548)
);

INVx2_ASAP7_75t_SL g550 ( 
.A(n_551),
.Y(n_550)
);

XNOR2xp5_ASAP7_75t_L g555 ( 
.A(n_556),
.B(n_563),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_556),
.B(n_564),
.C(n_565),
.Y(n_570)
);

INVxp67_ASAP7_75t_L g578 ( 
.A(n_557),
.Y(n_578)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_559),
.Y(n_558)
);

BUFx2_ASAP7_75t_SL g559 ( 
.A(n_560),
.Y(n_559)
);

XNOR2xp5_ASAP7_75t_L g563 ( 
.A(n_564),
.B(n_565),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_570),
.B(n_571),
.Y(n_569)
);

OR2x2_ASAP7_75t_L g611 ( 
.A(n_570),
.B(n_571),
.Y(n_611)
);

AOI21xp5_ASAP7_75t_L g573 ( 
.A1(n_574),
.A2(n_589),
.B(n_609),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_575),
.B(n_588),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_575),
.B(n_588),
.Y(n_609)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_577),
.Y(n_576)
);

INVxp67_ASAP7_75t_L g579 ( 
.A(n_580),
.Y(n_579)
);

OAI21xp5_ASAP7_75t_SL g592 ( 
.A1(n_580),
.A2(n_593),
.B(n_596),
.Y(n_592)
);

BUFx2_ASAP7_75t_L g581 ( 
.A(n_582),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_583),
.Y(n_582)
);

BUFx2_ASAP7_75t_SL g583 ( 
.A(n_584),
.Y(n_583)
);

INVx3_ASAP7_75t_L g585 ( 
.A(n_586),
.Y(n_585)
);

INVx5_ASAP7_75t_L g586 ( 
.A(n_587),
.Y(n_586)
);

OAI21xp5_ASAP7_75t_SL g589 ( 
.A1(n_590),
.A2(n_597),
.B(n_608),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_591),
.B(n_592),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_591),
.B(n_592),
.Y(n_608)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_594),
.Y(n_593)
);

BUFx2_ASAP7_75t_L g594 ( 
.A(n_595),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_598),
.B(n_599),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_SL g599 ( 
.A(n_600),
.B(n_605),
.Y(n_599)
);

BUFx6f_ASAP7_75t_L g601 ( 
.A(n_602),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_603),
.Y(n_602)
);

BUFx2_ASAP7_75t_L g603 ( 
.A(n_604),
.Y(n_603)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_606),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_607),
.Y(n_606)
);

NOR3xp33_ASAP7_75t_L g619 ( 
.A(n_620),
.B(n_674),
.C(n_689),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_621),
.B(n_665),
.Y(n_620)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_621),
.Y(n_697)
);

OAI21xp5_ASAP7_75t_L g621 ( 
.A1(n_622),
.A2(n_656),
.B(n_657),
.Y(n_621)
);

NOR3xp33_ASAP7_75t_L g702 ( 
.A(n_622),
.B(n_656),
.C(n_657),
.Y(n_702)
);

NOR2xp67_ASAP7_75t_L g622 ( 
.A(n_623),
.B(n_642),
.Y(n_622)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_623),
.B(n_642),
.Y(n_656)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_623),
.Y(n_677)
);

MAJIxp5_ASAP7_75t_L g623 ( 
.A(n_624),
.B(n_634),
.C(n_641),
.Y(n_623)
);

HB1xp67_ASAP7_75t_L g624 ( 
.A(n_625),
.Y(n_624)
);

OAI22xp5_ASAP7_75t_L g660 ( 
.A1(n_625),
.A2(n_641),
.B1(n_645),
.B2(n_661),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_625),
.Y(n_661)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_629),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_630),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_631),
.Y(n_630)
);

INVx3_ASAP7_75t_L g631 ( 
.A(n_632),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_633),
.Y(n_632)
);

XNOR2xp5_ASAP7_75t_L g642 ( 
.A(n_634),
.B(n_643),
.Y(n_642)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_634),
.Y(n_678)
);

BUFx2_ASAP7_75t_L g634 ( 
.A(n_635),
.Y(n_634)
);

XNOR2xp5_ASAP7_75t_L g659 ( 
.A(n_635),
.B(n_660),
.Y(n_659)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_636),
.Y(n_651)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_638),
.Y(n_637)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_640),
.Y(n_639)
);

AOI22xp5_ASAP7_75t_L g644 ( 
.A1(n_641),
.A2(n_645),
.B1(n_646),
.B2(n_649),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_641),
.Y(n_645)
);

INVxp33_ASAP7_75t_SL g679 ( 
.A(n_643),
.Y(n_679)
);

XOR2x2_ASAP7_75t_L g643 ( 
.A(n_644),
.B(n_650),
.Y(n_643)
);

MAJIxp5_ASAP7_75t_SL g681 ( 
.A(n_645),
.B(n_649),
.C(n_682),
.Y(n_681)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_646),
.Y(n_649)
);

HB1xp67_ASAP7_75t_L g682 ( 
.A(n_650),
.Y(n_682)
);

OAI22xp5_ASAP7_75t_L g650 ( 
.A1(n_651),
.A2(n_652),
.B1(n_653),
.B2(n_655),
.Y(n_650)
);

INVxp67_ASAP7_75t_L g686 ( 
.A(n_653),
.Y(n_686)
);

MAJIxp5_ASAP7_75t_L g657 ( 
.A(n_658),
.B(n_662),
.C(n_664),
.Y(n_657)
);

HB1xp67_ASAP7_75t_L g658 ( 
.A(n_659),
.Y(n_658)
);

OAI22xp5_ASAP7_75t_L g671 ( 
.A1(n_659),
.A2(n_664),
.B1(n_672),
.B2(n_673),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_659),
.Y(n_672)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_663),
.Y(n_662)
);

XNOR2xp5_ASAP7_75t_L g670 ( 
.A(n_663),
.B(n_671),
.Y(n_670)
);

INVxp67_ASAP7_75t_L g673 ( 
.A(n_664),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_666),
.B(n_670),
.Y(n_665)
);

NOR2xp67_ASAP7_75t_L g696 ( 
.A(n_666),
.B(n_670),
.Y(n_696)
);

MAJIxp5_ASAP7_75t_L g666 ( 
.A(n_667),
.B(n_668),
.C(n_669),
.Y(n_666)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_675),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_675),
.B(n_696),
.Y(n_695)
);

NAND3xp33_ASAP7_75t_L g701 ( 
.A(n_675),
.B(n_690),
.C(n_702),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_676),
.B(n_680),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_676),
.B(n_680),
.Y(n_699)
);

MAJIxp5_ASAP7_75t_L g676 ( 
.A(n_677),
.B(n_678),
.C(n_679),
.Y(n_676)
);

XNOR2xp5_ASAP7_75t_L g680 ( 
.A(n_681),
.B(n_683),
.Y(n_680)
);

MAJIxp5_ASAP7_75t_L g692 ( 
.A(n_681),
.B(n_685),
.C(n_687),
.Y(n_692)
);

AOI22xp5_ASAP7_75t_SL g683 ( 
.A1(n_684),
.A2(n_685),
.B1(n_687),
.B2(n_688),
.Y(n_683)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_684),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_685),
.Y(n_688)
);

OAI311xp33_ASAP7_75t_L g694 ( 
.A1(n_689),
.A2(n_695),
.A3(n_697),
.B1(n_698),
.C1(n_701),
.Y(n_694)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_690),
.Y(n_689)
);

AOI21xp33_ASAP7_75t_L g698 ( 
.A1(n_690),
.A2(n_699),
.B(n_700),
.Y(n_698)
);

NAND2x1_ASAP7_75t_L g690 ( 
.A(n_691),
.B(n_693),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_692),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_706),
.B(n_710),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_707),
.Y(n_706)
);

BUFx4f_ASAP7_75t_SL g707 ( 
.A(n_708),
.Y(n_707)
);

BUFx12f_ASAP7_75t_L g708 ( 
.A(n_709),
.Y(n_708)
);


endmodule