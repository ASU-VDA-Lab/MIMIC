module fake_netlist_6_1289_n_1782 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1782);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1782;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1371;
wire n_1285;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1517;
wire n_1393;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1757;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1373;
wire n_1292;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1721;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_59),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_77),
.Y(n_171)
);

BUFx10_ASAP7_75t_L g172 ( 
.A(n_118),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_124),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_32),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_110),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_145),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_104),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_26),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_120),
.Y(n_179)
);

CKINVDCx14_ASAP7_75t_R g180 ( 
.A(n_22),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_146),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_18),
.Y(n_182)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_160),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_116),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_14),
.Y(n_185)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_37),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_52),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_140),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_50),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_28),
.Y(n_190)
);

BUFx2_ASAP7_75t_L g191 ( 
.A(n_169),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_119),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_113),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_39),
.Y(n_194)
);

BUFx2_ASAP7_75t_L g195 ( 
.A(n_46),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_135),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_20),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_26),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_167),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_60),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_7),
.Y(n_201)
);

BUFx2_ASAP7_75t_L g202 ( 
.A(n_64),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_45),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_99),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_31),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_92),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_40),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_81),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_7),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_37),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_13),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_153),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_40),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_63),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_166),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_45),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_95),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_154),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_49),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_141),
.Y(n_220)
);

BUFx8_ASAP7_75t_SL g221 ( 
.A(n_71),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_16),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_53),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_122),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_158),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_91),
.Y(n_226)
);

BUFx10_ASAP7_75t_L g227 ( 
.A(n_164),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_80),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_3),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_32),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_96),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_121),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_25),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_105),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_75),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_168),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_100),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_5),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_58),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_18),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_3),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_111),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_163),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_74),
.Y(n_244)
);

BUFx10_ASAP7_75t_L g245 ( 
.A(n_107),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_38),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_94),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_13),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_1),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_129),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_34),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_23),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_123),
.Y(n_253)
);

BUFx2_ASAP7_75t_L g254 ( 
.A(n_127),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_47),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_43),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_76),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_33),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_6),
.Y(n_259)
);

INVx1_ASAP7_75t_SL g260 ( 
.A(n_97),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_131),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_41),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_62),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_108),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_70),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_98),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_149),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_67),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_165),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_39),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_15),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_61),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_1),
.Y(n_273)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_152),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_82),
.Y(n_275)
);

HB1xp67_ASAP7_75t_L g276 ( 
.A(n_73),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_69),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_12),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_25),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_85),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_4),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_29),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_21),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_87),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_34),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_115),
.Y(n_286)
);

INVx1_ASAP7_75t_SL g287 ( 
.A(n_52),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_159),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_157),
.Y(n_289)
);

INVx2_ASAP7_75t_SL g290 ( 
.A(n_30),
.Y(n_290)
);

INVx2_ASAP7_75t_SL g291 ( 
.A(n_24),
.Y(n_291)
);

INVx1_ASAP7_75t_SL g292 ( 
.A(n_6),
.Y(n_292)
);

INVx1_ASAP7_75t_SL g293 ( 
.A(n_144),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_36),
.Y(n_294)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_125),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_2),
.Y(n_296)
);

CKINVDCx14_ASAP7_75t_R g297 ( 
.A(n_84),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_11),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_143),
.Y(n_299)
);

BUFx2_ASAP7_75t_L g300 ( 
.A(n_53),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_132),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_51),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_43),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_78),
.Y(n_304)
);

BUFx2_ASAP7_75t_L g305 ( 
.A(n_150),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_29),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_24),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_35),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_9),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_27),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_156),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_48),
.Y(n_312)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_155),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_93),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_89),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_4),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_101),
.Y(n_317)
);

CKINVDCx11_ASAP7_75t_R g318 ( 
.A(n_109),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_138),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_44),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_137),
.Y(n_321)
);

BUFx10_ASAP7_75t_L g322 ( 
.A(n_20),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_5),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_14),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_128),
.Y(n_325)
);

INVx2_ASAP7_75t_SL g326 ( 
.A(n_57),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_88),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_21),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_103),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_86),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_55),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_114),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_79),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_117),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_130),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_48),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_35),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_193),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_203),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_204),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_203),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_221),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_203),
.Y(n_343)
);

INVxp67_ASAP7_75t_SL g344 ( 
.A(n_276),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_224),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_203),
.Y(n_346)
);

BUFx2_ASAP7_75t_L g347 ( 
.A(n_195),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_203),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_235),
.Y(n_349)
);

INVx1_ASAP7_75t_SL g350 ( 
.A(n_300),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_174),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_236),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_199),
.Y(n_353)
);

INVxp67_ASAP7_75t_SL g354 ( 
.A(n_191),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_318),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_263),
.Y(n_356)
);

HB1xp67_ASAP7_75t_L g357 ( 
.A(n_302),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_174),
.Y(n_358)
);

BUFx3_ASAP7_75t_L g359 ( 
.A(n_295),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_170),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_238),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_238),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_197),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g364 ( 
.A(n_186),
.Y(n_364)
);

CKINVDCx14_ASAP7_75t_R g365 ( 
.A(n_180),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_197),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_313),
.Y(n_367)
);

INVxp33_ASAP7_75t_SL g368 ( 
.A(n_207),
.Y(n_368)
);

CKINVDCx16_ASAP7_75t_R g369 ( 
.A(n_176),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_217),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_230),
.Y(n_371)
);

CKINVDCx16_ASAP7_75t_R g372 ( 
.A(n_297),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_218),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_228),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_234),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_230),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_248),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_182),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_243),
.Y(n_379)
);

INVxp33_ASAP7_75t_L g380 ( 
.A(n_223),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_185),
.Y(n_381)
);

HB1xp67_ASAP7_75t_L g382 ( 
.A(n_187),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_247),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_257),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_190),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_209),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_210),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_213),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_264),
.Y(n_389)
);

INVxp67_ASAP7_75t_SL g390 ( 
.A(n_202),
.Y(n_390)
);

INVxp33_ASAP7_75t_L g391 ( 
.A(n_240),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_241),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_252),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_255),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_256),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_265),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_266),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_267),
.Y(n_398)
);

BUFx3_ASAP7_75t_L g399 ( 
.A(n_295),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_271),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_279),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_281),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_268),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_282),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_272),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_283),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_322),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_280),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_310),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_323),
.Y(n_410)
);

BUFx2_ASAP7_75t_L g411 ( 
.A(n_187),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_286),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_290),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_289),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_205),
.Y(n_415)
);

INVx1_ASAP7_75t_SL g416 ( 
.A(n_246),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_290),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_291),
.Y(n_418)
);

INVxp33_ASAP7_75t_L g419 ( 
.A(n_254),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_291),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_353),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_SL g422 ( 
.A(n_350),
.B(n_172),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_353),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_370),
.B(n_326),
.Y(n_424)
);

AND2x4_ASAP7_75t_L g425 ( 
.A(n_339),
.B(n_183),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_359),
.B(n_305),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_339),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_419),
.B(n_326),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_353),
.Y(n_429)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_357),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_353),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_373),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_341),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_341),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_353),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_343),
.Y(n_436)
);

INVx3_ASAP7_75t_L g437 ( 
.A(n_343),
.Y(n_437)
);

BUFx3_ASAP7_75t_L g438 ( 
.A(n_359),
.Y(n_438)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_346),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_346),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_348),
.Y(n_441)
);

AND2x4_ASAP7_75t_L g442 ( 
.A(n_348),
.B(n_183),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_386),
.Y(n_443)
);

AND2x2_ASAP7_75t_L g444 ( 
.A(n_399),
.B(n_172),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_374),
.B(n_183),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_338),
.Y(n_446)
);

INVx4_ASAP7_75t_L g447 ( 
.A(n_375),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_351),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_379),
.B(n_184),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_351),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_358),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_381),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_340),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_345),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_358),
.Y(n_455)
);

INVx3_ASAP7_75t_L g456 ( 
.A(n_361),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_383),
.Y(n_457)
);

NAND2xp33_ASAP7_75t_L g458 ( 
.A(n_415),
.B(n_189),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_384),
.B(n_184),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_381),
.Y(n_460)
);

INVxp67_ASAP7_75t_L g461 ( 
.A(n_382),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_349),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_396),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_385),
.Y(n_464)
);

INVx6_ASAP7_75t_L g465 ( 
.A(n_399),
.Y(n_465)
);

AND2x4_ASAP7_75t_L g466 ( 
.A(n_363),
.B(n_261),
.Y(n_466)
);

OR2x2_ASAP7_75t_L g467 ( 
.A(n_411),
.B(n_178),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_361),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_385),
.Y(n_469)
);

HB1xp67_ASAP7_75t_L g470 ( 
.A(n_416),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_397),
.B(n_261),
.Y(n_471)
);

HB1xp67_ASAP7_75t_L g472 ( 
.A(n_365),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_387),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_387),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_362),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_388),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_388),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_408),
.B(n_284),
.Y(n_478)
);

HB1xp67_ASAP7_75t_L g479 ( 
.A(n_412),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_344),
.B(n_284),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_392),
.Y(n_481)
);

AND2x6_ASAP7_75t_L g482 ( 
.A(n_362),
.B(n_199),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g483 ( 
.A(n_392),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_342),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_393),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_R g486 ( 
.A(n_355),
.B(n_179),
.Y(n_486)
);

INVx3_ASAP7_75t_L g487 ( 
.A(n_394),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_394),
.Y(n_488)
);

INVx3_ASAP7_75t_L g489 ( 
.A(n_395),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_395),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_400),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_400),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_401),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_401),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_437),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_483),
.Y(n_496)
);

INVx3_ASAP7_75t_L g497 ( 
.A(n_421),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_437),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_445),
.B(n_369),
.Y(n_499)
);

INVx8_ASAP7_75t_L g500 ( 
.A(n_482),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_422),
.B(n_372),
.Y(n_501)
);

AND2x4_ASAP7_75t_L g502 ( 
.A(n_425),
.B(n_304),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_421),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_437),
.Y(n_504)
);

OAI21xp33_ASAP7_75t_L g505 ( 
.A1(n_480),
.A2(n_391),
.B(n_390),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_427),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_483),
.Y(n_507)
);

INVxp33_ASAP7_75t_L g508 ( 
.A(n_470),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_427),
.Y(n_509)
);

NAND3xp33_ASAP7_75t_L g510 ( 
.A(n_449),
.B(n_378),
.C(n_220),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_448),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_459),
.B(n_354),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_448),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_448),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_483),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g516 ( 
.A(n_421),
.Y(n_516)
);

INVx3_ASAP7_75t_L g517 ( 
.A(n_421),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_471),
.B(n_212),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_483),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_466),
.B(n_363),
.Y(n_520)
);

HB1xp67_ASAP7_75t_L g521 ( 
.A(n_438),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_483),
.Y(n_522)
);

AND2x4_ASAP7_75t_L g523 ( 
.A(n_425),
.B(n_304),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_448),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_448),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_421),
.Y(n_526)
);

INVx2_ASAP7_75t_SL g527 ( 
.A(n_444),
.Y(n_527)
);

BUFx6f_ASAP7_75t_SL g528 ( 
.A(n_447),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_448),
.Y(n_529)
);

NAND2xp33_ASAP7_75t_L g530 ( 
.A(n_424),
.B(n_199),
.Y(n_530)
);

INVx1_ASAP7_75t_SL g531 ( 
.A(n_446),
.Y(n_531)
);

INVx3_ASAP7_75t_L g532 ( 
.A(n_421),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_483),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_450),
.Y(n_534)
);

AO21x2_ASAP7_75t_L g535 ( 
.A1(n_478),
.A2(n_173),
.B(n_171),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_450),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_450),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_450),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_444),
.B(n_232),
.Y(n_539)
);

INVxp33_ASAP7_75t_L g540 ( 
.A(n_467),
.Y(n_540)
);

INVx3_ASAP7_75t_L g541 ( 
.A(n_423),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_433),
.Y(n_542)
);

OR2x6_ASAP7_75t_L g543 ( 
.A(n_447),
.B(n_175),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_466),
.B(n_366),
.Y(n_544)
);

BUFx6f_ASAP7_75t_L g545 ( 
.A(n_423),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_437),
.Y(n_546)
);

INVx2_ASAP7_75t_SL g547 ( 
.A(n_465),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_439),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_438),
.B(n_260),
.Y(n_549)
);

INVx4_ASAP7_75t_L g550 ( 
.A(n_440),
.Y(n_550)
);

INVx2_ASAP7_75t_SL g551 ( 
.A(n_465),
.Y(n_551)
);

AOI22xp33_ASAP7_75t_L g552 ( 
.A1(n_466),
.A2(n_368),
.B1(n_347),
.B2(n_364),
.Y(n_552)
);

OR2x6_ASAP7_75t_L g553 ( 
.A(n_447),
.B(n_177),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_434),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_434),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_436),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_436),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_441),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_439),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_439),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_441),
.Y(n_561)
);

AOI21x1_ASAP7_75t_L g562 ( 
.A1(n_425),
.A2(n_192),
.B(n_181),
.Y(n_562)
);

NOR2x1p5_ASAP7_75t_L g563 ( 
.A(n_447),
.B(n_189),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_487),
.Y(n_564)
);

INVxp67_ASAP7_75t_SL g565 ( 
.A(n_438),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_450),
.Y(n_566)
);

OAI22xp5_ASAP7_75t_L g567 ( 
.A1(n_461),
.A2(n_405),
.B1(n_414),
.B2(n_398),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_432),
.Y(n_568)
);

INVx4_ASAP7_75t_L g569 ( 
.A(n_440),
.Y(n_569)
);

AND2x2_ASAP7_75t_SL g570 ( 
.A(n_458),
.B(n_215),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_428),
.B(n_389),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_450),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_487),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_439),
.Y(n_574)
);

INVx3_ASAP7_75t_L g575 ( 
.A(n_423),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_440),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_440),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_426),
.B(n_274),
.Y(n_578)
);

NAND3xp33_ASAP7_75t_L g579 ( 
.A(n_466),
.B(n_376),
.C(n_371),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_440),
.Y(n_580)
);

INVx1_ASAP7_75t_SL g581 ( 
.A(n_453),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_465),
.B(n_403),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_457),
.B(n_360),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g584 ( 
.A(n_426),
.B(n_366),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_487),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_463),
.B(n_367),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_440),
.Y(n_587)
);

INVx2_ASAP7_75t_SL g588 ( 
.A(n_465),
.Y(n_588)
);

INVx3_ASAP7_75t_L g589 ( 
.A(n_423),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_425),
.B(n_293),
.Y(n_590)
);

INVx4_ASAP7_75t_L g591 ( 
.A(n_482),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_489),
.Y(n_592)
);

AOI21x1_ASAP7_75t_L g593 ( 
.A1(n_442),
.A2(n_208),
.B(n_206),
.Y(n_593)
);

INVx2_ASAP7_75t_SL g594 ( 
.A(n_467),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_430),
.B(n_380),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_423),
.Y(n_596)
);

OAI22xp33_ASAP7_75t_L g597 ( 
.A1(n_479),
.A2(n_292),
.B1(n_287),
.B2(n_347),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_423),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_489),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_435),
.Y(n_600)
);

INVx2_ASAP7_75t_SL g601 ( 
.A(n_442),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_456),
.Y(n_602)
);

BUFx3_ASAP7_75t_L g603 ( 
.A(n_442),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_456),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_472),
.B(n_411),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_489),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_456),
.Y(n_607)
);

OR2x6_ASAP7_75t_L g608 ( 
.A(n_493),
.B(n_214),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_442),
.B(n_225),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_456),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_489),
.B(n_226),
.Y(n_611)
);

INVx3_ASAP7_75t_L g612 ( 
.A(n_435),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_490),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_429),
.B(n_231),
.Y(n_614)
);

NAND2xp33_ASAP7_75t_L g615 ( 
.A(n_482),
.B(n_215),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_490),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_452),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_451),
.Y(n_618)
);

AOI22xp33_ASAP7_75t_SL g619 ( 
.A1(n_486),
.A2(n_262),
.B1(n_336),
.B2(n_356),
.Y(n_619)
);

NOR2x1p5_ASAP7_75t_L g620 ( 
.A(n_484),
.B(n_194),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_452),
.B(n_460),
.Y(n_621)
);

OAI22xp33_ASAP7_75t_L g622 ( 
.A1(n_460),
.A2(n_233),
.B1(n_211),
.B2(n_219),
.Y(n_622)
);

INVx2_ASAP7_75t_SL g623 ( 
.A(n_464),
.Y(n_623)
);

INVxp67_ASAP7_75t_SL g624 ( 
.A(n_435),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_451),
.Y(n_625)
);

HB1xp67_ASAP7_75t_L g626 ( 
.A(n_464),
.Y(n_626)
);

CKINVDCx6p67_ASAP7_75t_R g627 ( 
.A(n_454),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_451),
.Y(n_628)
);

BUFx4f_ASAP7_75t_L g629 ( 
.A(n_482),
.Y(n_629)
);

NOR2x1p5_ASAP7_75t_L g630 ( 
.A(n_469),
.B(n_194),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_469),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_473),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_429),
.B(n_237),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_473),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_474),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_476),
.Y(n_636)
);

AOI21x1_ASAP7_75t_L g637 ( 
.A1(n_429),
.A2(n_239),
.B(n_250),
.Y(n_637)
);

OAI21xp33_ASAP7_75t_SL g638 ( 
.A1(n_476),
.A2(n_377),
.B(n_418),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_435),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_477),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_435),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_623),
.B(n_431),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_495),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_623),
.B(n_431),
.Y(n_644)
);

AOI22xp33_ASAP7_75t_L g645 ( 
.A1(n_570),
.A2(n_317),
.B1(n_215),
.B2(n_325),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_512),
.B(n_407),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_518),
.B(n_179),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_570),
.B(n_431),
.Y(n_648)
);

AND2x4_ASAP7_75t_L g649 ( 
.A(n_565),
.B(n_477),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_570),
.B(n_269),
.Y(n_650)
);

NOR2xp67_ASAP7_75t_L g651 ( 
.A(n_567),
.B(n_494),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_495),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_603),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_527),
.B(n_275),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_540),
.B(n_352),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_527),
.B(n_277),
.Y(n_656)
);

BUFx2_ASAP7_75t_L g657 ( 
.A(n_594),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_495),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_603),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_601),
.B(n_288),
.Y(n_660)
);

INVx2_ASAP7_75t_SL g661 ( 
.A(n_584),
.Y(n_661)
);

OAI22xp33_ASAP7_75t_L g662 ( 
.A1(n_594),
.A2(n_312),
.B1(n_201),
.B2(n_294),
.Y(n_662)
);

HB1xp67_ASAP7_75t_L g663 ( 
.A(n_626),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_601),
.B(n_311),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_539),
.B(n_188),
.Y(n_665)
);

OR2x2_ASAP7_75t_L g666 ( 
.A(n_595),
.B(n_377),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_505),
.B(n_188),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_508),
.B(n_584),
.Y(n_668)
);

BUFx5_ASAP7_75t_L g669 ( 
.A(n_564),
.Y(n_669)
);

NOR2xp67_ASAP7_75t_L g670 ( 
.A(n_568),
.B(n_481),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_617),
.B(n_329),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_617),
.B(n_334),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_631),
.B(n_455),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_631),
.B(n_455),
.Y(n_674)
);

AND2x4_ASAP7_75t_L g675 ( 
.A(n_547),
.B(n_481),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_499),
.B(n_462),
.Y(n_676)
);

INVx5_ASAP7_75t_L g677 ( 
.A(n_500),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_498),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_498),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_632),
.B(n_455),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_578),
.B(n_505),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_549),
.B(n_196),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_632),
.B(n_468),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_634),
.B(n_468),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_634),
.B(n_468),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_603),
.Y(n_686)
);

INVx2_ASAP7_75t_SL g687 ( 
.A(n_630),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_571),
.B(n_196),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_621),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_635),
.B(n_636),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_635),
.B(n_475),
.Y(n_691)
);

OAI22xp5_ASAP7_75t_L g692 ( 
.A1(n_543),
.A2(n_301),
.B1(n_332),
.B2(n_335),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_582),
.B(n_200),
.Y(n_693)
);

BUFx6f_ASAP7_75t_L g694 ( 
.A(n_503),
.Y(n_694)
);

NAND2xp33_ASAP7_75t_SL g695 ( 
.A(n_563),
.B(n_630),
.Y(n_695)
);

INVxp67_ASAP7_75t_L g696 ( 
.A(n_520),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_621),
.Y(n_697)
);

A2O1A1Ixp33_ASAP7_75t_L g698 ( 
.A1(n_502),
.A2(n_523),
.B(n_573),
.C(n_564),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_636),
.B(n_475),
.Y(n_699)
);

BUFx3_ASAP7_75t_L g700 ( 
.A(n_627),
.Y(n_700)
);

NAND2xp33_ASAP7_75t_L g701 ( 
.A(n_590),
.B(n_215),
.Y(n_701)
);

AOI22xp5_ASAP7_75t_L g702 ( 
.A1(n_543),
.A2(n_200),
.B1(n_321),
.B2(n_319),
.Y(n_702)
);

INVx8_ASAP7_75t_L g703 ( 
.A(n_543),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_498),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_640),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_542),
.B(n_485),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_542),
.Y(n_707)
);

NAND2x1_ASAP7_75t_L g708 ( 
.A(n_591),
.B(n_435),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_521),
.B(n_510),
.Y(n_709)
);

INVxp67_ASAP7_75t_SL g710 ( 
.A(n_554),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_510),
.B(n_253),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_622),
.B(n_253),
.Y(n_712)
);

BUFx2_ASAP7_75t_L g713 ( 
.A(n_627),
.Y(n_713)
);

O2A1O1Ixp33_ASAP7_75t_L g714 ( 
.A1(n_638),
.A2(n_492),
.B(n_491),
.C(n_488),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_504),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_597),
.B(n_299),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_555),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_552),
.B(n_605),
.Y(n_718)
);

NOR2x1p5_ASAP7_75t_L g719 ( 
.A(n_579),
.B(n_198),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_555),
.B(n_556),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_501),
.B(n_299),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_544),
.B(n_301),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_556),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_504),
.Y(n_724)
);

INVxp67_ASAP7_75t_L g725 ( 
.A(n_544),
.Y(n_725)
);

NAND2xp33_ASAP7_75t_L g726 ( 
.A(n_547),
.B(n_215),
.Y(n_726)
);

BUFx6f_ASAP7_75t_SL g727 ( 
.A(n_543),
.Y(n_727)
);

INVxp67_ASAP7_75t_L g728 ( 
.A(n_579),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_557),
.Y(n_729)
);

AOI22xp33_ASAP7_75t_L g730 ( 
.A1(n_535),
.A2(n_242),
.B1(n_333),
.B2(n_327),
.Y(n_730)
);

NOR2xp67_ASAP7_75t_L g731 ( 
.A(n_583),
.B(n_488),
.Y(n_731)
);

NOR2xp67_ASAP7_75t_L g732 ( 
.A(n_586),
.B(n_551),
.Y(n_732)
);

INVx4_ASAP7_75t_L g733 ( 
.A(n_500),
.Y(n_733)
);

AND2x4_ASAP7_75t_L g734 ( 
.A(n_551),
.B(n_491),
.Y(n_734)
);

AOI22xp33_ASAP7_75t_L g735 ( 
.A1(n_535),
.A2(n_242),
.B1(n_244),
.B2(n_317),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_557),
.B(n_492),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_558),
.B(n_493),
.Y(n_737)
);

NOR3xp33_ASAP7_75t_L g738 ( 
.A(n_638),
.B(n_619),
.C(n_609),
.Y(n_738)
);

CKINVDCx20_ASAP7_75t_R g739 ( 
.A(n_531),
.Y(n_739)
);

INVxp67_ASAP7_75t_L g740 ( 
.A(n_535),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_561),
.B(n_443),
.Y(n_741)
);

INVxp67_ASAP7_75t_L g742 ( 
.A(n_502),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_561),
.Y(n_743)
);

INVx2_ASAP7_75t_SL g744 ( 
.A(n_563),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_504),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_502),
.B(n_314),
.Y(n_746)
);

INVx1_ASAP7_75t_SL g747 ( 
.A(n_581),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_585),
.B(n_315),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_546),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_585),
.B(n_482),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_592),
.B(n_482),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_592),
.B(n_482),
.Y(n_752)
);

NOR2xp67_ASAP7_75t_L g753 ( 
.A(n_588),
.B(n_413),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_599),
.B(n_242),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_599),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_606),
.B(n_242),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_606),
.B(n_242),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_523),
.B(n_244),
.Y(n_758)
);

AOI22xp5_ASAP7_75t_L g759 ( 
.A1(n_543),
.A2(n_335),
.B1(n_332),
.B2(n_315),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_546),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_523),
.B(n_244),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_523),
.B(n_244),
.Y(n_762)
);

HB1xp67_ASAP7_75t_L g763 ( 
.A(n_608),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_602),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_602),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_604),
.Y(n_766)
);

INVx2_ASAP7_75t_SL g767 ( 
.A(n_620),
.Y(n_767)
);

AOI21xp5_ASAP7_75t_L g768 ( 
.A1(n_624),
.A2(n_244),
.B(n_325),
.Y(n_768)
);

INVxp67_ASAP7_75t_L g769 ( 
.A(n_608),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_588),
.B(n_319),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_629),
.B(n_591),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_604),
.B(n_317),
.Y(n_772)
);

INVx2_ASAP7_75t_SL g773 ( 
.A(n_620),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_629),
.B(n_321),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_607),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_546),
.Y(n_776)
);

INVxp67_ASAP7_75t_L g777 ( 
.A(n_608),
.Y(n_777)
);

INVx2_ASAP7_75t_SL g778 ( 
.A(n_553),
.Y(n_778)
);

AOI22xp5_ASAP7_75t_L g779 ( 
.A1(n_553),
.A2(n_330),
.B1(n_331),
.B2(n_327),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_607),
.B(n_317),
.Y(n_780)
);

BUFx5_ASAP7_75t_L g781 ( 
.A(n_496),
.Y(n_781)
);

NOR4xp25_ASAP7_75t_SL g782 ( 
.A(n_528),
.B(n_306),
.C(n_198),
.D(n_201),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_528),
.B(n_330),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_629),
.B(n_331),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_610),
.B(n_574),
.Y(n_785)
);

OAI22xp33_ASAP7_75t_L g786 ( 
.A1(n_553),
.A2(n_308),
.B1(n_306),
.B2(n_307),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_610),
.Y(n_787)
);

AOI22xp33_ASAP7_75t_L g788 ( 
.A1(n_613),
.A2(n_317),
.B1(n_325),
.B2(n_327),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_553),
.B(n_216),
.Y(n_789)
);

AOI22xp5_ASAP7_75t_L g790 ( 
.A1(n_553),
.A2(n_325),
.B1(n_327),
.B2(n_333),
.Y(n_790)
);

HB1xp67_ASAP7_75t_L g791 ( 
.A(n_608),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_608),
.B(n_413),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_574),
.Y(n_793)
);

INVxp33_ASAP7_75t_L g794 ( 
.A(n_614),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_548),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_496),
.B(n_507),
.Y(n_796)
);

OR2x6_ASAP7_75t_L g797 ( 
.A(n_500),
.B(n_417),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_591),
.B(n_172),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_507),
.B(n_325),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_L g800 ( 
.A(n_528),
.B(n_222),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_548),
.Y(n_801)
);

BUFx6f_ASAP7_75t_L g802 ( 
.A(n_694),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_643),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_668),
.B(n_417),
.Y(n_804)
);

BUFx2_ASAP7_75t_L g805 ( 
.A(n_739),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_710),
.B(n_613),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_755),
.Y(n_807)
);

AND2x4_ASAP7_75t_L g808 ( 
.A(n_661),
.B(n_402),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_645),
.B(n_591),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_681),
.A2(n_611),
.B(n_500),
.Y(n_810)
);

INVx2_ASAP7_75t_SL g811 ( 
.A(n_657),
.Y(n_811)
);

BUFx3_ASAP7_75t_L g812 ( 
.A(n_700),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_710),
.B(n_616),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_705),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_652),
.Y(n_815)
);

OAI22xp5_ASAP7_75t_SL g816 ( 
.A1(n_676),
.A2(n_655),
.B1(n_646),
.B2(n_747),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_647),
.B(n_616),
.Y(n_817)
);

NAND2x1p5_ASAP7_75t_L g818 ( 
.A(n_677),
.B(n_550),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_713),
.Y(n_819)
);

OAI22xp5_ASAP7_75t_SL g820 ( 
.A1(n_646),
.A2(n_712),
.B1(n_688),
.B2(n_687),
.Y(n_820)
);

INVx3_ASAP7_75t_SL g821 ( 
.A(n_767),
.Y(n_821)
);

AOI22xp33_ASAP7_75t_L g822 ( 
.A1(n_645),
.A2(n_738),
.B1(n_730),
.B2(n_735),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_647),
.B(n_515),
.Y(n_823)
);

CKINVDCx6p67_ASAP7_75t_R g824 ( 
.A(n_727),
.Y(n_824)
);

BUFx2_ASAP7_75t_L g825 ( 
.A(n_663),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_707),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_649),
.B(n_515),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_649),
.B(n_519),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_717),
.B(n_519),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_658),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_723),
.Y(n_831)
);

AOI22xp5_ASAP7_75t_L g832 ( 
.A1(n_738),
.A2(n_522),
.B1(n_533),
.B2(n_530),
.Y(n_832)
);

AND2x4_ASAP7_75t_L g833 ( 
.A(n_689),
.B(n_402),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_718),
.B(n_522),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_677),
.B(n_548),
.Y(n_835)
);

NAND3xp33_ASAP7_75t_SL g836 ( 
.A(n_711),
.B(n_296),
.C(n_294),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_729),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_743),
.B(n_533),
.Y(n_838)
);

BUFx3_ASAP7_75t_L g839 ( 
.A(n_773),
.Y(n_839)
);

AND2x4_ASAP7_75t_L g840 ( 
.A(n_697),
.B(n_404),
.Y(n_840)
);

OAI22xp5_ASAP7_75t_L g841 ( 
.A1(n_742),
.A2(n_560),
.B1(n_559),
.B2(n_633),
.Y(n_841)
);

NAND2x1p5_ASAP7_75t_L g842 ( 
.A(n_677),
.B(n_550),
.Y(n_842)
);

BUFx6f_ASAP7_75t_L g843 ( 
.A(n_694),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_696),
.B(n_559),
.Y(n_844)
);

AND2x4_ASAP7_75t_L g845 ( 
.A(n_696),
.B(n_404),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_764),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_725),
.B(n_560),
.Y(n_847)
);

HB1xp67_ASAP7_75t_L g848 ( 
.A(n_663),
.Y(n_848)
);

INVx2_ASAP7_75t_SL g849 ( 
.A(n_719),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_677),
.B(n_560),
.Y(n_850)
);

AOI22xp33_ASAP7_75t_L g851 ( 
.A1(n_730),
.A2(n_735),
.B1(n_667),
.B2(n_650),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_765),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_725),
.B(n_497),
.Y(n_853)
);

BUFx3_ASAP7_75t_L g854 ( 
.A(n_744),
.Y(n_854)
);

BUFx3_ASAP7_75t_L g855 ( 
.A(n_792),
.Y(n_855)
);

NAND3xp33_ASAP7_75t_SL g856 ( 
.A(n_711),
.B(n_303),
.C(n_296),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_678),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_766),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_794),
.B(n_229),
.Y(n_859)
);

CKINVDCx11_ASAP7_75t_R g860 ( 
.A(n_703),
.Y(n_860)
);

INVx3_ASAP7_75t_L g861 ( 
.A(n_675),
.Y(n_861)
);

INVx5_ASAP7_75t_L g862 ( 
.A(n_797),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_690),
.B(n_497),
.Y(n_863)
);

NOR3xp33_ASAP7_75t_SL g864 ( 
.A(n_662),
.B(n_307),
.C(n_298),
.Y(n_864)
);

BUFx6f_ASAP7_75t_L g865 ( 
.A(n_694),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_679),
.Y(n_866)
);

AOI22xp33_ASAP7_75t_L g867 ( 
.A1(n_667),
.A2(n_628),
.B1(n_625),
.B2(n_618),
.Y(n_867)
);

HB1xp67_ASAP7_75t_SL g868 ( 
.A(n_763),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_775),
.Y(n_869)
);

AND2x4_ASAP7_75t_L g870 ( 
.A(n_732),
.B(n_406),
.Y(n_870)
);

NAND3xp33_ASAP7_75t_SL g871 ( 
.A(n_782),
.B(n_712),
.C(n_702),
.Y(n_871)
);

INVx4_ASAP7_75t_L g872 ( 
.A(n_694),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_787),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_704),
.Y(n_874)
);

BUFx3_ASAP7_75t_L g875 ( 
.A(n_675),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_793),
.Y(n_876)
);

BUFx6f_ASAP7_75t_L g877 ( 
.A(n_797),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_720),
.B(n_497),
.Y(n_878)
);

BUFx6f_ASAP7_75t_L g879 ( 
.A(n_703),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_669),
.B(n_511),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_728),
.B(n_497),
.Y(n_881)
);

INVx3_ASAP7_75t_L g882 ( 
.A(n_734),
.Y(n_882)
);

BUFx6f_ASAP7_75t_L g883 ( 
.A(n_703),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_795),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_L g885 ( 
.A(n_666),
.B(n_249),
.Y(n_885)
);

INVx5_ASAP7_75t_L g886 ( 
.A(n_733),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_801),
.Y(n_887)
);

AOI22xp33_ASAP7_75t_L g888 ( 
.A1(n_740),
.A2(n_628),
.B1(n_625),
.B2(n_618),
.Y(n_888)
);

NAND2xp33_ASAP7_75t_SL g889 ( 
.A(n_727),
.B(n_298),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_669),
.B(n_511),
.Y(n_890)
);

INVx3_ASAP7_75t_L g891 ( 
.A(n_734),
.Y(n_891)
);

BUFx3_ASAP7_75t_L g892 ( 
.A(n_654),
.Y(n_892)
);

AOI22xp33_ASAP7_75t_L g893 ( 
.A1(n_740),
.A2(n_509),
.B1(n_506),
.B2(n_333),
.Y(n_893)
);

INVx2_ASAP7_75t_SL g894 ( 
.A(n_656),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_653),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_659),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_686),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_800),
.Y(n_898)
);

AOI211xp5_ASAP7_75t_L g899 ( 
.A1(n_662),
.A2(n_309),
.B(n_328),
.C(n_324),
.Y(n_899)
);

HB1xp67_ASAP7_75t_L g900 ( 
.A(n_763),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_715),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_724),
.Y(n_902)
);

BUFx3_ASAP7_75t_L g903 ( 
.A(n_800),
.Y(n_903)
);

NAND3xp33_ASAP7_75t_L g904 ( 
.A(n_728),
.B(n_278),
.C(n_258),
.Y(n_904)
);

HB1xp67_ASAP7_75t_L g905 ( 
.A(n_791),
.Y(n_905)
);

BUFx6f_ASAP7_75t_L g906 ( 
.A(n_778),
.Y(n_906)
);

INVx1_ASAP7_75t_SL g907 ( 
.A(n_722),
.Y(n_907)
);

OAI22xp5_ASAP7_75t_L g908 ( 
.A1(n_648),
.A2(n_562),
.B1(n_593),
.B2(n_513),
.Y(n_908)
);

NOR2xp33_ASAP7_75t_R g909 ( 
.A(n_695),
.B(n_562),
.Y(n_909)
);

NOR2xp67_ASAP7_75t_L g910 ( 
.A(n_783),
.B(n_593),
.Y(n_910)
);

AND2x2_ASAP7_75t_L g911 ( 
.A(n_670),
.B(n_418),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_737),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_706),
.B(n_517),
.Y(n_913)
);

INVx3_ASAP7_75t_L g914 ( 
.A(n_745),
.Y(n_914)
);

CKINVDCx20_ASAP7_75t_R g915 ( 
.A(n_693),
.Y(n_915)
);

BUFx4f_ASAP7_75t_L g916 ( 
.A(n_749),
.Y(n_916)
);

BUFx4f_ASAP7_75t_L g917 ( 
.A(n_760),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_SL g918 ( 
.A(n_669),
.B(n_513),
.Y(n_918)
);

AND2x4_ASAP7_75t_L g919 ( 
.A(n_731),
.B(n_409),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_692),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_L g921 ( 
.A(n_709),
.B(n_251),
.Y(n_921)
);

OAI21xp33_ASAP7_75t_SL g922 ( 
.A1(n_771),
.A2(n_420),
.B(n_409),
.Y(n_922)
);

AOI22xp5_ASAP7_75t_L g923 ( 
.A1(n_651),
.A2(n_777),
.B1(n_769),
.B2(n_789),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_736),
.B(n_748),
.Y(n_924)
);

AOI22xp33_ASAP7_75t_L g925 ( 
.A1(n_786),
.A2(n_509),
.B1(n_506),
.B2(n_333),
.Y(n_925)
);

AND2x6_ASAP7_75t_SL g926 ( 
.A(n_789),
.B(n_420),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_776),
.Y(n_927)
);

AOI221xp5_ASAP7_75t_SL g928 ( 
.A1(n_714),
.A2(n_410),
.B1(n_615),
.B2(n_639),
.C(n_641),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_741),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_748),
.B(n_517),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_673),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_674),
.Y(n_932)
);

AND2x4_ASAP7_75t_L g933 ( 
.A(n_791),
.B(n_410),
.Y(n_933)
);

OAI21xp5_ASAP7_75t_L g934 ( 
.A1(n_698),
.A2(n_538),
.B(n_537),
.Y(n_934)
);

AND2x4_ASAP7_75t_L g935 ( 
.A(n_769),
.B(n_576),
.Y(n_935)
);

INVxp67_ASAP7_75t_SL g936 ( 
.A(n_669),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_669),
.B(n_517),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_669),
.B(n_517),
.Y(n_938)
);

HB1xp67_ASAP7_75t_L g939 ( 
.A(n_777),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_671),
.B(n_526),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_680),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_L g942 ( 
.A(n_786),
.B(n_259),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_785),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_665),
.B(n_322),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_683),
.Y(n_945)
);

AOI22xp5_ASAP7_75t_L g946 ( 
.A1(n_660),
.A2(n_529),
.B1(n_514),
.B2(n_524),
.Y(n_946)
);

BUFx6f_ASAP7_75t_L g947 ( 
.A(n_708),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_SL g948 ( 
.A(n_781),
.B(n_514),
.Y(n_948)
);

AND2x4_ASAP7_75t_L g949 ( 
.A(n_753),
.B(n_770),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_796),
.Y(n_950)
);

AOI22xp5_ASAP7_75t_L g951 ( 
.A1(n_664),
.A2(n_529),
.B1(n_524),
.B2(n_525),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_672),
.B(n_526),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_684),
.Y(n_953)
);

BUFx4f_ASAP7_75t_L g954 ( 
.A(n_746),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_716),
.B(n_721),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_685),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_691),
.Y(n_957)
);

BUFx6f_ASAP7_75t_L g958 ( 
.A(n_642),
.Y(n_958)
);

HB1xp67_ASAP7_75t_L g959 ( 
.A(n_644),
.Y(n_959)
);

INVx4_ASAP7_75t_L g960 ( 
.A(n_733),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_781),
.B(n_526),
.Y(n_961)
);

BUFx3_ASAP7_75t_L g962 ( 
.A(n_699),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_SL g963 ( 
.A(n_781),
.B(n_525),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_758),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_682),
.B(n_270),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_781),
.Y(n_966)
);

AND2x4_ASAP7_75t_L g967 ( 
.A(n_759),
.B(n_576),
.Y(n_967)
);

OR2x6_ASAP7_75t_L g968 ( 
.A(n_798),
.B(n_500),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_781),
.B(n_526),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_781),
.Y(n_970)
);

INVx5_ASAP7_75t_L g971 ( 
.A(n_726),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_761),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_762),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_SL g974 ( 
.A(n_779),
.B(n_534),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_754),
.Y(n_975)
);

AOI22xp33_ASAP7_75t_L g976 ( 
.A1(n_788),
.A2(n_333),
.B1(n_327),
.B2(n_322),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_772),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_774),
.Y(n_978)
);

NAND3xp33_ASAP7_75t_SL g979 ( 
.A(n_790),
.B(n_309),
.C(n_324),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_750),
.B(n_536),
.Y(n_980)
);

BUFx8_ASAP7_75t_L g981 ( 
.A(n_701),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_780),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_924),
.B(n_784),
.Y(n_983)
);

O2A1O1Ixp33_ASAP7_75t_L g984 ( 
.A1(n_836),
.A2(n_757),
.B(n_756),
.C(n_799),
.Y(n_984)
);

AOI21x1_ASAP7_75t_L g985 ( 
.A1(n_910),
.A2(n_751),
.B(n_752),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_L g986 ( 
.A(n_816),
.B(n_273),
.Y(n_986)
);

AOI22xp33_ASAP7_75t_L g987 ( 
.A1(n_836),
.A2(n_227),
.B1(n_245),
.B2(n_788),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_814),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_886),
.A2(n_550),
.B(n_569),
.Y(n_989)
);

OAI22xp5_ASAP7_75t_L g990 ( 
.A1(n_822),
.A2(n_328),
.B1(n_320),
.B2(n_316),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_914),
.Y(n_991)
);

AO21x1_ASAP7_75t_L g992 ( 
.A1(n_834),
.A2(n_768),
.B(n_637),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_914),
.Y(n_993)
);

AOI221xp5_ASAP7_75t_L g994 ( 
.A1(n_942),
.A2(n_308),
.B1(n_316),
.B2(n_312),
.C(n_320),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_826),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_929),
.B(n_596),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_831),
.Y(n_997)
);

O2A1O1Ixp33_ASAP7_75t_L g998 ( 
.A1(n_856),
.A2(n_572),
.B(n_536),
.C(n_537),
.Y(n_998)
);

O2A1O1Ixp33_ASAP7_75t_L g999 ( 
.A1(n_856),
.A2(n_572),
.B(n_538),
.C(n_566),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_837),
.Y(n_1000)
);

AOI22xp5_ASAP7_75t_L g1001 ( 
.A1(n_820),
.A2(n_566),
.B1(n_577),
.B2(n_580),
.Y(n_1001)
);

O2A1O1Ixp33_ASAP7_75t_L g1002 ( 
.A1(n_942),
.A2(n_580),
.B(n_587),
.C(n_641),
.Y(n_1002)
);

BUFx6f_ASAP7_75t_L g1003 ( 
.A(n_879),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_807),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_861),
.B(n_227),
.Y(n_1005)
);

OAI22xp5_ASAP7_75t_L g1006 ( 
.A1(n_822),
.A2(n_303),
.B1(n_285),
.B2(n_337),
.Y(n_1006)
);

A2O1A1Ixp33_ASAP7_75t_L g1007 ( 
.A1(n_851),
.A2(n_587),
.B(n_639),
.C(n_641),
.Y(n_1007)
);

AND2x2_ASAP7_75t_L g1008 ( 
.A(n_885),
.B(n_227),
.Y(n_1008)
);

CKINVDCx16_ASAP7_75t_R g1009 ( 
.A(n_805),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_884),
.Y(n_1010)
);

AOI21x1_ASAP7_75t_L g1011 ( 
.A1(n_930),
.A2(n_637),
.B(n_639),
.Y(n_1011)
);

INVx3_ASAP7_75t_SL g1012 ( 
.A(n_819),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_887),
.Y(n_1013)
);

BUFx6f_ASAP7_75t_L g1014 ( 
.A(n_879),
.Y(n_1014)
);

AOI22xp5_ASAP7_75t_L g1015 ( 
.A1(n_871),
.A2(n_612),
.B1(n_541),
.B2(n_532),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_844),
.Y(n_1016)
);

BUFx3_ASAP7_75t_L g1017 ( 
.A(n_825),
.Y(n_1017)
);

OR2x6_ASAP7_75t_L g1018 ( 
.A(n_879),
.B(n_569),
.Y(n_1018)
);

AND2x2_ASAP7_75t_L g1019 ( 
.A(n_885),
.B(n_245),
.Y(n_1019)
);

O2A1O1Ixp33_ASAP7_75t_SL g1020 ( 
.A1(n_809),
.A2(n_871),
.B(n_974),
.C(n_890),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_847),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_SL g1022 ( 
.A(n_861),
.B(n_245),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_SL g1023 ( 
.A(n_882),
.B(n_503),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_936),
.A2(n_503),
.B(n_516),
.Y(n_1024)
);

NAND3xp33_ASAP7_75t_SL g1025 ( 
.A(n_898),
.B(n_596),
.C(n_598),
.Y(n_1025)
);

NOR2xp33_ASAP7_75t_L g1026 ( 
.A(n_903),
.B(n_575),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_803),
.Y(n_1027)
);

O2A1O1Ixp33_ASAP7_75t_L g1028 ( 
.A1(n_899),
.A2(n_600),
.B(n_598),
.C(n_596),
.Y(n_1028)
);

AOI22xp5_ASAP7_75t_SL g1029 ( 
.A1(n_920),
.A2(n_0),
.B1(n_2),
.B2(n_8),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_846),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_852),
.Y(n_1031)
);

BUFx2_ASAP7_75t_L g1032 ( 
.A(n_848),
.Y(n_1032)
);

NOR2xp33_ASAP7_75t_L g1033 ( 
.A(n_894),
.B(n_589),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_858),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_815),
.Y(n_1035)
);

NAND3xp33_ASAP7_75t_L g1036 ( 
.A(n_921),
.B(n_600),
.C(n_598),
.Y(n_1036)
);

OAI22xp5_ASAP7_75t_L g1037 ( 
.A1(n_851),
.A2(n_600),
.B1(n_612),
.B2(n_589),
.Y(n_1037)
);

CKINVDCx20_ASAP7_75t_R g1038 ( 
.A(n_860),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_818),
.A2(n_503),
.B(n_516),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_SL g1040 ( 
.A(n_882),
.B(n_891),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_869),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_818),
.A2(n_503),
.B(n_516),
.Y(n_1042)
);

NOR2xp67_ASAP7_75t_L g1043 ( 
.A(n_904),
.B(n_66),
.Y(n_1043)
);

AND2x2_ASAP7_75t_SL g1044 ( 
.A(n_976),
.B(n_0),
.Y(n_1044)
);

BUFx6f_ASAP7_75t_L g1045 ( 
.A(n_879),
.Y(n_1045)
);

AND2x4_ASAP7_75t_L g1046 ( 
.A(n_855),
.B(n_612),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_L g1047 ( 
.A(n_848),
.B(n_575),
.Y(n_1047)
);

NOR2xp33_ASAP7_75t_L g1048 ( 
.A(n_892),
.B(n_575),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_842),
.A2(n_516),
.B(n_545),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_L g1050 ( 
.A(n_859),
.B(n_541),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_842),
.A2(n_545),
.B(n_532),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_961),
.A2(n_545),
.B(n_532),
.Y(n_1052)
);

BUFx2_ASAP7_75t_L g1053 ( 
.A(n_811),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_969),
.A2(n_545),
.B(n_532),
.Y(n_1054)
);

AND2x4_ASAP7_75t_L g1055 ( 
.A(n_875),
.B(n_162),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_830),
.Y(n_1056)
);

BUFx2_ASAP7_75t_L g1057 ( 
.A(n_900),
.Y(n_1057)
);

NAND2x2_ASAP7_75t_L g1058 ( 
.A(n_812),
.B(n_8),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_950),
.B(n_9),
.Y(n_1059)
);

O2A1O1Ixp33_ASAP7_75t_L g1060 ( 
.A1(n_921),
.A2(n_10),
.B(n_11),
.C(n_12),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_857),
.Y(n_1061)
);

BUFx6f_ASAP7_75t_L g1062 ( 
.A(n_883),
.Y(n_1062)
);

OR2x6_ASAP7_75t_L g1063 ( 
.A(n_883),
.B(n_56),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_912),
.B(n_15),
.Y(n_1064)
);

OAI22xp5_ASAP7_75t_L g1065 ( 
.A1(n_893),
.A2(n_17),
.B1(n_19),
.B2(n_22),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_937),
.A2(n_65),
.B(n_151),
.Y(n_1066)
);

INVx3_ASAP7_75t_L g1067 ( 
.A(n_802),
.Y(n_1067)
);

O2A1O1Ixp33_ASAP7_75t_L g1068 ( 
.A1(n_965),
.A2(n_17),
.B(n_19),
.C(n_23),
.Y(n_1068)
);

OAI22x1_ASAP7_75t_L g1069 ( 
.A1(n_923),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_1069)
);

INVx4_ASAP7_75t_L g1070 ( 
.A(n_883),
.Y(n_1070)
);

OA22x2_ASAP7_75t_L g1071 ( 
.A1(n_907),
.A2(n_31),
.B1(n_33),
.B2(n_36),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_931),
.B(n_38),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_938),
.A2(n_102),
.B(n_148),
.Y(n_1073)
);

A2O1A1Ixp33_ASAP7_75t_SL g1074 ( 
.A1(n_965),
.A2(n_90),
.B(n_147),
.C(n_142),
.Y(n_1074)
);

NAND3xp33_ASAP7_75t_L g1075 ( 
.A(n_864),
.B(n_41),
.C(n_42),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_810),
.A2(n_83),
.B(n_139),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_932),
.B(n_44),
.Y(n_1077)
);

INVx4_ASAP7_75t_L g1078 ( 
.A(n_802),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_866),
.Y(n_1079)
);

INVx3_ASAP7_75t_SL g1080 ( 
.A(n_824),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_810),
.A2(n_106),
.B(n_136),
.Y(n_1081)
);

AND2x4_ASAP7_75t_L g1082 ( 
.A(n_849),
.B(n_72),
.Y(n_1082)
);

OAI22xp5_ASAP7_75t_L g1083 ( 
.A1(n_893),
.A2(n_47),
.B1(n_50),
.B2(n_51),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_873),
.Y(n_1084)
);

OAI22xp5_ASAP7_75t_L g1085 ( 
.A1(n_976),
.A2(n_54),
.B1(n_68),
.B2(n_112),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_941),
.B(n_54),
.Y(n_1086)
);

AOI33xp33_ASAP7_75t_L g1087 ( 
.A1(n_804),
.A2(n_126),
.A3(n_133),
.B1(n_134),
.B2(n_161),
.B3(n_833),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_806),
.A2(n_813),
.B(n_971),
.Y(n_1088)
);

AND2x2_ASAP7_75t_L g1089 ( 
.A(n_859),
.B(n_845),
.Y(n_1089)
);

INVxp67_ASAP7_75t_SL g1090 ( 
.A(n_802),
.Y(n_1090)
);

AOI21x1_ASAP7_75t_L g1091 ( 
.A1(n_908),
.A2(n_890),
.B(n_880),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_874),
.Y(n_1092)
);

NAND2xp33_ASAP7_75t_SL g1093 ( 
.A(n_978),
.B(n_915),
.Y(n_1093)
);

O2A1O1Ixp33_ASAP7_75t_L g1094 ( 
.A1(n_864),
.A2(n_939),
.B(n_922),
.C(n_959),
.Y(n_1094)
);

NOR2xp33_ASAP7_75t_L g1095 ( 
.A(n_900),
.B(n_905),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_945),
.B(n_953),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_956),
.B(n_957),
.Y(n_1097)
);

OAI21xp33_ASAP7_75t_L g1098 ( 
.A1(n_845),
.A2(n_833),
.B(n_840),
.Y(n_1098)
);

BUFx6f_ASAP7_75t_L g1099 ( 
.A(n_802),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_971),
.A2(n_863),
.B(n_878),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_SL g1101 ( 
.A(n_954),
.B(n_955),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_876),
.Y(n_1102)
);

AOI22xp33_ASAP7_75t_L g1103 ( 
.A1(n_967),
.A2(n_979),
.B1(n_962),
.B2(n_935),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_959),
.B(n_943),
.Y(n_1104)
);

AOI22xp5_ASAP7_75t_L g1105 ( 
.A1(n_911),
.A2(n_870),
.B1(n_919),
.B2(n_967),
.Y(n_1105)
);

CKINVDCx8_ASAP7_75t_R g1106 ( 
.A(n_926),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_817),
.B(n_823),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_901),
.Y(n_1108)
);

OAI22xp5_ASAP7_75t_SL g1109 ( 
.A1(n_925),
.A2(n_821),
.B1(n_854),
.B2(n_839),
.Y(n_1109)
);

INVx5_ASAP7_75t_L g1110 ( 
.A(n_843),
.Y(n_1110)
);

INVxp67_ASAP7_75t_SL g1111 ( 
.A(n_843),
.Y(n_1111)
);

AO21x1_ASAP7_75t_L g1112 ( 
.A1(n_974),
.A2(n_832),
.B(n_973),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_895),
.Y(n_1113)
);

NOR2xp33_ASAP7_75t_L g1114 ( 
.A(n_868),
.B(n_944),
.Y(n_1114)
);

BUFx3_ASAP7_75t_L g1115 ( 
.A(n_821),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_971),
.A2(n_960),
.B(n_850),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_902),
.Y(n_1117)
);

INVx2_ASAP7_75t_SL g1118 ( 
.A(n_933),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_896),
.Y(n_1119)
);

OAI22xp5_ASAP7_75t_L g1120 ( 
.A1(n_925),
.A2(n_868),
.B1(n_867),
.B2(n_888),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_897),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_881),
.B(n_808),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_808),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_853),
.Y(n_1124)
);

OR2x2_ASAP7_75t_L g1125 ( 
.A(n_1104),
.B(n_1009),
.Y(n_1125)
);

AOI21xp33_ASAP7_75t_L g1126 ( 
.A1(n_1008),
.A2(n_827),
.B(n_828),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_988),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_1096),
.B(n_840),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_995),
.Y(n_1129)
);

OAI22xp5_ASAP7_75t_L g1130 ( 
.A1(n_1120),
.A2(n_1097),
.B1(n_1107),
.B2(n_1103),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_1012),
.Y(n_1131)
);

A2O1A1Ixp33_ASAP7_75t_L g1132 ( 
.A1(n_986),
.A2(n_949),
.B(n_964),
.C(n_917),
.Y(n_1132)
);

OAI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_983),
.A2(n_934),
.B(n_980),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_SL g1134 ( 
.A(n_1089),
.B(n_949),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1016),
.B(n_933),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_997),
.Y(n_1136)
);

AO31x2_ASAP7_75t_L g1137 ( 
.A1(n_1112),
.A2(n_975),
.A3(n_841),
.B(n_972),
.Y(n_1137)
);

BUFx2_ASAP7_75t_SL g1138 ( 
.A(n_1115),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1021),
.B(n_958),
.Y(n_1139)
);

OAI21x1_ASAP7_75t_SL g1140 ( 
.A1(n_1094),
.A2(n_829),
.B(n_838),
.Y(n_1140)
);

AOI211x1_ASAP7_75t_L g1141 ( 
.A1(n_1065),
.A2(n_979),
.B(n_913),
.C(n_927),
.Y(n_1141)
);

OAI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_1122),
.A2(n_980),
.B(n_940),
.Y(n_1142)
);

OAI21x1_ASAP7_75t_L g1143 ( 
.A1(n_1052),
.A2(n_1054),
.B(n_1011),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_1019),
.B(n_958),
.Y(n_1144)
);

NOR2xp33_ASAP7_75t_L g1145 ( 
.A(n_1114),
.B(n_906),
.Y(n_1145)
);

INVxp67_ASAP7_75t_L g1146 ( 
.A(n_1032),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_1124),
.B(n_958),
.Y(n_1147)
);

AO31x2_ASAP7_75t_L g1148 ( 
.A1(n_992),
.A2(n_982),
.A3(n_977),
.B(n_952),
.Y(n_1148)
);

AOI21x1_ASAP7_75t_SL g1149 ( 
.A1(n_1064),
.A2(n_935),
.B(n_928),
.Y(n_1149)
);

OAI22xp5_ASAP7_75t_SL g1150 ( 
.A1(n_1106),
.A2(n_877),
.B1(n_906),
.B2(n_862),
.Y(n_1150)
);

A2O1A1Ixp33_ASAP7_75t_L g1151 ( 
.A1(n_1098),
.A2(n_916),
.B(n_889),
.C(n_951),
.Y(n_1151)
);

OAI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_1020),
.A2(n_946),
.B(n_867),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_1088),
.A2(n_968),
.B(n_835),
.Y(n_1153)
);

AO31x2_ASAP7_75t_L g1154 ( 
.A1(n_1007),
.A2(n_970),
.A3(n_966),
.B(n_872),
.Y(n_1154)
);

BUFx6f_ASAP7_75t_L g1155 ( 
.A(n_1003),
.Y(n_1155)
);

OAI21x1_ASAP7_75t_L g1156 ( 
.A1(n_985),
.A2(n_918),
.B(n_880),
.Y(n_1156)
);

OAI21x1_ASAP7_75t_L g1157 ( 
.A1(n_1039),
.A2(n_918),
.B(n_948),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1000),
.Y(n_1158)
);

A2O1A1Ixp33_ASAP7_75t_L g1159 ( 
.A1(n_1098),
.A2(n_916),
.B(n_958),
.C(n_906),
.Y(n_1159)
);

OAI21x1_ASAP7_75t_L g1160 ( 
.A1(n_1042),
.A2(n_963),
.B(n_948),
.Y(n_1160)
);

AND2x2_ASAP7_75t_L g1161 ( 
.A(n_1123),
.B(n_906),
.Y(n_1161)
);

BUFx2_ASAP7_75t_L g1162 ( 
.A(n_1017),
.Y(n_1162)
);

NOR2xp67_ASAP7_75t_L g1163 ( 
.A(n_1105),
.B(n_862),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1100),
.A2(n_968),
.B(n_963),
.Y(n_1164)
);

A2O1A1Ixp33_ASAP7_75t_L g1165 ( 
.A1(n_1050),
.A2(n_877),
.B(n_888),
.C(n_947),
.Y(n_1165)
);

INVxp67_ASAP7_75t_L g1166 ( 
.A(n_1057),
.Y(n_1166)
);

OAI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_1036),
.A2(n_909),
.B(n_947),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1101),
.B(n_877),
.Y(n_1168)
);

NAND2x1_ASAP7_75t_L g1169 ( 
.A(n_1018),
.B(n_843),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1004),
.B(n_877),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_1013),
.Y(n_1171)
);

INVx3_ASAP7_75t_L g1172 ( 
.A(n_1018),
.Y(n_1172)
);

OA21x2_ASAP7_75t_L g1173 ( 
.A1(n_1036),
.A2(n_865),
.B(n_981),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1072),
.B(n_865),
.Y(n_1174)
);

OAI21xp33_ASAP7_75t_SL g1175 ( 
.A1(n_1044),
.A2(n_981),
.B(n_1065),
.Y(n_1175)
);

INVx2_ASAP7_75t_SL g1176 ( 
.A(n_1053),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1010),
.Y(n_1177)
);

NOR4xp25_ASAP7_75t_L g1178 ( 
.A(n_1068),
.B(n_1060),
.C(n_1075),
.D(n_1083),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1030),
.Y(n_1179)
);

BUFx6f_ASAP7_75t_L g1180 ( 
.A(n_1003),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_1038),
.Y(n_1181)
);

AOI21x1_ASAP7_75t_L g1182 ( 
.A1(n_1037),
.A2(n_1049),
.B(n_1081),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_1080),
.Y(n_1183)
);

INVx4_ASAP7_75t_L g1184 ( 
.A(n_1110),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1031),
.Y(n_1185)
);

OAI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_998),
.A2(n_999),
.B(n_1028),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1034),
.Y(n_1187)
);

AOI22xp5_ASAP7_75t_L g1188 ( 
.A1(n_1069),
.A2(n_1109),
.B1(n_1083),
.B2(n_1075),
.Y(n_1188)
);

OAI21x1_ASAP7_75t_L g1189 ( 
.A1(n_1051),
.A2(n_1024),
.B(n_1116),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1077),
.B(n_1086),
.Y(n_1190)
);

AOI21x1_ASAP7_75t_L g1191 ( 
.A1(n_1076),
.A2(n_1023),
.B(n_996),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_989),
.A2(n_984),
.B(n_996),
.Y(n_1192)
);

OR2x6_ASAP7_75t_L g1193 ( 
.A(n_1063),
.B(n_1003),
.Y(n_1193)
);

AOI221xp5_ASAP7_75t_L g1194 ( 
.A1(n_994),
.A2(n_1006),
.B1(n_990),
.B2(n_987),
.C(n_1085),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_1093),
.Y(n_1195)
);

INVx1_ASAP7_75t_SL g1196 ( 
.A(n_1095),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_1113),
.Y(n_1197)
);

OAI21x1_ASAP7_75t_L g1198 ( 
.A1(n_1002),
.A2(n_1015),
.B(n_1001),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1041),
.Y(n_1199)
);

AO31x2_ASAP7_75t_L g1200 ( 
.A1(n_1085),
.A2(n_1059),
.A3(n_1066),
.B(n_1073),
.Y(n_1200)
);

AO31x2_ASAP7_75t_L g1201 ( 
.A1(n_1006),
.A2(n_1033),
.A3(n_990),
.B(n_1047),
.Y(n_1201)
);

AO31x2_ASAP7_75t_L g1202 ( 
.A1(n_1084),
.A2(n_1102),
.A3(n_1048),
.B(n_1121),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1018),
.A2(n_1025),
.B(n_1111),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_SL g1204 ( 
.A(n_1118),
.B(n_1109),
.Y(n_1204)
);

NOR2xp67_ASAP7_75t_L g1205 ( 
.A(n_1070),
.B(n_1078),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1119),
.Y(n_1206)
);

AND2x2_ASAP7_75t_L g1207 ( 
.A(n_1055),
.B(n_1071),
.Y(n_1207)
);

INVx4_ASAP7_75t_L g1208 ( 
.A(n_1014),
.Y(n_1208)
);

AND2x6_ASAP7_75t_L g1209 ( 
.A(n_1014),
.B(n_1045),
.Y(n_1209)
);

AO31x2_ASAP7_75t_L g1210 ( 
.A1(n_991),
.A2(n_993),
.A3(n_1061),
.B(n_1117),
.Y(n_1210)
);

AOI22xp33_ASAP7_75t_L g1211 ( 
.A1(n_1040),
.A2(n_1055),
.B1(n_1022),
.B2(n_1005),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1026),
.B(n_1046),
.Y(n_1212)
);

AOI22xp5_ASAP7_75t_L g1213 ( 
.A1(n_1082),
.A2(n_1063),
.B1(n_1043),
.B2(n_1092),
.Y(n_1213)
);

A2O1A1Ixp33_ASAP7_75t_L g1214 ( 
.A1(n_1087),
.A2(n_1029),
.B(n_1027),
.C(n_1108),
.Y(n_1214)
);

AND2x4_ASAP7_75t_L g1215 ( 
.A(n_1046),
.B(n_1070),
.Y(n_1215)
);

OAI22xp5_ASAP7_75t_L g1216 ( 
.A1(n_1090),
.A2(n_1079),
.B1(n_1035),
.B2(n_1056),
.Y(n_1216)
);

INVxp67_ASAP7_75t_L g1217 ( 
.A(n_1029),
.Y(n_1217)
);

AO31x2_ASAP7_75t_L g1218 ( 
.A1(n_1078),
.A2(n_1074),
.A3(n_1067),
.B(n_1058),
.Y(n_1218)
);

AND2x2_ASAP7_75t_SL g1219 ( 
.A(n_1014),
.B(n_1045),
.Y(n_1219)
);

AO31x2_ASAP7_75t_L g1220 ( 
.A1(n_1062),
.A2(n_1112),
.A3(n_992),
.B(n_1007),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_988),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_988),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1088),
.A2(n_886),
.B(n_677),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1096),
.B(n_1097),
.Y(n_1224)
);

OAI21x1_ASAP7_75t_L g1225 ( 
.A1(n_1052),
.A2(n_934),
.B(n_1054),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1088),
.A2(n_886),
.B(n_677),
.Y(n_1226)
);

OAI22xp5_ASAP7_75t_L g1227 ( 
.A1(n_1120),
.A2(n_822),
.B1(n_851),
.B2(n_645),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_L g1228 ( 
.A1(n_1052),
.A2(n_934),
.B(n_1054),
.Y(n_1228)
);

AOI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1011),
.A2(n_1091),
.B(n_1100),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_1012),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1096),
.B(n_1097),
.Y(n_1231)
);

NOR2xp33_ASAP7_75t_L g1232 ( 
.A(n_1089),
.B(n_338),
.Y(n_1232)
);

INVx5_ASAP7_75t_L g1233 ( 
.A(n_1099),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1096),
.B(n_1097),
.Y(n_1234)
);

NAND2x1p5_ASAP7_75t_L g1235 ( 
.A(n_1070),
.B(n_1110),
.Y(n_1235)
);

AO31x2_ASAP7_75t_L g1236 ( 
.A1(n_1112),
.A2(n_992),
.A3(n_1007),
.B(n_908),
.Y(n_1236)
);

OAI21x1_ASAP7_75t_L g1237 ( 
.A1(n_1052),
.A2(n_934),
.B(n_1054),
.Y(n_1237)
);

AND2x2_ASAP7_75t_L g1238 ( 
.A(n_1089),
.B(n_668),
.Y(n_1238)
);

INVx1_ASAP7_75t_SL g1239 ( 
.A(n_1017),
.Y(n_1239)
);

INVx2_ASAP7_75t_SL g1240 ( 
.A(n_1115),
.Y(n_1240)
);

AO31x2_ASAP7_75t_L g1241 ( 
.A1(n_1112),
.A2(n_992),
.A3(n_1007),
.B(n_908),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_SL g1242 ( 
.A(n_1089),
.B(n_898),
.Y(n_1242)
);

INVx3_ASAP7_75t_SL g1243 ( 
.A(n_1012),
.Y(n_1243)
);

AOI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1088),
.A2(n_886),
.B(n_677),
.Y(n_1244)
);

O2A1O1Ixp5_ASAP7_75t_L g1245 ( 
.A1(n_1112),
.A2(n_1019),
.B(n_1008),
.C(n_1005),
.Y(n_1245)
);

OAI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_983),
.A2(n_851),
.B(n_740),
.Y(n_1246)
);

NOR4xp25_ASAP7_75t_L g1247 ( 
.A(n_1068),
.B(n_1060),
.C(n_856),
.D(n_836),
.Y(n_1247)
);

OAI22xp5_ASAP7_75t_L g1248 ( 
.A1(n_1120),
.A2(n_822),
.B1(n_851),
.B2(n_645),
.Y(n_1248)
);

CKINVDCx8_ASAP7_75t_R g1249 ( 
.A(n_1009),
.Y(n_1249)
);

AOI221x1_ASAP7_75t_L g1250 ( 
.A1(n_1120),
.A2(n_1083),
.B1(n_1065),
.B2(n_986),
.C(n_1069),
.Y(n_1250)
);

OAI22x1_ASAP7_75t_L g1251 ( 
.A1(n_986),
.A2(n_942),
.B1(n_920),
.B2(n_1114),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1096),
.B(n_1097),
.Y(n_1252)
);

NOR2xp33_ASAP7_75t_L g1253 ( 
.A(n_1089),
.B(n_338),
.Y(n_1253)
);

INVx2_ASAP7_75t_L g1254 ( 
.A(n_1013),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_988),
.Y(n_1255)
);

AOI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_1088),
.A2(n_886),
.B(n_677),
.Y(n_1256)
);

OAI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_983),
.A2(n_851),
.B(n_740),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1096),
.B(n_1097),
.Y(n_1258)
);

AOI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1088),
.A2(n_886),
.B(n_677),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1013),
.Y(n_1260)
);

AOI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_1088),
.A2(n_886),
.B(n_677),
.Y(n_1261)
);

OAI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1052),
.A2(n_934),
.B(n_1054),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_988),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1096),
.B(n_1097),
.Y(n_1264)
);

A2O1A1Ixp33_ASAP7_75t_L g1265 ( 
.A1(n_986),
.A2(n_822),
.B(n_851),
.C(n_688),
.Y(n_1265)
);

OAI21x1_ASAP7_75t_L g1266 ( 
.A1(n_1052),
.A2(n_934),
.B(n_1054),
.Y(n_1266)
);

AO31x2_ASAP7_75t_L g1267 ( 
.A1(n_1112),
.A2(n_992),
.A3(n_1007),
.B(n_908),
.Y(n_1267)
);

INVx2_ASAP7_75t_L g1268 ( 
.A(n_1197),
.Y(n_1268)
);

OAI22xp5_ASAP7_75t_L g1269 ( 
.A1(n_1265),
.A2(n_1234),
.B1(n_1264),
.B2(n_1258),
.Y(n_1269)
);

OR2x2_ASAP7_75t_L g1270 ( 
.A(n_1125),
.B(n_1196),
.Y(n_1270)
);

OAI21x1_ASAP7_75t_L g1271 ( 
.A1(n_1143),
.A2(n_1189),
.B(n_1229),
.Y(n_1271)
);

NAND2x1p5_ASAP7_75t_L g1272 ( 
.A(n_1172),
.B(n_1169),
.Y(n_1272)
);

BUFx3_ASAP7_75t_L g1273 ( 
.A(n_1162),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1224),
.B(n_1231),
.Y(n_1274)
);

OA21x2_ASAP7_75t_L g1275 ( 
.A1(n_1186),
.A2(n_1192),
.B(n_1198),
.Y(n_1275)
);

OAI22xp33_ASAP7_75t_L g1276 ( 
.A1(n_1227),
.A2(n_1248),
.B1(n_1250),
.B2(n_1188),
.Y(n_1276)
);

INVx2_ASAP7_75t_SL g1277 ( 
.A(n_1176),
.Y(n_1277)
);

INVx1_ASAP7_75t_SL g1278 ( 
.A(n_1239),
.Y(n_1278)
);

BUFx2_ASAP7_75t_SL g1279 ( 
.A(n_1249),
.Y(n_1279)
);

AO21x2_ASAP7_75t_L g1280 ( 
.A1(n_1164),
.A2(n_1153),
.B(n_1140),
.Y(n_1280)
);

OA21x2_ASAP7_75t_L g1281 ( 
.A1(n_1225),
.A2(n_1237),
.B(n_1228),
.Y(n_1281)
);

CKINVDCx6p67_ASAP7_75t_R g1282 ( 
.A(n_1243),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1252),
.B(n_1238),
.Y(n_1283)
);

NOR2xp67_ASAP7_75t_L g1284 ( 
.A(n_1146),
.B(n_1166),
.Y(n_1284)
);

OAI21x1_ASAP7_75t_L g1285 ( 
.A1(n_1262),
.A2(n_1266),
.B(n_1160),
.Y(n_1285)
);

OAI21x1_ASAP7_75t_L g1286 ( 
.A1(n_1157),
.A2(n_1226),
.B(n_1223),
.Y(n_1286)
);

AOI21xp33_ASAP7_75t_L g1287 ( 
.A1(n_1194),
.A2(n_1190),
.B(n_1251),
.Y(n_1287)
);

NAND2x1p5_ASAP7_75t_L g1288 ( 
.A(n_1172),
.B(n_1184),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_1127),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_1129),
.Y(n_1290)
);

AOI22xp33_ASAP7_75t_L g1291 ( 
.A1(n_1217),
.A2(n_1188),
.B1(n_1175),
.B2(n_1130),
.Y(n_1291)
);

OAI21x1_ASAP7_75t_L g1292 ( 
.A1(n_1244),
.A2(n_1259),
.B(n_1261),
.Y(n_1292)
);

OA21x2_ASAP7_75t_L g1293 ( 
.A1(n_1152),
.A2(n_1182),
.B(n_1133),
.Y(n_1293)
);

INVx2_ASAP7_75t_SL g1294 ( 
.A(n_1240),
.Y(n_1294)
);

AO31x2_ASAP7_75t_L g1295 ( 
.A1(n_1165),
.A2(n_1132),
.A3(n_1214),
.B(n_1256),
.Y(n_1295)
);

INVx4_ASAP7_75t_L g1296 ( 
.A(n_1233),
.Y(n_1296)
);

CKINVDCx11_ASAP7_75t_R g1297 ( 
.A(n_1193),
.Y(n_1297)
);

CKINVDCx16_ASAP7_75t_R g1298 ( 
.A(n_1138),
.Y(n_1298)
);

INVx5_ASAP7_75t_L g1299 ( 
.A(n_1209),
.Y(n_1299)
);

OAI21x1_ASAP7_75t_L g1300 ( 
.A1(n_1191),
.A2(n_1156),
.B(n_1149),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_1181),
.Y(n_1301)
);

AOI22xp5_ASAP7_75t_L g1302 ( 
.A1(n_1232),
.A2(n_1253),
.B1(n_1134),
.B2(n_1242),
.Y(n_1302)
);

AND2x4_ASAP7_75t_L g1303 ( 
.A(n_1163),
.B(n_1215),
.Y(n_1303)
);

INVx4_ASAP7_75t_L g1304 ( 
.A(n_1233),
.Y(n_1304)
);

NOR2xp33_ASAP7_75t_L g1305 ( 
.A(n_1128),
.B(n_1175),
.Y(n_1305)
);

OAI21x1_ASAP7_75t_L g1306 ( 
.A1(n_1203),
.A2(n_1167),
.B(n_1142),
.Y(n_1306)
);

INVxp67_ASAP7_75t_L g1307 ( 
.A(n_1145),
.Y(n_1307)
);

OAI22xp5_ASAP7_75t_L g1308 ( 
.A1(n_1213),
.A2(n_1211),
.B1(n_1204),
.B2(n_1193),
.Y(n_1308)
);

AOI22xp5_ASAP7_75t_L g1309 ( 
.A1(n_1213),
.A2(n_1163),
.B1(n_1195),
.B2(n_1207),
.Y(n_1309)
);

AO31x2_ASAP7_75t_L g1310 ( 
.A1(n_1159),
.A2(n_1151),
.A3(n_1216),
.B(n_1174),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1136),
.Y(n_1311)
);

NOR2xp33_ASAP7_75t_L g1312 ( 
.A(n_1135),
.B(n_1126),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1144),
.B(n_1139),
.Y(n_1313)
);

OAI21xp5_ASAP7_75t_L g1314 ( 
.A1(n_1245),
.A2(n_1247),
.B(n_1178),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1158),
.Y(n_1315)
);

OAI21x1_ASAP7_75t_L g1316 ( 
.A1(n_1246),
.A2(n_1257),
.B(n_1147),
.Y(n_1316)
);

AND2x4_ASAP7_75t_SL g1317 ( 
.A(n_1208),
.B(n_1180),
.Y(n_1317)
);

OAI21x1_ASAP7_75t_L g1318 ( 
.A1(n_1173),
.A2(n_1168),
.B(n_1170),
.Y(n_1318)
);

INVx1_ASAP7_75t_SL g1319 ( 
.A(n_1131),
.Y(n_1319)
);

INVx2_ASAP7_75t_SL g1320 ( 
.A(n_1230),
.Y(n_1320)
);

INVx1_ASAP7_75t_SL g1321 ( 
.A(n_1212),
.Y(n_1321)
);

BUFx3_ASAP7_75t_L g1322 ( 
.A(n_1219),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_1177),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_L g1324 ( 
.A1(n_1171),
.A2(n_1254),
.B1(n_1260),
.B2(n_1199),
.Y(n_1324)
);

OR2x6_ASAP7_75t_L g1325 ( 
.A(n_1150),
.B(n_1141),
.Y(n_1325)
);

NOR2xp67_ASAP7_75t_L g1326 ( 
.A(n_1208),
.B(n_1183),
.Y(n_1326)
);

OAI21x1_ASAP7_75t_L g1327 ( 
.A1(n_1173),
.A2(n_1206),
.B(n_1263),
.Y(n_1327)
);

AOI21xp33_ASAP7_75t_SL g1328 ( 
.A1(n_1179),
.A2(n_1222),
.B(n_1187),
.Y(n_1328)
);

OAI21x1_ASAP7_75t_L g1329 ( 
.A1(n_1185),
.A2(n_1255),
.B(n_1221),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1161),
.B(n_1201),
.Y(n_1330)
);

OR2x6_ASAP7_75t_L g1331 ( 
.A(n_1141),
.B(n_1235),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1210),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1210),
.Y(n_1333)
);

OAI21x1_ASAP7_75t_L g1334 ( 
.A1(n_1205),
.A2(n_1154),
.B(n_1220),
.Y(n_1334)
);

OAI21x1_ASAP7_75t_L g1335 ( 
.A1(n_1154),
.A2(n_1220),
.B(n_1241),
.Y(n_1335)
);

NOR2xp33_ASAP7_75t_L g1336 ( 
.A(n_1155),
.B(n_1180),
.Y(n_1336)
);

OAI21x1_ASAP7_75t_L g1337 ( 
.A1(n_1154),
.A2(n_1220),
.B(n_1241),
.Y(n_1337)
);

INVx1_ASAP7_75t_SL g1338 ( 
.A(n_1209),
.Y(n_1338)
);

AND2x4_ASAP7_75t_L g1339 ( 
.A(n_1218),
.B(n_1202),
.Y(n_1339)
);

AO21x2_ASAP7_75t_L g1340 ( 
.A1(n_1137),
.A2(n_1267),
.B(n_1241),
.Y(n_1340)
);

AO31x2_ASAP7_75t_L g1341 ( 
.A1(n_1236),
.A2(n_1267),
.A3(n_1137),
.B(n_1148),
.Y(n_1341)
);

OAI21xp5_ASAP7_75t_L g1342 ( 
.A1(n_1209),
.A2(n_1200),
.B(n_1201),
.Y(n_1342)
);

OAI21xp5_ASAP7_75t_L g1343 ( 
.A1(n_1200),
.A2(n_1202),
.B(n_1137),
.Y(n_1343)
);

A2O1A1Ixp33_ASAP7_75t_L g1344 ( 
.A1(n_1200),
.A2(n_1265),
.B(n_822),
.C(n_1248),
.Y(n_1344)
);

A2O1A1Ixp33_ASAP7_75t_L g1345 ( 
.A1(n_1265),
.A2(n_822),
.B(n_1248),
.C(n_1227),
.Y(n_1345)
);

OAI21x1_ASAP7_75t_L g1346 ( 
.A1(n_1143),
.A2(n_1189),
.B(n_1266),
.Y(n_1346)
);

OAI21x1_ASAP7_75t_L g1347 ( 
.A1(n_1143),
.A2(n_1189),
.B(n_1266),
.Y(n_1347)
);

OAI21xp5_ASAP7_75t_L g1348 ( 
.A1(n_1265),
.A2(n_1245),
.B(n_1019),
.Y(n_1348)
);

AOI22xp33_ASAP7_75t_L g1349 ( 
.A1(n_1194),
.A2(n_820),
.B1(n_1044),
.B2(n_856),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1224),
.B(n_1231),
.Y(n_1350)
);

AOI22xp33_ASAP7_75t_L g1351 ( 
.A1(n_1194),
.A2(n_820),
.B1(n_1044),
.B2(n_856),
.Y(n_1351)
);

OA21x2_ASAP7_75t_L g1352 ( 
.A1(n_1186),
.A2(n_1143),
.B(n_1192),
.Y(n_1352)
);

OA21x2_ASAP7_75t_L g1353 ( 
.A1(n_1186),
.A2(n_1143),
.B(n_1192),
.Y(n_1353)
);

AOI22xp5_ASAP7_75t_L g1354 ( 
.A1(n_1251),
.A2(n_676),
.B1(n_898),
.B2(n_816),
.Y(n_1354)
);

NOR2xp67_ASAP7_75t_L g1355 ( 
.A(n_1125),
.B(n_568),
.Y(n_1355)
);

OR2x2_ASAP7_75t_L g1356 ( 
.A(n_1125),
.B(n_1196),
.Y(n_1356)
);

OAI21x1_ASAP7_75t_L g1357 ( 
.A1(n_1143),
.A2(n_1189),
.B(n_1266),
.Y(n_1357)
);

AND2x4_ASAP7_75t_L g1358 ( 
.A(n_1163),
.B(n_1172),
.Y(n_1358)
);

OAI21x1_ASAP7_75t_L g1359 ( 
.A1(n_1143),
.A2(n_1189),
.B(n_1266),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1224),
.B(n_1231),
.Y(n_1360)
);

O2A1O1Ixp33_ASAP7_75t_SL g1361 ( 
.A1(n_1265),
.A2(n_1227),
.B(n_1248),
.C(n_1194),
.Y(n_1361)
);

OR2x2_ASAP7_75t_L g1362 ( 
.A(n_1125),
.B(n_1196),
.Y(n_1362)
);

INVxp67_ASAP7_75t_SL g1363 ( 
.A(n_1227),
.Y(n_1363)
);

AOI221xp5_ASAP7_75t_L g1364 ( 
.A1(n_1194),
.A2(n_986),
.B1(n_646),
.B2(n_942),
.C(n_1247),
.Y(n_1364)
);

CKINVDCx5p33_ASAP7_75t_R g1365 ( 
.A(n_1181),
.Y(n_1365)
);

OAI21x1_ASAP7_75t_L g1366 ( 
.A1(n_1143),
.A2(n_1189),
.B(n_1266),
.Y(n_1366)
);

OAI21x1_ASAP7_75t_L g1367 ( 
.A1(n_1143),
.A2(n_1189),
.B(n_1266),
.Y(n_1367)
);

CKINVDCx20_ASAP7_75t_R g1368 ( 
.A(n_1181),
.Y(n_1368)
);

INVxp67_ASAP7_75t_L g1369 ( 
.A(n_1196),
.Y(n_1369)
);

AND2x4_ASAP7_75t_L g1370 ( 
.A(n_1163),
.B(n_1172),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1197),
.Y(n_1371)
);

OA21x2_ASAP7_75t_L g1372 ( 
.A1(n_1186),
.A2(n_1143),
.B(n_1192),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1197),
.Y(n_1373)
);

AO21x2_ASAP7_75t_L g1374 ( 
.A1(n_1186),
.A2(n_1192),
.B(n_1164),
.Y(n_1374)
);

OAI21x1_ASAP7_75t_L g1375 ( 
.A1(n_1143),
.A2(n_1189),
.B(n_1266),
.Y(n_1375)
);

OAI21x1_ASAP7_75t_L g1376 ( 
.A1(n_1143),
.A2(n_1189),
.B(n_1266),
.Y(n_1376)
);

OAI22xp5_ASAP7_75t_L g1377 ( 
.A1(n_1265),
.A2(n_822),
.B1(n_851),
.B2(n_1224),
.Y(n_1377)
);

BUFx8_ASAP7_75t_L g1378 ( 
.A(n_1162),
.Y(n_1378)
);

INVx4_ASAP7_75t_L g1379 ( 
.A(n_1233),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1224),
.B(n_1231),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1197),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1197),
.Y(n_1382)
);

OAI21x1_ASAP7_75t_L g1383 ( 
.A1(n_1143),
.A2(n_1189),
.B(n_1266),
.Y(n_1383)
);

OAI21x1_ASAP7_75t_L g1384 ( 
.A1(n_1143),
.A2(n_1189),
.B(n_1266),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1224),
.B(n_1231),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_SL g1386 ( 
.A(n_1265),
.B(n_1194),
.Y(n_1386)
);

OAI222xp33_ASAP7_75t_L g1387 ( 
.A1(n_1188),
.A2(n_1248),
.B1(n_1227),
.B2(n_1029),
.C1(n_822),
.C2(n_1217),
.Y(n_1387)
);

OAI22xp5_ASAP7_75t_SL g1388 ( 
.A1(n_1251),
.A2(n_816),
.B1(n_1217),
.B2(n_898),
.Y(n_1388)
);

O2A1O1Ixp33_ASAP7_75t_SL g1389 ( 
.A1(n_1265),
.A2(n_1227),
.B(n_1248),
.C(n_1194),
.Y(n_1389)
);

A2O1A1Ixp33_ASAP7_75t_L g1390 ( 
.A1(n_1265),
.A2(n_822),
.B(n_1248),
.C(n_1227),
.Y(n_1390)
);

OAI21x1_ASAP7_75t_L g1391 ( 
.A1(n_1143),
.A2(n_1189),
.B(n_1266),
.Y(n_1391)
);

AOI221xp5_ASAP7_75t_L g1392 ( 
.A1(n_1364),
.A2(n_1276),
.B1(n_1349),
.B2(n_1351),
.C(n_1287),
.Y(n_1392)
);

CKINVDCx20_ASAP7_75t_R g1393 ( 
.A(n_1368),
.Y(n_1393)
);

AND2x4_ASAP7_75t_L g1394 ( 
.A(n_1358),
.B(n_1370),
.Y(n_1394)
);

AOI21xp5_ASAP7_75t_SL g1395 ( 
.A1(n_1269),
.A2(n_1377),
.B(n_1345),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_1368),
.Y(n_1396)
);

INVx3_ASAP7_75t_L g1397 ( 
.A(n_1334),
.Y(n_1397)
);

BUFx3_ASAP7_75t_L g1398 ( 
.A(n_1378),
.Y(n_1398)
);

O2A1O1Ixp5_ASAP7_75t_L g1399 ( 
.A1(n_1386),
.A2(n_1314),
.B(n_1348),
.C(n_1276),
.Y(n_1399)
);

O2A1O1Ixp33_ASAP7_75t_L g1400 ( 
.A1(n_1386),
.A2(n_1387),
.B(n_1351),
.C(n_1349),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1360),
.B(n_1380),
.Y(n_1401)
);

O2A1O1Ixp33_ASAP7_75t_L g1402 ( 
.A1(n_1387),
.A2(n_1361),
.B(n_1389),
.C(n_1390),
.Y(n_1402)
);

OR2x2_ASAP7_75t_L g1403 ( 
.A(n_1362),
.B(n_1321),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1363),
.B(n_1330),
.Y(n_1404)
);

OAI22xp5_ASAP7_75t_L g1405 ( 
.A1(n_1354),
.A2(n_1291),
.B1(n_1309),
.B2(n_1302),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1307),
.B(n_1283),
.Y(n_1406)
);

CKINVDCx5p33_ASAP7_75t_R g1407 ( 
.A(n_1301),
.Y(n_1407)
);

INVx3_ASAP7_75t_L g1408 ( 
.A(n_1339),
.Y(n_1408)
);

OAI22xp5_ASAP7_75t_L g1409 ( 
.A1(n_1291),
.A2(n_1385),
.B1(n_1388),
.B2(n_1369),
.Y(n_1409)
);

INVx1_ASAP7_75t_SL g1410 ( 
.A(n_1278),
.Y(n_1410)
);

A2O1A1Ixp33_ASAP7_75t_L g1411 ( 
.A1(n_1345),
.A2(n_1390),
.B(n_1344),
.C(n_1305),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1363),
.B(n_1342),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1313),
.B(n_1312),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1312),
.B(n_1305),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1322),
.B(n_1268),
.Y(n_1415)
);

CKINVDCx5p33_ASAP7_75t_R g1416 ( 
.A(n_1301),
.Y(n_1416)
);

INVx3_ASAP7_75t_L g1417 ( 
.A(n_1358),
.Y(n_1417)
);

OA21x2_ASAP7_75t_L g1418 ( 
.A1(n_1343),
.A2(n_1337),
.B(n_1335),
.Y(n_1418)
);

NOR2xp33_ASAP7_75t_L g1419 ( 
.A(n_1369),
.B(n_1308),
.Y(n_1419)
);

INVx1_ASAP7_75t_SL g1420 ( 
.A(n_1273),
.Y(n_1420)
);

OR2x2_ASAP7_75t_L g1421 ( 
.A(n_1289),
.B(n_1290),
.Y(n_1421)
);

OA21x2_ASAP7_75t_L g1422 ( 
.A1(n_1300),
.A2(n_1271),
.B(n_1306),
.Y(n_1422)
);

INVx8_ASAP7_75t_L g1423 ( 
.A(n_1299),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1371),
.B(n_1373),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1381),
.B(n_1382),
.Y(n_1425)
);

OA21x2_ASAP7_75t_L g1426 ( 
.A1(n_1271),
.A2(n_1306),
.B(n_1292),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1324),
.B(n_1323),
.Y(n_1427)
);

O2A1O1Ixp33_ASAP7_75t_L g1428 ( 
.A1(n_1361),
.A2(n_1389),
.B(n_1328),
.C(n_1325),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_1365),
.Y(n_1429)
);

OAI22xp5_ASAP7_75t_L g1430 ( 
.A1(n_1325),
.A2(n_1355),
.B1(n_1284),
.B2(n_1298),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1324),
.B(n_1303),
.Y(n_1431)
);

OAI22xp5_ASAP7_75t_L g1432 ( 
.A1(n_1325),
.A2(n_1273),
.B1(n_1277),
.B2(n_1331),
.Y(n_1432)
);

OAI22xp5_ASAP7_75t_L g1433 ( 
.A1(n_1331),
.A2(n_1294),
.B1(n_1279),
.B2(n_1303),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1303),
.B(n_1329),
.Y(n_1434)
);

INVx1_ASAP7_75t_SL g1435 ( 
.A(n_1297),
.Y(n_1435)
);

INVx1_ASAP7_75t_SL g1436 ( 
.A(n_1297),
.Y(n_1436)
);

AND2x4_ASAP7_75t_L g1437 ( 
.A(n_1327),
.B(n_1311),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1315),
.B(n_1336),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1316),
.B(n_1272),
.Y(n_1439)
);

NOR2xp67_ASAP7_75t_L g1440 ( 
.A(n_1320),
.B(n_1326),
.Y(n_1440)
);

INVx1_ASAP7_75t_SL g1441 ( 
.A(n_1319),
.Y(n_1441)
);

OR2x2_ASAP7_75t_L g1442 ( 
.A(n_1318),
.B(n_1310),
.Y(n_1442)
);

O2A1O1Ixp33_ASAP7_75t_L g1443 ( 
.A1(n_1374),
.A2(n_1331),
.B(n_1338),
.C(n_1275),
.Y(n_1443)
);

HB1xp67_ASAP7_75t_L g1444 ( 
.A(n_1332),
.Y(n_1444)
);

OAI22xp5_ASAP7_75t_L g1445 ( 
.A1(n_1299),
.A2(n_1288),
.B1(n_1282),
.B2(n_1365),
.Y(n_1445)
);

HB1xp67_ASAP7_75t_L g1446 ( 
.A(n_1333),
.Y(n_1446)
);

O2A1O1Ixp33_ASAP7_75t_L g1447 ( 
.A1(n_1275),
.A2(n_1280),
.B(n_1293),
.C(n_1352),
.Y(n_1447)
);

AOI221x1_ASAP7_75t_SL g1448 ( 
.A1(n_1378),
.A2(n_1295),
.B1(n_1275),
.B2(n_1341),
.C(n_1340),
.Y(n_1448)
);

OAI22xp5_ASAP7_75t_L g1449 ( 
.A1(n_1299),
.A2(n_1304),
.B1(n_1379),
.B2(n_1296),
.Y(n_1449)
);

O2A1O1Ixp33_ASAP7_75t_L g1450 ( 
.A1(n_1280),
.A2(n_1293),
.B(n_1352),
.C(n_1372),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1317),
.B(n_1310),
.Y(n_1451)
);

BUFx2_ASAP7_75t_L g1452 ( 
.A(n_1378),
.Y(n_1452)
);

AND2x4_ASAP7_75t_L g1453 ( 
.A(n_1296),
.B(n_1379),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1340),
.B(n_1293),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1341),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1281),
.Y(n_1456)
);

OA21x2_ASAP7_75t_L g1457 ( 
.A1(n_1346),
.A2(n_1366),
.B(n_1384),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1353),
.B(n_1372),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1353),
.B(n_1281),
.Y(n_1459)
);

O2A1O1Ixp33_ASAP7_75t_L g1460 ( 
.A1(n_1285),
.A2(n_1286),
.B(n_1347),
.C(n_1357),
.Y(n_1460)
);

AOI21xp5_ASAP7_75t_SL g1461 ( 
.A1(n_1359),
.A2(n_1367),
.B(n_1375),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1376),
.B(n_1383),
.Y(n_1462)
);

O2A1O1Ixp33_ASAP7_75t_L g1463 ( 
.A1(n_1391),
.A2(n_1364),
.B(n_1265),
.C(n_1287),
.Y(n_1463)
);

AOI21xp5_ASAP7_75t_L g1464 ( 
.A1(n_1269),
.A2(n_822),
.B(n_1265),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1274),
.B(n_1350),
.Y(n_1465)
);

AOI21xp5_ASAP7_75t_L g1466 ( 
.A1(n_1269),
.A2(n_822),
.B(n_1265),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1307),
.B(n_1321),
.Y(n_1467)
);

OAI22xp5_ASAP7_75t_L g1468 ( 
.A1(n_1349),
.A2(n_1351),
.B1(n_822),
.B2(n_1364),
.Y(n_1468)
);

AOI21xp5_ASAP7_75t_L g1469 ( 
.A1(n_1269),
.A2(n_822),
.B(n_1265),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1274),
.B(n_1350),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1363),
.B(n_1330),
.Y(n_1471)
);

OR2x2_ASAP7_75t_L g1472 ( 
.A(n_1270),
.B(n_1356),
.Y(n_1472)
);

O2A1O1Ixp33_ASAP7_75t_L g1473 ( 
.A1(n_1364),
.A2(n_1265),
.B(n_1287),
.C(n_1386),
.Y(n_1473)
);

AOI221xp5_ASAP7_75t_L g1474 ( 
.A1(n_1364),
.A2(n_986),
.B1(n_942),
.B2(n_1276),
.C(n_1194),
.Y(n_1474)
);

OAI22xp5_ASAP7_75t_L g1475 ( 
.A1(n_1349),
.A2(n_1351),
.B1(n_822),
.B2(n_1364),
.Y(n_1475)
);

AOI21xp5_ASAP7_75t_SL g1476 ( 
.A1(n_1269),
.A2(n_1265),
.B(n_1248),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1274),
.B(n_1350),
.Y(n_1477)
);

AOI221x1_ASAP7_75t_SL g1478 ( 
.A1(n_1287),
.A2(n_662),
.B1(n_899),
.B2(n_942),
.C(n_597),
.Y(n_1478)
);

OAI22xp5_ASAP7_75t_L g1479 ( 
.A1(n_1349),
.A2(n_1351),
.B1(n_822),
.B2(n_1364),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1274),
.B(n_1350),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1307),
.B(n_1321),
.Y(n_1481)
);

OAI22xp5_ASAP7_75t_L g1482 ( 
.A1(n_1349),
.A2(n_1351),
.B1(n_822),
.B2(n_1364),
.Y(n_1482)
);

HB1xp67_ASAP7_75t_L g1483 ( 
.A(n_1444),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1456),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1412),
.B(n_1404),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1404),
.B(n_1471),
.Y(n_1486)
);

OR2x2_ASAP7_75t_L g1487 ( 
.A(n_1454),
.B(n_1442),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1444),
.Y(n_1488)
);

BUFx2_ASAP7_75t_L g1489 ( 
.A(n_1437),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1408),
.B(n_1459),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1446),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1455),
.Y(n_1492)
);

BUFx12f_ASAP7_75t_L g1493 ( 
.A(n_1396),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1418),
.B(n_1437),
.Y(n_1494)
);

AND2x4_ASAP7_75t_L g1495 ( 
.A(n_1397),
.B(n_1462),
.Y(n_1495)
);

INVxp67_ASAP7_75t_SL g1496 ( 
.A(n_1443),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_1418),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1414),
.B(n_1413),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1421),
.Y(n_1499)
);

INVx5_ASAP7_75t_L g1500 ( 
.A(n_1423),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1422),
.Y(n_1501)
);

AND2x2_ASAP7_75t_SL g1502 ( 
.A(n_1474),
.B(n_1392),
.Y(n_1502)
);

OR2x2_ASAP7_75t_L g1503 ( 
.A(n_1458),
.B(n_1422),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1439),
.Y(n_1504)
);

HB1xp67_ASAP7_75t_L g1505 ( 
.A(n_1448),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_1457),
.Y(n_1506)
);

NOR2x1_ASAP7_75t_L g1507 ( 
.A(n_1395),
.B(n_1476),
.Y(n_1507)
);

AOI21x1_ASAP7_75t_L g1508 ( 
.A1(n_1457),
.A2(n_1426),
.B(n_1466),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1411),
.B(n_1434),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1411),
.B(n_1401),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1425),
.Y(n_1511)
);

NOR2xp33_ASAP7_75t_L g1512 ( 
.A(n_1405),
.B(n_1473),
.Y(n_1512)
);

OR2x6_ASAP7_75t_L g1513 ( 
.A(n_1395),
.B(n_1476),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1426),
.B(n_1451),
.Y(n_1514)
);

NOR2x1_ASAP7_75t_SL g1515 ( 
.A(n_1433),
.B(n_1432),
.Y(n_1515)
);

AOI21x1_ASAP7_75t_L g1516 ( 
.A1(n_1464),
.A2(n_1469),
.B(n_1479),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1424),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1447),
.B(n_1417),
.Y(n_1518)
);

OA21x2_ASAP7_75t_L g1519 ( 
.A1(n_1399),
.A2(n_1427),
.B(n_1475),
.Y(n_1519)
);

OAI21x1_ASAP7_75t_L g1520 ( 
.A1(n_1450),
.A2(n_1460),
.B(n_1461),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1417),
.B(n_1431),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1406),
.B(n_1438),
.Y(n_1522)
);

INVx3_ASAP7_75t_L g1523 ( 
.A(n_1394),
.Y(n_1523)
);

AND2x4_ASAP7_75t_L g1524 ( 
.A(n_1394),
.B(n_1415),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1463),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1428),
.Y(n_1526)
);

OA21x2_ASAP7_75t_L g1527 ( 
.A1(n_1468),
.A2(n_1482),
.B(n_1419),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1514),
.B(n_1419),
.Y(n_1528)
);

AOI22xp33_ASAP7_75t_L g1529 ( 
.A1(n_1502),
.A2(n_1512),
.B1(n_1507),
.B2(n_1527),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1496),
.B(n_1465),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1484),
.Y(n_1531)
);

BUFx3_ASAP7_75t_L g1532 ( 
.A(n_1495),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1514),
.B(n_1490),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1514),
.B(n_1481),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1506),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1496),
.B(n_1480),
.Y(n_1536)
);

AND2x4_ASAP7_75t_SL g1537 ( 
.A(n_1513),
.B(n_1453),
.Y(n_1537)
);

BUFx2_ASAP7_75t_L g1538 ( 
.A(n_1494),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1494),
.B(n_1467),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1487),
.B(n_1477),
.Y(n_1540)
);

HB1xp67_ASAP7_75t_L g1541 ( 
.A(n_1483),
.Y(n_1541)
);

OAI21xp5_ASAP7_75t_L g1542 ( 
.A1(n_1507),
.A2(n_1402),
.B(n_1400),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1504),
.B(n_1486),
.Y(n_1543)
);

BUFx6f_ASAP7_75t_L g1544 ( 
.A(n_1520),
.Y(n_1544)
);

AOI22xp33_ASAP7_75t_L g1545 ( 
.A1(n_1502),
.A2(n_1409),
.B1(n_1470),
.B2(n_1472),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1487),
.B(n_1478),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1497),
.B(n_1420),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1492),
.Y(n_1548)
);

OR2x2_ASAP7_75t_L g1549 ( 
.A(n_1503),
.B(n_1403),
.Y(n_1549)
);

OAI21xp5_ASAP7_75t_L g1550 ( 
.A1(n_1502),
.A2(n_1430),
.B(n_1445),
.Y(n_1550)
);

OR2x2_ASAP7_75t_L g1551 ( 
.A(n_1503),
.B(n_1410),
.Y(n_1551)
);

AOI221xp5_ASAP7_75t_L g1552 ( 
.A1(n_1529),
.A2(n_1512),
.B1(n_1542),
.B2(n_1546),
.C(n_1545),
.Y(n_1552)
);

OAI211xp5_ASAP7_75t_L g1553 ( 
.A1(n_1529),
.A2(n_1542),
.B(n_1545),
.C(n_1550),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1540),
.B(n_1504),
.Y(n_1554)
);

AOI22xp5_ASAP7_75t_L g1555 ( 
.A1(n_1542),
.A2(n_1502),
.B1(n_1513),
.B2(n_1527),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1540),
.B(n_1498),
.Y(n_1556)
);

AOI22xp33_ASAP7_75t_L g1557 ( 
.A1(n_1550),
.A2(n_1513),
.B1(n_1527),
.B2(n_1525),
.Y(n_1557)
);

OAI21x1_ASAP7_75t_L g1558 ( 
.A1(n_1535),
.A2(n_1520),
.B(n_1508),
.Y(n_1558)
);

OAI33xp33_ASAP7_75t_L g1559 ( 
.A1(n_1546),
.A2(n_1525),
.A3(n_1498),
.B1(n_1526),
.B2(n_1510),
.B3(n_1511),
.Y(n_1559)
);

OAI221xp5_ASAP7_75t_SL g1560 ( 
.A1(n_1546),
.A2(n_1513),
.B1(n_1510),
.B2(n_1525),
.C(n_1505),
.Y(n_1560)
);

AOI22xp33_ASAP7_75t_L g1561 ( 
.A1(n_1550),
.A2(n_1513),
.B1(n_1527),
.B2(n_1505),
.Y(n_1561)
);

NOR4xp25_ASAP7_75t_SL g1562 ( 
.A(n_1538),
.B(n_1396),
.C(n_1489),
.D(n_1416),
.Y(n_1562)
);

INVxp33_ASAP7_75t_L g1563 ( 
.A(n_1536),
.Y(n_1563)
);

BUFx3_ASAP7_75t_L g1564 ( 
.A(n_1551),
.Y(n_1564)
);

OAI211xp5_ASAP7_75t_SL g1565 ( 
.A1(n_1536),
.A2(n_1526),
.B(n_1441),
.C(n_1435),
.Y(n_1565)
);

BUFx3_ASAP7_75t_L g1566 ( 
.A(n_1551),
.Y(n_1566)
);

AOI221xp5_ASAP7_75t_L g1567 ( 
.A1(n_1530),
.A2(n_1509),
.B1(n_1511),
.B2(n_1499),
.C(n_1522),
.Y(n_1567)
);

AOI222xp33_ASAP7_75t_L g1568 ( 
.A1(n_1530),
.A2(n_1509),
.B1(n_1515),
.B2(n_1493),
.C1(n_1436),
.C2(n_1522),
.Y(n_1568)
);

AOI21xp5_ASAP7_75t_L g1569 ( 
.A1(n_1530),
.A2(n_1513),
.B(n_1527),
.Y(n_1569)
);

INVx2_ASAP7_75t_R g1570 ( 
.A(n_1531),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1533),
.B(n_1489),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1533),
.B(n_1485),
.Y(n_1572)
);

AOI221xp5_ASAP7_75t_L g1573 ( 
.A1(n_1540),
.A2(n_1509),
.B1(n_1499),
.B2(n_1522),
.C(n_1517),
.Y(n_1573)
);

HB1xp67_ASAP7_75t_L g1574 ( 
.A(n_1541),
.Y(n_1574)
);

NAND3xp33_ASAP7_75t_L g1575 ( 
.A(n_1551),
.B(n_1527),
.C(n_1513),
.Y(n_1575)
);

OAI31xp33_ASAP7_75t_SL g1576 ( 
.A1(n_1528),
.A2(n_1485),
.A3(n_1524),
.B(n_1521),
.Y(n_1576)
);

NAND3xp33_ASAP7_75t_L g1577 ( 
.A(n_1551),
.B(n_1519),
.C(n_1518),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1548),
.Y(n_1578)
);

NAND4xp25_ASAP7_75t_L g1579 ( 
.A(n_1549),
.B(n_1440),
.C(n_1487),
.D(n_1518),
.Y(n_1579)
);

AO21x1_ASAP7_75t_SL g1580 ( 
.A1(n_1543),
.A2(n_1491),
.B(n_1488),
.Y(n_1580)
);

INVx1_ASAP7_75t_SL g1581 ( 
.A(n_1549),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1548),
.Y(n_1582)
);

HB1xp67_ASAP7_75t_L g1583 ( 
.A(n_1541),
.Y(n_1583)
);

AND2x4_ASAP7_75t_L g1584 ( 
.A(n_1532),
.B(n_1523),
.Y(n_1584)
);

HB1xp67_ASAP7_75t_L g1585 ( 
.A(n_1574),
.Y(n_1585)
);

OA21x2_ASAP7_75t_L g1586 ( 
.A1(n_1558),
.A2(n_1497),
.B(n_1501),
.Y(n_1586)
);

INVx4_ASAP7_75t_SL g1587 ( 
.A(n_1564),
.Y(n_1587)
);

HB1xp67_ASAP7_75t_L g1588 ( 
.A(n_1583),
.Y(n_1588)
);

BUFx2_ASAP7_75t_L g1589 ( 
.A(n_1584),
.Y(n_1589)
);

NOR3xp33_ASAP7_75t_L g1590 ( 
.A(n_1553),
.B(n_1516),
.C(n_1452),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1563),
.B(n_1528),
.Y(n_1591)
);

INVx2_ASAP7_75t_SL g1592 ( 
.A(n_1584),
.Y(n_1592)
);

OR2x2_ASAP7_75t_L g1593 ( 
.A(n_1581),
.B(n_1549),
.Y(n_1593)
);

BUFx2_ASAP7_75t_L g1594 ( 
.A(n_1584),
.Y(n_1594)
);

INVx2_ASAP7_75t_SL g1595 ( 
.A(n_1578),
.Y(n_1595)
);

NAND3xp33_ASAP7_75t_SL g1596 ( 
.A(n_1552),
.B(n_1393),
.C(n_1407),
.Y(n_1596)
);

NAND3xp33_ASAP7_75t_SL g1597 ( 
.A(n_1555),
.B(n_1393),
.C(n_1407),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1578),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1582),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1582),
.Y(n_1600)
);

NOR2xp33_ASAP7_75t_L g1601 ( 
.A(n_1565),
.B(n_1493),
.Y(n_1601)
);

OR2x6_ASAP7_75t_L g1602 ( 
.A(n_1569),
.B(n_1544),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1572),
.B(n_1538),
.Y(n_1603)
);

INVx4_ASAP7_75t_L g1604 ( 
.A(n_1564),
.Y(n_1604)
);

BUFx3_ASAP7_75t_L g1605 ( 
.A(n_1566),
.Y(n_1605)
);

OR2x2_ASAP7_75t_L g1606 ( 
.A(n_1591),
.B(n_1577),
.Y(n_1606)
);

HB1xp67_ASAP7_75t_L g1607 ( 
.A(n_1595),
.Y(n_1607)
);

NOR2xp33_ASAP7_75t_L g1608 ( 
.A(n_1596),
.B(n_1493),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1585),
.B(n_1528),
.Y(n_1609)
);

CKINVDCx20_ASAP7_75t_R g1610 ( 
.A(n_1596),
.Y(n_1610)
);

OR2x2_ASAP7_75t_L g1611 ( 
.A(n_1591),
.B(n_1554),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_1586),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1585),
.B(n_1556),
.Y(n_1613)
);

NAND3xp33_ASAP7_75t_L g1614 ( 
.A(n_1590),
.B(n_1560),
.C(n_1561),
.Y(n_1614)
);

NOR2x1_ASAP7_75t_L g1615 ( 
.A(n_1604),
.B(n_1575),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1587),
.B(n_1576),
.Y(n_1616)
);

AND4x1_ASAP7_75t_L g1617 ( 
.A(n_1590),
.B(n_1559),
.C(n_1568),
.D(n_1557),
.Y(n_1617)
);

HB1xp67_ASAP7_75t_L g1618 ( 
.A(n_1595),
.Y(n_1618)
);

CKINVDCx20_ASAP7_75t_R g1619 ( 
.A(n_1601),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1587),
.B(n_1572),
.Y(n_1620)
);

NAND2x1_ASAP7_75t_L g1621 ( 
.A(n_1604),
.B(n_1538),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1587),
.B(n_1571),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1587),
.B(n_1571),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1587),
.B(n_1570),
.Y(n_1624)
);

OAI31xp33_ASAP7_75t_L g1625 ( 
.A1(n_1605),
.A2(n_1579),
.A3(n_1398),
.B(n_1566),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1588),
.B(n_1567),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1587),
.B(n_1533),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1598),
.Y(n_1628)
);

HB1xp67_ASAP7_75t_L g1629 ( 
.A(n_1595),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1588),
.B(n_1534),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1589),
.B(n_1570),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1599),
.Y(n_1632)
);

OAI31xp33_ASAP7_75t_L g1633 ( 
.A1(n_1605),
.A2(n_1398),
.A3(n_1537),
.B(n_1547),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1599),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1594),
.B(n_1534),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1594),
.B(n_1570),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1602),
.B(n_1592),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1602),
.B(n_1580),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1602),
.B(n_1580),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1628),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1628),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1623),
.B(n_1592),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1623),
.B(n_1604),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1632),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1631),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1632),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1622),
.B(n_1604),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1617),
.B(n_1614),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_SL g1649 ( 
.A(n_1625),
.B(n_1605),
.Y(n_1649)
);

NOR2xp33_ASAP7_75t_SL g1650 ( 
.A(n_1625),
.B(n_1597),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1617),
.B(n_1534),
.Y(n_1651)
);

NAND2x1p5_ASAP7_75t_L g1652 ( 
.A(n_1615),
.B(n_1500),
.Y(n_1652)
);

INVx1_ASAP7_75t_SL g1653 ( 
.A(n_1619),
.Y(n_1653)
);

INVx1_ASAP7_75t_SL g1654 ( 
.A(n_1610),
.Y(n_1654)
);

AOI22xp33_ASAP7_75t_SL g1655 ( 
.A1(n_1614),
.A2(n_1515),
.B1(n_1544),
.B2(n_1602),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1634),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1634),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1622),
.B(n_1603),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1622),
.B(n_1603),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1607),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1607),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1616),
.B(n_1603),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1618),
.Y(n_1663)
);

INVx1_ASAP7_75t_SL g1664 ( 
.A(n_1616),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1616),
.B(n_1602),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1618),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1620),
.B(n_1602),
.Y(n_1667)
);

AND2x4_ASAP7_75t_L g1668 ( 
.A(n_1620),
.B(n_1600),
.Y(n_1668)
);

INVxp67_ASAP7_75t_L g1669 ( 
.A(n_1608),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1626),
.B(n_1539),
.Y(n_1670)
);

OR2x6_ASAP7_75t_L g1671 ( 
.A(n_1615),
.B(n_1493),
.Y(n_1671)
);

INVxp67_ASAP7_75t_SL g1672 ( 
.A(n_1621),
.Y(n_1672)
);

OR2x2_ASAP7_75t_L g1673 ( 
.A(n_1613),
.B(n_1593),
.Y(n_1673)
);

NAND3xp33_ASAP7_75t_SL g1674 ( 
.A(n_1626),
.B(n_1562),
.C(n_1573),
.Y(n_1674)
);

OR2x2_ASAP7_75t_L g1675 ( 
.A(n_1613),
.B(n_1611),
.Y(n_1675)
);

BUFx3_ASAP7_75t_L g1676 ( 
.A(n_1660),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1643),
.B(n_1642),
.Y(n_1677)
);

OR2x2_ASAP7_75t_L g1678 ( 
.A(n_1673),
.B(n_1606),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_1658),
.Y(n_1679)
);

INVx1_ASAP7_75t_SL g1680 ( 
.A(n_1653),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1640),
.Y(n_1681)
);

BUFx12f_ASAP7_75t_L g1682 ( 
.A(n_1671),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1643),
.B(n_1620),
.Y(n_1683)
);

INVx4_ASAP7_75t_L g1684 ( 
.A(n_1671),
.Y(n_1684)
);

HB1xp67_ASAP7_75t_L g1685 ( 
.A(n_1660),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1640),
.Y(n_1686)
);

INVx1_ASAP7_75t_SL g1687 ( 
.A(n_1654),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_1645),
.Y(n_1688)
);

OAI22x1_ASAP7_75t_SL g1689 ( 
.A1(n_1664),
.A2(n_1416),
.B1(n_1429),
.B2(n_1633),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1658),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1641),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1642),
.B(n_1627),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1641),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1661),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1648),
.B(n_1635),
.Y(n_1695)
);

OR2x2_ASAP7_75t_L g1696 ( 
.A(n_1673),
.B(n_1606),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1661),
.Y(n_1697)
);

NOR2x1_ASAP7_75t_L g1698 ( 
.A(n_1671),
.B(n_1621),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1651),
.B(n_1635),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1666),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1666),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1685),
.Y(n_1702)
);

INVxp67_ASAP7_75t_L g1703 ( 
.A(n_1695),
.Y(n_1703)
);

NAND2x1_ASAP7_75t_SL g1704 ( 
.A(n_1698),
.B(n_1647),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1676),
.Y(n_1705)
);

HB1xp67_ASAP7_75t_L g1706 ( 
.A(n_1676),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1676),
.Y(n_1707)
);

OAI21xp5_ASAP7_75t_L g1708 ( 
.A1(n_1698),
.A2(n_1650),
.B(n_1655),
.Y(n_1708)
);

INVxp67_ASAP7_75t_L g1709 ( 
.A(n_1677),
.Y(n_1709)
);

NOR2xp33_ASAP7_75t_L g1710 ( 
.A(n_1687),
.B(n_1669),
.Y(n_1710)
);

NAND4xp25_ASAP7_75t_L g1711 ( 
.A(n_1680),
.B(n_1649),
.C(n_1674),
.D(n_1663),
.Y(n_1711)
);

AOI222xp33_ASAP7_75t_L g1712 ( 
.A1(n_1689),
.A2(n_1682),
.B1(n_1597),
.B2(n_1699),
.C1(n_1697),
.C2(n_1694),
.Y(n_1712)
);

INVx1_ASAP7_75t_SL g1713 ( 
.A(n_1677),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1683),
.B(n_1647),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1681),
.Y(n_1715)
);

AOI22xp33_ASAP7_75t_L g1716 ( 
.A1(n_1682),
.A2(n_1671),
.B1(n_1652),
.B2(n_1670),
.Y(n_1716)
);

INVx1_ASAP7_75t_SL g1717 ( 
.A(n_1678),
.Y(n_1717)
);

OAI21xp5_ASAP7_75t_L g1718 ( 
.A1(n_1678),
.A2(n_1652),
.B(n_1672),
.Y(n_1718)
);

NAND2x1_ASAP7_75t_SL g1719 ( 
.A(n_1683),
.B(n_1624),
.Y(n_1719)
);

OAI21xp5_ASAP7_75t_L g1720 ( 
.A1(n_1696),
.A2(n_1652),
.B(n_1665),
.Y(n_1720)
);

OR2x2_ASAP7_75t_L g1721 ( 
.A(n_1696),
.B(n_1675),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1719),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1706),
.Y(n_1723)
);

INVxp67_ASAP7_75t_L g1724 ( 
.A(n_1706),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1705),
.Y(n_1725)
);

NOR2xp33_ASAP7_75t_L g1726 ( 
.A(n_1717),
.B(n_1684),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1707),
.Y(n_1727)
);

INVx1_ASAP7_75t_SL g1728 ( 
.A(n_1704),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1713),
.B(n_1679),
.Y(n_1729)
);

INVx1_ASAP7_75t_SL g1730 ( 
.A(n_1721),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1710),
.B(n_1679),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1710),
.B(n_1690),
.Y(n_1732)
);

NAND2xp33_ASAP7_75t_L g1733 ( 
.A(n_1708),
.B(n_1690),
.Y(n_1733)
);

AOI21x1_ASAP7_75t_L g1734 ( 
.A1(n_1723),
.A2(n_1702),
.B(n_1715),
.Y(n_1734)
);

O2A1O1Ixp5_ASAP7_75t_SL g1735 ( 
.A1(n_1724),
.A2(n_1701),
.B(n_1700),
.C(n_1697),
.Y(n_1735)
);

O2A1O1Ixp33_ASAP7_75t_L g1736 ( 
.A1(n_1733),
.A2(n_1711),
.B(n_1712),
.C(n_1703),
.Y(n_1736)
);

NAND4xp25_ASAP7_75t_L g1737 ( 
.A(n_1726),
.B(n_1709),
.C(n_1716),
.D(n_1684),
.Y(n_1737)
);

AOI22xp5_ASAP7_75t_L g1738 ( 
.A1(n_1730),
.A2(n_1714),
.B1(n_1689),
.B2(n_1684),
.Y(n_1738)
);

OAI221xp5_ASAP7_75t_L g1739 ( 
.A1(n_1728),
.A2(n_1716),
.B1(n_1720),
.B2(n_1718),
.C(n_1684),
.Y(n_1739)
);

AOI31xp33_ASAP7_75t_L g1740 ( 
.A1(n_1726),
.A2(n_1700),
.A3(n_1694),
.B(n_1701),
.Y(n_1740)
);

OAI22xp5_ASAP7_75t_L g1741 ( 
.A1(n_1731),
.A2(n_1692),
.B1(n_1675),
.B2(n_1662),
.Y(n_1741)
);

OAI21xp33_ASAP7_75t_L g1742 ( 
.A1(n_1732),
.A2(n_1692),
.B(n_1662),
.Y(n_1742)
);

NOR3xp33_ASAP7_75t_L g1743 ( 
.A(n_1729),
.B(n_1693),
.C(n_1686),
.Y(n_1743)
);

AOI21xp5_ASAP7_75t_L g1744 ( 
.A1(n_1722),
.A2(n_1688),
.B(n_1686),
.Y(n_1744)
);

XNOR2xp5_ASAP7_75t_L g1745 ( 
.A(n_1738),
.B(n_1725),
.Y(n_1745)
);

OAI22xp5_ASAP7_75t_L g1746 ( 
.A1(n_1736),
.A2(n_1722),
.B1(n_1727),
.B2(n_1665),
.Y(n_1746)
);

OA22x2_ASAP7_75t_L g1747 ( 
.A1(n_1742),
.A2(n_1688),
.B1(n_1691),
.B2(n_1681),
.Y(n_1747)
);

O2A1O1Ixp33_ASAP7_75t_L g1748 ( 
.A1(n_1740),
.A2(n_1693),
.B(n_1691),
.C(n_1688),
.Y(n_1748)
);

NAND2xp33_ASAP7_75t_SL g1749 ( 
.A(n_1741),
.B(n_1429),
.Y(n_1749)
);

O2A1O1Ixp33_ASAP7_75t_L g1750 ( 
.A1(n_1739),
.A2(n_1646),
.B(n_1644),
.C(n_1656),
.Y(n_1750)
);

NOR3x1_ASAP7_75t_L g1751 ( 
.A(n_1737),
.B(n_1657),
.C(n_1609),
.Y(n_1751)
);

INVx1_ASAP7_75t_SL g1752 ( 
.A(n_1744),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1747),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1748),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1751),
.B(n_1734),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1750),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1745),
.B(n_1743),
.Y(n_1757)
);

INVx1_ASAP7_75t_SL g1758 ( 
.A(n_1752),
.Y(n_1758)
);

NAND2x1p5_ASAP7_75t_L g1759 ( 
.A(n_1749),
.B(n_1624),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1746),
.B(n_1735),
.Y(n_1760)
);

OAI22xp5_ASAP7_75t_L g1761 ( 
.A1(n_1759),
.A2(n_1645),
.B1(n_1668),
.B2(n_1629),
.Y(n_1761)
);

HB1xp67_ASAP7_75t_L g1762 ( 
.A(n_1759),
.Y(n_1762)
);

HB1xp67_ASAP7_75t_L g1763 ( 
.A(n_1758),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1753),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1755),
.B(n_1659),
.Y(n_1765)
);

OA22x2_ASAP7_75t_L g1766 ( 
.A1(n_1762),
.A2(n_1754),
.B1(n_1756),
.B2(n_1758),
.Y(n_1766)
);

INVx2_ASAP7_75t_SL g1767 ( 
.A(n_1763),
.Y(n_1767)
);

OAI221xp5_ASAP7_75t_L g1768 ( 
.A1(n_1765),
.A2(n_1760),
.B1(n_1757),
.B2(n_1667),
.C(n_1633),
.Y(n_1768)
);

XNOR2x1_ASAP7_75t_L g1769 ( 
.A(n_1766),
.B(n_1764),
.Y(n_1769)
);

OAI221xp5_ASAP7_75t_SL g1770 ( 
.A1(n_1769),
.A2(n_1768),
.B1(n_1767),
.B2(n_1761),
.C(n_1667),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1770),
.B(n_1668),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1770),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1771),
.Y(n_1773)
);

AOI22xp5_ASAP7_75t_L g1774 ( 
.A1(n_1772),
.A2(n_1668),
.B1(n_1659),
.B2(n_1637),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1773),
.Y(n_1775)
);

OAI21x1_ASAP7_75t_SL g1776 ( 
.A1(n_1774),
.A2(n_1609),
.B(n_1630),
.Y(n_1776)
);

INVx2_ASAP7_75t_L g1777 ( 
.A(n_1776),
.Y(n_1777)
);

NOR2xp33_ASAP7_75t_L g1778 ( 
.A(n_1777),
.B(n_1775),
.Y(n_1778)
);

OAI21xp5_ASAP7_75t_L g1779 ( 
.A1(n_1778),
.A2(n_1637),
.B(n_1629),
.Y(n_1779)
);

AOI22xp5_ASAP7_75t_L g1780 ( 
.A1(n_1779),
.A2(n_1637),
.B1(n_1636),
.B2(n_1631),
.Y(n_1780)
);

AOI221xp5_ASAP7_75t_L g1781 ( 
.A1(n_1780),
.A2(n_1624),
.B1(n_1639),
.B2(n_1638),
.C(n_1612),
.Y(n_1781)
);

AOI211xp5_ASAP7_75t_L g1782 ( 
.A1(n_1781),
.A2(n_1639),
.B(n_1638),
.C(n_1449),
.Y(n_1782)
);


endmodule