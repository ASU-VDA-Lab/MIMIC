module real_jpeg_28601_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_97, n_6, n_104, n_100, n_106, n_11, n_14, n_7, n_18, n_3, n_99, n_5, n_4, n_102, n_105, n_98, n_101, n_1, n_16, n_15, n_13, n_103, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_97;
input n_6;
input n_104;
input n_100;
input n_106;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_99;
input n_5;
input n_4;
input n_102;
input n_105;
input n_98;
input n_101;
input n_1;
input n_16;
input n_15;
input n_13;
input n_103;

output n_19;

wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_83;
wire n_78;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_27;
wire n_56;
wire n_48;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_44;
wire n_28;
wire n_62;
wire n_45;
wire n_42;
wire n_77;
wire n_39;
wire n_94;
wire n_26;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_92;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_85;
wire n_89;

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_0),
.Y(n_59)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_1),
.B(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_2),
.B(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_4),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_5),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_6),
.B(n_29),
.C(n_93),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_7),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_8),
.B(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_8),
.B(n_23),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_9),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_10),
.B(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_10),
.B(n_44),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_11),
.B(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_11),
.B(n_64),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_12),
.B(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_12),
.B(n_51),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_13),
.B(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_13),
.B(n_81),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_14),
.B(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_14),
.B(n_39),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_15),
.B(n_33),
.Y(n_32)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_15),
.B(n_33),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_16),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_17),
.B(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_17),
.B(n_90),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_18),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_28),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_27),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_25),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_25),
.B(n_40),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_25),
.B(n_76),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_25),
.B(n_86),
.Y(n_85)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_26),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g29 ( 
.A1(n_30),
.A2(n_89),
.B(n_92),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_SL g30 ( 
.A1(n_31),
.A2(n_84),
.B(n_88),
.Y(n_30)
);

A2O1A1Ixp33_ASAP7_75t_SL g31 ( 
.A1(n_32),
.A2(n_36),
.B(n_80),
.C(n_83),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_34),
.B(n_35),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_34),
.B(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_34),
.B(n_82),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_34),
.B(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_37),
.B(n_79),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_41),
.B(n_78),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_73),
.B(n_77),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_46),
.B(n_72),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_67),
.B(n_71),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_SL g47 ( 
.A1(n_48),
.A2(n_63),
.B(n_66),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_58),
.B(n_62),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_SL g49 ( 
.A1(n_50),
.A2(n_54),
.B(n_57),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_52),
.B(n_53),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_52),
.B(n_61),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_52),
.B(n_65),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_60),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_59),
.B(n_60),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_69),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_68),
.B(n_69),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_75),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_74),
.B(n_75),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_85),
.B(n_87),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_85),
.B(n_87),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_95),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_97),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_98),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_99),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_100),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_101),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_102),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_103),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_104),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_105),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_106),
.Y(n_82)
);


endmodule