module fake_jpeg_2394_n_453 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_453);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_453;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx10_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_12),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_11),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_16),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_0),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

CKINVDCx14_ASAP7_75t_R g47 ( 
.A(n_6),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_1),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_19),
.B(n_17),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_55),
.B(n_68),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_56),
.Y(n_123)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_57),
.Y(n_121)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_58),
.Y(n_128)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_59),
.Y(n_178)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

BUFx10_ASAP7_75t_L g174 ( 
.A(n_60),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_61),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_19),
.B(n_16),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_62),
.B(n_93),
.Y(n_132)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_63),
.Y(n_122)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_64),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_65),
.Y(n_120)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_66),
.Y(n_146)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g152 ( 
.A(n_67),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_31),
.B(n_15),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_69),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_70),
.Y(n_180)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_27),
.Y(n_71)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_71),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

INVx6_ASAP7_75t_L g187 ( 
.A(n_72),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

INVx6_ASAP7_75t_L g189 ( 
.A(n_73),
.Y(n_189)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_35),
.Y(n_74)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_74),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_75),
.Y(n_183)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_33),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_76),
.Y(n_185)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_27),
.Y(n_77)
);

INVx3_ASAP7_75t_SL g138 ( 
.A(n_77),
.Y(n_138)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_33),
.Y(n_78)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_78),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_31),
.B(n_15),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_79),
.B(n_80),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_36),
.B(n_11),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_36),
.B(n_11),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_81),
.B(n_85),
.Y(n_162)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_26),
.Y(n_82)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_82),
.Y(n_133)
);

BUFx12_ASAP7_75t_L g83 ( 
.A(n_35),
.Y(n_83)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_83),
.Y(n_140)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_33),
.Y(n_84)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_84),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_37),
.B(n_13),
.Y(n_85)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_35),
.Y(n_86)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_86),
.Y(n_148)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_28),
.Y(n_87)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_87),
.Y(n_135)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_28),
.Y(n_88)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_88),
.Y(n_149)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_27),
.Y(n_89)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_89),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_37),
.B(n_0),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_90),
.B(n_112),
.Y(n_163)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_91),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_38),
.Y(n_92)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_92),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_43),
.B(n_0),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_38),
.Y(n_94)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_94),
.Y(n_142)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_51),
.Y(n_95)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_95),
.Y(n_156)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_29),
.Y(n_96)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_96),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_51),
.Y(n_97)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_97),
.Y(n_167)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_30),
.Y(n_98)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_98),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_28),
.Y(n_99)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_99),
.Y(n_186)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_25),
.Y(n_100)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_100),
.Y(n_154)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_40),
.Y(n_101)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_101),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_45),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_102),
.B(n_105),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_40),
.B(n_1),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_103),
.B(n_104),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_43),
.B(n_1),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_25),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g106 ( 
.A(n_50),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_106),
.B(n_110),
.Y(n_151)
);

INVx13_ASAP7_75t_L g107 ( 
.A(n_47),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_107),
.Y(n_125)
);

INVx11_ASAP7_75t_L g108 ( 
.A(n_35),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_108),
.Y(n_158)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_30),
.B(n_1),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_109),
.B(n_111),
.Y(n_144)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_40),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g111 ( 
.A(n_24),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_45),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_46),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_113),
.B(n_114),
.Y(n_145)
);

OR2x2_ASAP7_75t_L g114 ( 
.A(n_46),
.B(n_2),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_54),
.B(n_8),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_115),
.B(n_2),
.Y(n_169)
);

BUFx12f_ASAP7_75t_L g116 ( 
.A(n_28),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_116),
.B(n_41),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_103),
.B(n_53),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_126),
.B(n_159),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_56),
.A2(n_45),
.B1(n_52),
.B2(n_47),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_130),
.A2(n_137),
.B1(n_191),
.B2(n_189),
.Y(n_238)
);

OAI21xp33_ASAP7_75t_L g134 ( 
.A1(n_109),
.A2(n_53),
.B(n_48),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_134),
.B(n_151),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_61),
.A2(n_45),
.B1(n_52),
.B2(n_20),
.Y(n_137)
);

OAI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_65),
.A2(n_52),
.B1(n_20),
.B2(n_41),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_150),
.A2(n_155),
.B1(n_73),
.B2(n_102),
.Y(n_196)
);

OAI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_69),
.A2(n_52),
.B1(n_20),
.B2(n_41),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_157),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_114),
.B(n_54),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_89),
.B(n_34),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_160),
.B(n_164),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_78),
.A2(n_48),
.B1(n_49),
.B2(n_42),
.Y(n_161)
);

OA22x2_ASAP7_75t_L g212 ( 
.A1(n_161),
.A2(n_168),
.B1(n_170),
.B2(n_5),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_60),
.B(n_34),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_60),
.B(n_32),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_165),
.B(n_171),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_84),
.A2(n_48),
.B1(n_49),
.B2(n_42),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_169),
.B(n_176),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_91),
.A2(n_39),
.B1(n_44),
.B2(n_21),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_111),
.B(n_21),
.Y(n_171)
);

NOR2x1_ASAP7_75t_L g173 ( 
.A(n_95),
.B(n_39),
.Y(n_173)
);

OR2x2_ASAP7_75t_L g241 ( 
.A(n_173),
.B(n_179),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_111),
.B(n_44),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_175),
.B(n_188),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_70),
.B(n_32),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_75),
.B(n_18),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_177),
.B(n_182),
.Y(n_210)
);

NOR2x1_ASAP7_75t_L g179 ( 
.A(n_59),
.B(n_18),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_97),
.B(n_18),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_116),
.B(n_2),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_107),
.B(n_99),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_190),
.B(n_138),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_72),
.A2(n_35),
.B1(n_50),
.B2(n_7),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_129),
.B(n_116),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_192),
.B(n_204),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_137),
.A2(n_130),
.B1(n_163),
.B2(n_92),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_194),
.A2(n_200),
.B1(n_203),
.B2(n_211),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_134),
.B(n_87),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g273 ( 
.A(n_195),
.B(n_214),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_196),
.A2(n_201),
.B1(n_226),
.B2(n_231),
.Y(n_257)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_119),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g256 ( 
.A(n_197),
.Y(n_256)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_135),
.Y(n_198)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_198),
.Y(n_269)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_141),
.Y(n_199)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_199),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_170),
.A2(n_112),
.B1(n_94),
.B2(n_88),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_144),
.A2(n_66),
.B1(n_67),
.B2(n_58),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_117),
.Y(n_202)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_202),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_179),
.A2(n_83),
.B1(n_86),
.B2(n_108),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_147),
.B(n_5),
.Y(n_204)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_149),
.Y(n_205)
);

INVx4_ASAP7_75t_SL g301 ( 
.A(n_205),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_173),
.A2(n_83),
.B(n_35),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_206),
.A2(n_254),
.B(n_249),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_162),
.B(n_5),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_207),
.B(n_220),
.Y(n_276)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_142),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_208),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_117),
.A2(n_74),
.B1(n_6),
.B2(n_7),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g274 ( 
.A(n_212),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_124),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_213),
.B(n_222),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_153),
.B(n_5),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_150),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_215)
);

OR2x2_ASAP7_75t_L g267 ( 
.A(n_215),
.B(n_229),
.Y(n_267)
);

AOI21xp33_ASAP7_75t_L g216 ( 
.A1(n_139),
.A2(n_7),
.B(n_145),
.Y(n_216)
);

AOI32xp33_ASAP7_75t_L g279 ( 
.A1(n_216),
.A2(n_152),
.A3(n_174),
.B1(n_195),
.B2(n_214),
.Y(n_279)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_156),
.Y(n_217)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_217),
.Y(n_265)
);

INVx6_ASAP7_75t_L g218 ( 
.A(n_123),
.Y(n_218)
);

BUFx3_ASAP7_75t_L g298 ( 
.A(n_218),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_132),
.B(n_125),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_154),
.Y(n_221)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_221),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_118),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_181),
.B(n_184),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_224),
.B(n_227),
.Y(n_277)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_186),
.Y(n_225)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_225),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_L g226 ( 
.A1(n_155),
.A2(n_133),
.B1(n_121),
.B2(n_122),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_120),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_120),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_228),
.B(n_230),
.Y(n_278)
);

OA22x2_ASAP7_75t_L g229 ( 
.A1(n_161),
.A2(n_168),
.B1(n_149),
.B2(n_143),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_127),
.B(n_143),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_L g231 ( 
.A1(n_172),
.A2(n_158),
.B1(n_123),
.B2(n_131),
.Y(n_231)
);

INVx6_ASAP7_75t_L g233 ( 
.A(n_131),
.Y(n_233)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_233),
.Y(n_284)
);

INVx6_ASAP7_75t_L g234 ( 
.A(n_178),
.Y(n_234)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_234),
.Y(n_290)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_180),
.Y(n_235)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_235),
.Y(n_295)
);

BUFx2_ASAP7_75t_L g236 ( 
.A(n_180),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_236),
.Y(n_289)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_172),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_237),
.B(n_239),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_238),
.A2(n_174),
.B1(n_194),
.B2(n_200),
.Y(n_282)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_166),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_127),
.B(n_140),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_240),
.B(n_247),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_151),
.A2(n_185),
.B1(n_136),
.B2(n_140),
.Y(n_242)
);

OAI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_242),
.A2(n_215),
.B1(n_241),
.B2(n_223),
.Y(n_283)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_167),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_244),
.B(n_248),
.Y(n_266)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_128),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_245),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_166),
.Y(n_246)
);

INVx6_ASAP7_75t_L g261 ( 
.A(n_246),
.Y(n_261)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_187),
.Y(n_247)
);

INVx4_ASAP7_75t_L g248 ( 
.A(n_128),
.Y(n_248)
);

A2O1A1Ixp33_ASAP7_75t_L g292 ( 
.A1(n_249),
.A2(n_203),
.B(n_241),
.C(n_211),
.Y(n_292)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_187),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_250),
.B(n_251),
.Y(n_280)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_189),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_146),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_252),
.B(n_253),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_183),
.B(n_178),
.Y(n_253)
);

NAND2xp33_ASAP7_75t_SL g254 ( 
.A(n_183),
.B(n_185),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_255),
.B(n_193),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_210),
.B(n_138),
.C(n_148),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_260),
.B(n_288),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_263),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_196),
.A2(n_148),
.B1(n_146),
.B2(n_152),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_270),
.A2(n_282),
.B1(n_303),
.B2(n_236),
.Y(n_312)
);

FAx1_ASAP7_75t_SL g272 ( 
.A(n_249),
.B(n_174),
.CI(n_152),
.CON(n_272),
.SN(n_272)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_272),
.B(n_286),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_279),
.B(n_288),
.Y(n_320)
);

INVxp33_ASAP7_75t_L g338 ( 
.A(n_283),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_209),
.B(n_223),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_287),
.B(n_291),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_202),
.B(n_243),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_206),
.B(n_253),
.Y(n_291)
);

A2O1A1Ixp33_ASAP7_75t_L g330 ( 
.A1(n_292),
.A2(n_259),
.B(n_262),
.C(n_272),
.Y(n_330)
);

OAI22xp33_ASAP7_75t_SL g294 ( 
.A1(n_229),
.A2(n_212),
.B1(n_205),
.B2(n_221),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_L g325 ( 
.A1(n_294),
.A2(n_300),
.B1(n_257),
.B2(n_260),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_219),
.B(n_232),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_296),
.B(n_297),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_225),
.B(n_244),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_198),
.B(n_212),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_300),
.B(n_267),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_212),
.A2(n_229),
.B1(n_251),
.B2(n_250),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_280),
.Y(n_304)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_304),
.Y(n_342)
);

NOR2x1_ASAP7_75t_L g305 ( 
.A(n_291),
.B(n_229),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_SL g367 ( 
.A1(n_305),
.A2(n_307),
.B(n_329),
.Y(n_367)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_280),
.Y(n_306)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_306),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_263),
.A2(n_254),
.B(n_217),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_274),
.A2(n_239),
.B1(n_247),
.B2(n_218),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_308),
.A2(n_312),
.B1(n_314),
.B2(n_316),
.Y(n_347)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_297),
.Y(n_310)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_310),
.Y(n_356)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_301),
.Y(n_311)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_311),
.Y(n_354)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_266),
.Y(n_313)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_313),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_282),
.A2(n_199),
.B1(n_208),
.B2(n_246),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_268),
.A2(n_252),
.B1(n_235),
.B2(n_245),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_281),
.B(n_248),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g361 ( 
.A(n_318),
.B(n_321),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_268),
.A2(n_233),
.B1(n_234),
.B2(n_303),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_319),
.A2(n_325),
.B1(n_290),
.B2(n_295),
.Y(n_348)
);

NOR3xp33_ASAP7_75t_L g359 ( 
.A(n_320),
.B(n_330),
.C(n_335),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_281),
.B(n_287),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_273),
.B(n_296),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_323),
.B(n_324),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_273),
.B(n_278),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_326),
.B(n_332),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_267),
.A2(n_262),
.B1(n_292),
.B2(n_286),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_328),
.A2(n_301),
.B1(n_284),
.B2(n_289),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_264),
.A2(n_299),
.B(n_277),
.Y(n_329)
);

OAI22xp33_ASAP7_75t_SL g331 ( 
.A1(n_270),
.A2(n_276),
.B1(n_266),
.B2(n_256),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_331),
.A2(n_328),
.B1(n_313),
.B2(n_317),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_271),
.B(n_275),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_271),
.Y(n_333)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_333),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_293),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_334),
.B(n_337),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_258),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_256),
.B(n_295),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_336),
.B(n_285),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_261),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_SL g339 ( 
.A(n_272),
.B(n_275),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_SL g346 ( 
.A(n_339),
.B(n_265),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_324),
.A2(n_284),
.B1(n_290),
.B2(n_261),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_343),
.B(n_308),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_327),
.B(n_265),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_344),
.B(n_353),
.C(n_365),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_346),
.B(n_330),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_348),
.A2(n_304),
.B1(n_306),
.B2(n_318),
.Y(n_380)
);

NAND4xp25_ASAP7_75t_L g386 ( 
.A(n_349),
.B(n_352),
.C(n_311),
.D(n_333),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_319),
.A2(n_301),
.B1(n_298),
.B2(n_302),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_350),
.A2(n_312),
.B1(n_316),
.B2(n_314),
.Y(n_368)
);

NOR3xp33_ASAP7_75t_SL g352 ( 
.A(n_320),
.B(n_298),
.C(n_269),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_327),
.B(n_269),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_332),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_355),
.B(n_363),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_L g358 ( 
.A1(n_309),
.A2(n_285),
.B(n_305),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_SL g385 ( 
.A1(n_358),
.A2(n_364),
.B(n_307),
.Y(n_385)
);

CKINVDCx14_ASAP7_75t_R g384 ( 
.A(n_360),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_322),
.B(n_321),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_315),
.B(n_326),
.C(n_323),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_315),
.B(n_339),
.C(n_322),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_366),
.B(n_317),
.C(n_365),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_368),
.A2(n_369),
.B1(n_348),
.B2(n_342),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_364),
.A2(n_305),
.B1(n_338),
.B2(n_310),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_351),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_370),
.B(n_378),
.Y(n_392)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_371),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_355),
.B(n_335),
.Y(n_373)
);

CKINVDCx14_ASAP7_75t_R g403 ( 
.A(n_373),
.Y(n_403)
);

INVx2_ASAP7_75t_SL g374 ( 
.A(n_362),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_374),
.B(n_376),
.Y(n_396)
);

OA21x2_ASAP7_75t_L g376 ( 
.A1(n_358),
.A2(n_367),
.B(n_349),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_356),
.B(n_329),
.Y(n_377)
);

AOI22xp33_ASAP7_75t_L g394 ( 
.A1(n_377),
.A2(n_381),
.B1(n_388),
.B2(n_362),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_343),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_361),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_379),
.B(n_383),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_380),
.B(n_387),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_356),
.B(n_336),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_382),
.B(n_389),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_361),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_L g395 ( 
.A1(n_385),
.A2(n_367),
.B(n_357),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_386),
.B(n_359),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_357),
.B(n_337),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_354),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_SL g413 ( 
.A1(n_393),
.A2(n_395),
.B(n_406),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_394),
.B(n_401),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_375),
.B(n_353),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_397),
.B(n_400),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_375),
.B(n_344),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_373),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_402),
.A2(n_378),
.B1(n_345),
.B2(n_371),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_389),
.B(n_366),
.C(n_346),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_404),
.B(n_405),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_382),
.B(n_341),
.C(n_342),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_L g406 ( 
.A1(n_376),
.A2(n_340),
.B(n_345),
.Y(n_406)
);

AOI321xp33_ASAP7_75t_L g407 ( 
.A1(n_398),
.A2(n_379),
.A3(n_383),
.B1(n_372),
.B2(n_385),
.C(n_377),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_L g421 ( 
.A1(n_407),
.A2(n_414),
.B(n_406),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_L g409 ( 
.A1(n_396),
.A2(n_376),
.B(n_369),
.Y(n_409)
);

AOI21xp5_ASAP7_75t_SL g424 ( 
.A1(n_409),
.A2(n_395),
.B(n_391),
.Y(n_424)
);

OAI22x1_ASAP7_75t_L g411 ( 
.A1(n_396),
.A2(n_376),
.B1(n_380),
.B2(n_386),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_411),
.A2(n_415),
.B1(n_390),
.B2(n_402),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_SL g412 ( 
.A(n_398),
.B(n_370),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_412),
.B(n_392),
.Y(n_422)
);

OA21x2_ASAP7_75t_SL g414 ( 
.A1(n_391),
.A2(n_372),
.B(n_341),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_405),
.B(n_340),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_416),
.B(n_401),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_397),
.B(n_381),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_418),
.B(n_419),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_403),
.A2(n_384),
.B1(n_368),
.B2(n_352),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_SL g435 ( 
.A(n_420),
.B(n_423),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_421),
.A2(n_427),
.B1(n_419),
.B2(n_409),
.Y(n_433)
);

NOR3xp33_ASAP7_75t_L g431 ( 
.A(n_422),
.B(n_428),
.C(n_413),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_413),
.B(n_392),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_424),
.B(n_429),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_417),
.B(n_418),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_426),
.B(n_410),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_408),
.B(n_387),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_410),
.B(n_400),
.Y(n_429)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_427),
.Y(n_430)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_430),
.Y(n_438)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_431),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_425),
.B(n_417),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_432),
.B(n_436),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_433),
.B(n_425),
.Y(n_441)
);

OAI221xp5_ASAP7_75t_L g442 ( 
.A1(n_434),
.A2(n_399),
.B1(n_404),
.B2(n_390),
.C(n_388),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_SL g436 ( 
.A1(n_424),
.A2(n_411),
.B(n_407),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_437),
.B(n_429),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_439),
.B(n_435),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_441),
.B(n_442),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_438),
.B(n_437),
.C(n_440),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_445),
.B(n_446),
.C(n_447),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_L g447 ( 
.A1(n_443),
.A2(n_430),
.B1(n_415),
.B2(n_399),
.Y(n_447)
);

A2O1A1Ixp33_ASAP7_75t_SL g448 ( 
.A1(n_445),
.A2(n_440),
.B(n_444),
.C(n_374),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_448),
.B(n_354),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_449),
.A2(n_444),
.B1(n_374),
.B2(n_347),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_450),
.B(n_451),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_452),
.B(n_350),
.Y(n_453)
);


endmodule