module fake_jpeg_31873_n_152 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_152);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_152;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_2),
.B(n_7),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx4f_ASAP7_75t_SL g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx14_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_29),
.Y(n_30)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_21),
.B(n_5),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_34),
.B(n_35),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_15),
.B(n_0),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx4_ASAP7_75t_SL g37 ( 
.A(n_18),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_42),
.Y(n_59)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_28),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_53),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_15),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_60),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_54),
.B(n_6),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_31),
.A2(n_25),
.B1(n_19),
.B2(n_14),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_55),
.A2(n_62),
.B1(n_63),
.B2(n_1),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_30),
.B(n_27),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_56),
.B(n_59),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_24),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_38),
.A2(n_26),
.B1(n_16),
.B2(n_19),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_43),
.A2(n_26),
.B1(n_16),
.B2(n_27),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_41),
.B(n_14),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_64),
.B(n_3),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_42),
.B(n_26),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_70),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_35),
.B(n_16),
.Y(n_70)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_74),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_0),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_77),
.B(n_58),
.C(n_68),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_78),
.B(n_88),
.Y(n_95)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g105 ( 
.A(n_80),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_59),
.A2(n_1),
.B(n_3),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_82),
.Y(n_104)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_84),
.B(n_87),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_85),
.B(n_90),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_47),
.B(n_4),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_10),
.Y(n_108)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_60),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_89),
.B(n_91),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_52),
.B(n_5),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_52),
.B(n_46),
.Y(n_91)
);

INVxp67_ASAP7_75t_SL g97 ( 
.A(n_92),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_73),
.B(n_65),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_93),
.B(n_87),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_75),
.A2(n_62),
.B1(n_67),
.B2(n_72),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_94),
.A2(n_78),
.B1(n_81),
.B2(n_76),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_75),
.B(n_9),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_101),
.B(n_106),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_102),
.B(n_108),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_77),
.B(n_79),
.C(n_89),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_102),
.B(n_79),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_113),
.Y(n_128)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_103),
.Y(n_111)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_111),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_112),
.A2(n_114),
.B1(n_95),
.B2(n_106),
.Y(n_124)
);

INVxp67_ASAP7_75t_SL g113 ( 
.A(n_107),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g114 ( 
.A(n_96),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_98),
.A2(n_88),
.B(n_86),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_115),
.B(n_121),
.C(n_95),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_74),
.Y(n_117)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_117),
.Y(n_127)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_104),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_118),
.Y(n_126)
);

NOR3xp33_ASAP7_75t_L g122 ( 
.A(n_119),
.B(n_120),
.C(n_108),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_93),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_98),
.A2(n_82),
.B(n_84),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_122),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_123),
.B(n_109),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_124),
.B(n_129),
.Y(n_134)
);

NOR2x1_ASAP7_75t_L g129 ( 
.A(n_112),
.B(n_97),
.Y(n_129)
);

AOI322xp5_ASAP7_75t_SL g130 ( 
.A1(n_120),
.A2(n_99),
.A3(n_53),
.B1(n_68),
.B2(n_54),
.C1(n_105),
.C2(n_67),
.Y(n_130)
);

BUFx24_ASAP7_75t_SL g131 ( 
.A(n_130),
.Y(n_131)
);

BUFx24_ASAP7_75t_SL g132 ( 
.A(n_128),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_132),
.B(n_136),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_133),
.B(n_137),
.C(n_116),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_123),
.B(n_110),
.C(n_109),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_127),
.B(n_115),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_134),
.A2(n_121),
.B(n_119),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_138),
.A2(n_118),
.B(n_83),
.Y(n_145)
);

OAI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_135),
.A2(n_127),
.B1(n_129),
.B2(n_125),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_140),
.A2(n_142),
.B1(n_126),
.B2(n_125),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_141),
.B(n_111),
.Y(n_143)
);

OAI21xp33_ASAP7_75t_SL g142 ( 
.A1(n_131),
.A2(n_117),
.B(n_126),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_143),
.B(n_144),
.Y(n_146)
);

INVxp33_ASAP7_75t_L g147 ( 
.A(n_145),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_146),
.B(n_139),
.Y(n_148)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_148),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_147),
.A2(n_100),
.B(n_80),
.Y(n_149)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_150),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_149),
.Y(n_152)
);


endmodule