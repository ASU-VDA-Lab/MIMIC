module fake_jpeg_23_n_434 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_434);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_434;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx8_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx14_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx16f_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

BUFx4f_ASAP7_75t_SL g48 ( 
.A(n_13),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_49),
.Y(n_137)
);

BUFx4f_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx2_ASAP7_75t_SL g143 ( 
.A(n_50),
.Y(n_143)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_51),
.Y(n_118)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

BUFx10_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_53),
.Y(n_105)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

INVx11_ASAP7_75t_L g119 ( 
.A(n_54),
.Y(n_119)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_55),
.Y(n_124)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_56),
.Y(n_141)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_57),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_58),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_22),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_59),
.B(n_62),
.Y(n_104)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_60),
.Y(n_108)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_61),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_22),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_63),
.Y(n_112)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_64),
.Y(n_128)
);

AND2x2_ASAP7_75t_SL g65 ( 
.A(n_25),
.B(n_0),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_65),
.B(n_3),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_22),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_66),
.B(n_71),
.Y(n_123)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

INVx11_ASAP7_75t_L g135 ( 
.A(n_67),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_21),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_68),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_26),
.B(n_14),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_69),
.B(n_77),
.Y(n_102)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_17),
.Y(n_70)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_70),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_23),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_16),
.Y(n_72)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_72),
.Y(n_136)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_25),
.Y(n_73)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_73),
.Y(n_113)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_16),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_74),
.B(n_79),
.Y(n_138)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_20),
.Y(n_75)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_75),
.Y(n_115)
);

INVx6_ASAP7_75t_SL g76 ( 
.A(n_48),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g134 ( 
.A(n_76),
.B(n_37),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_26),
.B(n_0),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_24),
.B(n_2),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_78),
.B(n_81),
.Y(n_103)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_28),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_23),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_80),
.B(n_85),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_27),
.B(n_2),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_29),
.Y(n_82)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_82),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_27),
.B(n_2),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_83),
.B(n_97),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_29),
.Y(n_84)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_84),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_35),
.B(n_2),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_29),
.Y(n_86)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_86),
.Y(n_130)
);

INVx13_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

INVx11_ASAP7_75t_L g154 ( 
.A(n_87),
.Y(n_154)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_28),
.Y(n_88)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_88),
.Y(n_110)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_18),
.Y(n_89)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_89),
.Y(n_144)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_25),
.Y(n_90)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_90),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_30),
.Y(n_91)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_19),
.Y(n_92)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_92),
.Y(n_117)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_15),
.Y(n_93)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_93),
.Y(n_120)
);

BUFx10_ASAP7_75t_L g94 ( 
.A(n_25),
.Y(n_94)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_94),
.Y(n_121)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_95),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_30),
.Y(n_96)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_96),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_35),
.B(n_13),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_48),
.Y(n_98)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_98),
.Y(n_145)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_32),
.Y(n_99)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_99),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_49),
.A2(n_23),
.B1(n_41),
.B2(n_30),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_100),
.A2(n_116),
.B1(n_139),
.B2(n_153),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_106),
.B(n_50),
.Y(n_159)
);

OAI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_96),
.A2(n_41),
.B1(n_15),
.B2(n_37),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_58),
.A2(n_41),
.B1(n_45),
.B2(n_44),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_125),
.A2(n_126),
.B1(n_146),
.B2(n_92),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_68),
.A2(n_86),
.B1(n_84),
.B2(n_82),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_63),
.A2(n_47),
.B1(n_40),
.B2(n_37),
.Y(n_132)
);

OA22x2_ASAP7_75t_L g166 ( 
.A1(n_132),
.A2(n_147),
.B1(n_89),
.B2(n_60),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_134),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_91),
.A2(n_15),
.B1(n_47),
.B2(n_40),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_76),
.B(n_32),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_140),
.B(n_142),
.Y(n_167)
);

OR2x2_ASAP7_75t_L g142 ( 
.A(n_70),
.B(n_33),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_51),
.A2(n_55),
.B1(n_93),
.B2(n_73),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_63),
.A2(n_47),
.B1(n_40),
.B2(n_33),
.Y(n_147)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_90),
.Y(n_150)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_150),
.Y(n_164)
);

OAI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_65),
.A2(n_39),
.B1(n_45),
.B2(n_44),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_138),
.B(n_57),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_156),
.B(n_169),
.Y(n_209)
);

OAI32xp33_ASAP7_75t_L g157 ( 
.A1(n_103),
.A2(n_65),
.A3(n_36),
.B1(n_34),
.B2(n_39),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_157),
.B(n_159),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_115),
.A2(n_54),
.B1(n_67),
.B2(n_34),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_158),
.Y(n_215)
);

INVx11_ASAP7_75t_L g160 ( 
.A(n_119),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_160),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_104),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_161),
.B(n_162),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_133),
.B(n_50),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_163),
.A2(n_166),
.B1(n_184),
.B2(n_191),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g165 ( 
.A(n_113),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_165),
.Y(n_234)
);

BUFx2_ASAP7_75t_L g168 ( 
.A(n_143),
.Y(n_168)
);

CKINVDCx14_ASAP7_75t_R g202 ( 
.A(n_168),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_129),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_110),
.Y(n_170)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_170),
.Y(n_206)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_149),
.Y(n_171)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_171),
.Y(n_214)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_112),
.Y(n_172)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_172),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_106),
.B(n_56),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_173),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_123),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_174),
.B(n_178),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_153),
.B(n_36),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_175),
.B(n_180),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_126),
.A2(n_94),
.B1(n_87),
.B2(n_52),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_176),
.A2(n_199),
.B1(n_101),
.B2(n_11),
.Y(n_229)
);

BUFx12_ASAP7_75t_L g177 ( 
.A(n_101),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_177),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_102),
.B(n_52),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_116),
.A2(n_94),
.B1(n_75),
.B2(n_46),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_179),
.A2(n_154),
.B1(n_119),
.B2(n_135),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_142),
.B(n_3),
.Y(n_180)
);

OR2x2_ASAP7_75t_L g181 ( 
.A(n_148),
.B(n_95),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_181),
.B(n_186),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_121),
.Y(n_182)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_182),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_134),
.B(n_5),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_183),
.B(n_188),
.Y(n_211)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_113),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_137),
.Y(n_185)
);

INVx6_ASAP7_75t_L g210 ( 
.A(n_185),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_122),
.Y(n_186)
);

OA22x2_ASAP7_75t_L g187 ( 
.A1(n_132),
.A2(n_125),
.B1(n_147),
.B2(n_130),
.Y(n_187)
);

AOI22x1_ASAP7_75t_L g213 ( 
.A1(n_187),
.A2(n_166),
.B1(n_199),
.B2(n_176),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_109),
.B(n_7),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_127),
.B(n_8),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_190),
.A2(n_144),
.B1(n_120),
.B2(n_155),
.Y(n_216)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_111),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_136),
.B(n_9),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_192),
.B(n_196),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_117),
.A2(n_46),
.B1(n_42),
.B2(n_19),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_194),
.A2(n_195),
.B1(n_198),
.B2(n_154),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_115),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_128),
.B(n_9),
.Y(n_196)
);

INVx6_ASAP7_75t_L g197 ( 
.A(n_137),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_197),
.B(n_10),
.Y(n_235)
);

BUFx2_ASAP7_75t_L g198 ( 
.A(n_143),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_131),
.A2(n_42),
.B1(n_11),
.B2(n_12),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_183),
.A2(n_108),
.B(n_144),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_200),
.A2(n_223),
.B(n_198),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_189),
.A2(n_124),
.B1(n_118),
.B2(n_151),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_201),
.A2(n_213),
.B1(n_219),
.B2(n_221),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_193),
.A2(n_175),
.B1(n_180),
.B2(n_167),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_203),
.A2(n_204),
.B1(n_164),
.B2(n_170),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_193),
.A2(n_105),
.B1(n_107),
.B2(n_130),
.Y(n_204)
);

FAx1_ASAP7_75t_SL g207 ( 
.A(n_162),
.B(n_145),
.CI(n_108),
.CON(n_207),
.SN(n_207)
);

OAI32xp33_ASAP7_75t_L g257 ( 
.A1(n_207),
.A2(n_164),
.A3(n_171),
.B1(n_169),
.B2(n_182),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_208),
.A2(n_160),
.B1(n_198),
.B2(n_168),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_216),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_178),
.A2(n_107),
.B1(n_114),
.B2(n_141),
.Y(n_219)
);

INVxp33_ASAP7_75t_L g263 ( 
.A(n_220),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_187),
.A2(n_114),
.B1(n_152),
.B2(n_135),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_183),
.A2(n_181),
.B(n_159),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_187),
.A2(n_152),
.B1(n_101),
.B2(n_12),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_226),
.A2(n_229),
.B1(n_194),
.B2(n_173),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_173),
.B(n_13),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_233),
.B(n_159),
.Y(n_236)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_235),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_236),
.B(n_233),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_203),
.B(n_188),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_237),
.B(n_240),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_239),
.A2(n_249),
.B1(n_251),
.B2(n_258),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_207),
.B(n_188),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_228),
.A2(n_166),
.B(n_187),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_241),
.A2(n_244),
.B(n_257),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_207),
.B(n_157),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_242),
.B(n_254),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_202),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_243),
.B(n_253),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_215),
.A2(n_166),
.B(n_195),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_200),
.Y(n_246)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_246),
.Y(n_267)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_206),
.Y(n_247)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_247),
.Y(n_275)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_206),
.Y(n_248)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_248),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_205),
.A2(n_163),
.B1(n_186),
.B2(n_174),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_224),
.A2(n_161),
.B1(n_197),
.B2(n_191),
.Y(n_251)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_252),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_209),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_211),
.B(n_192),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_214),
.Y(n_255)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_255),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_256),
.B(n_204),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_213),
.A2(n_185),
.B1(n_184),
.B2(n_172),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_210),
.Y(n_259)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_259),
.Y(n_273)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_210),
.Y(n_260)
);

INVx2_ASAP7_75t_SL g276 ( 
.A(n_260),
.Y(n_276)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_214),
.Y(n_261)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_261),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_262),
.A2(n_246),
.B(n_241),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_228),
.Y(n_264)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_264),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_268),
.B(n_257),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_264),
.A2(n_224),
.B1(n_213),
.B2(n_229),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_271),
.A2(n_238),
.B1(n_239),
.B2(n_244),
.Y(n_306)
);

O2A1O1Ixp33_ASAP7_75t_L g272 ( 
.A1(n_240),
.A2(n_221),
.B(n_226),
.C(n_215),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_272),
.B(n_291),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_274),
.A2(n_280),
.B(n_282),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_251),
.B(n_218),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_278),
.B(n_222),
.Y(n_307)
);

A2O1A1O1Ixp25_ASAP7_75t_L g282 ( 
.A1(n_237),
.A2(n_224),
.B(n_222),
.C(n_227),
.D(n_223),
.Y(n_282)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_247),
.Y(n_285)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_285),
.Y(n_296)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_248),
.Y(n_286)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_286),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_255),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_288),
.B(n_234),
.Y(n_315)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_261),
.Y(n_289)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_289),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_236),
.B(n_211),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_290),
.B(n_245),
.C(n_236),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_245),
.B(n_235),
.Y(n_291)
);

CKINVDCx14_ASAP7_75t_R g292 ( 
.A(n_277),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_292),
.A2(n_297),
.B1(n_306),
.B2(n_307),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_270),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_294),
.B(n_304),
.Y(n_322)
);

OR2x2_ASAP7_75t_L g295 ( 
.A(n_274),
.B(n_242),
.Y(n_295)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_295),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_284),
.A2(n_258),
.B1(n_238),
.B2(n_256),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_284),
.A2(n_269),
.B1(n_283),
.B2(n_265),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_298),
.A2(n_267),
.B1(n_291),
.B2(n_281),
.Y(n_319)
);

AOI21xp33_ASAP7_75t_L g299 ( 
.A1(n_265),
.A2(n_262),
.B(n_254),
.Y(n_299)
);

CKINVDCx14_ASAP7_75t_R g335 ( 
.A(n_299),
.Y(n_335)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_273),
.Y(n_300)
);

INVx1_ASAP7_75t_SL g328 ( 
.A(n_300),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_303),
.B(n_305),
.C(n_311),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_270),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_290),
.B(n_230),
.C(n_249),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_283),
.B(n_243),
.Y(n_308)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_308),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_279),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_309),
.B(n_313),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_SL g317 ( 
.A(n_310),
.B(n_266),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_268),
.B(n_256),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_279),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_269),
.A2(n_244),
.B(n_250),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_314),
.A2(n_216),
.B(n_219),
.Y(n_331)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_315),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_266),
.B(n_231),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_316),
.B(n_267),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_317),
.B(n_321),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_306),
.A2(n_272),
.B1(n_280),
.B2(n_271),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_318),
.B(n_330),
.Y(n_344)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_319),
.Y(n_346)
);

INVx4_ASAP7_75t_L g320 ( 
.A(n_300),
.Y(n_320)
);

INVx1_ASAP7_75t_SL g361 ( 
.A(n_320),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_303),
.B(n_282),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_323),
.B(n_310),
.C(n_293),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_298),
.A2(n_263),
.B1(n_289),
.B2(n_286),
.Y(n_324)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_324),
.Y(n_349)
);

XNOR2x1_ASAP7_75t_L g325 ( 
.A(n_311),
.B(n_287),
.Y(n_325)
);

XNOR2x1_ASAP7_75t_L g342 ( 
.A(n_325),
.B(n_305),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_308),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_329),
.B(n_338),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_302),
.A2(n_285),
.B1(n_275),
.B2(n_252),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g352 ( 
.A1(n_331),
.A2(n_314),
.B(n_293),
.Y(n_352)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_296),
.Y(n_333)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_333),
.Y(n_348)
);

INVxp33_ASAP7_75t_L g334 ( 
.A(n_302),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_334),
.B(n_304),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g338 ( 
.A(n_295),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_296),
.Y(n_339)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_339),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_342),
.B(n_324),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_327),
.B(n_307),
.Y(n_343)
);

NAND3xp33_ASAP7_75t_L g373 ( 
.A(n_343),
.B(n_355),
.C(n_357),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_345),
.B(n_337),
.Y(n_364)
);

BUFx24_ASAP7_75t_SL g347 ( 
.A(n_335),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_347),
.B(n_317),
.Y(n_366)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_322),
.Y(n_350)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_350),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_351),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_352),
.B(n_356),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_322),
.B(n_313),
.Y(n_354)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_354),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_326),
.B(n_316),
.Y(n_355)
);

NOR3xp33_ASAP7_75t_SL g356 ( 
.A(n_336),
.B(n_295),
.C(n_231),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_SL g357 ( 
.A(n_323),
.B(n_337),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_332),
.Y(n_358)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_358),
.Y(n_377)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_332),
.Y(n_359)
);

AOI22x1_ASAP7_75t_L g363 ( 
.A1(n_359),
.A2(n_340),
.B1(n_330),
.B2(n_318),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_346),
.A2(n_334),
.B1(n_336),
.B2(n_319),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_362),
.A2(n_351),
.B1(n_341),
.B2(n_297),
.Y(n_383)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_363),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_364),
.B(n_368),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_366),
.B(n_367),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_345),
.B(n_325),
.C(n_321),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_360),
.B(n_328),
.C(n_301),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_369),
.B(n_371),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_360),
.B(n_352),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_342),
.B(n_328),
.C(n_301),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_372),
.B(n_374),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_348),
.B(n_294),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_346),
.B(n_331),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_378),
.B(n_359),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_379),
.B(n_381),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_376),
.A2(n_358),
.B1(n_350),
.B2(n_349),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_380),
.A2(n_377),
.B1(n_375),
.B2(n_378),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_369),
.B(n_349),
.C(n_344),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_372),
.B(n_344),
.C(n_354),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_382),
.B(n_386),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_383),
.B(n_363),
.Y(n_395)
);

A2O1A1Ixp33_ASAP7_75t_SL g384 ( 
.A1(n_362),
.A2(n_356),
.B(n_312),
.C(n_309),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_384),
.A2(n_390),
.B1(n_276),
.B2(n_259),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_365),
.B(n_353),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_364),
.B(n_361),
.C(n_312),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_388),
.B(n_273),
.Y(n_401)
);

AOI22xp33_ASAP7_75t_SL g390 ( 
.A1(n_370),
.A2(n_361),
.B1(n_320),
.B2(n_276),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_388),
.B(n_367),
.C(n_368),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_393),
.B(n_396),
.Y(n_410)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_394),
.Y(n_405)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_395),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_381),
.B(n_373),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_387),
.B(n_371),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_397),
.B(n_399),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_382),
.B(n_260),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_401),
.B(n_402),
.C(n_384),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_391),
.B(n_389),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_403),
.A2(n_404),
.B1(n_384),
.B2(n_398),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_392),
.A2(n_276),
.B(n_212),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_393),
.B(n_385),
.C(n_390),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_406),
.B(n_407),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_400),
.B(n_384),
.C(n_232),
.Y(n_407)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_411),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_412),
.Y(n_416)
);

XNOR2x1_ASAP7_75t_SL g413 ( 
.A(n_395),
.B(n_208),
.Y(n_413)
);

OAI21x1_ASAP7_75t_L g418 ( 
.A1(n_413),
.A2(n_225),
.B(n_212),
.Y(n_418)
);

XOR2x2_ASAP7_75t_SL g414 ( 
.A(n_403),
.B(n_225),
.Y(n_414)
);

A2O1A1Ixp33_ASAP7_75t_SL g420 ( 
.A1(n_414),
.A2(n_217),
.B(n_177),
.C(n_234),
.Y(n_420)
);

NOR2x1_ASAP7_75t_L g417 ( 
.A(n_410),
.B(n_232),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_417),
.B(n_419),
.Y(n_422)
);

NAND2xp33_ASAP7_75t_SL g423 ( 
.A(n_418),
.B(n_407),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_409),
.B(n_232),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_L g426 ( 
.A1(n_420),
.A2(n_177),
.B(n_10),
.Y(n_426)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_423),
.Y(n_428)
);

OAI321xp33_ASAP7_75t_L g424 ( 
.A1(n_421),
.A2(n_408),
.A3(n_405),
.B1(n_414),
.B2(n_413),
.C(n_406),
.Y(n_424)
);

NAND3xp33_ASAP7_75t_L g427 ( 
.A(n_424),
.B(n_425),
.C(n_426),
.Y(n_427)
);

AOI31xp33_ASAP7_75t_L g425 ( 
.A1(n_415),
.A2(n_217),
.A3(n_177),
.B(n_11),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_422),
.B(n_416),
.C(n_420),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_429),
.B(n_10),
.C(n_428),
.Y(n_430)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_430),
.Y(n_432)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_427),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_432),
.B(n_431),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_433),
.B(n_10),
.Y(n_434)
);


endmodule