module fake_jpeg_3916_n_275 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_275);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_275;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_149;
wire n_48;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_140;
wire n_128;
wire n_82;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_8),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx4f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx2_ASAP7_75t_SL g31 ( 
.A(n_25),
.Y(n_31)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

INVx4_ASAP7_75t_SL g32 ( 
.A(n_25),
.Y(n_32)
);

HAxp5_ASAP7_75t_SL g51 ( 
.A(n_32),
.B(n_35),
.CON(n_51),
.SN(n_51)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_13),
.B(n_12),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_36),
.A2(n_22),
.B1(n_20),
.B2(n_24),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_36),
.A2(n_22),
.B1(n_26),
.B2(n_23),
.Y(n_38)
);

OAI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_38),
.A2(n_50),
.B1(n_53),
.B2(n_14),
.Y(n_73)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_40),
.B(n_31),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_41),
.Y(n_54)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_27),
.C(n_26),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_43),
.B(n_35),
.Y(n_72)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_36),
.A2(n_22),
.B1(n_27),
.B2(n_14),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_30),
.A2(n_19),
.B1(n_16),
.B2(n_23),
.Y(n_53)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_55),
.B(n_56),
.Y(n_80)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_47),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_57),
.B(n_58),
.Y(n_84)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_59),
.Y(n_93)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_40),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_60),
.B(n_62),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

CKINVDCx14_ASAP7_75t_R g63 ( 
.A(n_43),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_63),
.B(n_64),
.Y(n_87)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

AND2x2_ASAP7_75t_SL g66 ( 
.A(n_51),
.B(n_31),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_31),
.C(n_20),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_20),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_68),
.B(n_71),
.Y(n_92)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_69),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_52),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_72),
.A2(n_14),
.B(n_13),
.Y(n_81)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_73),
.Y(n_78)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_76),
.B(n_77),
.Y(n_97)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_85),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_81),
.B(n_60),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_83),
.B(n_71),
.C(n_24),
.Y(n_105)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_86),
.B(n_89),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_62),
.A2(n_46),
.B1(n_34),
.B2(n_33),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_88),
.A2(n_94),
.B1(n_54),
.B2(n_66),
.Y(n_96)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_70),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_44),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_64),
.A2(n_54),
.B1(n_66),
.B2(n_72),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_96),
.A2(n_112),
.B1(n_46),
.B2(n_70),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_74),
.A2(n_57),
.B1(n_65),
.B2(n_45),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_98),
.A2(n_75),
.B1(n_77),
.B2(n_85),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_87),
.B(n_92),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_99),
.B(n_100),
.Y(n_136)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_84),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_101),
.B(n_103),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_90),
.B(n_68),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_102),
.A2(n_104),
.B(n_115),
.Y(n_135)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_81),
.B(n_69),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_105),
.B(n_17),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_16),
.Y(n_131)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_108),
.Y(n_118)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_83),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_109),
.B(n_113),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_110),
.B(n_65),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_78),
.B(n_59),
.C(n_29),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_111),
.B(n_114),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_91),
.A2(n_46),
.B1(n_45),
.B2(n_39),
.Y(n_112)
);

OA21x2_ASAP7_75t_L g113 ( 
.A1(n_86),
.A2(n_33),
.B(n_34),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_59),
.C(n_29),
.Y(n_114)
);

O2A1O1Ixp33_ASAP7_75t_L g115 ( 
.A1(n_76),
.A2(n_33),
.B(n_34),
.C(n_37),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_116),
.A2(n_131),
.B(n_102),
.Y(n_142)
);

INVx1_ASAP7_75t_SL g117 ( 
.A(n_107),
.Y(n_117)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_117),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_119),
.B(n_122),
.Y(n_152)
);

INVx2_ASAP7_75t_SL g121 ( 
.A(n_113),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_121),
.B(n_132),
.Y(n_140)
);

NOR2xp67_ASAP7_75t_L g122 ( 
.A(n_96),
.B(n_59),
.Y(n_122)
);

BUFx2_ASAP7_75t_L g123 ( 
.A(n_95),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_123),
.B(n_128),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_125),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_106),
.B(n_28),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_126),
.B(n_127),
.C(n_133),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_99),
.B(n_28),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_107),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_129),
.B(n_126),
.Y(n_159)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_97),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_105),
.B(n_28),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_104),
.B(n_29),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_134),
.B(n_112),
.C(n_115),
.Y(n_155)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_95),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_137),
.B(n_89),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_135),
.A2(n_109),
.B(n_100),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_141),
.A2(n_154),
.B(n_156),
.Y(n_168)
);

NOR3xp33_ASAP7_75t_SL g182 ( 
.A(n_142),
.B(n_15),
.C(n_17),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_119),
.A2(n_111),
.B1(n_101),
.B2(n_103),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_143),
.A2(n_150),
.B1(n_158),
.B2(n_18),
.Y(n_178)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_136),
.Y(n_145)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_145),
.Y(n_176)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_120),
.Y(n_146)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_146),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_123),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_147),
.Y(n_167)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_127),
.Y(n_148)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_148),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_149),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_130),
.A2(n_45),
.B1(n_39),
.B2(n_113),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_118),
.B(n_113),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_151),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_135),
.A2(n_114),
.B(n_108),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_155),
.B(n_159),
.C(n_124),
.Y(n_164)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_128),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_134),
.B(n_75),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_157),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_121),
.A2(n_79),
.B1(n_115),
.B2(n_19),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_131),
.A2(n_16),
.B(n_19),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_160),
.B(n_133),
.Y(n_163)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_117),
.Y(n_161)
);

NOR3xp33_ASAP7_75t_L g177 ( 
.A(n_161),
.B(n_24),
.C(n_18),
.Y(n_177)
);

XNOR2x1_ASAP7_75t_SL g162 ( 
.A(n_141),
.B(n_131),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g191 ( 
.A(n_162),
.B(n_150),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_163),
.B(n_157),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_164),
.B(n_172),
.C(n_173),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_146),
.B(n_124),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_165),
.B(n_178),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_155),
.B(n_129),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_171),
.A2(n_139),
.B1(n_143),
.B2(n_140),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_144),
.B(n_121),
.C(n_37),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_144),
.B(n_37),
.C(n_39),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_149),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_174),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_141),
.B(n_15),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_175),
.B(n_179),
.Y(n_200)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_177),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_154),
.A2(n_13),
.B(n_18),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_138),
.A2(n_82),
.B1(n_15),
.B2(n_48),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_181),
.A2(n_161),
.B1(n_139),
.B2(n_140),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_182),
.B(n_151),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_148),
.B(n_48),
.C(n_82),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_184),
.B(n_153),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_185),
.B(n_15),
.C(n_17),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_162),
.A2(n_145),
.B1(n_147),
.B2(n_152),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_186),
.A2(n_191),
.B(n_171),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_187),
.B(n_182),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_181),
.Y(n_189)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_189),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_180),
.B(n_160),
.Y(n_192)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_192),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_178),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_194),
.B(n_198),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_176),
.B(n_142),
.Y(n_195)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_195),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_196),
.B(n_163),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_197),
.B(n_199),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_167),
.B(n_156),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_184),
.Y(n_202)
);

BUFx2_ASAP7_75t_L g206 ( 
.A(n_202),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_168),
.A2(n_158),
.B1(n_48),
.B2(n_15),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_203),
.A2(n_168),
.B1(n_183),
.B2(n_166),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_196),
.A2(n_195),
.B1(n_189),
.B2(n_169),
.Y(n_204)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_204),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_205),
.A2(n_211),
.B(n_215),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_201),
.A2(n_175),
.B1(n_170),
.B2(n_172),
.Y(n_207)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_207),
.Y(n_230)
);

XOR2x2_ASAP7_75t_L g222 ( 
.A(n_208),
.B(n_209),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_186),
.A2(n_164),
.B1(n_173),
.B2(n_171),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_210),
.B(n_198),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_190),
.B(n_179),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_212),
.B(n_217),
.C(n_218),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_191),
.A2(n_0),
.B(n_1),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_190),
.B(n_15),
.C(n_17),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_220),
.A2(n_187),
.B(n_203),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_223),
.A2(n_227),
.B(n_232),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_219),
.B(n_188),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_225),
.B(n_209),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_216),
.B(n_193),
.Y(n_226)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_226),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_205),
.B(n_200),
.Y(n_229)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_229),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g231 ( 
.A(n_206),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_231),
.B(n_1),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_213),
.B(n_200),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_208),
.B(n_17),
.C(n_1),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_233),
.B(n_217),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_214),
.B(n_0),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_234),
.B(n_215),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_222),
.B(n_211),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_235),
.B(n_17),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_236),
.B(n_243),
.Y(n_248)
);

OR2x2_ASAP7_75t_L g239 ( 
.A(n_222),
.B(n_223),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_239),
.B(n_240),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_228),
.B(n_206),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_241),
.A2(n_246),
.B(n_245),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_230),
.A2(n_209),
.B1(n_218),
.B2(n_212),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_242),
.B(n_244),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_233),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_246),
.B(n_238),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_237),
.B(n_224),
.C(n_221),
.Y(n_247)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_247),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_249),
.B(n_254),
.Y(n_258)
);

AOI21x1_ASAP7_75t_L g251 ( 
.A1(n_239),
.A2(n_221),
.B(n_224),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_251),
.A2(n_253),
.B(n_11),
.Y(n_259)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_252),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_235),
.B(n_2),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_238),
.B(n_12),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_256),
.B(n_3),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_248),
.B(n_12),
.Y(n_257)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_257),
.Y(n_265)
);

NAND3xp33_ASAP7_75t_L g268 ( 
.A(n_259),
.B(n_262),
.C(n_9),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_255),
.B(n_11),
.Y(n_260)
);

A2O1A1Ixp33_ASAP7_75t_SL g264 ( 
.A1(n_260),
.A2(n_250),
.B(n_247),
.C(n_8),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_264),
.A2(n_267),
.B(n_258),
.Y(n_270)
);

OAI21x1_ASAP7_75t_L g266 ( 
.A1(n_259),
.A2(n_252),
.B(n_9),
.Y(n_266)
);

NOR3xp33_ASAP7_75t_SL g269 ( 
.A(n_266),
.B(n_268),
.C(n_3),
.Y(n_269)
);

AO221x1_ASAP7_75t_L g267 ( 
.A1(n_261),
.A2(n_9),
.B1(n_4),
.B2(n_5),
.C(n_6),
.Y(n_267)
);

OAI221xp5_ASAP7_75t_L g271 ( 
.A1(n_269),
.A2(n_265),
.B1(n_4),
.B2(n_5),
.C(n_6),
.Y(n_271)
);

A2O1A1Ixp33_ASAP7_75t_L g272 ( 
.A1(n_270),
.A2(n_263),
.B(n_4),
.C(n_5),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_271),
.A2(n_272),
.B(n_3),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_273),
.B(n_6),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_274),
.B(n_6),
.Y(n_275)
);


endmodule