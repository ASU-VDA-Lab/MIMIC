module fake_jpeg_9715_n_253 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_253);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_253;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

BUFx3_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx24_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx4f_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx24_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx5_ASAP7_75t_SL g59 ( 
.A(n_36),
.Y(n_59)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_37),
.B(n_42),
.Y(n_60)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_27),
.B(n_0),
.Y(n_39)
);

OAI21xp33_ASAP7_75t_L g56 ( 
.A1(n_39),
.A2(n_40),
.B(n_1),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_14),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_45),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

BUFx24_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_38),
.A2(n_32),
.B1(n_25),
.B2(n_20),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_48),
.A2(n_52),
.B1(n_64),
.B2(n_73),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_38),
.A2(n_22),
.B1(n_32),
.B2(n_20),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_49),
.A2(n_50),
.B1(n_53),
.B2(n_21),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_L g50 ( 
.A1(n_46),
.A2(n_32),
.B1(n_25),
.B2(n_22),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_51),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_46),
.A2(n_25),
.B1(n_20),
.B2(n_22),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_L g53 ( 
.A1(n_42),
.A2(n_23),
.B1(n_21),
.B2(n_19),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_19),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_54),
.B(n_57),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_56),
.B(n_58),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_24),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_27),
.Y(n_58)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_62),
.B(n_66),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_63),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_41),
.A2(n_33),
.B1(n_23),
.B2(n_21),
.Y(n_64)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_31),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_67),
.B(n_72),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_36),
.B(n_24),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_69),
.B(n_47),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_36),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_41),
.A2(n_33),
.B1(n_30),
.B2(n_35),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_36),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_74),
.B(n_75),
.Y(n_100)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_54),
.A2(n_21),
.B1(n_28),
.B2(n_31),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_76),
.A2(n_86),
.B1(n_105),
.B2(n_106),
.Y(n_112)
);

OAI21xp33_ASAP7_75t_L g77 ( 
.A1(n_57),
.A2(n_1),
.B(n_2),
.Y(n_77)
);

NAND3xp33_ASAP7_75t_L g129 ( 
.A(n_77),
.B(n_92),
.C(n_107),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_74),
.Y(n_79)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_79),
.Y(n_109)
);

BUFx2_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_81),
.Y(n_124)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_82),
.B(n_87),
.Y(n_130)
);

OA22x2_ASAP7_75t_L g84 ( 
.A1(n_72),
.A2(n_71),
.B1(n_53),
.B2(n_50),
.Y(n_84)
);

OA22x2_ASAP7_75t_L g118 ( 
.A1(n_84),
.A2(n_68),
.B1(n_55),
.B2(n_18),
.Y(n_118)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_85),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_49),
.A2(n_21),
.B1(n_35),
.B2(n_30),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_64),
.Y(n_87)
);

AND2x2_ASAP7_75t_SL g89 ( 
.A(n_69),
.B(n_47),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_89),
.B(n_104),
.Y(n_116)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_90),
.B(n_94),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_58),
.B(n_47),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_60),
.A2(n_18),
.B(n_47),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_93),
.Y(n_126)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_51),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_51),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_95),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_59),
.Y(n_97)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_97),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_98),
.B(n_65),
.Y(n_114)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_55),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_101),
.A2(n_102),
.B1(n_5),
.B2(n_6),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_70),
.A2(n_28),
.B1(n_34),
.B2(n_26),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_61),
.B(n_34),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_103),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_66),
.B(n_26),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_70),
.A2(n_26),
.B1(n_24),
.B2(n_17),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_65),
.A2(n_26),
.B1(n_24),
.B2(n_17),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_59),
.B(n_36),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_75),
.B(n_68),
.Y(n_108)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_108),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_87),
.A2(n_83),
.B1(n_84),
.B2(n_85),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_110),
.A2(n_118),
.B1(n_123),
.B2(n_134),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_114),
.B(n_121),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_78),
.B(n_17),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_115),
.B(n_98),
.Y(n_140)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_104),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_120),
.B(n_128),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_78),
.B(n_18),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_80),
.B(n_1),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_122),
.B(n_125),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_84),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_123)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_86),
.B(n_13),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_127),
.Y(n_148)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_91),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_81),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_133),
.B(n_90),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_84),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_113),
.A2(n_92),
.B1(n_101),
.B2(n_89),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_135),
.Y(n_180)
);

INVxp33_ASAP7_75t_SL g137 ( 
.A(n_133),
.Y(n_137)
);

OA22x2_ASAP7_75t_L g167 ( 
.A1(n_137),
.A2(n_117),
.B1(n_109),
.B2(n_118),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_111),
.A2(n_113),
.B1(n_82),
.B2(n_96),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_138),
.A2(n_141),
.B(n_146),
.Y(n_165)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_131),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_139),
.B(n_142),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_140),
.B(n_119),
.C(n_112),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_114),
.B(n_89),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_131),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_110),
.A2(n_96),
.B1(n_94),
.B2(n_95),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_143),
.A2(n_117),
.B1(n_124),
.B2(n_128),
.Y(n_161)
);

OAI21xp33_ASAP7_75t_SL g145 ( 
.A1(n_123),
.A2(n_92),
.B(n_93),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_145),
.B(n_118),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_120),
.B(n_107),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_130),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_147),
.B(n_151),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_115),
.B(n_107),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_149),
.A2(n_157),
.B(n_160),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_122),
.Y(n_151)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_152),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_121),
.B(n_76),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_154),
.B(n_125),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_111),
.B(n_100),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_155),
.B(n_156),
.Y(n_164)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_116),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_126),
.A2(n_88),
.B(n_97),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_116),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_158),
.B(n_159),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_119),
.B(n_6),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_129),
.A2(n_79),
.B(n_8),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_161),
.A2(n_142),
.B1(n_148),
.B2(n_143),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_135),
.A2(n_118),
.B1(n_134),
.B2(n_112),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_163),
.A2(n_182),
.B1(n_150),
.B2(n_148),
.Y(n_184)
);

OAI21xp33_ASAP7_75t_SL g197 ( 
.A1(n_167),
.A2(n_168),
.B(n_141),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_139),
.B(n_118),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_170),
.B(n_179),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_171),
.B(n_176),
.C(n_178),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_172),
.B(n_163),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_147),
.B(n_109),
.Y(n_174)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_174),
.Y(n_185)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_136),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_175),
.B(n_177),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_140),
.B(n_124),
.C(n_132),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_153),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_156),
.B(n_125),
.C(n_99),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_153),
.B(n_7),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_150),
.A2(n_99),
.B1(n_8),
.B2(n_9),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_184),
.A2(n_196),
.B1(n_165),
.B2(n_181),
.Y(n_202)
);

INVxp33_ASAP7_75t_L g186 ( 
.A(n_166),
.Y(n_186)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_186),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_187),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_189),
.B(n_172),
.Y(n_201)
);

BUFx24_ASAP7_75t_SL g190 ( 
.A(n_175),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g204 ( 
.A(n_190),
.Y(n_204)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_166),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_191),
.B(n_195),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_165),
.B(n_149),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_192),
.B(n_183),
.C(n_171),
.Y(n_208)
);

INVxp33_ASAP7_75t_SL g193 ( 
.A(n_173),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_193),
.A2(n_197),
.B(n_198),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_180),
.A2(n_158),
.B1(n_154),
.B2(n_144),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_194),
.A2(n_199),
.B1(n_177),
.B2(n_168),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_173),
.B(n_144),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_162),
.Y(n_196)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_164),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_180),
.A2(n_141),
.B1(n_146),
.B2(n_149),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_201),
.B(n_206),
.C(n_209),
.Y(n_217)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_202),
.Y(n_220)
);

XNOR2x1_ASAP7_75t_L g203 ( 
.A(n_192),
.B(n_181),
.Y(n_203)
);

AOI21x1_ASAP7_75t_L g222 ( 
.A1(n_203),
.A2(n_186),
.B(n_146),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_183),
.B(n_176),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_208),
.B(n_206),
.C(n_201),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_199),
.B(n_178),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_184),
.A2(n_182),
.B1(n_167),
.B2(n_170),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_211),
.A2(n_213),
.B1(n_214),
.B2(n_168),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_188),
.A2(n_167),
.B1(n_157),
.B2(n_160),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_215),
.B(n_224),
.C(n_225),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_209),
.B(n_189),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_216),
.B(n_221),
.Y(n_228)
);

NOR3xp33_ASAP7_75t_L g218 ( 
.A(n_203),
.B(n_200),
.C(n_194),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_218),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_219),
.A2(n_223),
.B1(n_151),
.B2(n_8),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_208),
.B(n_200),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_222),
.B(n_226),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_210),
.A2(n_167),
.B1(n_185),
.B2(n_169),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_207),
.B(n_212),
.C(n_213),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_207),
.B(n_212),
.C(n_205),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_205),
.B(n_179),
.C(n_161),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_226),
.B(n_7),
.C(n_9),
.Y(n_232)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_229),
.Y(n_236)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_230),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_232),
.B(n_217),
.C(n_11),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_220),
.B(n_9),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_233),
.B(n_234),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_218),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_227),
.A2(n_217),
.B1(n_11),
.B2(n_13),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_235),
.B(n_237),
.Y(n_241)
);

OR2x2_ASAP7_75t_L g237 ( 
.A(n_227),
.B(n_10),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_238),
.B(n_237),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_242),
.B(n_243),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_235),
.B(n_232),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_240),
.A2(n_231),
.B(n_230),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_244),
.A2(n_238),
.B(n_228),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_236),
.B(n_231),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_245),
.B(n_228),
.C(n_241),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_247),
.B(n_248),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_246),
.A2(n_239),
.B(n_204),
.Y(n_250)
);

BUFx24_ASAP7_75t_SL g251 ( 
.A(n_250),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_251),
.B(n_249),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_252),
.A2(n_10),
.B(n_13),
.Y(n_253)
);


endmodule