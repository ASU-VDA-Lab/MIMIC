module fake_jpeg_31478_n_54 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_54);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_54;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_3),
.Y(n_7)
);

INVx3_ASAP7_75t_L g8 ( 
.A(n_6),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

INVx3_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

BUFx5_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_8),
.B(n_1),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_16),
.B(n_17),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_8),
.B(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_12),
.B(n_0),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_19),
.B(n_20),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_7),
.B(n_0),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_L g21 ( 
.A1(n_7),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_L g27 ( 
.A1(n_21),
.A2(n_23),
.B1(n_10),
.B2(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx10_ASAP7_75t_R g26 ( 
.A(n_22),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_9),
.B(n_0),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_27),
.A2(n_29),
.B1(n_19),
.B2(n_20),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_18),
.A2(n_15),
.B1(n_10),
.B2(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_26),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_30),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_33),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_32),
.A2(n_35),
.B1(n_25),
.B2(n_34),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_23),
.Y(n_33)
);

XOR2xp5_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_15),
.Y(n_34)
);

XNOR2xp5_ASAP7_75t_L g39 ( 
.A(n_34),
.B(n_32),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_24),
.B(n_25),
.Y(n_35)
);

XOR2xp5_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_39),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_35),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_27),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_36),
.B(n_30),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_41),
.B(n_42),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_38),
.B(n_28),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g44 ( 
.A1(n_43),
.A2(n_37),
.B(n_39),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_44),
.B(n_46),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_L g46 ( 
.A1(n_43),
.A2(n_28),
.B(n_31),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_47),
.B(n_22),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_45),
.B(n_4),
.Y(n_48)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_50),
.B(n_13),
.Y(n_52)
);

NOR3xp33_ASAP7_75t_L g53 ( 
.A(n_52),
.B(n_48),
.C(n_6),
.Y(n_53)
);

AOI321xp33_ASAP7_75t_L g54 ( 
.A1(n_53),
.A2(n_5),
.A3(n_49),
.B1(n_51),
.B2(n_45),
.C(n_52),
.Y(n_54)
);


endmodule