module fake_jpeg_460_n_497 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_497);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_497;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx24_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx14_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_13),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_14),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_14),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_12),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_3),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

BUFx16f_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_2),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_1),
.B(n_12),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_0),
.B(n_4),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_10),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_55),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_56),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_57),
.Y(n_124)
);

INVx4_ASAP7_75t_SL g58 ( 
.A(n_44),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_58),
.Y(n_161)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_59),
.Y(n_156)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_60),
.Y(n_128)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_61),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_62),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_63),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_8),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_64),
.B(n_65),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_53),
.B(n_8),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_66),
.Y(n_193)
);

CKINVDCx9p33_ASAP7_75t_R g67 ( 
.A(n_20),
.Y(n_67)
);

INVx13_ASAP7_75t_L g167 ( 
.A(n_67),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_68),
.Y(n_126)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_69),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_70),
.Y(n_138)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_28),
.Y(n_71)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_71),
.Y(n_142)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

INVx13_ASAP7_75t_L g198 ( 
.A(n_72),
.Y(n_198)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_73),
.Y(n_171)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_20),
.Y(n_74)
);

INVx5_ASAP7_75t_L g189 ( 
.A(n_74),
.Y(n_189)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_20),
.Y(n_75)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_75),
.Y(n_200)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_76),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_77),
.Y(n_147)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_23),
.Y(n_78)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_78),
.Y(n_157)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_79),
.Y(n_175)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_80),
.Y(n_136)
);

INVx2_ASAP7_75t_SL g81 ( 
.A(n_23),
.Y(n_81)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_81),
.Y(n_160)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

INVx11_ASAP7_75t_L g155 ( 
.A(n_82),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_50),
.B(n_21),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_83),
.B(n_89),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_84),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_50),
.B(n_8),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_85),
.B(n_115),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_51),
.Y(n_86)
);

INVx6_ASAP7_75t_L g176 ( 
.A(n_86),
.Y(n_176)
);

INVx13_ASAP7_75t_L g87 ( 
.A(n_23),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g190 ( 
.A(n_87),
.Y(n_190)
);

INVx13_ASAP7_75t_L g88 ( 
.A(n_23),
.Y(n_88)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_88),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_34),
.B(n_11),
.Y(n_89)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_27),
.Y(n_90)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_90),
.Y(n_143)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_91),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_30),
.Y(n_92)
);

INVx6_ASAP7_75t_L g177 ( 
.A(n_92),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_21),
.B(n_11),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_93),
.B(n_110),
.Y(n_134)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_94),
.Y(n_197)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

INVx11_ASAP7_75t_L g153 ( 
.A(n_95),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_46),
.Y(n_96)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_96),
.Y(n_145)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_30),
.Y(n_97)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_97),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_31),
.A2(n_11),
.B1(n_16),
.B2(n_12),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_98),
.A2(n_22),
.B1(n_18),
.B2(n_100),
.Y(n_152)
);

INVx3_ASAP7_75t_SL g99 ( 
.A(n_33),
.Y(n_99)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_99),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_31),
.Y(n_100)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_100),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_31),
.Y(n_101)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_101),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_24),
.Y(n_102)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_102),
.Y(n_163)
);

INVx3_ASAP7_75t_SL g103 ( 
.A(n_33),
.Y(n_103)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_103),
.Y(n_170)
);

BUFx12_ASAP7_75t_L g104 ( 
.A(n_26),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_104),
.B(n_107),
.Y(n_135)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_32),
.Y(n_105)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_105),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_24),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_106),
.B(n_108),
.Y(n_180)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_34),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_24),
.Y(n_108)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_19),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_109),
.B(n_45),
.Y(n_137)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_32),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_24),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_111),
.Y(n_150)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_43),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_112),
.B(n_114),
.Y(n_174)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_37),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_113),
.B(n_45),
.Y(n_139)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_43),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_35),
.B(n_16),
.Y(n_115)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_27),
.Y(n_116)
);

INVx2_ASAP7_75t_R g125 ( 
.A(n_116),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_37),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_117),
.Y(n_164)
);

INVx11_ASAP7_75t_L g118 ( 
.A(n_25),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_118),
.A2(n_49),
.B1(n_42),
.B2(n_22),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_38),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_119),
.B(n_2),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_56),
.A2(n_25),
.B1(n_42),
.B2(n_49),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_127),
.A2(n_141),
.B1(n_152),
.B2(n_185),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_129),
.Y(n_264)
);

CKINVDCx14_ASAP7_75t_R g244 ( 
.A(n_137),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_139),
.B(n_178),
.Y(n_226)
);

OAI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_57),
.A2(n_86),
.B1(n_77),
.B2(n_70),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_140),
.A2(n_179),
.B1(n_167),
.B2(n_150),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_85),
.A2(n_38),
.B1(n_40),
.B2(n_41),
.Y(n_141)
);

OR2x2_ASAP7_75t_SL g146 ( 
.A(n_104),
.B(n_41),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_146),
.B(n_191),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_115),
.B(n_40),
.C(n_36),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_148),
.B(n_134),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_81),
.A2(n_36),
.B1(n_35),
.B2(n_18),
.Y(n_151)
);

OA22x2_ASAP7_75t_L g210 ( 
.A1(n_151),
.A2(n_173),
.B1(n_181),
.B2(n_182),
.Y(n_210)
);

INVx2_ASAP7_75t_R g159 ( 
.A(n_72),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_159),
.Y(n_214)
);

OR2x2_ASAP7_75t_L g162 ( 
.A(n_58),
.B(n_29),
.Y(n_162)
);

CKINVDCx14_ASAP7_75t_R g265 ( 
.A(n_162),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_74),
.B(n_17),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_165),
.B(n_168),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_117),
.B(n_17),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_75),
.B(n_69),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_169),
.B(n_184),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_109),
.A2(n_91),
.B1(n_80),
.B2(n_97),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_92),
.A2(n_19),
.B1(n_29),
.B2(n_6),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_87),
.A2(n_19),
.B1(n_3),
.B2(n_6),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_88),
.A2(n_19),
.B1(n_6),
.B2(n_7),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_119),
.B(n_2),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_101),
.A2(n_19),
.B1(n_6),
.B2(n_7),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_99),
.B(n_2),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_186),
.B(n_187),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_102),
.B(n_7),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_106),
.B(n_7),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_188),
.B(n_196),
.Y(n_260)
);

OR2x2_ASAP7_75t_L g191 ( 
.A(n_108),
.B(n_111),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_103),
.B(n_62),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_68),
.B(n_63),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_199),
.B(n_140),
.Y(n_266)
);

OR2x2_ASAP7_75t_L g201 ( 
.A(n_66),
.B(n_83),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_201),
.B(n_133),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_121),
.Y(n_202)
);

INVx6_ASAP7_75t_L g318 ( 
.A(n_202),
.Y(n_318)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_189),
.Y(n_203)
);

INVx4_ASAP7_75t_L g310 ( 
.A(n_203),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_174),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_204),
.B(n_206),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_135),
.Y(n_206)
);

OR2x2_ASAP7_75t_L g306 ( 
.A(n_207),
.B(n_233),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_122),
.B(n_132),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_208),
.B(n_209),
.Y(n_280)
);

NAND2xp33_ASAP7_75t_SL g211 ( 
.A(n_162),
.B(n_191),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_211),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_145),
.A2(n_164),
.B1(n_192),
.B2(n_149),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_213),
.Y(n_274)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_154),
.Y(n_215)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_215),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_201),
.A2(n_127),
.B1(n_142),
.B2(n_128),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_216),
.A2(n_240),
.B1(n_251),
.B2(n_252),
.Y(n_282)
);

BUFx2_ASAP7_75t_L g217 ( 
.A(n_120),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g316 ( 
.A(n_217),
.Y(n_316)
);

INVx6_ASAP7_75t_L g218 ( 
.A(n_121),
.Y(n_218)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_218),
.Y(n_308)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_170),
.Y(n_219)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_219),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_L g221 ( 
.A1(n_140),
.A2(n_171),
.B1(n_172),
.B2(n_175),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_221),
.A2(n_232),
.B1(n_254),
.B2(n_257),
.Y(n_292)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_177),
.Y(n_222)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_222),
.Y(n_281)
);

INVx5_ASAP7_75t_L g224 ( 
.A(n_161),
.Y(n_224)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_224),
.Y(n_285)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_177),
.Y(n_225)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_225),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_143),
.B(n_161),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_227),
.B(n_241),
.Y(n_270)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_163),
.Y(n_228)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_228),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_166),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_229),
.B(n_236),
.Y(n_298)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_195),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_230),
.Y(n_276)
);

INVx2_ASAP7_75t_SL g231 ( 
.A(n_160),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_231),
.Y(n_291)
);

AOI21xp33_ASAP7_75t_L g233 ( 
.A1(n_125),
.A2(n_180),
.B(n_197),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_149),
.A2(n_190),
.B1(n_156),
.B2(n_157),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_234),
.Y(n_309)
);

BUFx4f_ASAP7_75t_SL g235 ( 
.A(n_190),
.Y(n_235)
);

BUFx8_ASAP7_75t_L g294 ( 
.A(n_235),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_198),
.Y(n_236)
);

INVx5_ASAP7_75t_L g237 ( 
.A(n_190),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_237),
.Y(n_271)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_195),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_239),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_151),
.A2(n_129),
.B1(n_173),
.B2(n_131),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_136),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_136),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_242),
.B(n_245),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_180),
.A2(n_158),
.B1(n_125),
.B2(n_181),
.Y(n_243)
);

MAJx2_ASAP7_75t_L g313 ( 
.A(n_243),
.B(n_269),
.C(n_255),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_158),
.B(n_200),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_130),
.B(n_194),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_246),
.B(n_247),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_194),
.B(n_159),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_126),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_248),
.Y(n_297)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_126),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_249),
.Y(n_302)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_138),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_250),
.Y(n_305)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_123),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_138),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_131),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_253),
.A2(n_255),
.B1(n_256),
.B2(n_258),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_147),
.A2(n_176),
.B1(n_182),
.B2(n_144),
.Y(n_254)
);

OA22x2_ASAP7_75t_L g255 ( 
.A1(n_147),
.A2(n_176),
.B1(n_124),
.B2(n_144),
.Y(n_255)
);

INVx3_ASAP7_75t_SL g256 ( 
.A(n_123),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_124),
.A2(n_183),
.B1(n_193),
.B2(n_153),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_183),
.Y(n_258)
);

A2O1A1Ixp33_ASAP7_75t_L g259 ( 
.A1(n_167),
.A2(n_198),
.B(n_153),
.C(n_155),
.Y(n_259)
);

A2O1A1Ixp33_ASAP7_75t_L g287 ( 
.A1(n_259),
.A2(n_211),
.B(n_214),
.C(n_267),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_193),
.A2(n_134),
.B(n_201),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_261),
.B(n_235),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_174),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_262),
.B(n_266),
.Y(n_300)
);

OA22x2_ASAP7_75t_L g263 ( 
.A1(n_181),
.A2(n_182),
.B1(n_173),
.B2(n_127),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_263),
.A2(n_240),
.B1(n_210),
.B2(n_251),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_159),
.B(n_174),
.Y(n_267)
);

XNOR2x1_ASAP7_75t_SL g283 ( 
.A(n_267),
.B(n_226),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_133),
.B(n_132),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_268),
.B(n_252),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_139),
.A2(n_179),
.B1(n_184),
.B2(n_174),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_269),
.A2(n_232),
.B1(n_264),
.B2(n_226),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_272),
.A2(n_277),
.B1(n_284),
.B2(n_299),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_264),
.A2(n_226),
.B1(n_265),
.B2(n_238),
.Y(n_277)
);

NAND2x1_ASAP7_75t_L g279 ( 
.A(n_267),
.B(n_223),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_279),
.B(n_287),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_283),
.B(n_290),
.C(n_301),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_243),
.A2(n_260),
.B1(n_216),
.B2(n_263),
.Y(n_284)
);

OA22x2_ASAP7_75t_L g356 ( 
.A1(n_289),
.A2(n_286),
.B1(n_294),
.B2(n_310),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_209),
.B(n_212),
.C(n_244),
.Y(n_290)
);

A2O1A1Ixp33_ASAP7_75t_L g296 ( 
.A1(n_220),
.A2(n_205),
.B(n_214),
.C(n_259),
.Y(n_296)
);

A2O1A1Ixp33_ASAP7_75t_L g335 ( 
.A1(n_296),
.A2(n_287),
.B(n_283),
.C(n_300),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_263),
.A2(n_210),
.B1(n_255),
.B2(n_250),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_SL g301 ( 
.A(n_210),
.B(n_263),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_210),
.B(n_249),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_303),
.B(n_319),
.C(n_202),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_304),
.B(n_315),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_255),
.A2(n_230),
.B1(n_248),
.B2(n_239),
.Y(n_312)
);

AO22x1_ASAP7_75t_SL g332 ( 
.A1(n_312),
.A2(n_292),
.B1(n_284),
.B2(n_277),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_313),
.B(n_272),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_222),
.B(n_225),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_317),
.B(n_218),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_231),
.B(n_217),
.Y(n_319)
);

NOR3xp33_ASAP7_75t_SL g320 ( 
.A(n_306),
.B(n_235),
.C(n_224),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_320),
.B(n_329),
.Y(n_377)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_317),
.Y(n_321)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_321),
.Y(n_383)
);

AO21x2_ASAP7_75t_SL g323 ( 
.A1(n_299),
.A2(n_301),
.B(n_303),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g372 ( 
.A(n_323),
.B(n_332),
.Y(n_372)
);

INVx4_ASAP7_75t_L g325 ( 
.A(n_294),
.Y(n_325)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_325),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_288),
.A2(n_237),
.B(n_256),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_326),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_328),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_290),
.B(n_203),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_330),
.B(n_335),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_331),
.B(n_334),
.Y(n_361)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_281),
.Y(n_333)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_333),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_304),
.B(n_300),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_315),
.B(n_280),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_336),
.B(n_339),
.Y(n_368)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_281),
.Y(n_338)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_338),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_275),
.B(n_319),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_293),
.Y(n_340)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_340),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_306),
.B(n_295),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_341),
.B(n_345),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_307),
.B(n_270),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_342),
.B(n_347),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_288),
.A2(n_296),
.B(n_279),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g386 ( 
.A1(n_343),
.A2(n_353),
.B(n_291),
.Y(n_386)
);

BUFx5_ASAP7_75t_L g344 ( 
.A(n_294),
.Y(n_344)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_344),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_298),
.B(n_313),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_293),
.Y(n_346)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_346),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_273),
.B(n_278),
.Y(n_347)
);

NAND2x1_ASAP7_75t_SL g348 ( 
.A(n_274),
.B(n_309),
.Y(n_348)
);

INVx1_ASAP7_75t_SL g364 ( 
.A(n_348),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_279),
.B(n_278),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_349),
.B(n_351),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_297),
.B(n_305),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_350),
.B(n_354),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_311),
.B(n_271),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_311),
.Y(n_352)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_352),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_282),
.A2(n_274),
.B(n_309),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_316),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_276),
.Y(n_355)
);

INVx1_ASAP7_75t_SL g378 ( 
.A(n_355),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_356),
.A2(n_285),
.B1(n_310),
.B2(n_314),
.Y(n_374)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_276),
.Y(n_357)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_357),
.Y(n_384)
);

CKINVDCx16_ASAP7_75t_R g363 ( 
.A(n_350),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_363),
.B(n_385),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_323),
.A2(n_312),
.B1(n_302),
.B2(n_308),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_L g397 ( 
.A1(n_365),
.A2(n_374),
.B1(n_379),
.B2(n_323),
.Y(n_397)
);

CKINVDCx12_ASAP7_75t_R g373 ( 
.A(n_344),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_373),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_337),
.A2(n_308),
.B1(n_318),
.B2(n_285),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_324),
.B(n_314),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_381),
.B(n_324),
.C(n_336),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_331),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_386),
.A2(n_364),
.B(n_371),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_388),
.B(n_389),
.C(n_390),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_381),
.B(n_345),
.C(n_327),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_360),
.B(n_382),
.C(n_368),
.Y(n_390)
);

CKINVDCx16_ASAP7_75t_R g391 ( 
.A(n_384),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_391),
.B(n_393),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_360),
.B(n_327),
.C(n_335),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_392),
.B(n_396),
.C(n_382),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_SL g393 ( 
.A(n_376),
.B(n_341),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_372),
.A2(n_323),
.B1(n_332),
.B2(n_343),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_394),
.A2(n_398),
.B1(n_411),
.B2(n_399),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_368),
.B(n_329),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_395),
.B(n_402),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_375),
.B(n_327),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_397),
.B(n_407),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_372),
.A2(n_332),
.B1(n_334),
.B2(n_337),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_387),
.Y(n_399)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_399),
.Y(n_414)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_387),
.Y(n_400)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_400),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_367),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g430 ( 
.A1(n_403),
.A2(n_405),
.B(n_406),
.Y(n_430)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_380),
.Y(n_404)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_404),
.Y(n_429)
);

AOI21xp5_ASAP7_75t_SL g405 ( 
.A1(n_372),
.A2(n_322),
.B(n_326),
.Y(n_405)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_380),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_361),
.B(n_321),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_408),
.Y(n_424)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_358),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_409),
.B(n_410),
.Y(n_423)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_358),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_365),
.A2(n_330),
.B1(n_322),
.B2(n_356),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_359),
.Y(n_412)
);

NAND2xp33_ASAP7_75t_R g433 ( 
.A(n_412),
.B(n_407),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_417),
.B(n_418),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_389),
.B(n_375),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_388),
.B(n_361),
.C(n_383),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_419),
.B(n_420),
.C(n_427),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_390),
.B(n_339),
.C(n_386),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_398),
.A2(n_371),
.B1(n_364),
.B2(n_377),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_421),
.A2(n_411),
.B1(n_403),
.B2(n_374),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_426),
.B(n_430),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_392),
.B(n_378),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_396),
.B(n_378),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_428),
.B(n_412),
.C(n_410),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_408),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_431),
.B(n_424),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_SL g432 ( 
.A(n_394),
.B(n_320),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_SL g442 ( 
.A(n_432),
.B(n_353),
.Y(n_442)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_433),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_434),
.B(n_446),
.Y(n_453)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_423),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_436),
.B(n_438),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_413),
.A2(n_400),
.B1(n_405),
.B2(n_393),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_437),
.A2(n_430),
.B1(n_421),
.B2(n_413),
.Y(n_458)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_423),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_419),
.B(n_401),
.Y(n_440)
);

CKINVDCx16_ASAP7_75t_R g462 ( 
.A(n_440),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_442),
.B(n_443),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_416),
.B(n_404),
.C(n_362),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_444),
.B(n_447),
.C(n_428),
.Y(n_459)
);

INVx1_ASAP7_75t_SL g446 ( 
.A(n_423),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_416),
.B(n_370),
.C(n_362),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_448),
.Y(n_452)
);

CKINVDCx16_ASAP7_75t_R g449 ( 
.A(n_425),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_449),
.B(n_402),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_439),
.B(n_427),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_451),
.B(n_454),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_439),
.B(n_418),
.Y(n_454)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_455),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_441),
.B(n_417),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_457),
.B(n_441),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_458),
.A2(n_434),
.B1(n_453),
.B2(n_445),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_459),
.B(n_460),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_447),
.B(n_420),
.C(n_426),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_SL g461 ( 
.A1(n_445),
.A2(n_413),
.B(n_432),
.Y(n_461)
);

CKINVDCx14_ASAP7_75t_R g472 ( 
.A(n_461),
.Y(n_472)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_463),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_464),
.B(n_465),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_451),
.B(n_444),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_454),
.B(n_443),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_466),
.B(n_471),
.Y(n_478)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_450),
.Y(n_470)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_470),
.Y(n_477)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_462),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_472),
.A2(n_458),
.B1(n_453),
.B2(n_452),
.Y(n_474)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_474),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_L g475 ( 
.A1(n_469),
.A2(n_437),
.B1(n_435),
.B2(n_422),
.Y(n_475)
);

INVxp67_ASAP7_75t_L g484 ( 
.A(n_475),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_L g479 ( 
.A1(n_468),
.A2(n_414),
.B1(n_415),
.B2(n_460),
.Y(n_479)
);

AOI21xp5_ASAP7_75t_L g485 ( 
.A1(n_479),
.A2(n_459),
.B(n_461),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_SL g480 ( 
.A(n_464),
.B(n_457),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_SL g481 ( 
.A(n_480),
.B(n_467),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_481),
.B(n_477),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_L g482 ( 
.A1(n_478),
.A2(n_466),
.B(n_465),
.Y(n_482)
);

AOI21xp5_ASAP7_75t_L g490 ( 
.A1(n_482),
.A2(n_485),
.B(n_486),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_L g486 ( 
.A1(n_474),
.A2(n_467),
.B(n_456),
.Y(n_486)
);

AOI21xp5_ASAP7_75t_SL g487 ( 
.A1(n_484),
.A2(n_477),
.B(n_476),
.Y(n_487)
);

HB1xp67_ASAP7_75t_L g492 ( 
.A(n_487),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_483),
.B(n_473),
.C(n_476),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_488),
.B(n_489),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_491),
.B(n_490),
.C(n_446),
.Y(n_493)
);

AOI321xp33_ASAP7_75t_L g495 ( 
.A1(n_493),
.A2(n_494),
.A3(n_429),
.B1(n_369),
.B2(n_354),
.C(n_366),
.Y(n_495)
);

AOI21xp5_ASAP7_75t_L g494 ( 
.A1(n_492),
.A2(n_456),
.B(n_401),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_495),
.B(n_369),
.C(n_359),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_496),
.B(n_370),
.Y(n_497)
);


endmodule