module fake_jpeg_9691_n_262 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_262);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_262;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

BUFx12_ASAP7_75t_L g13 ( 
.A(n_11),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx8_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_12),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_28),
.B(n_33),
.Y(n_54)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_29),
.B(n_32),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_13),
.B(n_0),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx3_ASAP7_75t_SL g48 ( 
.A(n_34),
.Y(n_48)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_40),
.B(n_41),
.Y(n_71)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_44),
.Y(n_56)
);

OA22x2_ASAP7_75t_L g45 ( 
.A1(n_34),
.A2(n_23),
.B1(n_17),
.B2(n_16),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_45),
.A2(n_52),
.B1(n_24),
.B2(n_21),
.Y(n_72)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_34),
.A2(n_18),
.B1(n_20),
.B2(n_17),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_58),
.B(n_62),
.Y(n_80)
);

NOR2x1_ASAP7_75t_R g59 ( 
.A(n_45),
.B(n_23),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_59),
.A2(n_65),
.B1(n_72),
.B2(n_24),
.Y(n_90)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_60),
.Y(n_76)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_51),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_63),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g65 ( 
.A(n_54),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g67 ( 
.A(n_44),
.Y(n_67)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_39),
.A2(n_34),
.B1(n_18),
.B2(n_20),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_69),
.A2(n_24),
.B1(n_21),
.B2(n_26),
.Y(n_91)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_73),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_59),
.A2(n_41),
.B1(n_39),
.B2(n_46),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_75),
.A2(n_86),
.B1(n_70),
.B2(n_49),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_57),
.B(n_42),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_77),
.B(n_81),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_72),
.B(n_45),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_61),
.A2(n_20),
.B1(n_18),
.B2(n_49),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_71),
.B(n_35),
.C(n_31),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_68),
.C(n_64),
.Y(n_104)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_85),
.B(n_87),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_58),
.A2(n_53),
.B1(n_35),
.B2(n_45),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_60),
.B(n_28),
.Y(n_87)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_89),
.Y(n_96)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_90),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_91),
.A2(n_22),
.B1(n_25),
.B2(n_26),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_66),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_92),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_94),
.B(n_103),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_81),
.A2(n_29),
.B(n_13),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_98),
.A2(n_110),
.B(n_22),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_33),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_SL g117 ( 
.A(n_99),
.B(n_31),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_101),
.Y(n_122)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_104),
.B(n_105),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_78),
.B(n_68),
.C(n_64),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_86),
.A2(n_66),
.B1(n_70),
.B2(n_73),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_106),
.A2(n_114),
.B1(n_76),
.B2(n_92),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_108),
.A2(n_111),
.B1(n_79),
.B2(n_89),
.Y(n_135)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_74),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_109),
.B(n_112),
.Y(n_133)
);

O2A1O1Ixp33_ASAP7_75t_SL g110 ( 
.A1(n_75),
.A2(n_26),
.B(n_22),
.C(n_25),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_78),
.A2(n_29),
.B1(n_37),
.B2(n_36),
.Y(n_111)
);

BUFx24_ASAP7_75t_SL g112 ( 
.A(n_77),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_88),
.Y(n_113)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_113),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_83),
.A2(n_29),
.B1(n_37),
.B2(n_36),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_115),
.A2(n_129),
.B1(n_108),
.B2(n_97),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_87),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_116),
.B(n_126),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_117),
.B(n_110),
.Y(n_139)
);

MAJx2_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_93),
.C(n_83),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_119),
.B(n_114),
.C(n_96),
.Y(n_143)
);

AOI32xp33_ASAP7_75t_L g121 ( 
.A1(n_100),
.A2(n_93),
.A3(n_76),
.B1(n_88),
.B2(n_33),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_121),
.A2(n_123),
.B(n_132),
.Y(n_151)
);

NOR2xp67_ASAP7_75t_SL g123 ( 
.A(n_101),
.B(n_93),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_102),
.A2(n_96),
.B1(n_109),
.B2(n_88),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_124),
.A2(n_127),
.B1(n_128),
.B2(n_130),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_107),
.B(n_104),
.Y(n_126)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_91),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_97),
.A2(n_79),
.B1(n_85),
.B2(n_89),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_105),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_98),
.B(n_74),
.Y(n_131)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_131),
.Y(n_141)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_111),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_95),
.B(n_74),
.Y(n_134)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_134),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_135),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_134),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_136),
.B(n_140),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_137),
.A2(n_27),
.B1(n_19),
.B2(n_23),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_125),
.B(n_126),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_138),
.B(n_143),
.C(n_152),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_139),
.B(n_128),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_131),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_129),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_144),
.B(n_147),
.Y(n_176)
);

INVxp33_ASAP7_75t_L g145 ( 
.A(n_115),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_145),
.B(n_154),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g147 ( 
.A(n_116),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_132),
.A2(n_110),
.B1(n_94),
.B2(n_113),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_150),
.A2(n_56),
.B1(n_19),
.B2(n_27),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_117),
.B(n_60),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_125),
.B(n_67),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_153),
.B(n_157),
.C(n_133),
.Y(n_170)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_120),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_130),
.B(n_0),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_155),
.A2(n_0),
.B(n_1),
.Y(n_178)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_135),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_156),
.B(n_127),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_119),
.B(n_67),
.C(n_56),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_159),
.B(n_175),
.Y(n_185)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_137),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_160),
.B(n_161),
.Y(n_180)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_142),
.Y(n_161)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_163),
.Y(n_188)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_155),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_164),
.B(n_173),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_148),
.A2(n_122),
.B1(n_118),
.B2(n_25),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_165),
.A2(n_166),
.B1(n_168),
.B2(n_171),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_141),
.A2(n_122),
.B1(n_118),
.B2(n_15),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_167),
.A2(n_146),
.B1(n_147),
.B2(n_150),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_144),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_170),
.B(n_172),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_145),
.A2(n_16),
.B1(n_15),
.B2(n_37),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_138),
.B(n_56),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_155),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_174),
.A2(n_149),
.B1(n_27),
.B2(n_19),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_152),
.B(n_23),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_153),
.B(n_27),
.C(n_19),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_177),
.B(n_139),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_178),
.B(n_151),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_158),
.Y(n_179)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_179),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_176),
.Y(n_181)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_181),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_182),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_165),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_183),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_162),
.A2(n_151),
.B1(n_143),
.B2(n_157),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_187),
.A2(n_195),
.B1(n_196),
.B2(n_13),
.Y(n_210)
);

CKINVDCx14_ASAP7_75t_R g212 ( 
.A(n_189),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_190),
.B(n_13),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_166),
.Y(n_191)
);

OAI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_191),
.A2(n_177),
.B1(n_172),
.B2(n_175),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_178),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_193),
.B(n_194),
.C(n_167),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_171),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_168),
.A2(n_149),
.B1(n_27),
.B2(n_19),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_185),
.B(n_159),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_SL g219 ( 
.A(n_197),
.B(n_205),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_199),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_200),
.B(n_210),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_184),
.B(n_169),
.C(n_187),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_203),
.B(n_204),
.C(n_208),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_184),
.B(n_169),
.C(n_170),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g205 ( 
.A(n_185),
.B(n_12),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_180),
.A2(n_11),
.B(n_10),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_206),
.A2(n_192),
.B(n_182),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_189),
.B(n_13),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_209),
.B(n_2),
.Y(n_225)
);

XOR2x2_ASAP7_75t_L g211 ( 
.A(n_190),
.B(n_10),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_211),
.A2(n_188),
.B(n_186),
.Y(n_213)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_213),
.Y(n_226)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_214),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_202),
.A2(n_191),
.B1(n_192),
.B2(n_2),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_216),
.B(n_223),
.C(n_207),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_201),
.B(n_10),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_218),
.B(n_222),
.Y(n_230)
);

NOR2xp67_ASAP7_75t_R g221 ( 
.A(n_211),
.B(n_0),
.Y(n_221)
);

XNOR2x2_ASAP7_75t_L g228 ( 
.A(n_221),
.B(n_223),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_206),
.B(n_9),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_212),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_198),
.B(n_2),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_224),
.B(n_3),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_225),
.B(n_205),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_227),
.B(n_236),
.Y(n_238)
);

AO21x1_ASAP7_75t_L g245 ( 
.A1(n_228),
.A2(n_231),
.B(n_4),
.Y(n_245)
);

NOR2xp67_ASAP7_75t_L g231 ( 
.A(n_217),
.B(n_200),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_232),
.B(n_234),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_215),
.B(n_203),
.Y(n_233)
);

OR2x2_ASAP7_75t_L g242 ( 
.A(n_233),
.B(n_235),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_215),
.B(n_220),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_219),
.B(n_197),
.C(n_208),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_229),
.A2(n_231),
.B(n_226),
.Y(n_237)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_237),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_230),
.B(n_216),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_239),
.B(n_240),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_230),
.B(n_225),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_232),
.B(n_219),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_241),
.B(n_4),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_230),
.B(n_4),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_244),
.B(n_245),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_238),
.B(n_4),
.C(n_5),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_247),
.B(n_248),
.Y(n_255)
);

OAI21x1_ASAP7_75t_L g250 ( 
.A1(n_242),
.A2(n_5),
.B(n_6),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_250),
.B(n_249),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_251),
.A2(n_243),
.B(n_244),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_252),
.B(n_253),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_246),
.A2(n_243),
.B(n_6),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_254),
.B(n_249),
.Y(n_257)
);

A2O1A1O1Ixp25_ASAP7_75t_L g258 ( 
.A1(n_257),
.A2(n_255),
.B(n_7),
.C(n_8),
.D(n_9),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_258),
.B(n_256),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_259),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_260),
.B(n_5),
.C(n_7),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_261),
.B(n_8),
.Y(n_262)
);


endmodule