module fake_jpeg_24263_n_79 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_79);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_79;

wire n_10;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_6),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_SL g12 ( 
.A(n_5),
.B(n_0),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx2_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx6_ASAP7_75t_SL g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_16),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_21),
.B(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_15),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_22),
.B(n_26),
.Y(n_33)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_16),
.B(n_1),
.C(n_2),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g37 ( 
.A1(n_24),
.A2(n_25),
.B(n_19),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g25 ( 
.A1(n_16),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_12),
.B(n_14),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_28),
.Y(n_34)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_30),
.A2(n_11),
.B1(n_13),
.B2(n_18),
.Y(n_39)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_15),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_32),
.B(n_35),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_21),
.B(n_12),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_19),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_10),
.C(n_14),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_37),
.A2(n_13),
.B1(n_11),
.B2(n_10),
.Y(n_40)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_39),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_43),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_35),
.A2(n_28),
.B1(n_23),
.B2(n_27),
.Y(n_41)
);

OAI32xp33_ASAP7_75t_L g48 ( 
.A1(n_41),
.A2(n_32),
.A3(n_37),
.B1(n_30),
.B2(n_25),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_33),
.B(n_20),
.Y(n_42)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_34),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_47),
.Y(n_55)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_48),
.A2(n_30),
.B1(n_28),
.B2(n_23),
.Y(n_62)
);

AND2x2_ASAP7_75t_SL g50 ( 
.A(n_46),
.B(n_32),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_44),
.C(n_45),
.Y(n_58)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_48),
.A2(n_46),
.B1(n_47),
.B2(n_41),
.Y(n_56)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_L g57 ( 
.A(n_50),
.B(n_36),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_58),
.C(n_62),
.Y(n_65)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_61),
.Y(n_63)
);

AO21x1_ASAP7_75t_L g64 ( 
.A1(n_59),
.A2(n_53),
.B(n_50),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_64),
.B(n_56),
.Y(n_70)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_66),
.B(n_49),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_68),
.A2(n_70),
.B(n_71),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_65),
.B(n_58),
.C(n_57),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_69),
.B(n_67),
.C(n_63),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_64),
.B(n_55),
.Y(n_71)
);

OAI21xp33_ASAP7_75t_L g76 ( 
.A1(n_72),
.A2(n_8),
.B(n_9),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_69),
.B(n_49),
.C(n_20),
.Y(n_74)
);

NOR3xp33_ASAP7_75t_L g75 ( 
.A(n_74),
.B(n_18),
.C(n_9),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_75),
.B(n_76),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_77),
.A2(n_73),
.B(n_29),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_78),
.B(n_29),
.Y(n_79)
);


endmodule