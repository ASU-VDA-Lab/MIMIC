module fake_jpeg_29203_n_167 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_167);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_167;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_14),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_11),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_50),
.Y(n_55)
);

CKINVDCx14_ASAP7_75t_R g56 ( 
.A(n_16),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_18),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_12),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_7),
.B(n_34),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_45),
.Y(n_63)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

BUFx4f_ASAP7_75t_L g65 ( 
.A(n_13),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_40),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_2),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

BUFx4f_ASAP7_75t_SL g71 ( 
.A(n_9),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_31),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_21),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_9),
.Y(n_74)
);

BUFx12_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_75),
.B(n_79),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

INVx2_ASAP7_75t_SL g96 ( 
.A(n_76),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_0),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_77),
.B(n_80),
.Y(n_84)
);

INVx3_ASAP7_75t_SL g78 ( 
.A(n_65),
.Y(n_78)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_73),
.Y(n_80)
);

AND2x2_ASAP7_75t_SL g81 ( 
.A(n_72),
.B(n_19),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_81),
.B(n_66),
.C(n_56),
.Y(n_86)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_62),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_61),
.B(n_23),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_83),
.B(n_0),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_83),
.B(n_53),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_94),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_86),
.B(n_92),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_78),
.A2(n_67),
.B1(n_74),
.B2(n_56),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_88),
.B(n_90),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_79),
.A2(n_73),
.B1(n_59),
.B2(n_60),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_89),
.A2(n_91),
.B1(n_98),
.B2(n_88),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_78),
.A2(n_52),
.B1(n_70),
.B2(n_54),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_80),
.A2(n_62),
.B1(n_68),
.B2(n_59),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_81),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_95),
.B(n_75),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_81),
.B(n_55),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_97),
.B(n_86),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_76),
.A2(n_82),
.B1(n_68),
.B2(n_64),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_96),
.Y(n_99)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_99),
.Y(n_122)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_96),
.Y(n_100)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_100),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_103),
.A2(n_113),
.B1(n_117),
.B2(n_7),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_104),
.B(n_8),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_91),
.A2(n_76),
.B1(n_71),
.B2(n_75),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_105),
.A2(n_109),
.B1(n_10),
.B2(n_11),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_6),
.Y(n_127)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_95),
.Y(n_107)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_107),
.Y(n_130)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_108),
.Y(n_131)
);

NAND2x1p5_ASAP7_75t_R g109 ( 
.A(n_89),
.B(n_71),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_84),
.B(n_57),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_111),
.B(n_5),
.Y(n_121)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_112),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_84),
.A2(n_76),
.B1(n_63),
.B2(n_58),
.Y(n_113)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_93),
.Y(n_114)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_115),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_89),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_116),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_94),
.A2(n_24),
.B1(n_44),
.B2(n_43),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_94),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_118),
.A2(n_8),
.B(n_10),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_110),
.B(n_25),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_119),
.B(n_126),
.C(n_28),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_120),
.A2(n_137),
.B1(n_12),
.B2(n_13),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_121),
.B(n_134),
.Y(n_141)
);

XNOR2x1_ASAP7_75t_SL g123 ( 
.A(n_101),
.B(n_26),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_123),
.B(n_14),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_114),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_124),
.B(n_127),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_106),
.B(n_27),
.C(n_42),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_128),
.A2(n_102),
.B1(n_116),
.B2(n_105),
.Y(n_140)
);

INVx13_ASAP7_75t_L g129 ( 
.A(n_115),
.Y(n_129)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_129),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_132),
.B(n_120),
.Y(n_150)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_99),
.Y(n_136)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_136),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_130),
.A2(n_101),
.B(n_113),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_138),
.A2(n_133),
.B(n_135),
.Y(n_153)
);

A2O1A1O1Ixp25_ASAP7_75t_L g157 ( 
.A1(n_140),
.A2(n_144),
.B(n_151),
.C(n_139),
.D(n_149),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_142),
.A2(n_149),
.B(n_126),
.Y(n_152)
);

AO22x1_ASAP7_75t_SL g144 ( 
.A1(n_131),
.A2(n_48),
.B1(n_15),
.B2(n_17),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_145),
.B(n_147),
.C(n_148),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_SL g148 ( 
.A(n_119),
.B(n_29),
.Y(n_148)
);

NOR2x1_ASAP7_75t_L g149 ( 
.A(n_128),
.B(n_32),
.Y(n_149)
);

NAND3xp33_ASAP7_75t_L g155 ( 
.A(n_150),
.B(n_38),
.C(n_41),
.Y(n_155)
);

OAI21xp33_ASAP7_75t_L g151 ( 
.A1(n_123),
.A2(n_33),
.B(n_37),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_152),
.A2(n_153),
.B1(n_155),
.B2(n_157),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_148),
.B(n_125),
.C(n_122),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_156),
.B(n_141),
.C(n_146),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_158),
.B(n_160),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_154),
.B(n_151),
.C(n_144),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_159),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_161),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_162),
.C(n_144),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_164),
.B(n_143),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_165),
.Y(n_166)
);

HB1xp67_ASAP7_75t_L g167 ( 
.A(n_166),
.Y(n_167)
);


endmodule