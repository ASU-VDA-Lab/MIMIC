module fake_jpeg_12275_n_526 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_526);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_526;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_SL g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

INVx11_ASAP7_75t_SL g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_0),
.B(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_13),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g44 ( 
.A(n_1),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_3),
.Y(n_46)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_49),
.Y(n_114)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

INVx11_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_51),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_52),
.Y(n_119)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_53),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g134 ( 
.A(n_54),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_55),
.Y(n_99)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_56),
.Y(n_105)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_57),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_58),
.Y(n_131)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_59),
.Y(n_117)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_60),
.Y(n_151)
);

BUFx10_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

INVxp67_ASAP7_75t_SL g120 ( 
.A(n_61),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_62),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_34),
.B(n_14),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_63),
.B(n_74),
.Y(n_118)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_21),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_64),
.Y(n_133)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_65),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_66),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_67),
.Y(n_147)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_68),
.Y(n_121)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_17),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g128 ( 
.A(n_69),
.Y(n_128)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g154 ( 
.A(n_70),
.Y(n_154)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_71),
.Y(n_122)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_72),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_34),
.B(n_14),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_73),
.B(n_82),
.Y(n_149)
);

AOI21xp33_ASAP7_75t_L g74 ( 
.A1(n_19),
.A2(n_14),
.B(n_12),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_20),
.Y(n_75)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_17),
.Y(n_76)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_76),
.Y(n_137)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_38),
.Y(n_77)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_77),
.Y(n_139)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_20),
.Y(n_78)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_78),
.Y(n_109)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_17),
.Y(n_79)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_79),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_37),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_80),
.B(n_94),
.Y(n_106)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_24),
.Y(n_81)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_81),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_19),
.B(n_14),
.Y(n_82)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_25),
.Y(n_83)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_83),
.Y(n_110)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_41),
.Y(n_84)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_84),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_24),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_85),
.Y(n_150)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_24),
.Y(n_86)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_86),
.Y(n_155)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_41),
.Y(n_87)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_87),
.Y(n_123)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_18),
.Y(n_88)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_44),
.B(n_11),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_89),
.B(n_37),
.Y(n_127)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_41),
.Y(n_90)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_90),
.Y(n_144)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_24),
.Y(n_91)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_91),
.Y(n_157)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_42),
.Y(n_92)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_92),
.Y(n_145)
);

BUFx4f_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_93),
.Y(n_153)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_18),
.Y(n_94)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_95),
.Y(n_115)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_23),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_96),
.B(n_26),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_28),
.Y(n_97)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_97),
.Y(n_135)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_28),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_98),
.B(n_35),
.Y(n_142)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_63),
.B(n_23),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_101),
.B(n_111),
.Y(n_168)
);

OAI22xp33_ASAP7_75t_L g107 ( 
.A1(n_53),
.A2(n_29),
.B1(n_39),
.B2(n_32),
.Y(n_107)
);

AO22x2_ASAP7_75t_L g202 ( 
.A1(n_107),
.A2(n_97),
.B1(n_67),
.B2(n_85),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_52),
.A2(n_29),
.B1(n_39),
.B2(n_32),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_L g197 ( 
.A1(n_108),
.A2(n_140),
.B1(n_29),
.B2(n_39),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_64),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_127),
.B(n_143),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_83),
.B(n_15),
.C(n_35),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_130),
.B(n_44),
.C(n_28),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_136),
.B(n_138),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_61),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_58),
.A2(n_48),
.B1(n_45),
.B2(n_42),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_142),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_89),
.B(n_33),
.Y(n_143)
);

OR2x2_ASAP7_75t_L g146 ( 
.A(n_61),
.B(n_43),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_146),
.B(n_156),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_55),
.B(n_33),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_148),
.B(n_15),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_66),
.A2(n_48),
.B1(n_45),
.B2(n_42),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_152),
.A2(n_39),
.B1(n_32),
.B2(n_29),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_55),
.B(n_31),
.Y(n_156)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_141),
.Y(n_158)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_158),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_120),
.A2(n_15),
.B1(n_35),
.B2(n_76),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_159),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_160),
.B(n_171),
.Y(n_223)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_144),
.Y(n_161)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_161),
.Y(n_215)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_155),
.Y(n_162)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_162),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_149),
.B(n_26),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_164),
.B(n_170),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_120),
.A2(n_49),
.B1(n_57),
.B2(n_51),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_165),
.Y(n_221)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_144),
.Y(n_166)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_166),
.Y(n_238)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_137),
.Y(n_167)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_167),
.Y(n_230)
);

INVx2_ASAP7_75t_SL g169 ( 
.A(n_110),
.Y(n_169)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_169),
.Y(n_209)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_103),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g171 ( 
.A(n_106),
.Y(n_171)
);

INVx6_ASAP7_75t_L g172 ( 
.A(n_119),
.Y(n_172)
);

INVx6_ASAP7_75t_L g226 ( 
.A(n_172),
.Y(n_226)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_109),
.Y(n_173)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_173),
.Y(n_211)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_119),
.Y(n_174)
);

INVx5_ASAP7_75t_L g210 ( 
.A(n_174),
.Y(n_210)
);

INVx5_ASAP7_75t_L g175 ( 
.A(n_115),
.Y(n_175)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_175),
.Y(n_235)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_157),
.Y(n_176)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_176),
.Y(n_227)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_122),
.Y(n_177)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_177),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_101),
.B(n_46),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_179),
.B(n_183),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_134),
.Y(n_180)
);

INVx13_ASAP7_75t_L g217 ( 
.A(n_180),
.Y(n_217)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_112),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_182),
.B(n_186),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_146),
.B(n_46),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_118),
.A2(n_54),
.B1(n_43),
.B2(n_30),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_184),
.Y(n_224)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_124),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_185),
.B(n_187),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_131),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_145),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_114),
.A2(n_30),
.B1(n_95),
.B2(n_62),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_188),
.A2(n_99),
.B1(n_114),
.B2(n_128),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_104),
.B(n_31),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_189),
.B(n_198),
.Y(n_244)
);

INVx6_ASAP7_75t_L g190 ( 
.A(n_131),
.Y(n_190)
);

INVxp33_ASAP7_75t_L g234 ( 
.A(n_190),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_134),
.Y(n_191)
);

CKINVDCx14_ASAP7_75t_R g241 ( 
.A(n_191),
.Y(n_241)
);

CKINVDCx12_ASAP7_75t_R g192 ( 
.A(n_102),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_192),
.Y(n_228)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_139),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_193),
.B(n_197),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_194),
.A2(n_202),
.B1(n_204),
.B2(n_107),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_154),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_196),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_121),
.B(n_133),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_199),
.B(n_154),
.C(n_128),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_134),
.Y(n_200)
);

NAND2xp33_ASAP7_75t_SL g236 ( 
.A(n_200),
.B(n_203),
.Y(n_236)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_116),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_201),
.B(n_205),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_153),
.Y(n_203)
);

OAI22xp33_ASAP7_75t_L g204 ( 
.A1(n_108),
.A2(n_28),
.B1(n_32),
.B2(n_48),
.Y(n_204)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_153),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_142),
.B(n_12),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_206),
.B(n_207),
.Y(n_214)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_129),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_208),
.A2(n_202),
.B1(n_150),
.B2(n_132),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_218),
.A2(n_123),
.B1(n_102),
.B2(n_200),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_199),
.B(n_178),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_220),
.B(n_229),
.C(n_232),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_168),
.B(n_100),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_225),
.B(n_176),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_163),
.B(n_105),
.C(n_151),
.Y(n_232)
);

OA21x2_ASAP7_75t_L g239 ( 
.A1(n_202),
.A2(n_105),
.B(n_117),
.Y(n_239)
);

O2A1O1Ixp33_ASAP7_75t_SL g250 ( 
.A1(n_239),
.A2(n_202),
.B(n_204),
.C(n_197),
.Y(n_250)
);

AND2x2_ASAP7_75t_SL g240 ( 
.A(n_169),
.B(n_99),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_240),
.Y(n_253)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_213),
.Y(n_246)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_246),
.Y(n_285)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_212),
.Y(n_247)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_247),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_225),
.B(n_181),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_248),
.B(n_251),
.Y(n_310)
);

OAI32xp33_ASAP7_75t_L g249 ( 
.A1(n_245),
.A2(n_195),
.A3(n_193),
.B1(n_177),
.B2(n_185),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_249),
.B(n_252),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_250),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_223),
.B(n_166),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_244),
.B(n_158),
.Y(n_252)
);

INVx13_ASAP7_75t_L g254 ( 
.A(n_217),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_254),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_255),
.A2(n_270),
.B1(n_218),
.B2(n_221),
.Y(n_284)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_213),
.Y(n_256)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_256),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_220),
.B(n_229),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_257),
.B(n_267),
.C(n_214),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_244),
.B(n_161),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_258),
.B(n_260),
.Y(n_299)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_209),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_259),
.B(n_265),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_232),
.B(n_242),
.Y(n_260)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_210),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_261),
.A2(n_263),
.B1(n_264),
.B2(n_266),
.Y(n_297)
);

OA22x2_ASAP7_75t_L g262 ( 
.A1(n_239),
.A2(n_207),
.B1(n_135),
.B2(n_115),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_262),
.A2(n_272),
.B(n_279),
.Y(n_292)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_212),
.Y(n_263)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_209),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_214),
.B(n_167),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_226),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_268),
.Y(n_302)
);

INVx6_ASAP7_75t_L g269 ( 
.A(n_226),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_269),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_239),
.A2(n_175),
.B1(n_126),
.B2(n_135),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_245),
.B(n_201),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g303 ( 
.A(n_271),
.B(n_216),
.Y(n_303)
);

AND2x6_ASAP7_75t_L g272 ( 
.A(n_224),
.B(n_125),
.Y(n_272)
);

INVx11_ASAP7_75t_L g273 ( 
.A(n_217),
.Y(n_273)
);

NAND2xp33_ASAP7_75t_SL g311 ( 
.A(n_273),
.B(n_277),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_242),
.B(n_203),
.Y(n_274)
);

MAJx2_ASAP7_75t_L g296 ( 
.A(n_274),
.B(n_275),
.C(n_278),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_228),
.B(n_191),
.Y(n_275)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_227),
.Y(n_277)
);

BUFx24_ASAP7_75t_SL g278 ( 
.A(n_211),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_230),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_281),
.B(n_301),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_257),
.B(n_211),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_283),
.B(n_287),
.C(n_298),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_284),
.A2(n_290),
.B1(n_291),
.B2(n_294),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_276),
.B(n_224),
.C(n_240),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_246),
.A2(n_239),
.B1(n_231),
.B2(n_208),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_288),
.A2(n_293),
.B1(n_305),
.B2(n_307),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_255),
.A2(n_231),
.B1(n_219),
.B2(n_233),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_270),
.A2(n_231),
.B1(n_172),
.B2(n_190),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_256),
.A2(n_240),
.B1(n_235),
.B2(n_234),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_250),
.A2(n_174),
.B1(n_226),
.B2(n_210),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_250),
.A2(n_276),
.B1(n_262),
.B2(n_253),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_295),
.B(n_306),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_267),
.B(n_240),
.C(n_228),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_252),
.B(n_216),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_303),
.B(n_247),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_271),
.B(n_216),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_304),
.B(n_308),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_253),
.A2(n_235),
.B1(n_237),
.B2(n_243),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_262),
.A2(n_186),
.B1(n_150),
.B2(n_132),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_262),
.A2(n_237),
.B1(n_243),
.B2(n_227),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_265),
.B(n_249),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_SL g309 ( 
.A(n_259),
.B(n_236),
.Y(n_309)
);

HAxp5_ASAP7_75t_SL g342 ( 
.A(n_309),
.B(n_217),
.CON(n_342),
.SN(n_342)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_272),
.A2(n_236),
.B(n_241),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_314),
.A2(n_125),
.B(n_273),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_299),
.B(n_310),
.Y(n_315)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_315),
.Y(n_357)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_312),
.Y(n_316)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_316),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_299),
.B(n_266),
.Y(n_317)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_317),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_318),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_285),
.B(n_277),
.Y(n_319)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_319),
.Y(n_367)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_285),
.Y(n_322)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_322),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_286),
.B(n_308),
.Y(n_323)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_323),
.Y(n_380)
);

INVx13_ASAP7_75t_L g324 ( 
.A(n_313),
.Y(n_324)
);

INVx2_ASAP7_75t_SL g366 ( 
.A(n_324),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_286),
.B(n_305),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_326),
.B(n_330),
.Y(n_356)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_293),
.B(n_261),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_327),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_300),
.A2(n_269),
.B1(n_268),
.B2(n_279),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_328),
.A2(n_334),
.B1(n_349),
.B2(n_123),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_287),
.B(n_268),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_329),
.B(n_335),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_307),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_280),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_331),
.B(n_332),
.Y(n_371)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_280),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_289),
.B(n_263),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_333),
.B(n_339),
.Y(n_373)
);

AOI22xp33_ASAP7_75t_SL g334 ( 
.A1(n_300),
.A2(n_238),
.B1(n_215),
.B2(n_254),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g335 ( 
.A(n_289),
.Y(n_335)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_304),
.Y(n_337)
);

INVx3_ASAP7_75t_L g350 ( 
.A(n_337),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_298),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_SL g377 ( 
.A(n_340),
.B(n_342),
.Y(n_377)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_311),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_343),
.B(n_347),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_SL g344 ( 
.A(n_296),
.B(n_222),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_344),
.B(n_346),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_288),
.A2(n_147),
.B1(n_126),
.B2(n_129),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_345),
.A2(n_306),
.B1(n_291),
.B2(n_282),
.Y(n_363)
);

CKINVDCx14_ASAP7_75t_R g346 ( 
.A(n_290),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_311),
.Y(n_347)
);

INVx4_ASAP7_75t_L g348 ( 
.A(n_302),
.Y(n_348)
);

AOI22xp33_ASAP7_75t_SL g353 ( 
.A1(n_348),
.A2(n_282),
.B1(n_215),
.B2(n_238),
.Y(n_353)
);

AO21x1_ASAP7_75t_L g349 ( 
.A1(n_295),
.A2(n_292),
.B(n_284),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_341),
.B(n_283),
.C(n_281),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_351),
.B(n_362),
.C(n_364),
.Y(n_391)
);

OAI22x1_ASAP7_75t_SL g352 ( 
.A1(n_320),
.A2(n_297),
.B1(n_292),
.B2(n_294),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_352),
.A2(n_378),
.B1(n_336),
.B2(n_327),
.Y(n_394)
);

HB1xp67_ASAP7_75t_L g413 ( 
.A(n_353),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_316),
.B(n_230),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_360),
.B(n_372),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_341),
.B(n_301),
.C(n_303),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_363),
.A2(n_369),
.B1(n_320),
.B2(n_321),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_325),
.B(n_309),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_336),
.A2(n_314),
.B1(n_296),
.B2(n_147),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_L g370 ( 
.A1(n_343),
.A2(n_180),
.B(n_222),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_370),
.B(n_381),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_344),
.B(n_205),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_325),
.B(n_151),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_374),
.B(n_375),
.C(n_379),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_338),
.B(n_117),
.C(n_100),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_338),
.B(n_113),
.C(n_93),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_319),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_SL g382 ( 
.A(n_329),
.B(n_10),
.C(n_113),
.Y(n_382)
);

MAJx2_ASAP7_75t_L g385 ( 
.A(n_382),
.B(n_317),
.C(n_327),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_337),
.B(n_116),
.C(n_90),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_383),
.B(n_374),
.C(n_375),
.Y(n_407)
);

AO22x1_ASAP7_75t_SL g384 ( 
.A1(n_380),
.A2(n_335),
.B1(n_349),
.B2(n_347),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_384),
.B(n_388),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_385),
.B(n_399),
.Y(n_415)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_367),
.Y(n_386)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_386),
.Y(n_416)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_359),
.Y(n_387)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_387),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_371),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_SL g389 ( 
.A(n_364),
.B(n_323),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_SL g423 ( 
.A(n_389),
.B(n_409),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_361),
.B(n_322),
.Y(n_390)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_390),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_371),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_392),
.B(n_397),
.Y(n_428)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_366),
.Y(n_393)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_393),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_394),
.A2(n_355),
.B1(n_352),
.B2(n_376),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_395),
.A2(n_405),
.B1(n_350),
.B2(n_370),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_356),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_368),
.Y(n_398)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_398),
.Y(n_433)
);

MAJx2_ASAP7_75t_L g399 ( 
.A(n_362),
.B(n_340),
.C(n_315),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_351),
.B(n_333),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_400),
.B(n_382),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_356),
.B(n_330),
.Y(n_401)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_401),
.Y(n_437)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_357),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g436 ( 
.A(n_402),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_373),
.B(n_348),
.Y(n_404)
);

NOR3xp33_ASAP7_75t_L g438 ( 
.A(n_404),
.B(n_411),
.C(n_45),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_369),
.A2(n_349),
.B1(n_321),
.B2(n_328),
.Y(n_405)
);

INVxp33_ASAP7_75t_SL g406 ( 
.A(n_373),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_406),
.B(n_407),
.C(n_408),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_379),
.B(n_318),
.C(n_326),
.Y(n_408)
);

XNOR2x1_ASAP7_75t_L g409 ( 
.A(n_377),
.B(n_345),
.Y(n_409)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_354),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_365),
.B(n_331),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_412),
.B(n_376),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_394),
.A2(n_363),
.B1(n_358),
.B2(n_365),
.Y(n_417)
);

BUFx2_ASAP7_75t_L g457 ( 
.A(n_417),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_419),
.A2(n_422),
.B1(n_42),
.B2(n_1),
.Y(n_458)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_421),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_401),
.A2(n_355),
.B1(n_350),
.B2(n_377),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_SL g425 ( 
.A(n_400),
.B(n_383),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_425),
.B(n_47),
.Y(n_459)
);

OAI22xp33_ASAP7_75t_SL g452 ( 
.A1(n_426),
.A2(n_438),
.B1(n_393),
.B2(n_384),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_427),
.B(n_399),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_391),
.B(n_396),
.C(n_407),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_430),
.B(n_432),
.Y(n_453)
);

NOR2xp67_ASAP7_75t_L g431 ( 
.A(n_391),
.B(n_332),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_431),
.B(n_434),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_L g432 ( 
.A1(n_413),
.A2(n_366),
.B1(n_324),
.B2(n_45),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_396),
.B(n_366),
.C(n_324),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_412),
.B(n_90),
.Y(n_435)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_435),
.Y(n_442)
);

BUFx12_ASAP7_75t_L g439 ( 
.A(n_434),
.Y(n_439)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_439),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_441),
.B(n_459),
.Y(n_477)
);

OAI21xp5_ASAP7_75t_L g443 ( 
.A1(n_414),
.A2(n_403),
.B(n_405),
.Y(n_443)
);

AOI21xp5_ASAP7_75t_SL g472 ( 
.A1(n_443),
.A2(n_423),
.B(n_1),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_SL g444 ( 
.A(n_430),
.B(n_390),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_444),
.B(n_455),
.Y(n_460)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_421),
.Y(n_446)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_446),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_418),
.B(n_408),
.Y(n_447)
);

NOR2xp67_ASAP7_75t_SL g469 ( 
.A(n_447),
.B(n_456),
.Y(n_469)
);

OAI21xp5_ASAP7_75t_SL g448 ( 
.A1(n_428),
.A2(n_384),
.B(n_385),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_448),
.B(n_452),
.Y(n_465)
);

INVx13_ASAP7_75t_L g449 ( 
.A(n_429),
.Y(n_449)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_449),
.Y(n_474)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_421),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_450),
.B(n_451),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_437),
.B(n_395),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_419),
.A2(n_409),
.B1(n_389),
.B2(n_410),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_454),
.A2(n_458),
.B1(n_426),
.B2(n_416),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_436),
.Y(n_455)
);

INVx13_ASAP7_75t_L g456 ( 
.A(n_424),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_459),
.B(n_418),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_462),
.B(n_0),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_464),
.A2(n_467),
.B1(n_442),
.B2(n_443),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_457),
.A2(n_422),
.B1(n_415),
.B2(n_427),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_447),
.B(n_425),
.C(n_415),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_468),
.B(n_471),
.Y(n_484)
);

OAI21xp5_ASAP7_75t_SL g470 ( 
.A1(n_440),
.A2(n_435),
.B(n_423),
.Y(n_470)
);

OR2x2_ASAP7_75t_L g483 ( 
.A(n_470),
.B(n_472),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_L g471 ( 
.A1(n_457),
.A2(n_433),
.B1(n_420),
.B2(n_435),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_445),
.B(n_47),
.C(n_1),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_473),
.B(n_475),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_453),
.B(n_441),
.C(n_439),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_439),
.B(n_47),
.C(n_2),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_476),
.B(n_2),
.C(n_4),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_477),
.B(n_462),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_478),
.B(n_489),
.Y(n_501)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_479),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_475),
.B(n_451),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_480),
.B(n_481),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_461),
.B(n_451),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_464),
.A2(n_440),
.B1(n_450),
.B2(n_446),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_SL g503 ( 
.A1(n_482),
.A2(n_463),
.B1(n_476),
.B2(n_477),
.Y(n_503)
);

CKINVDCx16_ASAP7_75t_R g485 ( 
.A(n_465),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_485),
.B(n_488),
.Y(n_500)
);

AOI21xp5_ASAP7_75t_L g486 ( 
.A1(n_469),
.A2(n_448),
.B(n_454),
.Y(n_486)
);

OAI21xp5_ASAP7_75t_L g502 ( 
.A1(n_486),
.A2(n_487),
.B(n_492),
.Y(n_502)
);

OAI21xp5_ASAP7_75t_SL g487 ( 
.A1(n_460),
.A2(n_442),
.B(n_456),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_474),
.B(n_458),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_L g489 ( 
.A1(n_466),
.A2(n_449),
.B1(n_47),
.B2(n_3),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_491),
.B(n_473),
.Y(n_494)
);

AOI221xp5_ASAP7_75t_L g492 ( 
.A1(n_467),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.C(n_5),
.Y(n_492)
);

HB1xp67_ASAP7_75t_L g495 ( 
.A(n_493),
.Y(n_495)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_494),
.Y(n_509)
);

AOI22xp33_ASAP7_75t_L g496 ( 
.A1(n_490),
.A2(n_463),
.B1(n_472),
.B2(n_470),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_496),
.B(n_498),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_484),
.B(n_468),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g506 ( 
.A(n_503),
.B(n_479),
.Y(n_506)
);

OAI21xp5_ASAP7_75t_L g504 ( 
.A1(n_486),
.A2(n_2),
.B(n_4),
.Y(n_504)
);

OAI21xp5_ASAP7_75t_L g510 ( 
.A1(n_504),
.A2(n_493),
.B(n_7),
.Y(n_510)
);

AOI22xp33_ASAP7_75t_SL g505 ( 
.A1(n_483),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_505),
.B(n_483),
.Y(n_508)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_506),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_499),
.B(n_478),
.C(n_482),
.Y(n_507)
);

INVxp33_ASAP7_75t_L g517 ( 
.A(n_507),
.Y(n_517)
);

AOI21xp5_ASAP7_75t_L g518 ( 
.A1(n_508),
.A2(n_510),
.B(n_6),
.Y(n_518)
);

AOI21x1_ASAP7_75t_L g511 ( 
.A1(n_502),
.A2(n_491),
.B(n_8),
.Y(n_511)
);

OAI21xp5_ASAP7_75t_L g514 ( 
.A1(n_511),
.A2(n_495),
.B(n_513),
.Y(n_514)
);

AOI322xp5_ASAP7_75t_L g512 ( 
.A1(n_497),
.A2(n_6),
.A3(n_8),
.B1(n_9),
.B2(n_500),
.C1(n_496),
.C2(n_501),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_L g515 ( 
.A1(n_512),
.A2(n_495),
.B1(n_509),
.B2(n_507),
.Y(n_515)
);

HB1xp67_ASAP7_75t_L g519 ( 
.A(n_514),
.Y(n_519)
);

NAND3xp33_ASAP7_75t_L g521 ( 
.A(n_515),
.B(n_518),
.C(n_8),
.Y(n_521)
);

NOR2x1_ASAP7_75t_L g520 ( 
.A(n_516),
.B(n_506),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_520),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_L g523 ( 
.A1(n_522),
.A2(n_519),
.B1(n_517),
.B2(n_521),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_523),
.B(n_8),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_524),
.B(n_9),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_525),
.B(n_9),
.Y(n_526)
);


endmodule