module fake_jpeg_14194_n_46 (n_3, n_2, n_1, n_0, n_4, n_5, n_46);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_46;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx20_ASAP7_75t_R g6 ( 
.A(n_2),
.Y(n_6)
);

INVx2_ASAP7_75t_L g7 ( 
.A(n_0),
.Y(n_7)
);

INVx8_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_4),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

INVx8_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

BUFx3_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_6),
.B(n_2),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_13),
.B(n_14),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_6),
.B(n_3),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_16),
.B(n_17),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_17),
.B(n_9),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_19),
.B(n_14),
.C(n_9),
.Y(n_23)
);

CKINVDCx14_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_23),
.B(n_18),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_L g25 ( 
.A1(n_22),
.A2(n_16),
.B1(n_15),
.B2(n_7),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_SL g28 ( 
.A1(n_25),
.A2(n_26),
.B(n_21),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_21),
.B(n_15),
.C(n_16),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_22),
.A2(n_8),
.B1(n_11),
.B2(n_12),
.Y(n_27)
);

OAI22x1_ASAP7_75t_L g31 ( 
.A1(n_27),
.A2(n_11),
.B1(n_8),
.B2(n_10),
.Y(n_31)
);

AOI21xp5_ASAP7_75t_L g35 ( 
.A1(n_28),
.A2(n_29),
.B(n_31),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_32),
.C(n_19),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_25),
.B(n_18),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_36),
.C(n_10),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_31),
.A2(n_20),
.B1(n_8),
.B2(n_11),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_34),
.Y(n_37)
);

MAJx2_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_5),
.C(n_4),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_38),
.B(n_39),
.C(n_10),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g39 ( 
.A1(n_35),
.A2(n_5),
.B(n_4),
.Y(n_39)
);

AOI22x1_ASAP7_75t_L g40 ( 
.A1(n_37),
.A2(n_36),
.B1(n_10),
.B2(n_5),
.Y(n_40)
);

AND2x2_ASAP7_75t_SL g42 ( 
.A(n_40),
.B(n_41),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_41),
.B(n_0),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_43),
.A2(n_8),
.B1(n_11),
.B2(n_42),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_44),
.B(n_12),
.C(n_0),
.Y(n_45)
);

AOI221xp5_ASAP7_75t_L g46 ( 
.A1(n_45),
.A2(n_0),
.B1(n_1),
.B2(n_12),
.C(n_20),
.Y(n_46)
);


endmodule