module fake_aes_10816_n_739 (n_117, n_44, n_133, n_149, n_81, n_69, n_185, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_125, n_9, n_161, n_10, n_177, n_130, n_103, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_154, n_7, n_29, n_165, n_146, n_45, n_85, n_181, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_139, n_16, n_13, n_169, n_152, n_113, n_95, n_124, n_156, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_38, n_64, n_142, n_184, n_46, n_31, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_12, n_86, n_143, n_182, n_166, n_162, n_186, n_75, n_163, n_105, n_159, n_174, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_67, n_77, n_20, n_2, n_147, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_150, n_168, n_3, n_18, n_110, n_66, n_134, n_1, n_164, n_82, n_106, n_175, n_15, n_173, n_145, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_96, n_39, n_739);
input n_117;
input n_44;
input n_133;
input n_149;
input n_81;
input n_69;
input n_185;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_125;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_103;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_154;
input n_7;
input n_29;
input n_165;
input n_146;
input n_45;
input n_85;
input n_181;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_139;
input n_16;
input n_13;
input n_169;
input n_152;
input n_113;
input n_95;
input n_124;
input n_156;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_38;
input n_64;
input n_142;
input n_184;
input n_46;
input n_31;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_12;
input n_86;
input n_143;
input n_182;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_105;
input n_159;
input n_174;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_67;
input n_77;
input n_20;
input n_2;
input n_147;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_150;
input n_168;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_1;
input n_164;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_145;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_96;
input n_39;
output n_739;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_607;
wire n_431;
wire n_484;
wire n_496;
wire n_667;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_202;
wire n_386;
wire n_432;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_678;
wire n_387;
wire n_434;
wire n_384;
wire n_227;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_489;
wire n_732;
wire n_199;
wire n_351;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_560;
wire n_517;
wire n_479;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_712;
wire n_447;
wire n_608;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_393;
wire n_247;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_329;
wire n_251;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_207;
wire n_565;
wire n_224;
wire n_219;
wire n_475;
wire n_578;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_673;
wire n_669;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_295;
wire n_654;
wire n_263;
wire n_495;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_449;
wire n_300;
wire n_734;
wire n_524;
wire n_584;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_602;
wire n_198;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_297;
wire n_410;
wire n_377;
wire n_510;
wire n_343;
wire n_675;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_375;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_521;
wire n_695;
wire n_650;
wire n_625;
wire n_469;
wire n_585;
wire n_713;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_736;
wire n_194;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_421;
wire n_709;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g189 ( .A(n_50), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_16), .Y(n_190) );
CKINVDCx5p33_ASAP7_75t_R g191 ( .A(n_75), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_168), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_147), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_41), .Y(n_194) );
BUFx3_ASAP7_75t_L g195 ( .A(n_83), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_82), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_181), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_109), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_169), .Y(n_199) );
BUFx6f_ASAP7_75t_L g200 ( .A(n_114), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_166), .Y(n_201) );
CKINVDCx5p33_ASAP7_75t_R g202 ( .A(n_127), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_129), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_176), .Y(n_204) );
CKINVDCx20_ASAP7_75t_R g205 ( .A(n_145), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_4), .Y(n_206) );
CKINVDCx5p33_ASAP7_75t_R g207 ( .A(n_3), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_175), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_52), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_105), .Y(n_210) );
BUFx6f_ASAP7_75t_L g211 ( .A(n_79), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_143), .Y(n_212) );
CKINVDCx5p33_ASAP7_75t_R g213 ( .A(n_136), .Y(n_213) );
INVxp67_ASAP7_75t_L g214 ( .A(n_31), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_163), .Y(n_215) );
CKINVDCx20_ASAP7_75t_R g216 ( .A(n_22), .Y(n_216) );
CKINVDCx16_ASAP7_75t_R g217 ( .A(n_111), .Y(n_217) );
CKINVDCx5p33_ASAP7_75t_R g218 ( .A(n_187), .Y(n_218) );
CKINVDCx5p33_ASAP7_75t_R g219 ( .A(n_100), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_164), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_86), .Y(n_221) );
CKINVDCx5p33_ASAP7_75t_R g222 ( .A(n_22), .Y(n_222) );
BUFx3_ASAP7_75t_L g223 ( .A(n_30), .Y(n_223) );
INVxp67_ASAP7_75t_L g224 ( .A(n_113), .Y(n_224) );
CKINVDCx5p33_ASAP7_75t_R g225 ( .A(n_16), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_43), .Y(n_226) );
CKINVDCx5p33_ASAP7_75t_R g227 ( .A(n_155), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_126), .Y(n_228) );
CKINVDCx5p33_ASAP7_75t_R g229 ( .A(n_148), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_99), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_69), .Y(n_231) );
CKINVDCx20_ASAP7_75t_R g232 ( .A(n_56), .Y(n_232) );
BUFx3_ASAP7_75t_L g233 ( .A(n_118), .Y(n_233) );
CKINVDCx5p33_ASAP7_75t_R g234 ( .A(n_123), .Y(n_234) );
CKINVDCx5p33_ASAP7_75t_R g235 ( .A(n_77), .Y(n_235) );
CKINVDCx5p33_ASAP7_75t_R g236 ( .A(n_2), .Y(n_236) );
NOR2xp67_ASAP7_75t_L g237 ( .A(n_133), .B(n_9), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_44), .Y(n_238) );
INVxp67_ASAP7_75t_SL g239 ( .A(n_146), .Y(n_239) );
CKINVDCx5p33_ASAP7_75t_R g240 ( .A(n_141), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_182), .Y(n_241) );
INVx2_ASAP7_75t_L g242 ( .A(n_74), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_53), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_48), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_1), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_24), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_94), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_179), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_49), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_68), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_64), .Y(n_251) );
CKINVDCx5p33_ASAP7_75t_R g252 ( .A(n_87), .Y(n_252) );
CKINVDCx5p33_ASAP7_75t_R g253 ( .A(n_85), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_170), .Y(n_254) );
CKINVDCx14_ASAP7_75t_R g255 ( .A(n_42), .Y(n_255) );
CKINVDCx20_ASAP7_75t_R g256 ( .A(n_89), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_93), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_177), .Y(n_258) );
CKINVDCx5p33_ASAP7_75t_R g259 ( .A(n_27), .Y(n_259) );
CKINVDCx5p33_ASAP7_75t_R g260 ( .A(n_122), .Y(n_260) );
CKINVDCx20_ASAP7_75t_R g261 ( .A(n_51), .Y(n_261) );
INVxp67_ASAP7_75t_SL g262 ( .A(n_185), .Y(n_262) );
BUFx3_ASAP7_75t_L g263 ( .A(n_90), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_183), .Y(n_264) );
BUFx6f_ASAP7_75t_L g265 ( .A(n_120), .Y(n_265) );
INVxp33_ASAP7_75t_L g266 ( .A(n_47), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_46), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_0), .Y(n_268) );
CKINVDCx5p33_ASAP7_75t_R g269 ( .A(n_32), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_62), .Y(n_270) );
CKINVDCx5p33_ASAP7_75t_R g271 ( .A(n_67), .Y(n_271) );
BUFx3_ASAP7_75t_L g272 ( .A(n_125), .Y(n_272) );
HB1xp67_ASAP7_75t_L g273 ( .A(n_149), .Y(n_273) );
INVx2_ASAP7_75t_L g274 ( .A(n_95), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_132), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_178), .Y(n_276) );
CKINVDCx5p33_ASAP7_75t_R g277 ( .A(n_11), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_165), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_25), .Y(n_279) );
BUFx6f_ASAP7_75t_L g280 ( .A(n_24), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_9), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_172), .Y(n_282) );
CKINVDCx20_ASAP7_75t_R g283 ( .A(n_19), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_58), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_116), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_142), .Y(n_286) );
CKINVDCx20_ASAP7_75t_R g287 ( .A(n_110), .Y(n_287) );
CKINVDCx5p33_ASAP7_75t_R g288 ( .A(n_76), .Y(n_288) );
AND2x2_ASAP7_75t_L g289 ( .A(n_266), .B(n_0), .Y(n_289) );
AND2x2_ASAP7_75t_L g290 ( .A(n_266), .B(n_1), .Y(n_290) );
BUFx8_ASAP7_75t_L g291 ( .A(n_280), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_212), .Y(n_292) );
AND2x4_ASAP7_75t_L g293 ( .A(n_273), .B(n_2), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_242), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_258), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_274), .Y(n_296) );
BUFx3_ASAP7_75t_L g297 ( .A(n_195), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_195), .Y(n_298) );
AND2x4_ASAP7_75t_L g299 ( .A(n_273), .B(n_3), .Y(n_299) );
HB1xp67_ASAP7_75t_L g300 ( .A(n_207), .Y(n_300) );
BUFx6f_ASAP7_75t_L g301 ( .A(n_200), .Y(n_301) );
INVx2_ASAP7_75t_SL g302 ( .A(n_223), .Y(n_302) );
INVx3_ASAP7_75t_L g303 ( .A(n_280), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_206), .Y(n_304) );
HB1xp67_ASAP7_75t_L g305 ( .A(n_222), .Y(n_305) );
INVx4_ASAP7_75t_L g306 ( .A(n_223), .Y(n_306) );
OAI22xp5_ASAP7_75t_R g307 ( .A1(n_225), .A2(n_4), .B1(n_5), .B2(n_6), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_189), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_190), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_233), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_245), .B(n_5), .Y(n_311) );
AOI22xp5_ASAP7_75t_L g312 ( .A1(n_217), .A2(n_6), .B1(n_7), .B2(n_8), .Y(n_312) );
CKINVDCx5p33_ASAP7_75t_R g313 ( .A(n_255), .Y(n_313) );
BUFx6f_ASAP7_75t_L g314 ( .A(n_200), .Y(n_314) );
AND2x2_ASAP7_75t_L g315 ( .A(n_255), .B(n_7), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_246), .B(n_8), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_301), .Y(n_317) );
NOR2xp33_ASAP7_75t_L g318 ( .A(n_308), .B(n_214), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_289), .Y(n_319) );
BUFx6f_ASAP7_75t_L g320 ( .A(n_301), .Y(n_320) );
INVx3_ASAP7_75t_L g321 ( .A(n_306), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_301), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_289), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_290), .Y(n_324) );
AND2x6_ASAP7_75t_L g325 ( .A(n_293), .B(n_233), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_300), .B(n_236), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_301), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_290), .Y(n_328) );
NAND3xp33_ASAP7_75t_L g329 ( .A(n_293), .B(n_299), .C(n_291), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_292), .Y(n_330) );
AND2x2_ASAP7_75t_L g331 ( .A(n_305), .B(n_277), .Y(n_331) );
NAND2xp5_ASAP7_75t_SL g332 ( .A(n_306), .B(n_192), .Y(n_332) );
INVx1_ASAP7_75t_SL g333 ( .A(n_315), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_306), .B(n_214), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_301), .Y(n_335) );
INVx4_ASAP7_75t_L g336 ( .A(n_293), .Y(n_336) );
NAND2xp5_ASAP7_75t_SL g337 ( .A(n_298), .B(n_193), .Y(n_337) );
BUFx2_ASAP7_75t_L g338 ( .A(n_313), .Y(n_338) );
AND2x2_ASAP7_75t_L g339 ( .A(n_313), .B(n_239), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_302), .B(n_224), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_319), .B(n_299), .Y(n_341) );
INVx2_ASAP7_75t_SL g342 ( .A(n_325), .Y(n_342) );
NAND2xp5_ASAP7_75t_SL g343 ( .A(n_329), .B(n_299), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_323), .B(n_315), .Y(n_344) );
NAND2xp5_ASAP7_75t_SL g345 ( .A(n_336), .B(n_194), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_324), .B(n_297), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_328), .B(n_309), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_318), .B(n_297), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_318), .B(n_302), .Y(n_349) );
OR2x2_ASAP7_75t_L g350 ( .A(n_326), .B(n_311), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_330), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_333), .B(n_294), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_336), .B(n_294), .Y(n_353) );
NOR2xp33_ASAP7_75t_L g354 ( .A(n_339), .B(n_304), .Y(n_354) );
INVxp67_ASAP7_75t_L g355 ( .A(n_331), .Y(n_355) );
AND2x2_ASAP7_75t_SL g356 ( .A(n_338), .B(n_312), .Y(n_356) );
NOR2xp33_ASAP7_75t_L g357 ( .A(n_340), .B(n_334), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_325), .B(n_295), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_325), .B(n_296), .Y(n_359) );
AOI22xp5_ASAP7_75t_L g360 ( .A1(n_325), .A2(n_232), .B1(n_256), .B2(n_205), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_325), .B(n_296), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_321), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_325), .B(n_316), .Y(n_363) );
NAND2xp5_ASAP7_75t_SL g364 ( .A(n_321), .B(n_196), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_321), .Y(n_365) );
BUFx6f_ASAP7_75t_L g366 ( .A(n_320), .Y(n_366) );
NAND2xp5_ASAP7_75t_SL g367 ( .A(n_342), .B(n_191), .Y(n_367) );
CKINVDCx5p33_ASAP7_75t_R g368 ( .A(n_360), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_362), .Y(n_369) );
BUFx3_ASAP7_75t_L g370 ( .A(n_347), .Y(n_370) );
AOI21xp5_ASAP7_75t_L g371 ( .A1(n_343), .A2(n_332), .B(n_337), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_357), .B(n_332), .Y(n_372) );
INVxp67_ASAP7_75t_L g373 ( .A(n_350), .Y(n_373) );
AOI22xp5_ASAP7_75t_L g374 ( .A1(n_355), .A2(n_261), .B1(n_287), .B2(n_337), .Y(n_374) );
OAI22xp5_ASAP7_75t_L g375 ( .A1(n_363), .A2(n_283), .B1(n_216), .B2(n_262), .Y(n_375) );
OAI21xp33_ASAP7_75t_SL g376 ( .A1(n_341), .A2(n_279), .B(n_268), .Y(n_376) );
O2A1O1Ixp33_ASAP7_75t_L g377 ( .A1(n_344), .A2(n_281), .B(n_310), .C(n_224), .Y(n_377) );
NOR2xp67_ASAP7_75t_L g378 ( .A(n_354), .B(n_10), .Y(n_378) );
AOI22x1_ASAP7_75t_L g379 ( .A1(n_362), .A2(n_310), .B1(n_314), .B2(n_317), .Y(n_379) );
AOI21xp5_ASAP7_75t_L g380 ( .A1(n_345), .A2(n_198), .B(n_197), .Y(n_380) );
NOR2xp67_ASAP7_75t_L g381 ( .A(n_347), .B(n_10), .Y(n_381) );
NOR2xp67_ASAP7_75t_L g382 ( .A(n_352), .B(n_11), .Y(n_382) );
OAI22xp5_ASAP7_75t_L g383 ( .A1(n_348), .A2(n_346), .B1(n_351), .B2(n_349), .Y(n_383) );
AOI22xp33_ASAP7_75t_SL g384 ( .A1(n_356), .A2(n_307), .B1(n_291), .B2(n_280), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_353), .B(n_291), .Y(n_385) );
AOI21x1_ASAP7_75t_L g386 ( .A1(n_364), .A2(n_322), .B(n_317), .Y(n_386) );
OAI22xp5_ASAP7_75t_L g387 ( .A1(n_356), .A2(n_237), .B1(n_201), .B2(n_203), .Y(n_387) );
O2A1O1Ixp33_ASAP7_75t_L g388 ( .A1(n_364), .A2(n_204), .B(n_208), .C(n_199), .Y(n_388) );
AO32x1_ASAP7_75t_L g389 ( .A1(n_342), .A2(n_249), .A3(n_209), .B1(n_210), .B2(n_215), .Y(n_389) );
AOI21xp5_ASAP7_75t_L g390 ( .A1(n_365), .A2(n_221), .B(n_220), .Y(n_390) );
AOI22x1_ASAP7_75t_L g391 ( .A1(n_365), .A2(n_314), .B1(n_327), .B2(n_322), .Y(n_391) );
NAND2xp5_ASAP7_75t_SL g392 ( .A(n_373), .B(n_358), .Y(n_392) );
OAI21xp5_ASAP7_75t_L g393 ( .A1(n_371), .A2(n_361), .B(n_359), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_370), .Y(n_394) );
A2O1A1Ixp33_ASAP7_75t_L g395 ( .A1(n_381), .A2(n_248), .B(n_250), .C(n_226), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_369), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_383), .B(n_280), .Y(n_397) );
AOI21xp5_ASAP7_75t_L g398 ( .A1(n_372), .A2(n_366), .B(n_228), .Y(n_398) );
AO31x2_ASAP7_75t_L g399 ( .A1(n_383), .A2(n_264), .A3(n_238), .B(n_241), .Y(n_399) );
NOR2xp33_ASAP7_75t_L g400 ( .A(n_368), .B(n_307), .Y(n_400) );
AOI21xp5_ASAP7_75t_L g401 ( .A1(n_385), .A2(n_366), .B(n_231), .Y(n_401) );
OAI22xp5_ASAP7_75t_L g402 ( .A1(n_382), .A2(n_259), .B1(n_202), .B2(n_218), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_376), .Y(n_403) );
A2O1A1Ixp33_ASAP7_75t_L g404 ( .A1(n_377), .A2(n_244), .B(n_267), .C(n_230), .Y(n_404) );
OAI21x1_ASAP7_75t_L g405 ( .A1(n_386), .A2(n_247), .B(n_243), .Y(n_405) );
BUFx6f_ASAP7_75t_L g406 ( .A(n_367), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g407 ( .A1(n_384), .A2(n_275), .B1(n_251), .B2(n_254), .Y(n_407) );
NAND2xp33_ASAP7_75t_L g408 ( .A(n_374), .B(n_213), .Y(n_408) );
OR2x6_ASAP7_75t_L g409 ( .A(n_375), .B(n_257), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_378), .Y(n_410) );
BUFx12f_ASAP7_75t_L g411 ( .A(n_387), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_387), .B(n_12), .Y(n_412) );
AOI21xp5_ASAP7_75t_SL g413 ( .A1(n_388), .A2(n_272), .B(n_263), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_379), .Y(n_414) );
OAI21xp5_ASAP7_75t_SL g415 ( .A1(n_380), .A2(n_276), .B(n_270), .Y(n_415) );
INVx3_ASAP7_75t_L g416 ( .A(n_390), .Y(n_416) );
INVxp67_ASAP7_75t_SL g417 ( .A(n_391), .Y(n_417) );
AOI221xp5_ASAP7_75t_L g418 ( .A1(n_389), .A2(n_278), .B1(n_282), .B2(n_284), .C(n_285), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_389), .Y(n_419) );
AOI221xp5_ASAP7_75t_SL g420 ( .A1(n_383), .A2(n_286), .B1(n_303), .B2(n_200), .C(n_265), .Y(n_420) );
BUFx6f_ASAP7_75t_L g421 ( .A(n_370), .Y(n_421) );
AOI22xp33_ASAP7_75t_L g422 ( .A1(n_411), .A2(n_200), .B1(n_211), .B2(n_265), .Y(n_422) );
OA21x2_ASAP7_75t_L g423 ( .A1(n_420), .A2(n_335), .B(n_327), .Y(n_423) );
AO21x2_ASAP7_75t_L g424 ( .A1(n_419), .A2(n_335), .B(n_314), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_409), .B(n_12), .Y(n_425) );
BUFx6f_ASAP7_75t_L g426 ( .A(n_421), .Y(n_426) );
AOI22xp33_ASAP7_75t_L g427 ( .A1(n_409), .A2(n_211), .B1(n_265), .B2(n_303), .Y(n_427) );
OA21x2_ASAP7_75t_L g428 ( .A1(n_420), .A2(n_227), .B(n_219), .Y(n_428) );
AO31x2_ASAP7_75t_L g429 ( .A1(n_397), .A2(n_314), .A3(n_265), .B(n_211), .Y(n_429) );
OA21x2_ASAP7_75t_L g430 ( .A1(n_405), .A2(n_234), .B(n_229), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_403), .Y(n_431) );
OAI22xp5_ASAP7_75t_L g432 ( .A1(n_409), .A2(n_211), .B1(n_303), .B2(n_288), .Y(n_432) );
NOR2xp33_ASAP7_75t_L g433 ( .A(n_400), .B(n_235), .Y(n_433) );
BUFx6f_ASAP7_75t_L g434 ( .A(n_406), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_394), .Y(n_435) );
AO31x2_ASAP7_75t_L g436 ( .A1(n_414), .A2(n_314), .A3(n_320), .B(n_15), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_412), .B(n_13), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_396), .Y(n_438) );
NOR2xp33_ASAP7_75t_L g439 ( .A(n_407), .B(n_240), .Y(n_439) );
AOI21xp5_ASAP7_75t_L g440 ( .A1(n_398), .A2(n_253), .B(n_252), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_404), .B(n_13), .Y(n_441) );
OAI21x1_ASAP7_75t_L g442 ( .A1(n_416), .A2(n_104), .B(n_188), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_416), .Y(n_443) );
AND2x4_ASAP7_75t_L g444 ( .A(n_410), .B(n_14), .Y(n_444) );
OAI22xp5_ASAP7_75t_L g445 ( .A1(n_415), .A2(n_271), .B1(n_269), .B2(n_260), .Y(n_445) );
INVx2_ASAP7_75t_SL g446 ( .A(n_406), .Y(n_446) );
HB1xp67_ASAP7_75t_L g447 ( .A(n_399), .Y(n_447) );
INVx3_ASAP7_75t_L g448 ( .A(n_406), .Y(n_448) );
OAI21x1_ASAP7_75t_L g449 ( .A1(n_393), .A2(n_102), .B(n_186), .Y(n_449) );
AO21x2_ASAP7_75t_L g450 ( .A1(n_395), .A2(n_101), .B(n_184), .Y(n_450) );
HB1xp67_ASAP7_75t_L g451 ( .A(n_399), .Y(n_451) );
INVx2_ASAP7_75t_SL g452 ( .A(n_392), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_408), .B(n_15), .Y(n_453) );
AOI21xp33_ASAP7_75t_L g454 ( .A1(n_402), .A2(n_17), .B(n_18), .Y(n_454) );
NAND2x1p5_ASAP7_75t_L g455 ( .A(n_401), .B(n_20), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_418), .A2(n_20), .B1(n_21), .B2(n_23), .Y(n_456) );
AOI21xp5_ASAP7_75t_L g457 ( .A1(n_413), .A2(n_106), .B(n_180), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_403), .Y(n_458) );
AO31x2_ASAP7_75t_L g459 ( .A1(n_419), .A2(n_21), .A3(n_23), .B(n_25), .Y(n_459) );
AOI21xp5_ASAP7_75t_L g460 ( .A1(n_417), .A2(n_107), .B(n_28), .Y(n_460) );
OR2x2_ASAP7_75t_L g461 ( .A(n_409), .B(n_26), .Y(n_461) );
NOR2xp33_ASAP7_75t_L g462 ( .A(n_411), .B(n_29), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_403), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_403), .Y(n_464) );
OA21x2_ASAP7_75t_L g465 ( .A1(n_420), .A2(n_33), .B(n_34), .Y(n_465) );
OA21x2_ASAP7_75t_L g466 ( .A1(n_420), .A2(n_35), .B(n_36), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_424), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_435), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_438), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_431), .Y(n_470) );
INVx3_ASAP7_75t_L g471 ( .A(n_426), .Y(n_471) );
INVx2_ASAP7_75t_SL g472 ( .A(n_426), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_458), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_437), .B(n_37), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_463), .Y(n_475) );
AO21x2_ASAP7_75t_L g476 ( .A1(n_424), .A2(n_38), .B(n_39), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_461), .B(n_40), .Y(n_477) );
OR2x2_ASAP7_75t_L g478 ( .A(n_425), .B(n_174), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_464), .B(n_45), .Y(n_479) );
HB1xp67_ASAP7_75t_L g480 ( .A(n_447), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_443), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_444), .Y(n_482) );
AO21x2_ASAP7_75t_L g483 ( .A1(n_451), .A2(n_54), .B(n_55), .Y(n_483) );
HB1xp67_ASAP7_75t_L g484 ( .A(n_429), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_459), .Y(n_485) );
INVx3_ASAP7_75t_L g486 ( .A(n_434), .Y(n_486) );
INVx2_ASAP7_75t_L g487 ( .A(n_423), .Y(n_487) );
AO21x2_ASAP7_75t_L g488 ( .A1(n_449), .A2(n_57), .B(n_59), .Y(n_488) );
OAI21x1_ASAP7_75t_L g489 ( .A1(n_442), .A2(n_60), .B(n_61), .Y(n_489) );
INVx2_ASAP7_75t_SL g490 ( .A(n_434), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_459), .Y(n_491) );
AND2x4_ASAP7_75t_L g492 ( .A(n_446), .B(n_63), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_459), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_429), .Y(n_494) );
OR2x6_ASAP7_75t_L g495 ( .A(n_432), .B(n_65), .Y(n_495) );
INVxp67_ASAP7_75t_SL g496 ( .A(n_423), .Y(n_496) );
INVx2_ASAP7_75t_L g497 ( .A(n_429), .Y(n_497) );
OAI22xp33_ASAP7_75t_L g498 ( .A1(n_432), .A2(n_66), .B1(n_70), .B2(n_71), .Y(n_498) );
INVx3_ASAP7_75t_L g499 ( .A(n_434), .Y(n_499) );
OR2x2_ASAP7_75t_L g500 ( .A(n_448), .B(n_72), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_436), .Y(n_501) );
OR2x6_ASAP7_75t_L g502 ( .A(n_452), .B(n_73), .Y(n_502) );
OR2x2_ASAP7_75t_L g503 ( .A(n_448), .B(n_78), .Y(n_503) );
HB1xp67_ASAP7_75t_L g504 ( .A(n_428), .Y(n_504) );
HB1xp67_ASAP7_75t_L g505 ( .A(n_428), .Y(n_505) );
AOI21x1_ASAP7_75t_L g506 ( .A1(n_465), .A2(n_173), .B(n_80), .Y(n_506) );
INVx2_ASAP7_75t_L g507 ( .A(n_436), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_455), .Y(n_508) );
AND2x4_ASAP7_75t_L g509 ( .A(n_450), .B(n_81), .Y(n_509) );
OA21x2_ASAP7_75t_L g510 ( .A1(n_457), .A2(n_84), .B(n_88), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_441), .Y(n_511) );
BUFx4f_ASAP7_75t_SL g512 ( .A(n_462), .Y(n_512) );
AO21x2_ASAP7_75t_L g513 ( .A1(n_453), .A2(n_91), .B(n_92), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_436), .Y(n_514) );
INVx3_ASAP7_75t_L g515 ( .A(n_430), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_456), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_465), .B(n_96), .Y(n_517) );
NAND2xp33_ASAP7_75t_R g518 ( .A(n_466), .B(n_97), .Y(n_518) );
BUFx4f_ASAP7_75t_L g519 ( .A(n_466), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_450), .Y(n_520) );
OR2x2_ASAP7_75t_L g521 ( .A(n_445), .B(n_171), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_454), .Y(n_522) );
BUFx4f_ASAP7_75t_SL g523 ( .A(n_422), .Y(n_523) );
BUFx3_ASAP7_75t_L g524 ( .A(n_445), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_427), .Y(n_525) );
AO21x2_ASAP7_75t_L g526 ( .A1(n_460), .A2(n_98), .B(n_103), .Y(n_526) );
BUFx6f_ASAP7_75t_L g527 ( .A(n_439), .Y(n_527) );
OR2x2_ASAP7_75t_L g528 ( .A(n_433), .B(n_167), .Y(n_528) );
AO21x2_ASAP7_75t_L g529 ( .A1(n_440), .A2(n_108), .B(n_112), .Y(n_529) );
AND2x4_ASAP7_75t_L g530 ( .A(n_426), .B(n_115), .Y(n_530) );
BUFx6f_ASAP7_75t_L g531 ( .A(n_426), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_437), .B(n_117), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_435), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_435), .Y(n_534) );
HB1xp67_ASAP7_75t_L g535 ( .A(n_480), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_470), .B(n_119), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_468), .Y(n_537) );
INVx2_ASAP7_75t_L g538 ( .A(n_481), .Y(n_538) );
HB1xp67_ASAP7_75t_L g539 ( .A(n_480), .Y(n_539) );
HB1xp67_ASAP7_75t_L g540 ( .A(n_484), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_533), .B(n_121), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_534), .B(n_124), .Y(n_542) );
INVxp67_ASAP7_75t_SL g543 ( .A(n_484), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_474), .B(n_128), .Y(n_544) );
OR2x2_ASAP7_75t_L g545 ( .A(n_469), .B(n_130), .Y(n_545) );
HB1xp67_ASAP7_75t_L g546 ( .A(n_497), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_473), .Y(n_547) );
INVx2_ASAP7_75t_L g548 ( .A(n_497), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_475), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_511), .B(n_131), .Y(n_550) );
OR2x2_ASAP7_75t_L g551 ( .A(n_524), .B(n_134), .Y(n_551) );
HB1xp67_ASAP7_75t_L g552 ( .A(n_494), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_532), .B(n_135), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_482), .Y(n_554) );
AOI22xp33_ASAP7_75t_SL g555 ( .A1(n_524), .A2(n_137), .B1(n_138), .B2(n_139), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_479), .Y(n_556) );
AND2x4_ASAP7_75t_L g557 ( .A(n_495), .B(n_140), .Y(n_557) );
INVx2_ASAP7_75t_L g558 ( .A(n_487), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_477), .B(n_144), .Y(n_559) );
INVx2_ASAP7_75t_L g560 ( .A(n_487), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_485), .Y(n_561) );
INVx3_ASAP7_75t_L g562 ( .A(n_495), .Y(n_562) );
BUFx2_ASAP7_75t_L g563 ( .A(n_495), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_522), .B(n_150), .Y(n_564) );
HB1xp67_ASAP7_75t_L g565 ( .A(n_467), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_527), .B(n_151), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_491), .Y(n_567) );
AND2x4_ASAP7_75t_L g568 ( .A(n_486), .B(n_152), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_493), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_527), .B(n_153), .Y(n_570) );
OR2x2_ASAP7_75t_L g571 ( .A(n_527), .B(n_154), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_508), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_502), .Y(n_573) );
INVx2_ASAP7_75t_SL g574 ( .A(n_531), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_516), .B(n_156), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_492), .B(n_157), .Y(n_576) );
INVx2_ASAP7_75t_SL g577 ( .A(n_531), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_500), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_503), .Y(n_579) );
HB1xp67_ASAP7_75t_L g580 ( .A(n_467), .Y(n_580) );
OR2x2_ASAP7_75t_L g581 ( .A(n_472), .B(n_162), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_492), .B(n_158), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_525), .B(n_159), .Y(n_583) );
INVx2_ASAP7_75t_L g584 ( .A(n_501), .Y(n_584) );
AND2x4_ASAP7_75t_L g585 ( .A(n_486), .B(n_160), .Y(n_585) );
OR2x2_ASAP7_75t_L g586 ( .A(n_478), .B(n_490), .Y(n_586) );
AND2x4_ASAP7_75t_L g587 ( .A(n_499), .B(n_161), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_515), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_515), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_501), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_507), .Y(n_591) );
INVx4_ASAP7_75t_L g592 ( .A(n_531), .Y(n_592) );
AND2x2_ASAP7_75t_L g593 ( .A(n_521), .B(n_471), .Y(n_593) );
HB1xp67_ASAP7_75t_L g594 ( .A(n_507), .Y(n_594) );
INVx2_ASAP7_75t_L g595 ( .A(n_514), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_514), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_499), .B(n_471), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_504), .B(n_505), .Y(n_598) );
AND2x2_ASAP7_75t_L g599 ( .A(n_528), .B(n_530), .Y(n_599) );
INVx2_ASAP7_75t_SL g600 ( .A(n_512), .Y(n_600) );
AND2x4_ASAP7_75t_L g601 ( .A(n_509), .B(n_504), .Y(n_601) );
AND2x2_ASAP7_75t_L g602 ( .A(n_561), .B(n_520), .Y(n_602) );
AND2x2_ASAP7_75t_L g603 ( .A(n_567), .B(n_496), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_569), .B(n_496), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_537), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_538), .B(n_483), .Y(n_606) );
OR2x2_ASAP7_75t_L g607 ( .A(n_535), .B(n_483), .Y(n_607) );
INVx2_ASAP7_75t_L g608 ( .A(n_558), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_547), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_549), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_554), .Y(n_611) );
NOR2x1_ASAP7_75t_L g612 ( .A(n_557), .B(n_498), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_572), .B(n_523), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_535), .Y(n_614) );
AND2x2_ASAP7_75t_L g615 ( .A(n_588), .B(n_509), .Y(n_615) );
HB1xp67_ASAP7_75t_L g616 ( .A(n_539), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_539), .Y(n_617) );
OR2x2_ASAP7_75t_L g618 ( .A(n_563), .B(n_476), .Y(n_618) );
AND2x2_ASAP7_75t_L g619 ( .A(n_589), .B(n_476), .Y(n_619) );
AND2x4_ASAP7_75t_L g620 ( .A(n_562), .B(n_513), .Y(n_620) );
INVx2_ASAP7_75t_SL g621 ( .A(n_592), .Y(n_621) );
HB1xp67_ASAP7_75t_L g622 ( .A(n_540), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_573), .Y(n_623) );
AND2x2_ASAP7_75t_L g624 ( .A(n_591), .B(n_519), .Y(n_624) );
AND2x2_ASAP7_75t_L g625 ( .A(n_596), .B(n_519), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_548), .B(n_513), .Y(n_626) );
INVx2_ASAP7_75t_L g627 ( .A(n_560), .Y(n_627) );
AND2x2_ASAP7_75t_L g628 ( .A(n_584), .B(n_529), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_578), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_556), .B(n_517), .Y(n_630) );
BUFx2_ASAP7_75t_L g631 ( .A(n_562), .Y(n_631) );
INVx3_ASAP7_75t_L g632 ( .A(n_601), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_579), .Y(n_633) );
AND2x2_ASAP7_75t_L g634 ( .A(n_590), .B(n_595), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_586), .B(n_488), .Y(n_635) );
NAND2x1p5_ASAP7_75t_L g636 ( .A(n_557), .B(n_489), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_597), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_599), .B(n_526), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_540), .Y(n_639) );
OR2x2_ASAP7_75t_L g640 ( .A(n_598), .B(n_526), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_593), .B(n_510), .Y(n_641) );
AND2x2_ASAP7_75t_L g642 ( .A(n_565), .B(n_506), .Y(n_642) );
HB1xp67_ASAP7_75t_L g643 ( .A(n_565), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_598), .Y(n_644) );
HB1xp67_ASAP7_75t_L g645 ( .A(n_580), .Y(n_645) );
INVx2_ASAP7_75t_L g646 ( .A(n_580), .Y(n_646) );
INVx1_ASAP7_75t_SL g647 ( .A(n_600), .Y(n_647) );
AND2x2_ASAP7_75t_L g648 ( .A(n_601), .B(n_510), .Y(n_648) );
AND2x2_ASAP7_75t_L g649 ( .A(n_601), .B(n_518), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_583), .B(n_542), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_605), .Y(n_651) );
OR2x2_ASAP7_75t_L g652 ( .A(n_644), .B(n_543), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_629), .B(n_543), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_633), .B(n_546), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_609), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_610), .Y(n_656) );
AND2x2_ASAP7_75t_L g657 ( .A(n_623), .B(n_546), .Y(n_657) );
INVx2_ASAP7_75t_L g658 ( .A(n_643), .Y(n_658) );
OR2x2_ASAP7_75t_L g659 ( .A(n_616), .B(n_552), .Y(n_659) );
AOI22xp5_ASAP7_75t_L g660 ( .A1(n_612), .A2(n_555), .B1(n_582), .B2(n_576), .Y(n_660) );
AND2x2_ASAP7_75t_L g661 ( .A(n_632), .B(n_577), .Y(n_661) );
AOI21xp5_ASAP7_75t_L g662 ( .A1(n_636), .A2(n_552), .B(n_574), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_611), .Y(n_663) );
AND2x2_ASAP7_75t_L g664 ( .A(n_632), .B(n_594), .Y(n_664) );
AND2x2_ASAP7_75t_L g665 ( .A(n_649), .B(n_594), .Y(n_665) );
AND2x2_ASAP7_75t_L g666 ( .A(n_649), .B(n_570), .Y(n_666) );
AND2x2_ASAP7_75t_L g667 ( .A(n_631), .B(n_566), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_614), .Y(n_668) );
AND2x2_ASAP7_75t_L g669 ( .A(n_631), .B(n_592), .Y(n_669) );
OR2x6_ASAP7_75t_L g670 ( .A(n_636), .B(n_551), .Y(n_670) );
OR2x2_ASAP7_75t_L g671 ( .A(n_617), .B(n_545), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_637), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_639), .Y(n_673) );
INVx2_ASAP7_75t_SL g674 ( .A(n_647), .Y(n_674) );
OR2x2_ASAP7_75t_L g675 ( .A(n_645), .B(n_571), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_622), .B(n_575), .Y(n_676) );
OR2x2_ASAP7_75t_L g677 ( .A(n_646), .B(n_608), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_602), .B(n_564), .Y(n_678) );
AND2x4_ASAP7_75t_L g679 ( .A(n_615), .B(n_568), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_602), .Y(n_680) );
AND2x4_ASAP7_75t_L g681 ( .A(n_615), .B(n_568), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_634), .B(n_541), .Y(n_682) );
BUFx2_ASAP7_75t_L g683 ( .A(n_621), .Y(n_683) );
INVx2_ASAP7_75t_L g684 ( .A(n_677), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_651), .Y(n_685) );
INVx1_ASAP7_75t_SL g686 ( .A(n_683), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_680), .B(n_646), .Y(n_687) );
OR2x2_ASAP7_75t_L g688 ( .A(n_658), .B(n_638), .Y(n_688) );
AND2x2_ASAP7_75t_L g689 ( .A(n_665), .B(n_648), .Y(n_689) );
INVx1_ASAP7_75t_SL g690 ( .A(n_674), .Y(n_690) );
OAI322xp33_ASAP7_75t_L g691 ( .A1(n_660), .A2(n_618), .A3(n_640), .B1(n_607), .B2(n_635), .C1(n_613), .C2(n_641), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_655), .Y(n_692) );
INVxp67_ASAP7_75t_L g693 ( .A(n_659), .Y(n_693) );
AND2x2_ASAP7_75t_L g694 ( .A(n_666), .B(n_624), .Y(n_694) );
OR2x2_ASAP7_75t_L g695 ( .A(n_654), .B(n_640), .Y(n_695) );
INVx2_ASAP7_75t_L g696 ( .A(n_656), .Y(n_696) );
HB1xp67_ASAP7_75t_L g697 ( .A(n_654), .Y(n_697) );
AND2x4_ASAP7_75t_L g698 ( .A(n_664), .B(n_620), .Y(n_698) );
INVx2_ASAP7_75t_L g699 ( .A(n_663), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_668), .Y(n_700) );
AND2x2_ASAP7_75t_L g701 ( .A(n_661), .B(n_648), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_673), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_672), .Y(n_703) );
AND2x2_ASAP7_75t_L g704 ( .A(n_701), .B(n_669), .Y(n_704) );
INVxp67_ASAP7_75t_SL g705 ( .A(n_697), .Y(n_705) );
NOR2xp33_ASAP7_75t_L g706 ( .A(n_690), .B(n_686), .Y(n_706) );
OAI22xp5_ASAP7_75t_L g707 ( .A1(n_693), .A2(n_681), .B1(n_679), .B2(n_670), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_697), .Y(n_708) );
OAI211xp5_ASAP7_75t_L g709 ( .A1(n_695), .A2(n_676), .B(n_653), .C(n_662), .Y(n_709) );
OAI221xp5_ASAP7_75t_L g710 ( .A1(n_685), .A2(n_676), .B1(n_678), .B2(n_670), .C(n_671), .Y(n_710) );
INVx1_ASAP7_75t_L g711 ( .A(n_696), .Y(n_711) );
OAI21xp5_ASAP7_75t_L g712 ( .A1(n_696), .A2(n_621), .B(n_620), .Y(n_712) );
INVx1_ASAP7_75t_L g713 ( .A(n_699), .Y(n_713) );
AOI22xp5_ASAP7_75t_L g714 ( .A1(n_698), .A2(n_667), .B1(n_682), .B2(n_620), .Y(n_714) );
NAND2x1p5_ASAP7_75t_L g715 ( .A(n_706), .B(n_568), .Y(n_715) );
AOI22xp33_ASAP7_75t_SL g716 ( .A1(n_709), .A2(n_698), .B1(n_694), .B2(n_689), .Y(n_716) );
AOI22xp5_ASAP7_75t_L g717 ( .A1(n_710), .A2(n_689), .B1(n_703), .B2(n_702), .Y(n_717) );
AOI22xp5_ASAP7_75t_L g718 ( .A1(n_707), .A2(n_700), .B1(n_692), .B2(n_699), .Y(n_718) );
AOI22xp5_ASAP7_75t_L g719 ( .A1(n_714), .A2(n_684), .B1(n_687), .B2(n_688), .Y(n_719) );
OAI31xp33_ASAP7_75t_L g720 ( .A1(n_705), .A2(n_652), .A3(n_657), .B(n_675), .Y(n_720) );
AOI211x1_ASAP7_75t_L g721 ( .A1(n_712), .A2(n_650), .B(n_691), .C(n_544), .Y(n_721) );
INVx2_ASAP7_75t_L g722 ( .A(n_711), .Y(n_722) );
AOI221xp5_ASAP7_75t_L g723 ( .A1(n_708), .A2(n_619), .B1(n_630), .B2(n_604), .C(n_603), .Y(n_723) );
AOI211xp5_ASAP7_75t_L g724 ( .A1(n_704), .A2(n_553), .B(n_559), .C(n_625), .Y(n_724) );
NOR2xp33_ASAP7_75t_L g725 ( .A(n_713), .B(n_536), .Y(n_725) );
OAI211xp5_ASAP7_75t_L g726 ( .A1(n_721), .A2(n_716), .B(n_717), .C(n_718), .Y(n_726) );
NOR2xp33_ASAP7_75t_SL g727 ( .A(n_720), .B(n_715), .Y(n_727) );
INVxp67_ASAP7_75t_L g728 ( .A(n_725), .Y(n_728) );
AOI21xp5_ASAP7_75t_L g729 ( .A1(n_726), .A2(n_724), .B(n_722), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_728), .B(n_719), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_729), .B(n_727), .Y(n_731) );
NOR3xp33_ASAP7_75t_L g732 ( .A(n_730), .B(n_550), .C(n_723), .Y(n_732) );
INVx2_ASAP7_75t_L g733 ( .A(n_731), .Y(n_733) );
OAI22x1_ASAP7_75t_L g734 ( .A1(n_733), .A2(n_732), .B1(n_585), .B2(n_587), .Y(n_734) );
AOI21xp33_ASAP7_75t_SL g735 ( .A1(n_734), .A2(n_585), .B(n_587), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_735), .B(n_642), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_736), .B(n_581), .Y(n_737) );
OR2x6_ASAP7_75t_L g738 ( .A(n_737), .B(n_627), .Y(n_738) );
AOI22xp33_ASAP7_75t_L g739 ( .A1(n_738), .A2(n_628), .B1(n_606), .B2(n_626), .Y(n_739) );
endmodule