module fake_jpeg_23739_n_265 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_265);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_265;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx12_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_39),
.Y(n_51)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_41),
.Y(n_81)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_47),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_17),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_17),
.B(n_0),
.Y(n_45)
);

AOI21xp33_ASAP7_75t_L g82 ( 
.A1(n_45),
.A2(n_48),
.B(n_1),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_22),
.B(n_0),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_17),
.B(n_0),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_50),
.B(n_52),
.Y(n_95)
);

CKINVDCx12_ASAP7_75t_R g52 ( 
.A(n_44),
.Y(n_52)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_54),
.B(n_57),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_40),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_55),
.A2(n_63),
.B1(n_72),
.B2(n_76),
.Y(n_91)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_31),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_60),
.B(n_67),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_61),
.B(n_69),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx3_ASAP7_75t_SL g116 ( 
.A(n_62),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_40),
.A2(n_20),
.B1(n_19),
.B2(n_21),
.Y(n_63)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_64),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_47),
.B(n_31),
.Y(n_65)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_65),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_45),
.B(n_18),
.Y(n_66)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_66),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_48),
.Y(n_67)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_70),
.B(n_71),
.Y(n_109)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_48),
.A2(n_20),
.B1(n_19),
.B2(n_27),
.Y(n_72)
);

CKINVDCx12_ASAP7_75t_R g73 ( 
.A(n_44),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_73),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_38),
.B(n_21),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_74),
.B(n_78),
.Y(n_101)
);

CKINVDCx12_ASAP7_75t_R g75 ( 
.A(n_40),
.Y(n_75)
);

OR2x2_ASAP7_75t_SL g115 ( 
.A(n_75),
.B(n_82),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_40),
.A2(n_27),
.B1(n_19),
.B2(n_26),
.Y(n_76)
);

OA22x2_ASAP7_75t_L g77 ( 
.A1(n_37),
.A2(n_25),
.B1(n_33),
.B2(n_26),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_77),
.A2(n_86),
.B1(n_32),
.B2(n_24),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_38),
.B(n_27),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_79),
.Y(n_93)
);

BUFx8_ASAP7_75t_L g80 ( 
.A(n_39),
.Y(n_80)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_41),
.Y(n_83)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_83),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_41),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_84),
.B(n_85),
.Y(n_90)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_41),
.Y(n_85)
);

OA22x2_ASAP7_75t_L g86 ( 
.A1(n_43),
.A2(n_25),
.B1(n_33),
.B2(n_30),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_39),
.Y(n_87)
);

O2A1O1Ixp33_ASAP7_75t_L g112 ( 
.A1(n_87),
.A2(n_36),
.B(n_30),
.C(n_29),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_96),
.A2(n_99),
.B1(n_114),
.B2(n_110),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_59),
.B(n_42),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_98),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_51),
.A2(n_42),
.B(n_32),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_87),
.B(n_43),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_104),
.B(n_105),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_80),
.B(n_86),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_80),
.B(n_86),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_106),
.B(n_107),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_77),
.B(n_43),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_77),
.B(n_43),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_108),
.B(n_113),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_68),
.A2(n_18),
.B1(n_35),
.B2(n_34),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_110),
.A2(n_76),
.B1(n_63),
.B2(n_24),
.Y(n_118)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_112),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_49),
.B(n_17),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_49),
.B(n_35),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_117),
.B(n_58),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_118),
.A2(n_127),
.B1(n_116),
.B2(n_81),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_117),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_119),
.Y(n_160)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_103),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_120),
.B(n_130),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_101),
.B(n_55),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_122),
.B(n_128),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_88),
.B(n_114),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_123),
.B(n_125),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_97),
.B(n_50),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_124),
.B(n_2),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_94),
.B(n_61),
.Y(n_125)
);

AOI32xp33_ASAP7_75t_L g126 ( 
.A1(n_115),
.A2(n_53),
.A3(n_56),
.B1(n_29),
.B2(n_36),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_SL g165 ( 
.A(n_126),
.B(n_13),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_94),
.B(n_34),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_102),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_129),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_99),
.B(n_92),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_112),
.B(n_1),
.Y(n_131)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_131),
.Y(n_154)
);

OAI22xp33_ASAP7_75t_L g132 ( 
.A1(n_107),
.A2(n_84),
.B1(n_83),
.B2(n_62),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_132),
.A2(n_93),
.B1(n_89),
.B2(n_111),
.Y(n_156)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_95),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_134),
.Y(n_167)
);

OAI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_108),
.A2(n_96),
.B1(n_91),
.B2(n_105),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_135),
.A2(n_90),
.B1(n_81),
.B2(n_68),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_113),
.B(n_16),
.Y(n_136)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_136),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g137 ( 
.A(n_103),
.Y(n_137)
);

INVxp33_ASAP7_75t_L g149 ( 
.A(n_137),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_98),
.B(n_15),
.Y(n_138)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_138),
.Y(n_176)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_89),
.Y(n_139)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_139),
.Y(n_151)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_111),
.Y(n_142)
);

INVx13_ASAP7_75t_L g152 ( 
.A(n_142),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_100),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_143),
.B(n_145),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_106),
.B(n_1),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_144),
.A2(n_2),
.B(n_3),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_109),
.Y(n_145)
);

OAI32xp33_ASAP7_75t_L g147 ( 
.A1(n_91),
.A2(n_115),
.A3(n_92),
.B1(n_104),
.B2(n_90),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_147),
.B(n_148),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_153),
.A2(n_156),
.B1(n_163),
.B2(n_168),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_155),
.B(n_139),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_157),
.A2(n_158),
.B(n_169),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_140),
.A2(n_93),
.B(n_116),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_124),
.B(n_116),
.C(n_15),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_162),
.B(n_165),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_133),
.A2(n_141),
.B1(n_140),
.B2(n_147),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_166),
.B(n_171),
.Y(n_188)
);

AO22x1_ASAP7_75t_SL g168 ( 
.A1(n_132),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_141),
.A2(n_5),
.B(n_7),
.Y(n_169)
);

INVx13_ASAP7_75t_L g170 ( 
.A(n_137),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_170),
.B(n_142),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_121),
.B(n_146),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_133),
.A2(n_146),
.B1(n_119),
.B2(n_148),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_173),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_160),
.B(n_144),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_177),
.B(n_178),
.Y(n_205)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_150),
.Y(n_178)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_150),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_180),
.B(n_186),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_172),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_181),
.B(n_182),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_161),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_184),
.B(n_185),
.Y(n_210)
);

BUFx24_ASAP7_75t_SL g185 ( 
.A(n_159),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_169),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_174),
.A2(n_121),
.B1(n_144),
.B2(n_118),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_187),
.A2(n_168),
.B1(n_154),
.B2(n_167),
.Y(n_208)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_156),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_189),
.B(n_191),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_190),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_157),
.B(n_158),
.Y(n_191)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_155),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_193),
.B(n_194),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_164),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_149),
.B(n_151),
.Y(n_195)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_195),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_174),
.A2(n_129),
.B(n_145),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_197),
.B(n_167),
.Y(n_212)
);

OAI322xp33_ASAP7_75t_L g198 ( 
.A1(n_188),
.A2(n_171),
.A3(n_166),
.B1(n_165),
.B2(n_162),
.C1(n_168),
.C2(n_176),
.Y(n_198)
);

AOI31xp33_ASAP7_75t_L g227 ( 
.A1(n_198),
.A2(n_179),
.A3(n_177),
.B(n_191),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_188),
.B(n_143),
.C(n_176),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_201),
.B(n_204),
.C(n_214),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_197),
.B(n_175),
.C(n_151),
.Y(n_204)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_181),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_207),
.B(n_182),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_208),
.B(n_212),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_189),
.Y(n_209)
);

INVxp67_ASAP7_75t_SL g217 ( 
.A(n_209),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_186),
.B(n_170),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_213),
.A2(n_206),
.B(n_199),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_187),
.B(n_175),
.C(n_149),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_199),
.A2(n_193),
.B1(n_180),
.B2(n_178),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_216),
.A2(n_223),
.B1(n_8),
.B2(n_10),
.Y(n_238)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_218),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_214),
.B(n_183),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_219),
.B(n_224),
.C(n_200),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_203),
.B(n_194),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_220),
.B(n_221),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_202),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_L g223 ( 
.A1(n_213),
.A2(n_183),
.B1(n_152),
.B2(n_154),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_209),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_225),
.Y(n_239)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_202),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_226),
.B(n_213),
.Y(n_233)
);

OAI322xp33_ASAP7_75t_L g229 ( 
.A1(n_227),
.A2(n_205),
.A3(n_211),
.B1(n_212),
.B2(n_201),
.C1(n_179),
.C2(n_204),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_210),
.B(n_196),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_228),
.B(n_120),
.Y(n_236)
);

MAJx2_ASAP7_75t_L g247 ( 
.A(n_229),
.B(n_234),
.C(n_240),
.Y(n_247)
);

FAx1_ASAP7_75t_SL g230 ( 
.A(n_215),
.B(n_208),
.CI(n_196),
.CON(n_230),
.SN(n_230)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_230),
.B(n_236),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_232),
.B(n_8),
.C(n_11),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_233),
.A2(n_237),
.B(n_224),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_219),
.B(n_192),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_226),
.B(n_152),
.Y(n_237)
);

AOI21x1_ASAP7_75t_SL g241 ( 
.A1(n_238),
.A2(n_217),
.B(n_11),
.Y(n_241)
);

XOR2x2_ASAP7_75t_SL g240 ( 
.A(n_215),
.B(n_8),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_241),
.A2(n_243),
.B1(n_233),
.B2(n_240),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_242),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_231),
.A2(n_216),
.B1(n_222),
.B2(n_14),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_235),
.B(n_222),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_244),
.B(n_245),
.Y(n_249)
);

INVx11_ASAP7_75t_L g245 ( 
.A(n_239),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_248),
.A2(n_237),
.B(n_232),
.Y(n_250)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_250),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_246),
.B(n_234),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_251),
.B(n_254),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_252),
.B(n_230),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_242),
.A2(n_230),
.B(n_12),
.Y(n_254)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_255),
.Y(n_259)
);

OAI21xp33_ASAP7_75t_L g256 ( 
.A1(n_253),
.A2(n_247),
.B(n_241),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_256),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_257),
.B(n_258),
.C(n_249),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_260),
.B(n_249),
.C(n_248),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_262),
.B(n_263),
.C(n_259),
.Y(n_264)
);

NOR4xp25_ASAP7_75t_L g263 ( 
.A(n_261),
.B(n_256),
.C(n_247),
.D(n_245),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_264),
.B(n_12),
.Y(n_265)
);


endmodule