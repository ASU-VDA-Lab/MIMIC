module fake_jpeg_26370_n_229 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_229);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_229;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_2),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_19),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_24),
.B(n_26),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

NAND2xp33_ASAP7_75t_SL g40 ( 
.A(n_27),
.B(n_21),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g28 ( 
.A1(n_13),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_28),
.A2(n_23),
.B1(n_20),
.B2(n_17),
.Y(n_39)
);

INVx1_ASAP7_75t_SL g29 ( 
.A(n_19),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_29),
.B(n_31),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_13),
.B(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_32),
.B(n_14),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_L g33 ( 
.A1(n_24),
.A2(n_15),
.B1(n_16),
.B2(n_19),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_33),
.A2(n_29),
.B1(n_12),
.B2(n_23),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_32),
.B(n_21),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_35),
.B(n_38),
.Y(n_51)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_39),
.A2(n_20),
.B1(n_23),
.B2(n_17),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_27),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_43),
.Y(n_44)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_32),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_46),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_41),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_27),
.C(n_30),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_47),
.A2(n_48),
.B1(n_53),
.B2(n_59),
.Y(n_77)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_41),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_50),
.B(n_55),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_38),
.A2(n_29),
.B1(n_24),
.B2(n_18),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

AO22x2_ASAP7_75t_L g53 ( 
.A1(n_39),
.A2(n_27),
.B1(n_30),
.B2(n_26),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

CKINVDCx9p33_ASAP7_75t_R g56 ( 
.A(n_33),
.Y(n_56)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_60),
.Y(n_76)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_53),
.A2(n_43),
.B1(n_37),
.B2(n_39),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_62),
.A2(n_53),
.B1(n_57),
.B2(n_58),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_44),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_68),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_36),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_51),
.Y(n_80)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_69),
.B(n_72),
.Y(n_94)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_53),
.A2(n_56),
.B1(n_46),
.B2(n_50),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_75),
.A2(n_53),
.B1(n_43),
.B2(n_37),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_77),
.B(n_47),
.C(n_55),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_79),
.B(n_84),
.C(n_85),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_80),
.B(n_86),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_81),
.A2(n_89),
.B1(n_74),
.B2(n_78),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_77),
.B(n_47),
.C(n_57),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_77),
.B(n_57),
.C(n_60),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_67),
.B(n_45),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_65),
.B(n_48),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_88),
.B(n_91),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_76),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_90),
.Y(n_98)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_62),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_63),
.B(n_48),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_92),
.B(n_93),
.Y(n_107)
);

AO22x1_ASAP7_75t_SL g93 ( 
.A1(n_74),
.A2(n_59),
.B1(n_52),
.B2(n_37),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_61),
.A2(n_36),
.B(n_52),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_95),
.A2(n_92),
.B(n_88),
.Y(n_99)
);

OAI32xp33_ASAP7_75t_L g96 ( 
.A1(n_91),
.A2(n_63),
.A3(n_73),
.B1(n_68),
.B2(n_75),
.Y(n_96)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_96),
.Y(n_118)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_94),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_97),
.B(n_104),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_99),
.A2(n_100),
.B(n_83),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_81),
.A2(n_95),
.B(n_62),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_103),
.A2(n_87),
.B1(n_78),
.B2(n_93),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_76),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_94),
.Y(n_105)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_105),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_82),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_106),
.Y(n_121)
);

AOI22x1_ASAP7_75t_SL g108 ( 
.A1(n_85),
.A2(n_70),
.B1(n_78),
.B2(n_73),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_108),
.A2(n_110),
.B1(n_87),
.B2(n_93),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_82),
.B(n_64),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_109),
.Y(n_122)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_89),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_86),
.B(n_64),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_112),
.B(n_83),
.Y(n_113)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_113),
.Y(n_134)
);

BUFx12_ASAP7_75t_L g114 ( 
.A(n_108),
.Y(n_114)
);

INVx11_ASAP7_75t_L g149 ( 
.A(n_114),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_102),
.B(n_79),
.C(n_84),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_115),
.B(n_111),
.C(n_101),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_116),
.A2(n_117),
.B1(n_71),
.B2(n_26),
.Y(n_146)
);

OAI21xp33_ASAP7_75t_L g119 ( 
.A1(n_108),
.A2(n_98),
.B(n_106),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_119),
.A2(n_121),
.B1(n_131),
.B2(n_118),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g120 ( 
.A(n_102),
.B(n_79),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_SL g133 ( 
.A(n_120),
.B(n_128),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_110),
.A2(n_85),
.B1(n_93),
.B2(n_80),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_123),
.A2(n_127),
.B1(n_129),
.B2(n_71),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_38),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_124),
.B(n_26),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_107),
.A2(n_72),
.B(n_66),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_126),
.A2(n_130),
.B(n_98),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_107),
.A2(n_28),
.B1(n_66),
.B2(n_69),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_101),
.A2(n_69),
.B1(n_71),
.B2(n_18),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_99),
.A2(n_0),
.B(n_1),
.Y(n_130)
);

OAI22x1_ASAP7_75t_L g132 ( 
.A1(n_114),
.A2(n_103),
.B1(n_96),
.B2(n_100),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_132),
.A2(n_141),
.B1(n_148),
.B2(n_18),
.Y(n_166)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_113),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_135),
.B(n_142),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_136),
.B(n_139),
.C(n_144),
.Y(n_153)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_137),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_120),
.B(n_111),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_138),
.B(n_140),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_112),
.C(n_105),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_124),
.B(n_97),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_128),
.B(n_104),
.Y(n_142)
);

MAJx2_ASAP7_75t_L g143 ( 
.A(n_114),
.B(n_109),
.C(n_27),
.Y(n_143)
);

A2O1A1O1Ixp25_ASAP7_75t_L g165 ( 
.A1(n_143),
.A2(n_145),
.B(n_22),
.C(n_25),
.D(n_19),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_123),
.B(n_27),
.C(n_30),
.Y(n_144)
);

XNOR2x2_ASAP7_75t_SL g145 ( 
.A(n_126),
.B(n_22),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_146),
.A2(n_113),
.B1(n_117),
.B2(n_116),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_121),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_147),
.B(n_150),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_125),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_151),
.B(n_25),
.C(n_15),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_136),
.B(n_118),
.Y(n_154)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_154),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_141),
.B(n_131),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_155),
.B(n_156),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_139),
.B(n_122),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_157),
.B(n_159),
.Y(n_176)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_144),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_158),
.B(n_168),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_132),
.Y(n_159)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_149),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_161),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_149),
.A2(n_114),
.B1(n_130),
.B2(n_12),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_164),
.A2(n_166),
.B1(n_20),
.B2(n_17),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_165),
.B(n_143),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_167),
.B(n_133),
.Y(n_170)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_151),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_162),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_169),
.B(n_173),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_170),
.B(n_181),
.Y(n_185)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_171),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_160),
.B(n_138),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_160),
.B(n_133),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_177),
.B(n_178),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_153),
.B(n_140),
.C(n_134),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_163),
.B(n_14),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_180),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_153),
.B(n_145),
.C(n_42),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_182),
.A2(n_152),
.B1(n_167),
.B2(n_165),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_155),
.B(n_14),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_183),
.B(n_174),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_176),
.A2(n_152),
.B(n_157),
.Y(n_184)
);

O2A1O1Ixp33_ASAP7_75t_SL g202 ( 
.A1(n_184),
.A2(n_193),
.B(n_16),
.C(n_15),
.Y(n_202)
);

OA21x2_ASAP7_75t_SL g186 ( 
.A1(n_169),
.A2(n_178),
.B(n_179),
.Y(n_186)
);

OR2x2_ASAP7_75t_L g198 ( 
.A(n_186),
.B(n_42),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_189),
.B(n_194),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_170),
.B(n_164),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_192),
.B(n_195),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_175),
.A2(n_161),
.B(n_159),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_172),
.B(n_12),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_187),
.A2(n_174),
.B1(n_181),
.B2(n_11),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_196),
.B(n_198),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_195),
.B(n_16),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_199),
.B(n_202),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_191),
.B(n_22),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_200),
.B(n_201),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_188),
.A2(n_0),
.B(n_1),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_184),
.B(n_193),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_203),
.B(n_15),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_190),
.A2(n_22),
.B(n_16),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_205),
.B(n_194),
.C(n_185),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_197),
.B(n_185),
.C(n_192),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_206),
.B(n_42),
.C(n_4),
.Y(n_217)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_207),
.Y(n_216)
);

OAI21x1_ASAP7_75t_L g208 ( 
.A1(n_204),
.A2(n_201),
.B(n_22),
.Y(n_208)
);

AOI322xp5_ASAP7_75t_L g214 ( 
.A1(n_208),
.A2(n_211),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_7),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_209),
.B(n_42),
.Y(n_219)
);

OAI21x1_ASAP7_75t_L g211 ( 
.A1(n_198),
.A2(n_2),
.B(n_3),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_214),
.A2(n_215),
.B1(n_220),
.B2(n_9),
.Y(n_224)
);

AOI322xp5_ASAP7_75t_L g215 ( 
.A1(n_210),
.A2(n_3),
.A3(n_4),
.B1(n_6),
.B2(n_7),
.C1(n_8),
.C2(n_9),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_217),
.B(n_218),
.C(n_212),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_213),
.B(n_3),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_219),
.Y(n_222)
);

AOI322xp5_ASAP7_75t_L g220 ( 
.A1(n_206),
.A2(n_6),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.C1(n_10),
.C2(n_42),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_221),
.Y(n_227)
);

NAND3xp33_ASAP7_75t_L g223 ( 
.A(n_216),
.B(n_6),
.C(n_7),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_223),
.A2(n_224),
.B(n_225),
.Y(n_226)
);

OA21x2_ASAP7_75t_SL g225 ( 
.A1(n_217),
.A2(n_9),
.B(n_10),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_227),
.B(n_222),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_228),
.B(n_226),
.Y(n_229)
);


endmodule