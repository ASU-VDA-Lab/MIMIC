module real_jpeg_20850_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_83;
wire n_78;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_44;
wire n_28;
wire n_62;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

AOI22xp33_ASAP7_75t_SL g28 ( 
.A1(n_0),
.A2(n_20),
.B1(n_21),
.B2(n_29),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_0),
.A2(n_24),
.B1(n_25),
.B2(n_29),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_1),
.A2(n_24),
.B1(n_25),
.B2(n_43),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_1),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_2),
.A2(n_24),
.B1(n_25),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_2),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_2),
.A2(n_20),
.B1(n_21),
.B2(n_39),
.Y(n_64)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_3),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_4),
.A2(n_24),
.B1(n_25),
.B2(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_4),
.Y(n_48)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_7),
.A2(n_20),
.B1(n_21),
.B2(n_27),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_7),
.A2(n_27),
.B1(n_50),
.B2(n_51),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_7),
.A2(n_24),
.B1(n_25),
.B2(n_27),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_8),
.A2(n_20),
.B1(n_21),
.B2(n_34),
.Y(n_33)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

OAI32xp33_ASAP7_75t_L g49 ( 
.A1(n_8),
.A2(n_21),
.A3(n_50),
.B1(n_52),
.B2(n_53),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_9),
.B(n_32),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_9),
.Y(n_54)
);

AOI21xp33_ASAP7_75t_L g59 ( 
.A1(n_9),
.A2(n_50),
.B(n_60),
.Y(n_59)
);

AOI21xp33_ASAP7_75t_L g80 ( 
.A1(n_9),
.A2(n_10),
.B(n_24),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_9),
.A2(n_20),
.B1(n_21),
.B2(n_54),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_9),
.A2(n_36),
.B1(n_37),
.B2(n_88),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_L g19 ( 
.A1(n_10),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_19)
);

INVx6_ASAP7_75t_SL g22 ( 
.A(n_10),
.Y(n_22)
);

OA22x2_ASAP7_75t_L g23 ( 
.A1(n_10),
.A2(n_22),
.B1(n_24),
.B2(n_25),
.Y(n_23)
);

BUFx3_ASAP7_75t_SL g21 ( 
.A(n_11),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_69),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_68),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_44),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_16),
.B(n_44),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_30),
.C(n_35),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_17),
.A2(n_30),
.B1(n_31),
.B2(n_100),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_17),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_23),
.B1(n_26),
.B2(n_28),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_18),
.A2(n_23),
.B1(n_28),
.B2(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_18),
.A2(n_23),
.B1(n_26),
.B2(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_23),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_20),
.B(n_34),
.Y(n_52)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

A2O1A1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_21),
.A2(n_22),
.B(n_54),
.C(n_80),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_23),
.B(n_54),
.Y(n_86)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_24),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_25),
.B(n_91),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_33),
.A2(n_57),
.B1(n_59),
.B2(n_61),
.Y(n_56)
);

A2O1A1Ixp33_ASAP7_75t_L g57 ( 
.A1(n_33),
.A2(n_34),
.B(n_51),
.C(n_58),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_34),
.B(n_51),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_35),
.B(n_99),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_38),
.B1(n_40),
.B2(n_42),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_36),
.A2(n_37),
.B1(n_42),
.B2(n_47),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_36),
.A2(n_37),
.B1(n_75),
.B2(n_88),
.Y(n_87)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_38),
.Y(n_76)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_41),
.A2(n_73),
.B1(n_74),
.B2(n_76),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_55),
.B1(n_66),
.B2(n_67),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_45),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_49),
.Y(n_45)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_51),
.B(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_53),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_54),
.B(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_62),
.B1(n_63),
.B2(n_65),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_56),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_SL g69 ( 
.A1(n_70),
.A2(n_96),
.B(n_101),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_84),
.B(n_95),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_77),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_72),
.B(n_77),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_79),
.B1(n_81),
.B2(n_82),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_79),
.B(n_81),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_85),
.A2(n_89),
.B(n_94),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_87),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_86),
.B(n_87),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_93),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_98),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_97),
.B(n_98),
.Y(n_101)
);


endmodule