module fake_jpeg_16329_n_334 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_334);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_334;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_SL g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_6),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx4f_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

BUFx10_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

BUFx24_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

INVx3_ASAP7_75t_SL g98 ( 
.A(n_43),
.Y(n_98)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_45),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_17),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_46),
.B(n_58),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_16),
.B(n_6),
.Y(n_47)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_47),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_16),
.B(n_8),
.Y(n_48)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_49),
.Y(n_90)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_50),
.Y(n_96)
);

BUFx4f_ASAP7_75t_SL g51 ( 
.A(n_40),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g81 ( 
.A(n_51),
.Y(n_81)
);

INVx6_ASAP7_75t_SL g52 ( 
.A(n_23),
.Y(n_52)
);

INVx6_ASAP7_75t_SL g111 ( 
.A(n_52),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_53),
.Y(n_126)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_54),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_55),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_56),
.Y(n_115)
);

INVx3_ASAP7_75t_SL g57 ( 
.A(n_37),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_57),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_17),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_59),
.B(n_61),
.Y(n_93)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_60),
.B(n_64),
.Y(n_85)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_22),
.B(n_0),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_63),
.B(n_76),
.Y(n_118)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_65),
.B(n_66),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_21),
.B(n_8),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_21),
.B(n_5),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_67),
.B(n_68),
.Y(n_107)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_69),
.B(n_70),
.Y(n_121)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

CKINVDCx12_ASAP7_75t_R g71 ( 
.A(n_23),
.Y(n_71)
);

CKINVDCx12_ASAP7_75t_R g88 ( 
.A(n_71),
.Y(n_88)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_25),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_73),
.B(n_75),
.Y(n_109)
);

CKINVDCx9p33_ASAP7_75t_R g74 ( 
.A(n_41),
.Y(n_74)
);

CKINVDCx9p33_ASAP7_75t_R g97 ( 
.A(n_74),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_24),
.B(n_5),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_22),
.B(n_26),
.Y(n_76)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_77),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_24),
.B(n_5),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_78),
.B(n_70),
.Y(n_123)
);

INVx2_ASAP7_75t_SL g79 ( 
.A(n_23),
.Y(n_79)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_79),
.Y(n_101)
);

INVx2_ASAP7_75t_SL g80 ( 
.A(n_29),
.Y(n_80)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_80),
.Y(n_104)
);

OA22x2_ASAP7_75t_L g91 ( 
.A1(n_57),
.A2(n_74),
.B1(n_72),
.B2(n_80),
.Y(n_91)
);

OAI32xp33_ASAP7_75t_L g136 ( 
.A1(n_91),
.A2(n_117),
.A3(n_51),
.B1(n_50),
.B2(n_56),
.Y(n_136)
);

OR2x4_ASAP7_75t_L g94 ( 
.A(n_76),
.B(n_41),
.Y(n_94)
);

OR2x4_ASAP7_75t_L g162 ( 
.A(n_94),
.B(n_117),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_43),
.A2(n_30),
.B1(n_42),
.B2(n_27),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_99),
.A2(n_100),
.B1(n_102),
.B2(n_112),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_54),
.A2(n_30),
.B1(n_57),
.B2(n_61),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_65),
.A2(n_25),
.B1(n_36),
.B2(n_27),
.Y(n_102)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_79),
.Y(n_105)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_105),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_46),
.A2(n_28),
.B1(n_31),
.B2(n_35),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_106),
.A2(n_108),
.B1(n_114),
.B2(n_113),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_68),
.A2(n_28),
.B1(n_31),
.B2(n_35),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_58),
.B(n_36),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_110),
.B(n_116),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_44),
.A2(n_77),
.B1(n_26),
.B2(n_32),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_73),
.A2(n_34),
.B1(n_32),
.B2(n_38),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_60),
.B(n_34),
.Y(n_116)
);

OA22x2_ASAP7_75t_L g117 ( 
.A1(n_79),
.A2(n_41),
.B1(n_33),
.B2(n_29),
.Y(n_117)
);

CKINVDCx9p33_ASAP7_75t_R g119 ( 
.A(n_51),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_119),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_64),
.B(n_38),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_120),
.B(n_15),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_63),
.B(n_0),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_122),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_123),
.B(n_127),
.Y(n_167)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_80),
.Y(n_124)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_124),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_69),
.B(n_29),
.Y(n_127)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_45),
.Y(n_129)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_129),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_52),
.A2(n_41),
.B1(n_38),
.B2(n_12),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_130),
.A2(n_133),
.B1(n_98),
.B2(n_84),
.Y(n_172)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_62),
.Y(n_131)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_131),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_53),
.A2(n_33),
.B1(n_29),
.B2(n_11),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_132),
.A2(n_113),
.B1(n_98),
.B2(n_129),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_55),
.A2(n_11),
.B1(n_15),
.B2(n_13),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_94),
.B(n_59),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_135),
.B(n_143),
.Y(n_184)
);

AO22x1_ASAP7_75t_L g208 ( 
.A1(n_136),
.A2(n_148),
.B1(n_142),
.B2(n_138),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_118),
.B(n_1),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_137),
.B(n_138),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_1),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_97),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_139),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_85),
.B(n_49),
.C(n_33),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_141),
.B(n_142),
.C(n_178),
.Y(n_212)
);

AND2x2_ASAP7_75t_SL g142 ( 
.A(n_121),
.B(n_33),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_118),
.B(n_1),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_117),
.B(n_2),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_146),
.Y(n_187)
);

CKINVDCx14_ASAP7_75t_R g193 ( 
.A(n_147),
.Y(n_193)
);

OR2x2_ASAP7_75t_L g148 ( 
.A(n_97),
.B(n_3),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_148),
.B(n_153),
.Y(n_191)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_151),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_82),
.B(n_15),
.Y(n_152)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_152),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_122),
.B(n_10),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_109),
.B(n_12),
.Y(n_154)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_154),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_107),
.B(n_103),
.Y(n_155)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_155),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_87),
.B(n_89),
.Y(n_156)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_156),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_122),
.B(n_93),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_158),
.B(n_163),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_92),
.B(n_105),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_159),
.B(n_161),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_81),
.B(n_111),
.Y(n_160)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_160),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_81),
.B(n_111),
.Y(n_161)
);

FAx1_ASAP7_75t_SL g202 ( 
.A(n_162),
.B(n_179),
.CI(n_163),
.CON(n_202),
.SN(n_202)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_92),
.B(n_104),
.Y(n_163)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_164),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_165),
.A2(n_144),
.B1(n_171),
.B2(n_179),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_95),
.A2(n_128),
.B1(n_126),
.B2(n_131),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_166),
.A2(n_174),
.B1(n_86),
.B2(n_146),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_83),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_168),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_101),
.B(n_104),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_169),
.B(n_170),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_101),
.B(n_124),
.Y(n_170)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_83),
.Y(n_171)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_171),
.Y(n_181)
);

OAI22x1_ASAP7_75t_L g198 ( 
.A1(n_172),
.A2(n_174),
.B1(n_146),
.B2(n_147),
.Y(n_198)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_90),
.Y(n_173)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_173),
.Y(n_190)
);

OA22x2_ASAP7_75t_L g174 ( 
.A1(n_117),
.A2(n_91),
.B1(n_119),
.B2(n_84),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_115),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_175),
.B(n_176),
.Y(n_186)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_125),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_125),
.Y(n_177)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_177),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_91),
.B(n_88),
.C(n_96),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_95),
.B(n_126),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_96),
.B(n_91),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_180),
.B(n_139),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_162),
.A2(n_86),
.B1(n_128),
.B2(n_157),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_185),
.A2(n_189),
.B1(n_194),
.B2(n_204),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_L g219 ( 
.A1(n_188),
.A2(n_199),
.B1(n_205),
.B2(n_208),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_178),
.A2(n_136),
.B1(n_143),
.B2(n_135),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_135),
.A2(n_158),
.B1(n_174),
.B2(n_141),
.Y(n_194)
);

BUFx2_ASAP7_75t_L g197 ( 
.A(n_177),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_197),
.B(n_195),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_198),
.A2(n_176),
.B1(n_149),
.B2(n_173),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_202),
.B(n_148),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_174),
.A2(n_153),
.B1(n_144),
.B2(n_150),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_137),
.A2(n_138),
.B1(n_142),
.B2(n_166),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_211),
.A2(n_149),
.B(n_168),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_150),
.A2(n_137),
.B1(n_134),
.B2(n_140),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_L g241 ( 
.A1(n_215),
.A2(n_216),
.B1(n_193),
.B2(n_209),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_167),
.A2(n_145),
.B1(n_175),
.B2(n_140),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_217),
.B(n_227),
.C(n_232),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_202),
.B(n_167),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_218),
.B(n_221),
.Y(n_247)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_181),
.Y(n_220)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_220),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_202),
.B(n_134),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_222),
.A2(n_233),
.B(n_223),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_223),
.A2(n_225),
.B(n_230),
.Y(n_257)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_181),
.Y(n_224)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_224),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_187),
.A2(n_198),
.B(n_188),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_212),
.B(n_168),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_201),
.B(n_139),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_228),
.B(n_236),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_191),
.B(n_201),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_229),
.B(n_234),
.Y(n_246)
);

AND2x4_ASAP7_75t_L g230 ( 
.A(n_208),
.B(n_185),
.Y(n_230)
);

AO22x1_ASAP7_75t_L g231 ( 
.A1(n_204),
.A2(n_208),
.B1(n_215),
.B2(n_209),
.Y(n_231)
);

OA21x2_ASAP7_75t_L g249 ( 
.A1(n_231),
.A2(n_206),
.B(n_221),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_212),
.B(n_194),
.C(n_189),
.Y(n_232)
);

AND2x4_ASAP7_75t_L g233 ( 
.A(n_205),
.B(n_184),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_207),
.B(n_182),
.Y(n_234)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_235),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_184),
.B(n_191),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_186),
.B(n_203),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_237),
.B(n_239),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_214),
.B(n_200),
.Y(n_238)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_238),
.Y(n_264)
);

INVxp33_ASAP7_75t_L g239 ( 
.A(n_197),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_210),
.B(n_183),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_240),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_241),
.A2(n_222),
.B1(n_225),
.B2(n_243),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_214),
.B(n_190),
.Y(n_242)
);

NOR4xp25_ASAP7_75t_L g254 ( 
.A(n_242),
.B(n_243),
.C(n_228),
.D(n_230),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_214),
.B(n_190),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_192),
.A2(n_196),
.B(n_195),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_244),
.A2(n_217),
.B(n_220),
.Y(n_262)
);

NOR3xp33_ASAP7_75t_L g245 ( 
.A(n_233),
.B(n_213),
.C(n_206),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_245),
.B(n_249),
.Y(n_270)
);

NOR2x1_ASAP7_75t_L g248 ( 
.A(n_233),
.B(n_213),
.Y(n_248)
);

NOR2x1_ASAP7_75t_L g268 ( 
.A(n_248),
.B(n_244),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_230),
.A2(n_233),
.B1(n_219),
.B2(n_231),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_250),
.A2(n_260),
.B1(n_265),
.B2(n_249),
.Y(n_282)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_254),
.Y(n_271)
);

AOI221xp5_ASAP7_75t_L g274 ( 
.A1(n_255),
.A2(n_261),
.B1(n_262),
.B2(n_245),
.C(n_248),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_230),
.A2(n_232),
.B(n_242),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_SL g286 ( 
.A(n_256),
.B(n_267),
.Y(n_286)
);

OA21x2_ASAP7_75t_L g258 ( 
.A1(n_230),
.A2(n_231),
.B(n_218),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_258),
.B(n_249),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_226),
.A2(n_238),
.B1(n_227),
.B2(n_229),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_236),
.A2(n_226),
.B(n_224),
.Y(n_265)
);

XNOR2x1_ASAP7_75t_SL g287 ( 
.A(n_268),
.B(n_275),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_253),
.B(n_247),
.Y(n_269)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_269),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_267),
.B(n_256),
.C(n_260),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_272),
.B(n_276),
.C(n_286),
.Y(n_289)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_251),
.Y(n_273)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_273),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_274),
.A2(n_277),
.B(n_279),
.Y(n_296)
);

OAI322xp33_ASAP7_75t_L g275 ( 
.A1(n_247),
.A2(n_253),
.A3(n_248),
.B1(n_254),
.B2(n_264),
.C1(n_258),
.C2(n_256),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_267),
.B(n_265),
.C(n_262),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_246),
.B(n_264),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_251),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_278),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_246),
.B(n_255),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_280),
.B(n_281),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_261),
.B(n_263),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_282),
.B(n_285),
.Y(n_288)
);

INVx13_ASAP7_75t_L g283 ( 
.A(n_252),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_283),
.B(n_284),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_250),
.A2(n_249),
.B1(n_258),
.B2(n_257),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_263),
.B(n_257),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_277),
.B(n_259),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_290),
.B(n_280),
.Y(n_301)
);

A2O1A1O1Ixp25_ASAP7_75t_L g292 ( 
.A1(n_275),
.A2(n_258),
.B(n_266),
.C(n_259),
.D(n_252),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_292),
.A2(n_291),
.B(n_296),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_286),
.B(n_266),
.C(n_272),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_294),
.B(n_295),
.C(n_300),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_276),
.B(n_281),
.C(n_271),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_271),
.B(n_285),
.C(n_269),
.Y(n_300)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_301),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_293),
.B(n_283),
.Y(n_302)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_302),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_287),
.A2(n_268),
.B1(n_284),
.B2(n_282),
.Y(n_304)
);

AOI21x1_ASAP7_75t_SL g317 ( 
.A1(n_304),
.A2(n_288),
.B(n_295),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_299),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_305),
.B(n_306),
.Y(n_315)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_298),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_287),
.A2(n_279),
.B1(n_270),
.B2(n_268),
.Y(n_307)
);

OR2x2_ASAP7_75t_L g318 ( 
.A(n_307),
.B(n_310),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_308),
.B(n_309),
.C(n_311),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_297),
.B(n_283),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_292),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_300),
.B(n_273),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_289),
.B(n_278),
.C(n_294),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_312),
.B(n_303),
.C(n_308),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_317),
.A2(n_319),
.B(n_318),
.Y(n_325)
);

OAI21xp33_ASAP7_75t_L g319 ( 
.A1(n_304),
.A2(n_289),
.B(n_307),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_320),
.B(n_303),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_313),
.B(n_312),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_321),
.B(n_322),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_314),
.B(n_305),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_323),
.B(n_316),
.C(n_317),
.Y(n_326)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_315),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_324),
.B(n_318),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_325),
.B(n_319),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_326),
.B(n_327),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_328),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_330),
.A2(n_327),
.B(n_323),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_331),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_330),
.Y(n_334)
);


endmodule