module fake_jpeg_19182_n_266 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_266);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_266;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

BUFx5_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_SL g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_4),
.B(n_14),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx4f_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_12),
.B(n_0),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_0),
.B(n_3),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_42),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx4_ASAP7_75t_SL g42 ( 
.A(n_25),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_7),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_45),
.Y(n_52)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_47),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_7),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_45),
.A2(n_38),
.B1(n_46),
.B2(n_19),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_49),
.A2(n_55),
.B1(n_64),
.B2(n_42),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_50),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_30),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_53),
.B(n_37),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_45),
.A2(n_19),
.B1(n_20),
.B2(n_34),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_34),
.Y(n_57)
);

FAx1_ASAP7_75t_SL g90 ( 
.A(n_57),
.B(n_33),
.CI(n_16),
.CON(n_90),
.SN(n_90)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_47),
.B(n_28),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_59),
.B(n_21),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_42),
.A2(n_19),
.B1(n_20),
.B2(n_24),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_48),
.A2(n_20),
.B1(n_24),
.B2(n_21),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_65),
.A2(n_62),
.B1(n_33),
.B2(n_16),
.Y(n_102)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_69),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_58),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_70),
.B(n_71),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_52),
.B(n_28),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

INVxp33_ASAP7_75t_L g121 ( 
.A(n_72),
.Y(n_121)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_73),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_58),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_74),
.B(n_75),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_67),
.A2(n_48),
.B1(n_42),
.B2(n_44),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_76),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_77),
.B(n_90),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_52),
.A2(n_44),
.B1(n_41),
.B2(n_36),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_78),
.A2(n_82),
.B1(n_87),
.B2(n_88),
.Y(n_123)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_79),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_57),
.A2(n_51),
.B(n_55),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_80),
.A2(n_104),
.B(n_1),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_81),
.B(n_91),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_49),
.A2(n_41),
.B1(n_36),
.B2(n_39),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_37),
.C(n_30),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_83),
.B(n_93),
.C(n_109),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_63),
.B(n_17),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_84),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_58),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_85),
.B(n_89),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_57),
.A2(n_53),
.B1(n_61),
.B2(n_66),
.Y(n_87)
);

OA22x2_ASAP7_75t_L g88 ( 
.A1(n_61),
.A2(n_39),
.B1(n_35),
.B2(n_22),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_59),
.B(n_31),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_69),
.B(n_18),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_67),
.B(n_31),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_92),
.B(n_94),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_54),
.B(n_23),
.C(n_26),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_56),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_50),
.B(n_29),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_95),
.B(n_96),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_50),
.B(n_29),
.Y(n_96)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_68),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_0),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_60),
.B(n_27),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_98),
.B(n_6),
.Y(n_127)
);

OAI32xp33_ASAP7_75t_L g99 ( 
.A1(n_60),
.A2(n_27),
.A3(n_22),
.B1(n_33),
.B2(n_16),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_99),
.B(n_100),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_62),
.B(n_18),
.Y(n_100)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_68),
.Y(n_101)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_101),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_102),
.A2(n_4),
.B1(n_8),
.B2(n_9),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_56),
.A2(n_26),
.B1(n_23),
.B2(n_35),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_103),
.A2(n_82),
.B1(n_77),
.B2(n_72),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_57),
.A2(n_33),
.B(n_15),
.Y(n_104)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_60),
.Y(n_105)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_105),
.Y(n_115)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_61),
.Y(n_107)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_107),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_63),
.A2(n_26),
.B1(n_23),
.B2(n_33),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_108),
.A2(n_110),
.B1(n_14),
.B2(n_5),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_63),
.B(n_15),
.C(n_8),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_63),
.A2(n_6),
.B1(n_13),
.B2(n_11),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_117),
.B(n_127),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_119),
.B(n_88),
.Y(n_150)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_107),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_124),
.B(n_129),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_100),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_130),
.A2(n_114),
.B1(n_119),
.B2(n_128),
.Y(n_146)
);

AO21x1_ASAP7_75t_SL g153 ( 
.A1(n_132),
.A2(n_123),
.B(n_128),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_84),
.B(n_1),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_133),
.B(n_119),
.Y(n_149)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_86),
.Y(n_136)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_136),
.Y(n_152)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_86),
.Y(n_138)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_138),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_139),
.B(n_93),
.Y(n_162)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_91),
.Y(n_141)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_141),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_105),
.A2(n_99),
.B1(n_97),
.B2(n_101),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g160 ( 
.A(n_142),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_137),
.B(n_81),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_143),
.B(n_158),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_136),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_144),
.B(n_149),
.Y(n_171)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_140),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_145),
.B(n_168),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_146),
.A2(n_153),
.B1(n_112),
.B2(n_132),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_150),
.B(n_167),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_137),
.B(n_83),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_151),
.A2(n_166),
.B(n_150),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_122),
.B(n_109),
.Y(n_156)
);

CKINVDCx14_ASAP7_75t_R g188 ( 
.A(n_156),
.Y(n_188)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_140),
.Y(n_157)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_157),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_126),
.B(n_80),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_126),
.B(n_104),
.C(n_84),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_159),
.B(n_164),
.C(n_90),
.Y(n_179)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_140),
.Y(n_161)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_161),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_162),
.B(n_133),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_138),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_163),
.B(n_165),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_139),
.B(n_90),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_122),
.B(n_79),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_114),
.A2(n_85),
.B(n_70),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_135),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_135),
.Y(n_168)
);

OR2x2_ASAP7_75t_L g169 ( 
.A(n_148),
.B(n_129),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_169),
.B(n_181),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_155),
.B(n_116),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_172),
.B(n_180),
.Y(n_200)
);

XOR2x2_ASAP7_75t_L g174 ( 
.A(n_153),
.B(n_134),
.Y(n_174)
);

OAI322xp33_ASAP7_75t_L g201 ( 
.A1(n_174),
.A2(n_178),
.A3(n_189),
.B1(n_180),
.B2(n_177),
.C1(n_169),
.C2(n_179),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_177),
.B(n_179),
.Y(n_209)
);

NAND3xp33_ASAP7_75t_L g178 ( 
.A(n_155),
.B(n_141),
.C(n_131),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_164),
.B(n_121),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_143),
.B(n_112),
.C(n_134),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_182),
.A2(n_88),
.B1(n_168),
.B2(n_163),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_158),
.B(n_125),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_183),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_151),
.B(n_112),
.C(n_123),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_185),
.B(n_186),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_151),
.B(n_120),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_159),
.B(n_117),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_190),
.B(n_152),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_174),
.A2(n_160),
.B1(n_146),
.B2(n_150),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_191),
.A2(n_195),
.B1(n_203),
.B2(n_190),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_189),
.A2(n_162),
.B1(n_147),
.B2(n_166),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_196),
.B(n_197),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_184),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_170),
.Y(n_198)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_198),
.Y(n_215)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_175),
.Y(n_199)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_199),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_201),
.A2(n_208),
.B1(n_185),
.B2(n_111),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_186),
.Y(n_202)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_202),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_182),
.A2(n_144),
.B1(n_167),
.B2(n_154),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_175),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_204),
.B(n_205),
.Y(n_218)
);

AOI221xp5_ASAP7_75t_L g205 ( 
.A1(n_188),
.A2(n_154),
.B1(n_152),
.B2(n_88),
.C(n_74),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_206),
.A2(n_106),
.B(n_124),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_171),
.B(n_161),
.Y(n_207)
);

INVxp33_ASAP7_75t_L g224 ( 
.A(n_207),
.Y(n_224)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_176),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_209),
.B(n_173),
.C(n_181),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_210),
.B(n_214),
.C(n_217),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_211),
.A2(n_208),
.B1(n_192),
.B2(n_199),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_206),
.A2(n_176),
.B(n_173),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_212),
.A2(n_201),
.B(n_200),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_213),
.B(n_191),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_209),
.B(n_194),
.C(n_195),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_193),
.B(n_187),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_193),
.B(n_187),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_220),
.B(n_221),
.C(n_204),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_194),
.B(n_157),
.C(n_106),
.Y(n_221)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_222),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_217),
.B(n_197),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_225),
.B(n_227),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_223),
.B(n_207),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_228),
.B(n_234),
.Y(n_239)
);

AOI221xp5_ASAP7_75t_L g229 ( 
.A1(n_218),
.A2(n_200),
.B1(n_203),
.B2(n_192),
.C(n_196),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_229),
.B(n_231),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_220),
.B(n_198),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_230),
.B(n_233),
.Y(n_243)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_215),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_235),
.A2(n_222),
.B1(n_224),
.B2(n_213),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_221),
.B(n_115),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_236),
.A2(n_237),
.B(n_219),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_216),
.A2(n_113),
.B(n_118),
.Y(n_237)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_240),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_241),
.B(n_244),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_228),
.A2(n_214),
.B1(n_211),
.B2(n_224),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_232),
.A2(n_210),
.B1(n_145),
.B2(n_115),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_245),
.B(n_231),
.C(n_226),
.Y(n_251)
);

OAI31xp33_ASAP7_75t_L g246 ( 
.A1(n_232),
.A2(n_118),
.A3(n_113),
.B(n_111),
.Y(n_246)
);

NAND2xp33_ASAP7_75t_L g248 ( 
.A(n_246),
.B(n_73),
.Y(n_248)
);

AOI31xp67_ASAP7_75t_SL g247 ( 
.A1(n_243),
.A2(n_235),
.A3(n_227),
.B(n_237),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_247),
.B(n_252),
.Y(n_256)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_248),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_251),
.A2(n_239),
.B1(n_246),
.B2(n_10),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_245),
.A2(n_226),
.B(n_8),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_242),
.B(n_10),
.C(n_2),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_253),
.B(n_238),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_249),
.B(n_242),
.C(n_240),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_255),
.B(n_257),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_258),
.B(n_10),
.Y(n_261)
);

AOI21xp33_ASAP7_75t_L g260 ( 
.A1(n_256),
.A2(n_249),
.B(n_250),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_260),
.B(n_261),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_259),
.Y(n_263)
);

AOI21xp33_ASAP7_75t_L g264 ( 
.A1(n_263),
.A2(n_254),
.B(n_258),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_264),
.A2(n_262),
.B(n_255),
.Y(n_265)
);

NAND2x1p5_ASAP7_75t_SL g266 ( 
.A(n_265),
.B(n_239),
.Y(n_266)
);


endmodule