module fake_ibex_1436_n_1543 (n_151, n_85, n_84, n_64, n_171, n_103, n_204, n_274, n_130, n_177, n_76, n_273, n_309, n_9, n_293, n_124, n_37, n_256, n_193, n_108, n_165, n_86, n_70, n_255, n_175, n_59, n_28, n_125, n_304, n_191, n_5, n_62, n_71, n_153, n_194, n_249, n_239, n_94, n_134, n_88, n_142, n_226, n_258, n_40, n_90, n_17, n_74, n_176, n_58, n_43, n_216, n_33, n_166, n_163, n_114, n_236, n_34, n_15, n_24, n_189, n_280, n_105, n_187, n_1, n_154, n_182, n_196, n_89, n_50, n_144, n_170, n_270, n_113, n_117, n_265, n_158, n_259, n_276, n_210, n_220, n_91, n_287, n_54, n_243, n_19, n_228, n_147, n_251, n_244, n_73, n_310, n_143, n_106, n_8, n_224, n_183, n_67, n_110, n_306, n_47, n_169, n_10, n_21, n_242, n_278, n_16, n_60, n_7, n_109, n_127, n_121, n_48, n_57, n_301, n_296, n_120, n_168, n_155, n_13, n_122, n_116, n_0, n_289, n_12, n_150, n_286, n_133, n_51, n_215, n_279, n_49, n_235, n_22, n_136, n_261, n_30, n_221, n_102, n_52, n_99, n_269, n_156, n_126, n_25, n_104, n_45, n_141, n_222, n_186, n_295, n_230, n_96, n_185, n_290, n_174, n_157, n_219, n_246, n_31, n_146, n_207, n_167, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_205, n_139, n_275, n_98, n_129, n_267, n_245, n_229, n_209, n_82, n_263, n_27, n_299, n_87, n_262, n_75, n_137, n_173, n_180, n_201, n_14, n_257, n_77, n_44, n_66, n_305, n_307, n_192, n_140, n_4, n_6, n_100, n_179, n_206, n_26, n_188, n_200, n_199, n_308, n_135, n_283, n_111, n_36, n_18, n_53, n_227, n_115, n_11, n_248, n_92, n_101, n_190, n_138, n_214, n_238, n_211, n_218, n_132, n_277, n_225, n_272, n_23, n_223, n_95, n_285, n_288, n_247, n_55, n_291, n_63, n_161, n_237, n_29, n_203, n_268, n_148, n_2, n_233, n_118, n_164, n_38, n_198, n_264, n_217, n_78, n_20, n_69, n_39, n_178, n_303, n_93, n_162, n_240, n_282, n_61, n_266, n_42, n_294, n_112, n_46, n_284, n_80, n_172, n_250, n_119, n_72, n_195, n_212, n_97, n_197, n_181, n_131, n_123, n_260, n_302, n_297, n_41, n_252, n_83, n_32, n_107, n_149, n_254, n_213, n_271, n_241, n_68, n_292, n_79, n_81, n_35, n_159, n_202, n_231, n_298, n_160, n_184, n_56, n_232, n_281, n_1543);

input n_151;
input n_85;
input n_84;
input n_64;
input n_171;
input n_103;
input n_204;
input n_274;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_9;
input n_293;
input n_124;
input n_37;
input n_256;
input n_193;
input n_108;
input n_165;
input n_86;
input n_70;
input n_255;
input n_175;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_5;
input n_62;
input n_71;
input n_153;
input n_194;
input n_249;
input n_239;
input n_94;
input n_134;
input n_88;
input n_142;
input n_226;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_166;
input n_163;
input n_114;
input n_236;
input n_34;
input n_15;
input n_24;
input n_189;
input n_280;
input n_105;
input n_187;
input n_1;
input n_154;
input n_182;
input n_196;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_113;
input n_117;
input n_265;
input n_158;
input n_259;
input n_276;
input n_210;
input n_220;
input n_91;
input n_287;
input n_54;
input n_243;
input n_19;
input n_228;
input n_147;
input n_251;
input n_244;
input n_73;
input n_310;
input n_143;
input n_106;
input n_8;
input n_224;
input n_183;
input n_67;
input n_110;
input n_306;
input n_47;
input n_169;
input n_10;
input n_21;
input n_242;
input n_278;
input n_16;
input n_60;
input n_7;
input n_109;
input n_127;
input n_121;
input n_48;
input n_57;
input n_301;
input n_296;
input n_120;
input n_168;
input n_155;
input n_13;
input n_122;
input n_116;
input n_0;
input n_289;
input n_12;
input n_150;
input n_286;
input n_133;
input n_51;
input n_215;
input n_279;
input n_49;
input n_235;
input n_22;
input n_136;
input n_261;
input n_30;
input n_221;
input n_102;
input n_52;
input n_99;
input n_269;
input n_156;
input n_126;
input n_25;
input n_104;
input n_45;
input n_141;
input n_222;
input n_186;
input n_295;
input n_230;
input n_96;
input n_185;
input n_290;
input n_174;
input n_157;
input n_219;
input n_246;
input n_31;
input n_146;
input n_207;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_205;
input n_139;
input n_275;
input n_98;
input n_129;
input n_267;
input n_245;
input n_229;
input n_209;
input n_82;
input n_263;
input n_27;
input n_299;
input n_87;
input n_262;
input n_75;
input n_137;
input n_173;
input n_180;
input n_201;
input n_14;
input n_257;
input n_77;
input n_44;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_4;
input n_6;
input n_100;
input n_179;
input n_206;
input n_26;
input n_188;
input n_200;
input n_199;
input n_308;
input n_135;
input n_283;
input n_111;
input n_36;
input n_18;
input n_53;
input n_227;
input n_115;
input n_11;
input n_248;
input n_92;
input n_101;
input n_190;
input n_138;
input n_214;
input n_238;
input n_211;
input n_218;
input n_132;
input n_277;
input n_225;
input n_272;
input n_23;
input n_223;
input n_95;
input n_285;
input n_288;
input n_247;
input n_55;
input n_291;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_148;
input n_2;
input n_233;
input n_118;
input n_164;
input n_38;
input n_198;
input n_264;
input n_217;
input n_78;
input n_20;
input n_69;
input n_39;
input n_178;
input n_303;
input n_93;
input n_162;
input n_240;
input n_282;
input n_61;
input n_266;
input n_42;
input n_294;
input n_112;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_119;
input n_72;
input n_195;
input n_212;
input n_97;
input n_197;
input n_181;
input n_131;
input n_123;
input n_260;
input n_302;
input n_297;
input n_41;
input n_252;
input n_83;
input n_32;
input n_107;
input n_149;
input n_254;
input n_213;
input n_271;
input n_241;
input n_68;
input n_292;
input n_79;
input n_81;
input n_35;
input n_159;
input n_202;
input n_231;
input n_298;
input n_160;
input n_184;
input n_56;
input n_232;
input n_281;

output n_1543;

wire n_1084;
wire n_1474;
wire n_1295;
wire n_507;
wire n_992;
wire n_766;
wire n_1110;
wire n_1382;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_446;
wire n_452;
wire n_1234;
wire n_773;
wire n_1469;
wire n_821;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_957;
wire n_678;
wire n_969;
wire n_1125;
wire n_733;
wire n_312;
wire n_622;
wire n_1226;
wire n_1034;
wire n_872;
wire n_457;
wire n_494;
wire n_930;
wire n_1044;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_911;
wire n_652;
wire n_781;
wire n_475;
wire n_802;
wire n_1233;
wire n_1045;
wire n_500;
wire n_963;
wire n_376;
wire n_531;
wire n_1308;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_375;
wire n_1391;
wire n_667;
wire n_884;
wire n_850;
wire n_879;
wire n_723;
wire n_1144;
wire n_346;
wire n_1392;
wire n_1268;
wire n_739;
wire n_853;
wire n_504;
wire n_948;
wire n_1338;
wire n_875;
wire n_1307;
wire n_1327;
wire n_481;
wire n_876;
wire n_497;
wire n_711;
wire n_671;
wire n_989;
wire n_829;
wire n_825;
wire n_1480;
wire n_1463;
wire n_939;
wire n_655;
wire n_550;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_496;
wire n_434;
wire n_1258;
wire n_1344;
wire n_835;
wire n_1195;
wire n_824;
wire n_441;
wire n_694;
wire n_523;
wire n_787;
wire n_614;
wire n_431;
wire n_1130;
wire n_1228;
wire n_321;
wire n_1081;
wire n_374;
wire n_538;
wire n_1155;
wire n_1292;
wire n_459;
wire n_518;
wire n_852;
wire n_1427;
wire n_1133;
wire n_904;
wire n_355;
wire n_448;
wire n_646;
wire n_466;
wire n_1030;
wire n_1094;
wire n_1496;
wire n_715;
wire n_530;
wire n_1214;
wire n_1274;
wire n_420;
wire n_769;
wire n_1509;
wire n_857;
wire n_765;
wire n_1070;
wire n_777;
wire n_331;
wire n_917;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_1493;
wire n_1313;
wire n_352;
wire n_558;
wire n_666;
wire n_1071;
wire n_1449;
wire n_793;
wire n_937;
wire n_973;
wire n_1038;
wire n_618;
wire n_1269;
wire n_662;
wire n_979;
wire n_1309;
wire n_1316;
wire n_1215;
wire n_629;
wire n_1445;
wire n_573;
wire n_359;
wire n_1466;
wire n_1412;
wire n_433;
wire n_439;
wire n_1007;
wire n_643;
wire n_1276;
wire n_841;
wire n_772;
wire n_810;
wire n_338;
wire n_1401;
wire n_369;
wire n_1301;
wire n_869;
wire n_718;
wire n_553;
wire n_554;
wire n_1078;
wire n_1219;
wire n_713;
wire n_1252;
wire n_1170;
wire n_605;
wire n_539;
wire n_630;
wire n_567;
wire n_745;
wire n_447;
wire n_564;
wire n_562;
wire n_1322;
wire n_1305;
wire n_795;
wire n_592;
wire n_1248;
wire n_762;
wire n_1388;
wire n_800;
wire n_706;
wire n_784;
wire n_684;
wire n_1375;
wire n_397;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_709;
wire n_1296;
wire n_499;
wire n_702;
wire n_971;
wire n_1326;
wire n_451;
wire n_1350;
wire n_906;
wire n_1093;
wire n_978;
wire n_579;
wire n_899;
wire n_1019;
wire n_902;
wire n_1250;
wire n_1190;
wire n_1304;
wire n_744;
wire n_314;
wire n_563;
wire n_1506;
wire n_881;
wire n_734;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_382;
wire n_1423;
wire n_1239;
wire n_1370;
wire n_1209;
wire n_379;
wire n_551;
wire n_729;
wire n_1434;
wire n_603;
wire n_422;
wire n_324;
wire n_391;
wire n_820;
wire n_805;
wire n_670;
wire n_1132;
wire n_892;
wire n_390;
wire n_1467;
wire n_544;
wire n_1281;
wire n_1447;
wire n_695;
wire n_639;
wire n_1531;
wire n_1332;
wire n_482;
wire n_1424;
wire n_870;
wire n_1298;
wire n_1387;
wire n_609;
wire n_1040;
wire n_476;
wire n_1159;
wire n_1368;
wire n_1154;
wire n_345;
wire n_455;
wire n_1243;
wire n_1121;
wire n_693;
wire n_406;
wire n_606;
wire n_737;
wire n_462;
wire n_1407;
wire n_1235;
wire n_1003;
wire n_889;
wire n_435;
wire n_396;
wire n_816;
wire n_1058;
wire n_399;
wire n_823;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1441;
wire n_657;
wire n_1156;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1394;
wire n_1347;
wire n_819;
wire n_822;
wire n_1042;
wire n_743;
wire n_754;
wire n_395;
wire n_1319;
wire n_389;
wire n_1041;
wire n_1090;
wire n_1196;
wire n_330;
wire n_1182;
wire n_1271;
wire n_1031;
wire n_372;
wire n_981;
wire n_350;
wire n_398;
wire n_583;
wire n_1409;
wire n_1015;
wire n_663;
wire n_1377;
wire n_1521;
wire n_1152;
wire n_371;
wire n_1036;
wire n_974;
wire n_608;
wire n_864;
wire n_412;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_449;
wire n_1452;
wire n_1318;
wire n_1508;
wire n_421;
wire n_738;
wire n_1217;
wire n_1189;
wire n_761;
wire n_748;
wire n_901;
wire n_340;
wire n_1255;
wire n_1218;
wire n_1181;
wire n_1140;
wire n_1056;
wire n_1283;
wire n_1446;
wire n_1487;
wire n_840;
wire n_1203;
wire n_1421;
wire n_561;
wire n_846;
wire n_471;
wire n_1237;
wire n_859;
wire n_1109;
wire n_965;
wire n_384;
wire n_1051;
wire n_1008;
wire n_458;
wire n_1498;
wire n_1053;
wire n_1207;
wire n_1076;
wire n_1032;
wire n_936;
wire n_469;
wire n_1210;
wire n_591;
wire n_1510;
wire n_1201;
wire n_1246;
wire n_732;
wire n_1236;
wire n_832;
wire n_316;
wire n_590;
wire n_325;
wire n_1184;
wire n_1477;
wire n_1364;
wire n_1540;
wire n_1013;
wire n_929;
wire n_315;
wire n_637;
wire n_1136;
wire n_1075;
wire n_1249;
wire n_574;
wire n_515;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_907;
wire n_1179;
wire n_1153;
wire n_669;
wire n_521;
wire n_1117;
wire n_1273;
wire n_1083;
wire n_1014;
wire n_724;
wire n_437;
wire n_938;
wire n_1178;
wire n_474;
wire n_878;
wire n_594;
wire n_1464;
wire n_944;
wire n_623;
wire n_585;
wire n_1334;
wire n_483;
wire n_1418;
wire n_1137;
wire n_660;
wire n_524;
wire n_1200;
wire n_1120;
wire n_576;
wire n_388;
wire n_1522;
wire n_1279;
wire n_931;
wire n_607;
wire n_827;
wire n_1064;
wire n_1408;
wire n_1028;
wire n_1264;
wire n_1146;
wire n_358;
wire n_488;
wire n_705;
wire n_429;
wire n_1009;
wire n_1260;
wire n_589;
wire n_472;
wire n_347;
wire n_847;
wire n_1436;
wire n_413;
wire n_1069;
wire n_1485;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_679;
wire n_1345;
wire n_696;
wire n_837;
wire n_640;
wire n_954;
wire n_363;
wire n_725;
wire n_596;
wire n_351;
wire n_456;
wire n_1471;
wire n_1115;
wire n_998;
wire n_1395;
wire n_801;
wire n_1479;
wire n_1046;
wire n_882;
wire n_942;
wire n_1431;
wire n_651;
wire n_721;
wire n_365;
wire n_814;
wire n_943;
wire n_1086;
wire n_1523;
wire n_1470;
wire n_444;
wire n_986;
wire n_495;
wire n_1420;
wire n_411;
wire n_927;
wire n_615;
wire n_803;
wire n_1087;
wire n_757;
wire n_1400;
wire n_712;
wire n_1539;
wire n_650;
wire n_409;
wire n_332;
wire n_1448;
wire n_517;
wire n_817;
wire n_555;
wire n_337;
wire n_951;
wire n_468;
wire n_780;
wire n_502;
wire n_633;
wire n_726;
wire n_532;
wire n_1439;
wire n_863;
wire n_597;
wire n_1128;
wire n_1266;
wire n_1300;
wire n_318;
wire n_807;
wire n_741;
wire n_430;
wire n_486;
wire n_1405;
wire n_997;
wire n_1428;
wire n_891;
wire n_1528;
wire n_1495;
wire n_717;
wire n_1357;
wire n_1512;
wire n_668;
wire n_871;
wire n_1339;
wire n_1426;
wire n_485;
wire n_1315;
wire n_1413;
wire n_811;
wire n_808;
wire n_945;
wire n_460;
wire n_1461;
wire n_461;
wire n_903;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_1378;
wire n_1048;
wire n_774;
wire n_588;
wire n_1430;
wire n_1251;
wire n_1247;
wire n_528;
wire n_836;
wire n_1475;
wire n_1263;
wire n_443;
wire n_1185;
wire n_344;
wire n_436;
wire n_1122;
wire n_890;
wire n_628;
wire n_874;
wire n_1505;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_916;
wire n_503;
wire n_895;
wire n_687;
wire n_1035;
wire n_1535;
wire n_751;
wire n_1127;
wire n_932;
wire n_380;
wire n_1004;
wire n_947;
wire n_831;
wire n_778;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1104;
wire n_1011;
wire n_1437;
wire n_529;
wire n_626;
wire n_1497;
wire n_1143;
wire n_328;
wire n_418;
wire n_510;
wire n_972;
wire n_601;
wire n_610;
wire n_1444;
wire n_920;
wire n_664;
wire n_1067;
wire n_994;
wire n_545;
wire n_887;
wire n_1162;
wire n_334;
wire n_634;
wire n_961;
wire n_991;
wire n_1223;
wire n_1349;
wire n_1331;
wire n_1323;
wire n_578;
wire n_432;
wire n_403;
wire n_1353;
wire n_423;
wire n_357;
wire n_1429;
wire n_1432;
wire n_1320;
wire n_996;
wire n_915;
wire n_1174;
wire n_1286;
wire n_542;
wire n_1294;
wire n_900;
wire n_1351;
wire n_377;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_317;
wire n_1458;
wire n_1460;
wire n_326;
wire n_1340;
wire n_339;
wire n_348;
wire n_674;
wire n_552;
wire n_1112;
wire n_1267;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_703;
wire n_426;
wire n_1172;
wire n_1099;
wire n_598;
wire n_1422;
wire n_508;
wire n_453;
wire n_1527;
wire n_400;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_404;
wire n_1177;
wire n_1025;
wire n_1517;
wire n_690;
wire n_1225;
wire n_982;
wire n_785;
wire n_604;
wire n_977;
wire n_719;
wire n_370;
wire n_1491;
wire n_716;
wire n_923;
wire n_642;
wire n_933;
wire n_1037;
wire n_464;
wire n_1348;
wire n_838;
wire n_1289;
wire n_1021;
wire n_746;
wire n_1188;
wire n_742;
wire n_1191;
wire n_1503;
wire n_1052;
wire n_789;
wire n_656;
wire n_602;
wire n_842;
wire n_767;
wire n_636;
wire n_1259;
wire n_407;
wire n_490;
wire n_595;
wire n_1001;
wire n_570;
wire n_1396;
wire n_1224;
wire n_356;
wire n_1538;
wire n_487;
wire n_349;
wire n_454;
wire n_1017;
wire n_730;
wire n_1456;
wire n_625;
wire n_619;
wire n_1124;
wire n_611;
wire n_922;
wire n_851;
wire n_993;
wire n_1135;
wire n_541;
wire n_613;
wire n_659;
wire n_1494;
wire n_1066;
wire n_1169;
wire n_571;
wire n_648;
wire n_830;
wire n_473;
wire n_1241;
wire n_445;
wire n_1072;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_353;
wire n_826;
wire n_1337;
wire n_839;
wire n_768;
wire n_1278;
wire n_796;
wire n_797;
wire n_1006;
wire n_402;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1063;
wire n_1270;
wire n_834;
wire n_1476;
wire n_935;
wire n_925;
wire n_1054;
wire n_722;
wire n_1406;
wire n_1489;
wire n_804;
wire n_484;
wire n_1455;
wire n_480;
wire n_354;
wire n_1057;
wire n_1473;
wire n_516;
wire n_1403;
wire n_329;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_506;
wire n_868;
wire n_1202;
wire n_1065;
wire n_1457;
wire n_905;
wire n_975;
wire n_675;
wire n_463;
wire n_624;
wire n_520;
wire n_934;
wire n_775;
wire n_950;
wire n_512;
wire n_685;
wire n_1222;
wire n_1198;
wire n_1311;
wire n_1261;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_1282;
wire n_1321;
wire n_700;
wire n_360;
wire n_1107;
wire n_525;
wire n_815;
wire n_919;
wire n_535;
wire n_681;
wire n_415;
wire n_320;
wire n_1411;
wire n_1139;
wire n_858;
wire n_1018;
wire n_385;
wire n_1324;
wire n_1501;
wire n_782;
wire n_616;
wire n_833;
wire n_1343;
wire n_1371;
wire n_1513;
wire n_728;
wire n_786;
wire n_362;
wire n_505;
wire n_1342;
wire n_501;
wire n_752;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1221;
wire n_1047;
wire n_1515;
wire n_1374;
wire n_1435;
wire n_792;
wire n_1314;
wire n_1433;
wire n_575;
wire n_313;
wire n_1242;
wire n_1119;
wire n_1085;
wire n_419;
wire n_885;
wire n_1530;
wire n_513;
wire n_877;
wire n_311;
wire n_1088;
wire n_896;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_393;
wire n_428;
wire n_697;
wire n_1105;
wire n_1459;
wire n_912;
wire n_424;
wire n_701;
wire n_995;
wire n_1000;
wire n_1256;
wire n_587;
wire n_1303;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_855;
wire n_812;
wire n_1050;
wire n_599;
wire n_1060;
wire n_1372;
wire n_756;
wire n_1257;
wire n_387;
wire n_688;
wire n_1542;
wire n_946;
wire n_707;
wire n_1362;
wire n_1097;
wire n_341;
wire n_621;
wire n_956;
wire n_790;
wire n_1541;
wire n_586;
wire n_1330;
wire n_638;
wire n_593;
wire n_1212;
wire n_1199;
wire n_1443;
wire n_478;
wire n_336;
wire n_861;
wire n_1389;
wire n_1131;
wire n_547;
wire n_727;
wire n_1077;
wire n_1481;
wire n_828;
wire n_1438;
wire n_753;
wire n_645;
wire n_747;
wire n_1147;
wire n_1363;
wire n_1098;
wire n_584;
wire n_1366;
wire n_1518;
wire n_1361;
wire n_1187;
wire n_698;
wire n_1061;
wire n_682;
wire n_1373;
wire n_327;
wire n_1302;
wire n_383;
wire n_886;
wire n_1010;
wire n_883;
wire n_417;
wire n_755;
wire n_1029;
wire n_470;
wire n_770;
wire n_941;
wire n_1245;
wire n_1317;
wire n_632;
wire n_1329;
wire n_373;
wire n_854;
wire n_343;
wire n_714;
wire n_1297;
wire n_1369;
wire n_323;
wire n_740;
wire n_386;
wire n_549;
wire n_533;
wire n_928;
wire n_898;
wire n_333;
wire n_1285;
wire n_967;
wire n_736;
wire n_1529;
wire n_1381;
wire n_1103;
wire n_1161;
wire n_465;
wire n_1486;
wire n_1068;
wire n_617;
wire n_914;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1197;
wire n_1168;
wire n_865;
wire n_569;
wire n_600;
wire n_1192;
wire n_1290;
wire n_987;
wire n_750;
wire n_1299;
wire n_665;
wire n_1101;
wire n_367;
wire n_880;
wire n_654;
wire n_731;
wire n_1336;
wire n_758;
wire n_1166;
wire n_720;
wire n_710;
wire n_1390;
wire n_1023;
wire n_568;
wire n_1358;
wire n_813;
wire n_1211;
wire n_1397;
wire n_1284;
wire n_1359;
wire n_1116;
wire n_791;
wire n_1532;
wire n_1419;
wire n_543;
wire n_580;
wire n_1082;
wire n_1213;
wire n_1193;
wire n_980;
wire n_849;
wire n_1488;
wire n_1074;
wire n_759;
wire n_1379;
wire n_953;
wire n_1180;
wire n_1462;
wire n_536;
wire n_1220;
wire n_467;
wire n_1398;
wire n_427;
wire n_1262;
wire n_442;
wire n_438;
wire n_1012;
wire n_689;
wire n_960;
wire n_1022;
wire n_676;
wire n_1240;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_771;
wire n_999;
wire n_514;
wire n_1092;
wire n_560;
wire n_1386;
wire n_910;
wire n_635;
wire n_844;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1385;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_335;
wire n_1499;
wire n_1500;
wire n_966;
wire n_949;
wire n_704;
wire n_924;
wire n_477;
wire n_699;
wire n_368;
wire n_918;
wire n_672;
wire n_1039;
wire n_401;
wire n_1043;
wire n_1402;
wire n_735;
wire n_1450;
wire n_566;
wire n_416;
wire n_581;
wire n_1472;
wire n_1365;
wire n_1089;
wire n_392;
wire n_1536;
wire n_1049;
wire n_548;
wire n_1158;
wire n_763;
wire n_940;
wire n_1404;
wire n_546;
wire n_788;
wire n_410;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1216;
wire n_1026;
wire n_366;
wire n_1454;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_322;
wire n_888;
wire n_1325;
wire n_582;
wire n_1483;
wire n_653;
wire n_1205;
wire n_843;
wire n_1059;
wire n_799;
wire n_691;
wire n_522;
wire n_479;
wire n_534;
wire n_511;
wire n_381;
wire n_1414;
wire n_1002;
wire n_1111;
wire n_1341;
wire n_405;
wire n_1310;
wire n_612;
wire n_955;
wire n_440;
wire n_1333;
wire n_342;
wire n_414;
wire n_378;
wire n_952;
wire n_1145;
wire n_1533;
wire n_1511;
wire n_537;
wire n_1113;
wire n_1468;
wire n_913;
wire n_509;
wire n_1164;
wire n_1354;
wire n_1277;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_856;
wire n_779;
wire n_1280;
wire n_493;
wire n_1335;
wire n_519;
wire n_408;
wire n_361;
wire n_319;
wire n_1091;
wire n_1287;
wire n_1482;
wire n_860;
wire n_1525;
wire n_661;
wire n_848;
wire n_683;
wire n_1150;
wire n_1194;
wire n_620;
wire n_1399;
wire n_450;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_577;
wire n_970;
wire n_491;
wire n_921;
wire n_489;
wire n_1534;
wire n_908;
wire n_1346;
wire n_565;
wire n_1123;
wire n_1272;
wire n_1393;
wire n_984;
wire n_394;
wire n_364;
wire n_1410;
wire n_988;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_492;
wire n_649;
wire n_866;
wire n_559;
wire n_425;

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_117),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_6),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_2),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_225),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_192),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_173),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_232),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_219),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_239),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_69),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_269),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_64),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_201),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_22),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_242),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_258),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_38),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_260),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_246),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_119),
.Y(n_330)
);

CKINVDCx14_ASAP7_75t_R g331 ( 
.A(n_296),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_130),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_82),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_282),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_274),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_196),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_247),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_113),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_280),
.Y(n_339)
);

INVx2_ASAP7_75t_SL g340 ( 
.A(n_255),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_248),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_216),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_307),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_281),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_291),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_98),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_297),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_253),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_157),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_283),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_301),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_287),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_276),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_302),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_256),
.Y(n_355)
);

BUFx10_ASAP7_75t_L g356 ( 
.A(n_124),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_303),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_251),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_179),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_208),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_146),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_306),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_150),
.Y(n_363)
);

BUFx10_ASAP7_75t_L g364 ( 
.A(n_217),
.Y(n_364)
);

INVx1_ASAP7_75t_SL g365 ( 
.A(n_295),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_125),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_263),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_226),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_262),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_69),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_259),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_300),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_268),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_308),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_136),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_170),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_61),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_95),
.Y(n_378)
);

BUFx10_ASAP7_75t_L g379 ( 
.A(n_40),
.Y(n_379)
);

BUFx5_ASAP7_75t_L g380 ( 
.A(n_310),
.Y(n_380)
);

INVx1_ASAP7_75t_SL g381 ( 
.A(n_178),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_14),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_168),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_165),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_215),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_257),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_71),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_285),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_305),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_23),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_250),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_233),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_309),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_205),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_36),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_74),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_19),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_266),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_65),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_293),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_227),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_131),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_167),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_41),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_22),
.Y(n_405)
);

CKINVDCx16_ASAP7_75t_R g406 ( 
.A(n_265),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_84),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_60),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_30),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_55),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_166),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_174),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_289),
.Y(n_413)
);

INVx2_ASAP7_75t_SL g414 ( 
.A(n_207),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_16),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_3),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_206),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_202),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_198),
.Y(n_419)
);

BUFx10_ASAP7_75t_L g420 ( 
.A(n_241),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_264),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_111),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_175),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_102),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_74),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_31),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_12),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_243),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_186),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_237),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_286),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_98),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_171),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_223),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_31),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_46),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_244),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_70),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_267),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_138),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_272),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_16),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_236),
.Y(n_443)
);

INVx1_ASAP7_75t_SL g444 ( 
.A(n_144),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_123),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_230),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_77),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_229),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_261),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_240),
.Y(n_450)
);

INVx1_ASAP7_75t_SL g451 ( 
.A(n_10),
.Y(n_451)
);

CKINVDCx16_ASAP7_75t_R g452 ( 
.A(n_163),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_252),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_190),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_145),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_78),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_92),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_96),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_210),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_86),
.Y(n_460)
);

CKINVDCx16_ASAP7_75t_R g461 ( 
.A(n_177),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_23),
.Y(n_462)
);

BUFx10_ASAP7_75t_L g463 ( 
.A(n_102),
.Y(n_463)
);

BUFx3_ASAP7_75t_L g464 ( 
.A(n_15),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_249),
.Y(n_465)
);

BUFx3_ASAP7_75t_L g466 ( 
.A(n_273),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_43),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_200),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_299),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_182),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_140),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_7),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_21),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_7),
.Y(n_474)
);

INVxp67_ASAP7_75t_L g475 ( 
.A(n_169),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_277),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_197),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_112),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_78),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_235),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_148),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_84),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_172),
.Y(n_483)
);

BUFx2_ASAP7_75t_L g484 ( 
.A(n_161),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_73),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_304),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_224),
.Y(n_487)
);

CKINVDCx16_ASAP7_75t_R g488 ( 
.A(n_43),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_55),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_81),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_30),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_122),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_220),
.Y(n_493)
);

BUFx2_ASAP7_75t_R g494 ( 
.A(n_94),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_228),
.Y(n_495)
);

INVx2_ASAP7_75t_SL g496 ( 
.A(n_290),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_176),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_107),
.Y(n_498)
);

HB1xp67_ASAP7_75t_L g499 ( 
.A(n_222),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_254),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_3),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_189),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_294),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_61),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_6),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_38),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_155),
.Y(n_507)
);

INVx1_ASAP7_75t_SL g508 ( 
.A(n_164),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_142),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_37),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_187),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_238),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_91),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_284),
.Y(n_514)
);

CKINVDCx16_ASAP7_75t_R g515 ( 
.A(n_270),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_4),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_245),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_234),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_183),
.Y(n_519)
);

HB1xp67_ASAP7_75t_L g520 ( 
.A(n_279),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_54),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_298),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_5),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_153),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_275),
.Y(n_525)
);

BUFx5_ASAP7_75t_L g526 ( 
.A(n_15),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_288),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_90),
.Y(n_528)
);

BUFx6f_ASAP7_75t_L g529 ( 
.A(n_139),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_48),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_89),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_25),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_5),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_212),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_271),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_94),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_292),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_278),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_4),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_231),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_96),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_128),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_108),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_54),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_499),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_520),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_484),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_464),
.Y(n_548)
);

CKINVDCx20_ASAP7_75t_R g549 ( 
.A(n_488),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_323),
.Y(n_550)
);

HB1xp67_ASAP7_75t_L g551 ( 
.A(n_464),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_521),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_340),
.B(n_414),
.Y(n_553)
);

CKINVDCx20_ASAP7_75t_R g554 ( 
.A(n_324),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_329),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_521),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_539),
.Y(n_557)
);

INVxp67_ASAP7_75t_SL g558 ( 
.A(n_539),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_541),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_541),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_526),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_526),
.Y(n_562)
);

HB1xp67_ASAP7_75t_L g563 ( 
.A(n_312),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_526),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_344),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_367),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_369),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_526),
.Y(n_568)
);

CKINVDCx20_ASAP7_75t_R g569 ( 
.A(n_382),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_526),
.Y(n_570)
);

INVxp67_ASAP7_75t_SL g571 ( 
.A(n_370),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_526),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_389),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_413),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_387),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_430),
.Y(n_576)
);

CKINVDCx20_ASAP7_75t_R g577 ( 
.A(n_396),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_395),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_405),
.Y(n_579)
);

CKINVDCx20_ASAP7_75t_R g580 ( 
.A(n_440),
.Y(n_580)
);

CKINVDCx20_ASAP7_75t_R g581 ( 
.A(n_441),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_465),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_408),
.Y(n_583)
);

INVxp67_ASAP7_75t_SL g584 ( 
.A(n_409),
.Y(n_584)
);

INVxp67_ASAP7_75t_SL g585 ( 
.A(n_415),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_416),
.Y(n_586)
);

CKINVDCx20_ASAP7_75t_R g587 ( 
.A(n_477),
.Y(n_587)
);

INVxp67_ASAP7_75t_L g588 ( 
.A(n_424),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_435),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_483),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_438),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_493),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_447),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_456),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_462),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_380),
.Y(n_596)
);

CKINVDCx20_ASAP7_75t_R g597 ( 
.A(n_514),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_519),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_406),
.Y(n_599)
);

CKINVDCx20_ASAP7_75t_R g600 ( 
.A(n_452),
.Y(n_600)
);

CKINVDCx20_ASAP7_75t_R g601 ( 
.A(n_461),
.Y(n_601)
);

BUFx3_ASAP7_75t_L g602 ( 
.A(n_466),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_515),
.Y(n_603)
);

BUFx2_ASAP7_75t_SL g604 ( 
.A(n_356),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_474),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_491),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_501),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_331),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_380),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_R g610 ( 
.A(n_331),
.B(n_104),
.Y(n_610)
);

CKINVDCx20_ASAP7_75t_R g611 ( 
.A(n_379),
.Y(n_611)
);

NOR2xp67_ASAP7_75t_L g612 ( 
.A(n_505),
.B(n_0),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_313),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_510),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_320),
.Y(n_615)
);

HB1xp67_ASAP7_75t_L g616 ( 
.A(n_322),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_327),
.Y(n_617)
);

HB1xp67_ASAP7_75t_L g618 ( 
.A(n_333),
.Y(n_618)
);

CKINVDCx20_ASAP7_75t_R g619 ( 
.A(n_379),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_528),
.Y(n_620)
);

INVxp67_ASAP7_75t_SL g621 ( 
.A(n_530),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_536),
.Y(n_622)
);

BUFx6f_ASAP7_75t_L g623 ( 
.A(n_568),
.Y(n_623)
);

CKINVDCx20_ASAP7_75t_R g624 ( 
.A(n_569),
.Y(n_624)
);

BUFx6f_ASAP7_75t_L g625 ( 
.A(n_568),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_548),
.B(n_496),
.Y(n_626)
);

AND2x4_ASAP7_75t_L g627 ( 
.A(n_545),
.B(n_346),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_551),
.Y(n_628)
);

INVx3_ASAP7_75t_L g629 ( 
.A(n_602),
.Y(n_629)
);

CKINVDCx20_ASAP7_75t_R g630 ( 
.A(n_569),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_602),
.Y(n_631)
);

CKINVDCx20_ASAP7_75t_R g632 ( 
.A(n_577),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_553),
.B(n_377),
.Y(n_633)
);

AND3x2_ASAP7_75t_L g634 ( 
.A(n_563),
.B(n_494),
.C(n_475),
.Y(n_634)
);

CKINVDCx20_ASAP7_75t_R g635 ( 
.A(n_577),
.Y(n_635)
);

BUFx6f_ASAP7_75t_L g636 ( 
.A(n_596),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_546),
.B(n_378),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_558),
.B(n_316),
.Y(n_638)
);

BUFx6f_ASAP7_75t_L g639 ( 
.A(n_596),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_616),
.B(n_463),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_618),
.B(n_463),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_561),
.Y(n_642)
);

AND2x4_ASAP7_75t_L g643 ( 
.A(n_547),
.B(n_571),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_555),
.Y(n_644)
);

AND2x4_ASAP7_75t_L g645 ( 
.A(n_584),
.B(n_346),
.Y(n_645)
);

HB1xp67_ASAP7_75t_L g646 ( 
.A(n_613),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_562),
.Y(n_647)
);

BUFx2_ASAP7_75t_L g648 ( 
.A(n_615),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_608),
.B(n_617),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_565),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_564),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_570),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_572),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_566),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_588),
.B(n_356),
.Y(n_655)
);

BUFx6f_ASAP7_75t_L g656 ( 
.A(n_609),
.Y(n_656)
);

INVx3_ASAP7_75t_L g657 ( 
.A(n_609),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_567),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_575),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_578),
.B(n_316),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_R g661 ( 
.A(n_600),
.B(n_311),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_579),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_583),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_552),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_573),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_586),
.Y(n_666)
);

HB1xp67_ASAP7_75t_L g667 ( 
.A(n_599),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_589),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_591),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_574),
.Y(n_670)
);

BUFx2_ASAP7_75t_L g671 ( 
.A(n_603),
.Y(n_671)
);

CKINVDCx20_ASAP7_75t_R g672 ( 
.A(n_554),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_593),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_604),
.B(n_364),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_594),
.Y(n_675)
);

INVx4_ASAP7_75t_L g676 ( 
.A(n_595),
.Y(n_676)
);

BUFx6f_ASAP7_75t_L g677 ( 
.A(n_556),
.Y(n_677)
);

CKINVDCx20_ASAP7_75t_R g678 ( 
.A(n_580),
.Y(n_678)
);

BUFx6f_ASAP7_75t_L g679 ( 
.A(n_557),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_605),
.B(n_390),
.Y(n_680)
);

BUFx6f_ASAP7_75t_L g681 ( 
.A(n_559),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_576),
.Y(n_682)
);

AND2x4_ASAP7_75t_L g683 ( 
.A(n_585),
.B(n_346),
.Y(n_683)
);

INVxp67_ASAP7_75t_L g684 ( 
.A(n_582),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_606),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_607),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_622),
.B(n_614),
.Y(n_687)
);

CKINVDCx20_ASAP7_75t_R g688 ( 
.A(n_580),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_620),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_560),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_R g691 ( 
.A(n_600),
.B(n_314),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_590),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_621),
.Y(n_693)
);

INVx3_ASAP7_75t_L g694 ( 
.A(n_612),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_592),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_598),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_610),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_581),
.Y(n_698)
);

NOR2xp67_ASAP7_75t_L g699 ( 
.A(n_611),
.B(n_317),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_581),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_611),
.Y(n_701)
);

AND2x2_ASAP7_75t_L g702 ( 
.A(n_619),
.B(n_364),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_619),
.B(n_385),
.Y(n_703)
);

CKINVDCx20_ASAP7_75t_R g704 ( 
.A(n_587),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_601),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_601),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_549),
.Y(n_707)
);

INVx3_ASAP7_75t_L g708 ( 
.A(n_549),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_587),
.B(n_420),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_597),
.B(n_397),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_597),
.Y(n_711)
);

BUFx6f_ASAP7_75t_L g712 ( 
.A(n_568),
.Y(n_712)
);

HB1xp67_ASAP7_75t_L g713 ( 
.A(n_616),
.Y(n_713)
);

BUFx6f_ASAP7_75t_L g714 ( 
.A(n_568),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_551),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_550),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_551),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_551),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_551),
.Y(n_719)
);

HB1xp67_ASAP7_75t_L g720 ( 
.A(n_616),
.Y(n_720)
);

CKINVDCx20_ASAP7_75t_R g721 ( 
.A(n_569),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_550),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_547),
.B(n_315),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_551),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_550),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_551),
.Y(n_726)
);

INVx3_ASAP7_75t_L g727 ( 
.A(n_602),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_602),
.Y(n_728)
);

HB1xp67_ASAP7_75t_L g729 ( 
.A(n_616),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_551),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_551),
.Y(n_731)
);

INVx6_ASAP7_75t_L g732 ( 
.A(n_602),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_602),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_602),
.Y(n_734)
);

CKINVDCx20_ASAP7_75t_R g735 ( 
.A(n_569),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_551),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_548),
.B(n_385),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_551),
.Y(n_738)
);

BUFx6f_ASAP7_75t_L g739 ( 
.A(n_568),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_548),
.B(n_429),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_551),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_553),
.B(n_399),
.Y(n_742)
);

CKINVDCx20_ASAP7_75t_R g743 ( 
.A(n_569),
.Y(n_743)
);

HB1xp67_ASAP7_75t_L g744 ( 
.A(n_616),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_602),
.Y(n_745)
);

OAI21x1_ASAP7_75t_L g746 ( 
.A1(n_596),
.A2(n_437),
.B(n_429),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_548),
.B(n_437),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_608),
.B(n_420),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_602),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_551),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_550),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_551),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_551),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_R g754 ( 
.A(n_600),
.B(n_319),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_551),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_551),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_550),
.Y(n_757)
);

BUFx6f_ASAP7_75t_L g758 ( 
.A(n_568),
.Y(n_758)
);

CKINVDCx16_ASAP7_75t_R g759 ( 
.A(n_600),
.Y(n_759)
);

AND2x6_ASAP7_75t_L g760 ( 
.A(n_674),
.B(n_466),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_627),
.Y(n_761)
);

INVx5_ASAP7_75t_L g762 ( 
.A(n_732),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_627),
.Y(n_763)
);

INVx1_ASAP7_75t_SL g764 ( 
.A(n_720),
.Y(n_764)
);

INVx5_ASAP7_75t_L g765 ( 
.A(n_732),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_645),
.Y(n_766)
);

INVx3_ASAP7_75t_L g767 ( 
.A(n_645),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_629),
.Y(n_768)
);

BUFx6f_ASAP7_75t_L g769 ( 
.A(n_677),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_633),
.B(n_742),
.Y(n_770)
);

AND2x4_ASAP7_75t_L g771 ( 
.A(n_655),
.B(n_451),
.Y(n_771)
);

INVx2_ASAP7_75t_SL g772 ( 
.A(n_729),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_629),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_727),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_683),
.Y(n_775)
);

AND2x4_ASAP7_75t_L g776 ( 
.A(n_643),
.B(n_404),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_727),
.Y(n_777)
);

INVx1_ASAP7_75t_SL g778 ( 
.A(n_744),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_693),
.B(n_365),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_683),
.Y(n_780)
);

INVx3_ASAP7_75t_L g781 ( 
.A(n_677),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_677),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_679),
.Y(n_783)
);

BUFx3_ASAP7_75t_L g784 ( 
.A(n_648),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_690),
.Y(n_785)
);

AND2x2_ASAP7_75t_L g786 ( 
.A(n_640),
.B(n_407),
.Y(n_786)
);

AND2x6_ASAP7_75t_L g787 ( 
.A(n_643),
.B(n_318),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_679),
.Y(n_788)
);

AND2x2_ASAP7_75t_L g789 ( 
.A(n_641),
.B(n_410),
.Y(n_789)
);

AND2x2_ASAP7_75t_SL g790 ( 
.A(n_759),
.B(n_346),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_664),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_679),
.Y(n_792)
);

INVx4_ASAP7_75t_L g793 ( 
.A(n_676),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_L g794 ( 
.A(n_637),
.B(n_381),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_628),
.B(n_425),
.Y(n_795)
);

BUFx6f_ASAP7_75t_L g796 ( 
.A(n_681),
.Y(n_796)
);

BUFx6f_ASAP7_75t_L g797 ( 
.A(n_681),
.Y(n_797)
);

HB1xp67_ASAP7_75t_L g798 ( 
.A(n_646),
.Y(n_798)
);

OAI22xp33_ASAP7_75t_L g799 ( 
.A1(n_715),
.A2(n_427),
.B1(n_432),
.B2(n_426),
.Y(n_799)
);

INVx4_ASAP7_75t_SL g800 ( 
.A(n_717),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_659),
.B(n_326),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_718),
.B(n_444),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_680),
.B(n_330),
.Y(n_803)
);

INVx5_ASAP7_75t_L g804 ( 
.A(n_681),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_662),
.B(n_663),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_631),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_L g807 ( 
.A(n_719),
.B(n_508),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_666),
.Y(n_808)
);

BUFx2_ASAP7_75t_L g809 ( 
.A(n_661),
.Y(n_809)
);

AOI22xp5_ASAP7_75t_L g810 ( 
.A1(n_724),
.A2(n_544),
.B1(n_442),
.B2(n_457),
.Y(n_810)
);

INVx2_ASAP7_75t_SL g811 ( 
.A(n_726),
.Y(n_811)
);

INVx1_ASAP7_75t_SL g812 ( 
.A(n_691),
.Y(n_812)
);

AND2x2_ASAP7_75t_L g813 ( 
.A(n_730),
.B(n_436),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_668),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_669),
.B(n_337),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_673),
.Y(n_816)
);

INVx1_ASAP7_75t_SL g817 ( 
.A(n_754),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_675),
.B(n_338),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_728),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_731),
.B(n_339),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_733),
.Y(n_821)
);

INVx3_ASAP7_75t_L g822 ( 
.A(n_694),
.Y(n_822)
);

BUFx3_ASAP7_75t_L g823 ( 
.A(n_671),
.Y(n_823)
);

AOI22xp33_ASAP7_75t_L g824 ( 
.A1(n_736),
.A2(n_328),
.B1(n_332),
.B2(n_321),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_685),
.B(n_341),
.Y(n_825)
);

AND2x6_ASAP7_75t_L g826 ( 
.A(n_738),
.B(n_334),
.Y(n_826)
);

INVx4_ASAP7_75t_SL g827 ( 
.A(n_741),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_750),
.B(n_343),
.Y(n_828)
);

BUFx3_ASAP7_75t_L g829 ( 
.A(n_734),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_686),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_745),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_752),
.B(n_458),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_689),
.B(n_345),
.Y(n_833)
);

AOI22xp33_ASAP7_75t_L g834 ( 
.A1(n_753),
.A2(n_335),
.B1(n_342),
.B2(n_336),
.Y(n_834)
);

OR2x2_ASAP7_75t_L g835 ( 
.A(n_710),
.B(n_460),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_672),
.Y(n_836)
);

OR2x2_ASAP7_75t_L g837 ( 
.A(n_703),
.B(n_467),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_749),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_624),
.Y(n_839)
);

INVx4_ASAP7_75t_L g840 ( 
.A(n_657),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_755),
.B(n_347),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_636),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_636),
.Y(n_843)
);

BUFx2_ASAP7_75t_L g844 ( 
.A(n_684),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_636),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_638),
.Y(n_846)
);

AND2x2_ASAP7_75t_SL g847 ( 
.A(n_702),
.B(n_351),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_639),
.Y(n_848)
);

INVx3_ASAP7_75t_L g849 ( 
.A(n_746),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_756),
.B(n_703),
.Y(n_850)
);

OR2x2_ASAP7_75t_L g851 ( 
.A(n_707),
.B(n_472),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_638),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_SL g853 ( 
.A(n_687),
.B(n_348),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_737),
.Y(n_854)
);

NAND3xp33_ASAP7_75t_L g855 ( 
.A(n_723),
.B(n_647),
.C(n_642),
.Y(n_855)
);

AND2x6_ASAP7_75t_L g856 ( 
.A(n_737),
.B(n_352),
.Y(n_856)
);

BUFx3_ASAP7_75t_L g857 ( 
.A(n_644),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_639),
.Y(n_858)
);

INVx5_ASAP7_75t_L g859 ( 
.A(n_639),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_740),
.Y(n_860)
);

BUFx6f_ASAP7_75t_L g861 ( 
.A(n_656),
.Y(n_861)
);

INVx3_ASAP7_75t_L g862 ( 
.A(n_657),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_740),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_630),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_660),
.B(n_350),
.Y(n_865)
);

NAND2x1p5_ASAP7_75t_L g866 ( 
.A(n_699),
.B(n_355),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_747),
.Y(n_867)
);

OAI21xp33_ASAP7_75t_L g868 ( 
.A1(n_660),
.A2(n_626),
.B(n_747),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_L g869 ( 
.A(n_748),
.B(n_353),
.Y(n_869)
);

CKINVDCx20_ASAP7_75t_R g870 ( 
.A(n_632),
.Y(n_870)
);

INVx3_ASAP7_75t_L g871 ( 
.A(n_623),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_635),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_626),
.B(n_354),
.Y(n_873)
);

AND2x6_ASAP7_75t_L g874 ( 
.A(n_709),
.B(n_357),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_651),
.Y(n_875)
);

AND2x4_ASAP7_75t_L g876 ( 
.A(n_699),
.B(n_473),
.Y(n_876)
);

BUFx8_ASAP7_75t_SL g877 ( 
.A(n_721),
.Y(n_877)
);

OR2x2_ASAP7_75t_L g878 ( 
.A(n_705),
.B(n_479),
.Y(n_878)
);

AOI22xp5_ASAP7_75t_L g879 ( 
.A1(n_649),
.A2(n_485),
.B1(n_489),
.B2(n_482),
.Y(n_879)
);

AOI22xp33_ASAP7_75t_L g880 ( 
.A1(n_652),
.A2(n_363),
.B1(n_371),
.B2(n_358),
.Y(n_880)
);

BUFx4f_ASAP7_75t_L g881 ( 
.A(n_701),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_653),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_L g883 ( 
.A(n_667),
.B(n_359),
.Y(n_883)
);

INVx4_ASAP7_75t_L g884 ( 
.A(n_758),
.Y(n_884)
);

INVx4_ASAP7_75t_SL g885 ( 
.A(n_634),
.Y(n_885)
);

BUFx2_ASAP7_75t_L g886 ( 
.A(n_650),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_623),
.Y(n_887)
);

AO22x2_ASAP7_75t_L g888 ( 
.A1(n_711),
.A2(n_375),
.B1(n_376),
.B2(n_374),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_625),
.Y(n_889)
);

INVx3_ASAP7_75t_L g890 ( 
.A(n_625),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_625),
.B(n_360),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_712),
.Y(n_892)
);

AND2x2_ASAP7_75t_L g893 ( 
.A(n_654),
.B(n_490),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_712),
.B(n_361),
.Y(n_894)
);

INVx3_ASAP7_75t_L g895 ( 
.A(n_658),
.Y(n_895)
);

XOR2xp5_ASAP7_75t_L g896 ( 
.A(n_735),
.B(n_504),
.Y(n_896)
);

BUFx6f_ASAP7_75t_L g897 ( 
.A(n_714),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_714),
.Y(n_898)
);

INVx4_ASAP7_75t_L g899 ( 
.A(n_714),
.Y(n_899)
);

INVx3_ASAP7_75t_L g900 ( 
.A(n_665),
.Y(n_900)
);

INVx4_ASAP7_75t_L g901 ( 
.A(n_758),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_739),
.B(n_362),
.Y(n_902)
);

INVx3_ASAP7_75t_L g903 ( 
.A(n_739),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_739),
.Y(n_904)
);

INVx5_ASAP7_75t_L g905 ( 
.A(n_758),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_706),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_743),
.Y(n_907)
);

NAND2x1p5_ASAP7_75t_L g908 ( 
.A(n_670),
.B(n_384),
.Y(n_908)
);

INVx3_ASAP7_75t_L g909 ( 
.A(n_682),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_692),
.Y(n_910)
);

INVx1_ASAP7_75t_SL g911 ( 
.A(n_695),
.Y(n_911)
);

AND2x4_ASAP7_75t_L g912 ( 
.A(n_696),
.B(n_506),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_716),
.Y(n_913)
);

INVx3_ASAP7_75t_L g914 ( 
.A(n_722),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_725),
.B(n_366),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_751),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_757),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_698),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_L g919 ( 
.A(n_700),
.B(n_368),
.Y(n_919)
);

INVx3_ASAP7_75t_L g920 ( 
.A(n_704),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_L g921 ( 
.A(n_678),
.B(n_372),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_688),
.B(n_373),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_L g923 ( 
.A(n_633),
.B(n_383),
.Y(n_923)
);

BUFx6f_ASAP7_75t_L g924 ( 
.A(n_677),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_SL g925 ( 
.A(n_676),
.B(n_386),
.Y(n_925)
);

BUFx6f_ASAP7_75t_L g926 ( 
.A(n_677),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_SL g927 ( 
.A(n_676),
.B(n_388),
.Y(n_927)
);

OR2x2_ASAP7_75t_L g928 ( 
.A(n_713),
.B(n_513),
.Y(n_928)
);

INVx6_ASAP7_75t_L g929 ( 
.A(n_627),
.Y(n_929)
);

INVx4_ASAP7_75t_L g930 ( 
.A(n_732),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_L g931 ( 
.A(n_633),
.B(n_394),
.Y(n_931)
);

BUFx3_ASAP7_75t_L g932 ( 
.A(n_648),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_629),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_629),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_SL g935 ( 
.A(n_676),
.B(n_398),
.Y(n_935)
);

AND2x4_ASAP7_75t_L g936 ( 
.A(n_674),
.B(n_516),
.Y(n_936)
);

BUFx3_ASAP7_75t_L g937 ( 
.A(n_648),
.Y(n_937)
);

AND2x2_ASAP7_75t_L g938 ( 
.A(n_713),
.B(n_523),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_627),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_627),
.Y(n_940)
);

NAND2xp33_ASAP7_75t_SL g941 ( 
.A(n_661),
.B(n_531),
.Y(n_941)
);

BUFx6f_ASAP7_75t_L g942 ( 
.A(n_677),
.Y(n_942)
);

OR2x2_ASAP7_75t_L g943 ( 
.A(n_713),
.B(n_532),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_629),
.Y(n_944)
);

NAND2xp33_ASAP7_75t_L g945 ( 
.A(n_697),
.B(n_380),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_SL g946 ( 
.A(n_676),
.B(n_400),
.Y(n_946)
);

BUFx10_ASAP7_75t_L g947 ( 
.A(n_667),
.Y(n_947)
);

AND2x6_ASAP7_75t_L g948 ( 
.A(n_674),
.B(n_391),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_SL g949 ( 
.A(n_676),
.B(n_402),
.Y(n_949)
);

INVx1_ASAP7_75t_SL g950 ( 
.A(n_713),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_676),
.B(n_403),
.Y(n_951)
);

INVx2_ASAP7_75t_SL g952 ( 
.A(n_713),
.Y(n_952)
);

OR2x2_ASAP7_75t_L g953 ( 
.A(n_713),
.B(n_533),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_SL g954 ( 
.A(n_676),
.B(n_411),
.Y(n_954)
);

OR2x6_ASAP7_75t_L g955 ( 
.A(n_708),
.B(n_392),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_676),
.B(n_412),
.Y(n_956)
);

INVx4_ASAP7_75t_SL g957 ( 
.A(n_732),
.Y(n_957)
);

INVx4_ASAP7_75t_L g958 ( 
.A(n_732),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_676),
.B(n_417),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_627),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_SL g961 ( 
.A(n_676),
.B(n_418),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_846),
.B(n_419),
.Y(n_962)
);

AND2x2_ASAP7_75t_L g963 ( 
.A(n_764),
.B(n_0),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_852),
.B(n_422),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_854),
.B(n_423),
.Y(n_965)
);

INVx3_ASAP7_75t_L g966 ( 
.A(n_840),
.Y(n_966)
);

AND2x6_ASAP7_75t_SL g967 ( 
.A(n_921),
.B(n_393),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_860),
.B(n_439),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_863),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_769),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_867),
.B(n_868),
.Y(n_971)
);

INVxp67_ASAP7_75t_SL g972 ( 
.A(n_784),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_769),
.Y(n_973)
);

AOI22xp33_ASAP7_75t_L g974 ( 
.A1(n_787),
.A2(n_401),
.B1(n_428),
.B2(n_421),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_770),
.B(n_443),
.Y(n_975)
);

AOI22xp33_ASAP7_75t_L g976 ( 
.A1(n_787),
.A2(n_431),
.B1(n_434),
.B2(n_433),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_766),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_L g978 ( 
.A(n_772),
.B(n_445),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_793),
.B(n_446),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_793),
.B(n_448),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_775),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_780),
.Y(n_982)
);

INVxp67_ASAP7_75t_L g983 ( 
.A(n_778),
.Y(n_983)
);

AND2x6_ASAP7_75t_L g984 ( 
.A(n_808),
.B(n_450),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_769),
.Y(n_985)
);

BUFx3_ASAP7_75t_L g986 ( 
.A(n_823),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_787),
.B(n_449),
.Y(n_987)
);

HB1xp67_ASAP7_75t_L g988 ( 
.A(n_950),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_796),
.Y(n_989)
);

AOI22xp33_ASAP7_75t_L g990 ( 
.A1(n_787),
.A2(n_455),
.B1(n_481),
.B2(n_468),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_826),
.B(n_453),
.Y(n_991)
);

AOI22xp5_ASAP7_75t_L g992 ( 
.A1(n_952),
.A2(n_507),
.B1(n_509),
.B2(n_486),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_877),
.Y(n_993)
);

A2O1A1Ixp33_ASAP7_75t_SL g994 ( 
.A1(n_794),
.A2(n_497),
.B(n_522),
.C(n_517),
.Y(n_994)
);

INVx2_ASAP7_75t_SL g995 ( 
.A(n_932),
.Y(n_995)
);

NOR2xp33_ASAP7_75t_L g996 ( 
.A(n_837),
.B(n_454),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_SL g997 ( 
.A(n_811),
.B(n_543),
.Y(n_997)
);

O2A1O1Ixp5_ASAP7_75t_L g998 ( 
.A1(n_803),
.A2(n_497),
.B(n_537),
.C(n_380),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_826),
.B(n_459),
.Y(n_999)
);

OR2x2_ASAP7_75t_L g1000 ( 
.A(n_937),
.B(n_1),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_826),
.B(n_469),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_796),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_876),
.B(n_470),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_767),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_876),
.B(n_542),
.Y(n_1005)
);

NAND2xp33_ASAP7_75t_L g1006 ( 
.A(n_826),
.B(n_380),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_805),
.B(n_814),
.Y(n_1007)
);

O2A1O1Ixp33_ASAP7_75t_L g1008 ( 
.A1(n_850),
.A2(n_8),
.B(n_1),
.C(n_2),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_816),
.B(n_830),
.Y(n_1009)
);

A2O1A1Ixp33_ASAP7_75t_L g1010 ( 
.A1(n_875),
.A2(n_349),
.B(n_529),
.C(n_325),
.Y(n_1010)
);

A2O1A1Ixp33_ASAP7_75t_L g1011 ( 
.A1(n_855),
.A2(n_349),
.B(n_529),
.C(n_325),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_SL g1012 ( 
.A(n_844),
.B(n_471),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_796),
.Y(n_1013)
);

AOI22xp33_ASAP7_75t_L g1014 ( 
.A1(n_856),
.A2(n_380),
.B1(n_478),
.B2(n_476),
.Y(n_1014)
);

NOR2xp33_ASAP7_75t_L g1015 ( 
.A(n_936),
.B(n_480),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_856),
.B(n_487),
.Y(n_1016)
);

AOI22xp33_ASAP7_75t_L g1017 ( 
.A1(n_856),
.A2(n_495),
.B1(n_498),
.B2(n_492),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_L g1018 ( 
.A(n_936),
.B(n_500),
.Y(n_1018)
);

AOI22xp33_ASAP7_75t_L g1019 ( 
.A1(n_856),
.A2(n_503),
.B1(n_511),
.B2(n_502),
.Y(n_1019)
);

BUFx6f_ASAP7_75t_L g1020 ( 
.A(n_797),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_SL g1021 ( 
.A(n_947),
.B(n_865),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_SL g1022 ( 
.A(n_947),
.B(n_540),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_785),
.B(n_512),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_761),
.Y(n_1024)
);

AOI22xp5_ASAP7_75t_L g1025 ( 
.A1(n_776),
.A2(n_771),
.B1(n_789),
.B2(n_786),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_798),
.B(n_538),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_763),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_939),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_779),
.B(n_518),
.Y(n_1029)
);

OAI22xp5_ASAP7_75t_L g1030 ( 
.A1(n_847),
.A2(n_525),
.B1(n_527),
.B2(n_524),
.Y(n_1030)
);

NOR2xp33_ASAP7_75t_L g1031 ( 
.A(n_776),
.B(n_534),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_SL g1032 ( 
.A(n_771),
.B(n_840),
.Y(n_1032)
);

NOR2xp33_ASAP7_75t_SL g1033 ( 
.A(n_911),
.B(n_535),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_948),
.B(n_8),
.Y(n_1034)
);

AOI22xp33_ASAP7_75t_L g1035 ( 
.A1(n_888),
.A2(n_349),
.B1(n_529),
.B2(n_325),
.Y(n_1035)
);

INVx2_ASAP7_75t_SL g1036 ( 
.A(n_881),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_873),
.B(n_9),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_791),
.B(n_795),
.Y(n_1038)
);

INVx3_ASAP7_75t_L g1039 ( 
.A(n_862),
.Y(n_1039)
);

AOI22xp33_ASAP7_75t_L g1040 ( 
.A1(n_888),
.A2(n_529),
.B1(n_12),
.B2(n_10),
.Y(n_1040)
);

NAND3xp33_ASAP7_75t_L g1041 ( 
.A(n_880),
.B(n_834),
.C(n_824),
.Y(n_1041)
);

INVx3_ASAP7_75t_L g1042 ( 
.A(n_862),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_813),
.B(n_11),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_836),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_832),
.B(n_11),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_760),
.B(n_13),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_849),
.A2(n_106),
.B(n_105),
.Y(n_1047)
);

AND2x6_ASAP7_75t_SL g1048 ( 
.A(n_955),
.B(n_13),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_760),
.B(n_14),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_797),
.Y(n_1050)
);

NOR2xp33_ASAP7_75t_L g1051 ( 
.A(n_928),
.B(n_943),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_760),
.B(n_17),
.Y(n_1052)
);

OR2x6_ASAP7_75t_L g1053 ( 
.A(n_886),
.B(n_18),
.Y(n_1053)
);

INVxp67_ASAP7_75t_L g1054 ( 
.A(n_938),
.Y(n_1054)
);

INVx3_ASAP7_75t_L g1055 ( 
.A(n_884),
.Y(n_1055)
);

INVx2_ASAP7_75t_SL g1056 ( 
.A(n_955),
.Y(n_1056)
);

AND2x6_ASAP7_75t_L g1057 ( 
.A(n_909),
.B(n_109),
.Y(n_1057)
);

AOI22xp5_ASAP7_75t_L g1058 ( 
.A1(n_874),
.A2(n_20),
.B1(n_18),
.B2(n_19),
.Y(n_1058)
);

AND2x2_ASAP7_75t_SL g1059 ( 
.A(n_790),
.B(n_20),
.Y(n_1059)
);

AOI22xp33_ASAP7_75t_L g1060 ( 
.A1(n_874),
.A2(n_25),
.B1(n_21),
.B2(n_24),
.Y(n_1060)
);

OR2x2_ASAP7_75t_L g1061 ( 
.A(n_953),
.B(n_24),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_923),
.B(n_26),
.Y(n_1062)
);

O2A1O1Ixp33_ASAP7_75t_L g1063 ( 
.A1(n_906),
.A2(n_28),
.B(n_26),
.C(n_27),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_SL g1064 ( 
.A(n_951),
.B(n_27),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_940),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_931),
.B(n_28),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_797),
.Y(n_1067)
);

INVx1_ASAP7_75t_SL g1068 ( 
.A(n_896),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_924),
.Y(n_1069)
);

AOI22xp33_ASAP7_75t_L g1070 ( 
.A1(n_874),
.A2(n_33),
.B1(n_29),
.B2(n_32),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_960),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_924),
.Y(n_1072)
);

OAI22xp5_ASAP7_75t_SL g1073 ( 
.A1(n_870),
.A2(n_33),
.B1(n_29),
.B2(n_32),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_929),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_929),
.Y(n_1075)
);

AOI22xp33_ASAP7_75t_L g1076 ( 
.A1(n_874),
.A2(n_36),
.B1(n_34),
.B2(n_35),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_L g1077 ( 
.A(n_835),
.B(n_922),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_882),
.Y(n_1078)
);

BUFx3_ASAP7_75t_L g1079 ( 
.A(n_857),
.Y(n_1079)
);

NOR2xp33_ASAP7_75t_L g1080 ( 
.A(n_851),
.B(n_35),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_L g1081 ( 
.A(n_878),
.B(n_39),
.Y(n_1081)
);

NOR3xp33_ASAP7_75t_SL g1082 ( 
.A(n_839),
.B(n_39),
.C(n_40),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_802),
.B(n_807),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_801),
.B(n_41),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_SL g1085 ( 
.A(n_956),
.B(n_42),
.Y(n_1085)
);

AOI22xp5_ASAP7_75t_SL g1086 ( 
.A1(n_896),
.A2(n_45),
.B1(n_42),
.B2(n_44),
.Y(n_1086)
);

OR2x6_ASAP7_75t_L g1087 ( 
.A(n_809),
.B(n_44),
.Y(n_1087)
);

NOR2xp33_ASAP7_75t_SL g1088 ( 
.A(n_812),
.B(n_46),
.Y(n_1088)
);

NOR2xp33_ASAP7_75t_L g1089 ( 
.A(n_918),
.B(n_47),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_815),
.B(n_47),
.Y(n_1090)
);

AOI22xp33_ASAP7_75t_L g1091 ( 
.A1(n_829),
.A2(n_50),
.B1(n_48),
.B2(n_49),
.Y(n_1091)
);

NOR2xp33_ASAP7_75t_L g1092 ( 
.A(n_820),
.B(n_828),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_833),
.B(n_49),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_768),
.Y(n_1094)
);

NOR2x1p5_ASAP7_75t_L g1095 ( 
.A(n_895),
.B(n_900),
.Y(n_1095)
);

NAND2x1p5_ASAP7_75t_L g1096 ( 
.A(n_817),
.B(n_50),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_864),
.Y(n_1097)
);

NOR2x2_ASAP7_75t_L g1098 ( 
.A(n_916),
.B(n_51),
.Y(n_1098)
);

A2O1A1Ixp33_ASAP7_75t_L g1099 ( 
.A1(n_841),
.A2(n_53),
.B(n_51),
.C(n_52),
.Y(n_1099)
);

O2A1O1Ixp5_ASAP7_75t_L g1100 ( 
.A1(n_961),
.A2(n_114),
.B(n_115),
.C(n_110),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_959),
.B(n_52),
.Y(n_1101)
);

BUFx12f_ASAP7_75t_L g1102 ( 
.A(n_872),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_810),
.B(n_53),
.Y(n_1103)
);

AND2x2_ASAP7_75t_L g1104 ( 
.A(n_893),
.B(n_56),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_SL g1105 ( 
.A(n_799),
.B(n_56),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_773),
.Y(n_1106)
);

NOR2xp33_ASAP7_75t_L g1107 ( 
.A(n_912),
.B(n_57),
.Y(n_1107)
);

HB1xp67_ASAP7_75t_L g1108 ( 
.A(n_907),
.Y(n_1108)
);

OAI221xp5_ASAP7_75t_L g1109 ( 
.A1(n_879),
.A2(n_57),
.B1(n_58),
.B2(n_59),
.C(n_60),
.Y(n_1109)
);

NAND2x1p5_ASAP7_75t_L g1110 ( 
.A(n_804),
.B(n_58),
.Y(n_1110)
);

AND2x2_ASAP7_75t_SL g1111 ( 
.A(n_912),
.B(n_59),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_774),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_883),
.B(n_62),
.Y(n_1113)
);

O2A1O1Ixp5_ASAP7_75t_L g1114 ( 
.A1(n_925),
.A2(n_927),
.B(n_946),
.C(n_935),
.Y(n_1114)
);

AND2x4_ASAP7_75t_L g1115 ( 
.A(n_800),
.B(n_62),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_822),
.B(n_63),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_949),
.B(n_64),
.Y(n_1117)
);

AOI22xp33_ASAP7_75t_L g1118 ( 
.A1(n_806),
.A2(n_67),
.B1(n_65),
.B2(n_66),
.Y(n_1118)
);

AOI22xp33_ASAP7_75t_L g1119 ( 
.A1(n_819),
.A2(n_821),
.B1(n_838),
.B2(n_831),
.Y(n_1119)
);

AO22x1_ASAP7_75t_L g1120 ( 
.A1(n_909),
.A2(n_68),
.B1(n_66),
.B2(n_67),
.Y(n_1120)
);

HB1xp67_ASAP7_75t_L g1121 ( 
.A(n_914),
.Y(n_1121)
);

INVx3_ASAP7_75t_L g1122 ( 
.A(n_884),
.Y(n_1122)
);

NAND2x1p5_ASAP7_75t_L g1123 ( 
.A(n_804),
.B(n_68),
.Y(n_1123)
);

OAI221xp5_ASAP7_75t_L g1124 ( 
.A1(n_908),
.A2(n_70),
.B1(n_71),
.B2(n_72),
.C(n_73),
.Y(n_1124)
);

AOI22xp5_ASAP7_75t_L g1125 ( 
.A1(n_941),
.A2(n_76),
.B1(n_72),
.B2(n_75),
.Y(n_1125)
);

OAI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_910),
.A2(n_77),
.B1(n_75),
.B2(n_76),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_926),
.Y(n_1127)
);

AOI22xp5_ASAP7_75t_L g1128 ( 
.A1(n_913),
.A2(n_81),
.B1(n_79),
.B2(n_80),
.Y(n_1128)
);

NOR2xp33_ASAP7_75t_SL g1129 ( 
.A(n_914),
.B(n_79),
.Y(n_1129)
);

HB1xp67_ASAP7_75t_L g1130 ( 
.A(n_800),
.Y(n_1130)
);

OR2x6_ASAP7_75t_L g1131 ( 
.A(n_917),
.B(n_80),
.Y(n_1131)
);

HB1xp67_ASAP7_75t_L g1132 ( 
.A(n_988),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_969),
.Y(n_1133)
);

AO22x1_ASAP7_75t_L g1134 ( 
.A1(n_1115),
.A2(n_920),
.B1(n_919),
.B2(n_885),
.Y(n_1134)
);

INVx5_ASAP7_75t_L g1135 ( 
.A(n_1053),
.Y(n_1135)
);

XNOR2x2_ASAP7_75t_SL g1136 ( 
.A(n_1098),
.B(n_885),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_1024),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_1007),
.B(n_827),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_971),
.A2(n_945),
.B(n_853),
.Y(n_1139)
);

CKINVDCx16_ASAP7_75t_R g1140 ( 
.A(n_1102),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1038),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_1027),
.Y(n_1142)
);

INVxp67_ASAP7_75t_L g1143 ( 
.A(n_983),
.Y(n_1143)
);

INVx3_ASAP7_75t_L g1144 ( 
.A(n_986),
.Y(n_1144)
);

OR2x6_ASAP7_75t_L g1145 ( 
.A(n_1053),
.B(n_866),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_1051),
.B(n_827),
.Y(n_1146)
);

OR2x6_ASAP7_75t_L g1147 ( 
.A(n_1053),
.B(n_930),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1077),
.B(n_954),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1009),
.Y(n_1149)
);

INVx1_ASAP7_75t_SL g1150 ( 
.A(n_995),
.Y(n_1150)
);

OR2x6_ASAP7_75t_L g1151 ( 
.A(n_1131),
.B(n_958),
.Y(n_1151)
);

NOR2xp33_ASAP7_75t_L g1152 ( 
.A(n_1025),
.B(n_1054),
.Y(n_1152)
);

OAI22xp5_ASAP7_75t_L g1153 ( 
.A1(n_1083),
.A2(n_933),
.B1(n_934),
.B2(n_777),
.Y(n_1153)
);

BUFx2_ASAP7_75t_L g1154 ( 
.A(n_972),
.Y(n_1154)
);

NAND3xp33_ASAP7_75t_L g1155 ( 
.A(n_1092),
.B(n_915),
.C(n_869),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1041),
.B(n_1104),
.Y(n_1156)
);

BUFx3_ASAP7_75t_L g1157 ( 
.A(n_1079),
.Y(n_1157)
);

CKINVDCx20_ASAP7_75t_R g1158 ( 
.A(n_993),
.Y(n_1158)
);

AND2x2_ASAP7_75t_L g1159 ( 
.A(n_1111),
.B(n_930),
.Y(n_1159)
);

INVx5_ASAP7_75t_L g1160 ( 
.A(n_1057),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1078),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_1028),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_984),
.B(n_818),
.Y(n_1163)
);

INVxp67_ASAP7_75t_L g1164 ( 
.A(n_1033),
.Y(n_1164)
);

NOR2xp33_ASAP7_75t_R g1165 ( 
.A(n_1044),
.B(n_762),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_1097),
.Y(n_1166)
);

NOR3xp33_ASAP7_75t_SL g1167 ( 
.A(n_1073),
.B(n_1124),
.C(n_1022),
.Y(n_1167)
);

BUFx6f_ASAP7_75t_L g1168 ( 
.A(n_1020),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1065),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1071),
.Y(n_1170)
);

AND2x4_ASAP7_75t_L g1171 ( 
.A(n_1095),
.B(n_957),
.Y(n_1171)
);

OR2x6_ASAP7_75t_L g1172 ( 
.A(n_1131),
.B(n_958),
.Y(n_1172)
);

INVx1_ASAP7_75t_SL g1173 ( 
.A(n_1000),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_984),
.B(n_825),
.Y(n_1174)
);

INVx3_ASAP7_75t_L g1175 ( 
.A(n_1056),
.Y(n_1175)
);

NOR3xp33_ASAP7_75t_SL g1176 ( 
.A(n_1073),
.B(n_894),
.C(n_891),
.Y(n_1176)
);

BUFx8_ASAP7_75t_L g1177 ( 
.A(n_1115),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_977),
.Y(n_1178)
);

CKINVDCx20_ASAP7_75t_R g1179 ( 
.A(n_1108),
.Y(n_1179)
);

INVxp67_ASAP7_75t_SL g1180 ( 
.A(n_1020),
.Y(n_1180)
);

AND2x4_ASAP7_75t_L g1181 ( 
.A(n_1036),
.B(n_1021),
.Y(n_1181)
);

NOR2xp33_ASAP7_75t_L g1182 ( 
.A(n_1032),
.B(n_762),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_981),
.Y(n_1183)
);

NOR3xp33_ASAP7_75t_SL g1184 ( 
.A(n_1107),
.B(n_902),
.C(n_889),
.Y(n_1184)
);

BUFx2_ASAP7_75t_L g1185 ( 
.A(n_984),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_982),
.Y(n_1186)
);

BUFx6f_ASAP7_75t_L g1187 ( 
.A(n_966),
.Y(n_1187)
);

BUFx10_ASAP7_75t_L g1188 ( 
.A(n_1048),
.Y(n_1188)
);

OR2x2_ASAP7_75t_L g1189 ( 
.A(n_1068),
.B(n_944),
.Y(n_1189)
);

INVx1_ASAP7_75t_SL g1190 ( 
.A(n_963),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_1094),
.Y(n_1191)
);

BUFx3_ASAP7_75t_L g1192 ( 
.A(n_1121),
.Y(n_1192)
);

BUFx4f_ASAP7_75t_L g1193 ( 
.A(n_1087),
.Y(n_1193)
);

INVx4_ASAP7_75t_L g1194 ( 
.A(n_1087),
.Y(n_1194)
);

NOR3xp33_ASAP7_75t_SL g1195 ( 
.A(n_1003),
.B(n_892),
.C(n_887),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_1106),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_1112),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1004),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_R g1199 ( 
.A(n_1059),
.B(n_1048),
.Y(n_1199)
);

BUFx3_ASAP7_75t_L g1200 ( 
.A(n_1087),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_SL g1201 ( 
.A(n_1129),
.B(n_765),
.Y(n_1201)
);

AND2x2_ASAP7_75t_L g1202 ( 
.A(n_1061),
.B(n_899),
.Y(n_1202)
);

INVx4_ASAP7_75t_L g1203 ( 
.A(n_1057),
.Y(n_1203)
);

INVx2_ASAP7_75t_SL g1204 ( 
.A(n_1130),
.Y(n_1204)
);

BUFx3_ASAP7_75t_L g1205 ( 
.A(n_1110),
.Y(n_1205)
);

A2O1A1Ixp33_ASAP7_75t_L g1206 ( 
.A1(n_1080),
.A2(n_1081),
.B(n_1063),
.C(n_1089),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_1123),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1043),
.Y(n_1208)
);

BUFx3_ASAP7_75t_L g1209 ( 
.A(n_1123),
.Y(n_1209)
);

BUFx3_ASAP7_75t_L g1210 ( 
.A(n_1074),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1045),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_984),
.B(n_859),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_975),
.B(n_859),
.Y(n_1213)
);

CKINVDCx20_ASAP7_75t_R g1214 ( 
.A(n_1086),
.Y(n_1214)
);

NOR3xp33_ASAP7_75t_SL g1215 ( 
.A(n_1005),
.B(n_904),
.C(n_82),
.Y(n_1215)
);

OR2x6_ASAP7_75t_L g1216 ( 
.A(n_1120),
.B(n_899),
.Y(n_1216)
);

INVx4_ASAP7_75t_L g1217 ( 
.A(n_1057),
.Y(n_1217)
);

OR2x2_ASAP7_75t_L g1218 ( 
.A(n_1030),
.B(n_901),
.Y(n_1218)
);

BUFx6f_ASAP7_75t_L g1219 ( 
.A(n_966),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_996),
.B(n_905),
.Y(n_1220)
);

NAND2xp33_ASAP7_75t_SL g1221 ( 
.A(n_1034),
.B(n_901),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_992),
.B(n_905),
.Y(n_1222)
);

INVx3_ASAP7_75t_L g1223 ( 
.A(n_1075),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1116),
.Y(n_1224)
);

BUFx6f_ASAP7_75t_L g1225 ( 
.A(n_1057),
.Y(n_1225)
);

NOR3xp33_ASAP7_75t_SL g1226 ( 
.A(n_1031),
.B(n_83),
.C(n_85),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1117),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1103),
.B(n_905),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1128),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1084),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_962),
.B(n_781),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_SL g1232 ( 
.A(n_978),
.B(n_926),
.Y(n_1232)
);

NOR2xp33_ASAP7_75t_L g1233 ( 
.A(n_1015),
.B(n_781),
.Y(n_1233)
);

AND2x6_ASAP7_75t_L g1234 ( 
.A(n_1058),
.B(n_942),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_SL g1235 ( 
.A(n_991),
.B(n_942),
.Y(n_1235)
);

AND2x4_ASAP7_75t_L g1236 ( 
.A(n_1039),
.B(n_782),
.Y(n_1236)
);

INVx5_ASAP7_75t_L g1237 ( 
.A(n_1055),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_1055),
.Y(n_1238)
);

INVx2_ASAP7_75t_SL g1239 ( 
.A(n_1096),
.Y(n_1239)
);

NOR2xp33_ASAP7_75t_R g1240 ( 
.A(n_1006),
.B(n_83),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1090),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_1086),
.B(n_942),
.Y(n_1242)
);

AND2x2_ASAP7_75t_L g1243 ( 
.A(n_1018),
.B(n_85),
.Y(n_1243)
);

NOR3xp33_ASAP7_75t_SL g1244 ( 
.A(n_1126),
.B(n_86),
.C(n_87),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_964),
.B(n_783),
.Y(n_1245)
);

AND3x1_ASAP7_75t_SL g1246 ( 
.A(n_1109),
.B(n_87),
.C(n_88),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1093),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1037),
.Y(n_1248)
);

HB1xp67_ASAP7_75t_L g1249 ( 
.A(n_1122),
.Y(n_1249)
);

BUFx6f_ASAP7_75t_L g1250 ( 
.A(n_1122),
.Y(n_1250)
);

AOI221xp5_ASAP7_75t_L g1251 ( 
.A1(n_1105),
.A2(n_788),
.B1(n_792),
.B2(n_903),
.C(n_871),
.Y(n_1251)
);

AO22x1_ASAP7_75t_L g1252 ( 
.A1(n_1046),
.A2(n_90),
.B1(n_88),
.B2(n_89),
.Y(n_1252)
);

BUFx6f_ASAP7_75t_L g1253 ( 
.A(n_970),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_965),
.B(n_871),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_1133),
.Y(n_1255)
);

NOR2xp33_ASAP7_75t_L g1256 ( 
.A(n_1152),
.B(n_967),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1149),
.B(n_974),
.Y(n_1257)
);

A2O1A1Ixp33_ASAP7_75t_L g1258 ( 
.A1(n_1206),
.A2(n_1008),
.B(n_1066),
.C(n_1062),
.Y(n_1258)
);

AOI21xp33_ASAP7_75t_L g1259 ( 
.A1(n_1156),
.A2(n_994),
.B(n_1113),
.Y(n_1259)
);

OAI21x1_ASAP7_75t_L g1260 ( 
.A1(n_1207),
.A2(n_1047),
.B(n_1100),
.Y(n_1260)
);

OAI21x1_ASAP7_75t_L g1261 ( 
.A1(n_1235),
.A2(n_1127),
.B(n_985),
.Y(n_1261)
);

OAI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1148),
.A2(n_1114),
.B(n_968),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1141),
.B(n_1229),
.Y(n_1263)
);

BUFx6f_ASAP7_75t_L g1264 ( 
.A(n_1168),
.Y(n_1264)
);

OAI21x1_ASAP7_75t_L g1265 ( 
.A1(n_1139),
.A2(n_989),
.B(n_973),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1161),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1169),
.Y(n_1267)
);

OA21x2_ASAP7_75t_L g1268 ( 
.A1(n_1248),
.A2(n_1011),
.B(n_1010),
.Y(n_1268)
);

AOI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1230),
.A2(n_1101),
.B(n_998),
.Y(n_1269)
);

OAI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1155),
.A2(n_990),
.B(n_976),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1154),
.B(n_1040),
.Y(n_1271)
);

AOI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1241),
.A2(n_1085),
.B(n_1064),
.Y(n_1272)
);

BUFx6f_ASAP7_75t_L g1273 ( 
.A(n_1168),
.Y(n_1273)
);

NOR2xp67_ASAP7_75t_L g1274 ( 
.A(n_1135),
.B(n_1026),
.Y(n_1274)
);

CKINVDCx16_ASAP7_75t_R g1275 ( 
.A(n_1140),
.Y(n_1275)
);

BUFx6f_ASAP7_75t_L g1276 ( 
.A(n_1168),
.Y(n_1276)
);

AOI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_1247),
.A2(n_1013),
.B(n_1002),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_1158),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1154),
.B(n_967),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1170),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1178),
.B(n_1023),
.Y(n_1281)
);

OAI21x1_ASAP7_75t_L g1282 ( 
.A1(n_1180),
.A2(n_1067),
.B(n_1050),
.Y(n_1282)
);

AND2x4_ASAP7_75t_L g1283 ( 
.A(n_1135),
.B(n_1203),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1183),
.B(n_1082),
.Y(n_1284)
);

INVxp67_ASAP7_75t_L g1285 ( 
.A(n_1132),
.Y(n_1285)
);

BUFx6f_ASAP7_75t_L g1286 ( 
.A(n_1225),
.Y(n_1286)
);

O2A1O1Ixp5_ASAP7_75t_L g1287 ( 
.A1(n_1201),
.A2(n_1052),
.B(n_1049),
.C(n_1099),
.Y(n_1287)
);

AND2x2_ASAP7_75t_L g1288 ( 
.A(n_1159),
.B(n_1012),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1186),
.B(n_1029),
.Y(n_1289)
);

A2O1A1Ixp33_ASAP7_75t_L g1290 ( 
.A1(n_1208),
.A2(n_1125),
.B(n_1035),
.C(n_1070),
.Y(n_1290)
);

OAI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1211),
.A2(n_1227),
.B(n_1224),
.Y(n_1291)
);

AOI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1245),
.A2(n_1072),
.B(n_1069),
.Y(n_1292)
);

BUFx3_ASAP7_75t_L g1293 ( 
.A(n_1157),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1137),
.B(n_997),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1142),
.Y(n_1295)
);

AO21x2_ASAP7_75t_L g1296 ( 
.A1(n_1228),
.A2(n_1016),
.B(n_1001),
.Y(n_1296)
);

BUFx2_ASAP7_75t_L g1297 ( 
.A(n_1179),
.Y(n_1297)
);

AO21x1_ASAP7_75t_L g1298 ( 
.A1(n_1217),
.A2(n_1088),
.B(n_999),
.Y(n_1298)
);

OAI21xp5_ASAP7_75t_L g1299 ( 
.A1(n_1153),
.A2(n_1014),
.B(n_1119),
.Y(n_1299)
);

OAI22xp5_ASAP7_75t_L g1300 ( 
.A1(n_1151),
.A2(n_1076),
.B1(n_1060),
.B2(n_1091),
.Y(n_1300)
);

AOI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1232),
.A2(n_1042),
.B(n_1039),
.Y(n_1301)
);

OAI22xp5_ASAP7_75t_L g1302 ( 
.A1(n_1151),
.A2(n_1118),
.B1(n_1017),
.B2(n_1019),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1162),
.B(n_979),
.Y(n_1303)
);

AOI22xp5_ASAP7_75t_L g1304 ( 
.A1(n_1214),
.A2(n_987),
.B1(n_980),
.B2(n_890),
.Y(n_1304)
);

BUFx2_ASAP7_75t_SL g1305 ( 
.A(n_1135),
.Y(n_1305)
);

OR2x2_ASAP7_75t_L g1306 ( 
.A(n_1143),
.B(n_91),
.Y(n_1306)
);

BUFx2_ASAP7_75t_L g1307 ( 
.A(n_1177),
.Y(n_1307)
);

NAND3xp33_ASAP7_75t_L g1308 ( 
.A(n_1226),
.B(n_897),
.C(n_861),
.Y(n_1308)
);

AO31x2_ASAP7_75t_L g1309 ( 
.A1(n_1185),
.A2(n_843),
.A3(n_845),
.B(n_842),
.Y(n_1309)
);

INVx1_ASAP7_75t_SL g1310 ( 
.A(n_1150),
.Y(n_1310)
);

OAI21x1_ASAP7_75t_L g1311 ( 
.A1(n_1212),
.A2(n_858),
.B(n_848),
.Y(n_1311)
);

OA22x2_ASAP7_75t_L g1312 ( 
.A1(n_1147),
.A2(n_95),
.B1(n_92),
.B2(n_93),
.Y(n_1312)
);

AOI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1254),
.A2(n_898),
.B(n_897),
.Y(n_1313)
);

AO21x2_ASAP7_75t_L g1314 ( 
.A1(n_1184),
.A2(n_897),
.B(n_861),
.Y(n_1314)
);

OAI21x1_ASAP7_75t_L g1315 ( 
.A1(n_1213),
.A2(n_118),
.B(n_116),
.Y(n_1315)
);

AOI21xp5_ASAP7_75t_L g1316 ( 
.A1(n_1231),
.A2(n_121),
.B(n_120),
.Y(n_1316)
);

OAI21x1_ASAP7_75t_SL g1317 ( 
.A1(n_1194),
.A2(n_93),
.B(n_97),
.Y(n_1317)
);

AOI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1138),
.A2(n_127),
.B(n_126),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1191),
.Y(n_1319)
);

OAI21x1_ASAP7_75t_L g1320 ( 
.A1(n_1220),
.A2(n_132),
.B(n_129),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1190),
.B(n_97),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1196),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1199),
.B(n_99),
.Y(n_1323)
);

OAI21xp33_ASAP7_75t_L g1324 ( 
.A1(n_1167),
.A2(n_99),
.B(n_100),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1197),
.Y(n_1325)
);

OAI22xp5_ASAP7_75t_L g1326 ( 
.A1(n_1172),
.A2(n_100),
.B1(n_101),
.B2(n_103),
.Y(n_1326)
);

NAND3xp33_ASAP7_75t_L g1327 ( 
.A(n_1244),
.B(n_101),
.C(n_103),
.Y(n_1327)
);

CKINVDCx14_ASAP7_75t_R g1328 ( 
.A(n_1307),
.Y(n_1328)
);

AO31x2_ASAP7_75t_L g1329 ( 
.A1(n_1258),
.A2(n_1185),
.A3(n_1198),
.B(n_1174),
.Y(n_1329)
);

OAI21x1_ASAP7_75t_L g1330 ( 
.A1(n_1260),
.A2(n_1242),
.B(n_1238),
.Y(n_1330)
);

OAI21x1_ASAP7_75t_L g1331 ( 
.A1(n_1311),
.A2(n_1163),
.B(n_1218),
.Y(n_1331)
);

AND2x4_ASAP7_75t_L g1332 ( 
.A(n_1283),
.B(n_1160),
.Y(n_1332)
);

CKINVDCx20_ASAP7_75t_R g1333 ( 
.A(n_1275),
.Y(n_1333)
);

OAI21x1_ASAP7_75t_L g1334 ( 
.A1(n_1265),
.A2(n_1251),
.B(n_1222),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1319),
.B(n_1176),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1266),
.Y(n_1336)
);

NOR2xp33_ASAP7_75t_L g1337 ( 
.A(n_1256),
.B(n_1145),
.Y(n_1337)
);

HB1xp67_ASAP7_75t_L g1338 ( 
.A(n_1285),
.Y(n_1338)
);

AND2x4_ASAP7_75t_L g1339 ( 
.A(n_1283),
.B(n_1160),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1266),
.Y(n_1340)
);

INVx4_ASAP7_75t_L g1341 ( 
.A(n_1286),
.Y(n_1341)
);

AND3x1_ASAP7_75t_L g1342 ( 
.A(n_1323),
.B(n_1136),
.C(n_1215),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1280),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_1280),
.Y(n_1344)
);

OAI21x1_ASAP7_75t_L g1345 ( 
.A1(n_1320),
.A2(n_1146),
.B(n_1202),
.Y(n_1345)
);

INVx2_ASAP7_75t_L g1346 ( 
.A(n_1255),
.Y(n_1346)
);

OAI21x1_ASAP7_75t_L g1347 ( 
.A1(n_1315),
.A2(n_1182),
.B(n_1223),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1263),
.B(n_1173),
.Y(n_1348)
);

INVx1_ASAP7_75t_SL g1349 ( 
.A(n_1310),
.Y(n_1349)
);

OR2x6_ASAP7_75t_L g1350 ( 
.A(n_1305),
.B(n_1172),
.Y(n_1350)
);

OR2x2_ASAP7_75t_L g1351 ( 
.A(n_1279),
.B(n_1147),
.Y(n_1351)
);

NOR2xp33_ASAP7_75t_L g1352 ( 
.A(n_1297),
.B(n_1145),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1295),
.B(n_1216),
.Y(n_1353)
);

OAI21x1_ASAP7_75t_L g1354 ( 
.A1(n_1282),
.A2(n_1243),
.B(n_1249),
.Y(n_1354)
);

OAI21x1_ASAP7_75t_L g1355 ( 
.A1(n_1261),
.A2(n_1233),
.B(n_1221),
.Y(n_1355)
);

OAI22xp5_ASAP7_75t_L g1356 ( 
.A1(n_1304),
.A2(n_1193),
.B1(n_1216),
.B2(n_1200),
.Y(n_1356)
);

NOR2xp33_ASAP7_75t_L g1357 ( 
.A(n_1288),
.B(n_1164),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_1264),
.Y(n_1358)
);

OAI21x1_ASAP7_75t_L g1359 ( 
.A1(n_1269),
.A2(n_1175),
.B(n_1144),
.Y(n_1359)
);

BUFx6f_ASAP7_75t_L g1360 ( 
.A(n_1264),
.Y(n_1360)
);

BUFx2_ASAP7_75t_SL g1361 ( 
.A(n_1293),
.Y(n_1361)
);

OA21x2_ASAP7_75t_L g1362 ( 
.A1(n_1259),
.A2(n_1195),
.B(n_1236),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1267),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_1264),
.Y(n_1364)
);

NAND2x1_ASAP7_75t_L g1365 ( 
.A(n_1344),
.B(n_1273),
.Y(n_1365)
);

INVx2_ASAP7_75t_SL g1366 ( 
.A(n_1350),
.Y(n_1366)
);

AOI22xp33_ASAP7_75t_L g1367 ( 
.A1(n_1335),
.A2(n_1327),
.B1(n_1324),
.B2(n_1300),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1335),
.B(n_1322),
.Y(n_1368)
);

AOI222xp33_ASAP7_75t_L g1369 ( 
.A1(n_1356),
.A2(n_1177),
.B1(n_1188),
.B2(n_1291),
.C1(n_1284),
.C2(n_1326),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1344),
.Y(n_1370)
);

INVx1_ASAP7_75t_SL g1371 ( 
.A(n_1361),
.Y(n_1371)
);

CKINVDCx6p67_ASAP7_75t_R g1372 ( 
.A(n_1333),
.Y(n_1372)
);

INVx4_ASAP7_75t_L g1373 ( 
.A(n_1332),
.Y(n_1373)
);

AOI22xp33_ASAP7_75t_L g1374 ( 
.A1(n_1357),
.A2(n_1312),
.B1(n_1302),
.B2(n_1234),
.Y(n_1374)
);

AOI21xp33_ASAP7_75t_L g1375 ( 
.A1(n_1362),
.A2(n_1298),
.B(n_1239),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1336),
.Y(n_1376)
);

INVx3_ASAP7_75t_L g1377 ( 
.A(n_1360),
.Y(n_1377)
);

BUFx2_ASAP7_75t_L g1378 ( 
.A(n_1360),
.Y(n_1378)
);

BUFx2_ASAP7_75t_L g1379 ( 
.A(n_1360),
.Y(n_1379)
);

INVx4_ASAP7_75t_L g1380 ( 
.A(n_1332),
.Y(n_1380)
);

BUFx12f_ASAP7_75t_L g1381 ( 
.A(n_1350),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1340),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1343),
.Y(n_1383)
);

BUFx12f_ASAP7_75t_L g1384 ( 
.A(n_1350),
.Y(n_1384)
);

INVx3_ASAP7_75t_L g1385 ( 
.A(n_1360),
.Y(n_1385)
);

OR2x6_ASAP7_75t_L g1386 ( 
.A(n_1350),
.B(n_1205),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1346),
.Y(n_1387)
);

AND2x4_ASAP7_75t_L g1388 ( 
.A(n_1330),
.B(n_1314),
.Y(n_1388)
);

HB1xp67_ASAP7_75t_L g1389 ( 
.A(n_1338),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1346),
.B(n_1325),
.Y(n_1390)
);

OAI21x1_ASAP7_75t_L g1391 ( 
.A1(n_1359),
.A2(n_1287),
.B(n_1318),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1363),
.B(n_1271),
.Y(n_1392)
);

BUFx6f_ASAP7_75t_L g1393 ( 
.A(n_1378),
.Y(n_1393)
);

AOI22xp33_ASAP7_75t_L g1394 ( 
.A1(n_1374),
.A2(n_1234),
.B1(n_1317),
.B2(n_1353),
.Y(n_1394)
);

OAI22xp5_ASAP7_75t_L g1395 ( 
.A1(n_1367),
.A2(n_1328),
.B1(n_1342),
.B2(n_1351),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1390),
.B(n_1349),
.Y(n_1396)
);

BUFx4f_ASAP7_75t_SL g1397 ( 
.A(n_1372),
.Y(n_1397)
);

OAI211xp5_ASAP7_75t_SL g1398 ( 
.A1(n_1369),
.A2(n_1351),
.B(n_1328),
.C(n_1371),
.Y(n_1398)
);

OAI21xp5_ASAP7_75t_L g1399 ( 
.A1(n_1375),
.A2(n_1262),
.B(n_1290),
.Y(n_1399)
);

OAI22xp33_ASAP7_75t_L g1400 ( 
.A1(n_1381),
.A2(n_1209),
.B1(n_1348),
.B2(n_1333),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1382),
.Y(n_1401)
);

INVx2_ASAP7_75t_L g1402 ( 
.A(n_1390),
.Y(n_1402)
);

NOR2xp33_ASAP7_75t_L g1403 ( 
.A(n_1372),
.B(n_1337),
.Y(n_1403)
);

AOI22xp33_ASAP7_75t_L g1404 ( 
.A1(n_1381),
.A2(n_1353),
.B1(n_1270),
.B2(n_1352),
.Y(n_1404)
);

OAI22xp33_ASAP7_75t_L g1405 ( 
.A1(n_1384),
.A2(n_1306),
.B1(n_1257),
.B2(n_1274),
.Y(n_1405)
);

AOI22xp33_ASAP7_75t_L g1406 ( 
.A1(n_1384),
.A2(n_1240),
.B1(n_1188),
.B2(n_1296),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1389),
.B(n_1329),
.Y(n_1407)
);

INVx3_ASAP7_75t_L g1408 ( 
.A(n_1373),
.Y(n_1408)
);

AOI22xp33_ASAP7_75t_L g1409 ( 
.A1(n_1366),
.A2(n_1368),
.B1(n_1380),
.B2(n_1373),
.Y(n_1409)
);

HB1xp67_ASAP7_75t_L g1410 ( 
.A(n_1370),
.Y(n_1410)
);

AOI22xp33_ASAP7_75t_L g1411 ( 
.A1(n_1366),
.A2(n_1299),
.B1(n_1362),
.B2(n_1272),
.Y(n_1411)
);

AOI211xp5_ASAP7_75t_L g1412 ( 
.A1(n_1392),
.A2(n_1134),
.B(n_1252),
.C(n_1321),
.Y(n_1412)
);

AOI22xp5_ASAP7_75t_L g1413 ( 
.A1(n_1386),
.A2(n_1246),
.B1(n_1289),
.B2(n_1281),
.Y(n_1413)
);

OAI21xp5_ASAP7_75t_SL g1414 ( 
.A1(n_1386),
.A2(n_1339),
.B(n_1332),
.Y(n_1414)
);

INVx3_ASAP7_75t_L g1415 ( 
.A(n_1373),
.Y(n_1415)
);

AOI221xp5_ASAP7_75t_L g1416 ( 
.A1(n_1382),
.A2(n_1294),
.B1(n_1303),
.B2(n_1181),
.C(n_1192),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1383),
.Y(n_1417)
);

INVxp67_ASAP7_75t_SL g1418 ( 
.A(n_1410),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1396),
.B(n_1383),
.Y(n_1419)
);

OR2x2_ASAP7_75t_L g1420 ( 
.A(n_1402),
.B(n_1410),
.Y(n_1420)
);

BUFx2_ASAP7_75t_L g1421 ( 
.A(n_1393),
.Y(n_1421)
);

HB1xp67_ASAP7_75t_L g1422 ( 
.A(n_1393),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1401),
.B(n_1376),
.Y(n_1423)
);

AND2x2_ASAP7_75t_SL g1424 ( 
.A(n_1408),
.B(n_1373),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_1417),
.Y(n_1425)
);

AOI21xp33_ASAP7_75t_L g1426 ( 
.A1(n_1395),
.A2(n_1398),
.B(n_1405),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1407),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1408),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1415),
.B(n_1376),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1415),
.B(n_1370),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1393),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1393),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1411),
.B(n_1388),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1409),
.B(n_1387),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1399),
.B(n_1388),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1414),
.B(n_1388),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1404),
.B(n_1387),
.Y(n_1437)
);

HB1xp67_ASAP7_75t_L g1438 ( 
.A(n_1397),
.Y(n_1438)
);

AOI22xp33_ASAP7_75t_L g1439 ( 
.A1(n_1426),
.A2(n_1394),
.B1(n_1405),
.B2(n_1413),
.Y(n_1439)
);

AOI211xp5_ASAP7_75t_L g1440 ( 
.A1(n_1435),
.A2(n_1400),
.B(n_1403),
.C(n_1412),
.Y(n_1440)
);

AOI222xp33_ASAP7_75t_L g1441 ( 
.A1(n_1435),
.A2(n_1400),
.B1(n_1416),
.B2(n_1406),
.C1(n_1380),
.C2(n_1210),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1425),
.Y(n_1442)
);

AOI221x1_ASAP7_75t_SL g1443 ( 
.A1(n_1419),
.A2(n_1339),
.B1(n_1388),
.B2(n_1181),
.C(n_1171),
.Y(n_1443)
);

AOI221xp5_ASAP7_75t_L g1444 ( 
.A1(n_1427),
.A2(n_1437),
.B1(n_1434),
.B2(n_1436),
.C(n_1433),
.Y(n_1444)
);

AOI22xp33_ASAP7_75t_L g1445 ( 
.A1(n_1433),
.A2(n_1386),
.B1(n_1380),
.B2(n_1362),
.Y(n_1445)
);

HB1xp67_ASAP7_75t_L g1446 ( 
.A(n_1418),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1425),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1420),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1420),
.Y(n_1449)
);

AO21x2_ASAP7_75t_L g1450 ( 
.A1(n_1431),
.A2(n_1359),
.B(n_1391),
.Y(n_1450)
);

INVxp67_ASAP7_75t_L g1451 ( 
.A(n_1438),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1446),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1448),
.B(n_1436),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1446),
.Y(n_1454)
);

NAND2x1p5_ASAP7_75t_L g1455 ( 
.A(n_1442),
.B(n_1424),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1449),
.Y(n_1456)
);

INVx1_ASAP7_75t_SL g1457 ( 
.A(n_1447),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1444),
.B(n_1427),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1451),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1445),
.B(n_1429),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1443),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1450),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1440),
.B(n_1429),
.Y(n_1463)
);

NOR2xp33_ASAP7_75t_L g1464 ( 
.A(n_1439),
.B(n_1422),
.Y(n_1464)
);

OR2x2_ASAP7_75t_L g1465 ( 
.A(n_1445),
.B(n_1423),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1441),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1452),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1456),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1453),
.B(n_1460),
.Y(n_1469)
);

OR2x2_ASAP7_75t_L g1470 ( 
.A(n_1454),
.B(n_1430),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1454),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1453),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1459),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1468),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1470),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1471),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1473),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_L g1478 ( 
.A1(n_1475),
.A2(n_1466),
.B1(n_1461),
.B2(n_1464),
.Y(n_1478)
);

OAI21xp5_ASAP7_75t_SL g1479 ( 
.A1(n_1477),
.A2(n_1464),
.B(n_1455),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1474),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1480),
.Y(n_1481)
);

AND2x4_ASAP7_75t_SL g1482 ( 
.A(n_1478),
.B(n_1380),
.Y(n_1482)
);

CKINVDCx16_ASAP7_75t_R g1483 ( 
.A(n_1479),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1478),
.B(n_1458),
.Y(n_1484)
);

OAI211xp5_ASAP7_75t_L g1485 ( 
.A1(n_1484),
.A2(n_1278),
.B(n_1166),
.C(n_1165),
.Y(n_1485)
);

NOR2x1_ASAP7_75t_L g1486 ( 
.A(n_1481),
.B(n_1474),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1482),
.Y(n_1487)
);

OAI22xp5_ASAP7_75t_L g1488 ( 
.A1(n_1483),
.A2(n_1463),
.B1(n_1469),
.B2(n_1476),
.Y(n_1488)
);

NOR2xp33_ASAP7_75t_L g1489 ( 
.A(n_1483),
.B(n_1467),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1488),
.B(n_1460),
.Y(n_1490)
);

AOI21xp5_ASAP7_75t_L g1491 ( 
.A1(n_1485),
.A2(n_1462),
.B(n_1472),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1486),
.Y(n_1492)
);

A2O1A1Ixp33_ASAP7_75t_L g1493 ( 
.A1(n_1487),
.A2(n_1462),
.B(n_1465),
.C(n_1457),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1489),
.B(n_1428),
.Y(n_1494)
);

OAI21xp33_ASAP7_75t_SL g1495 ( 
.A1(n_1489),
.A2(n_1386),
.B(n_1431),
.Y(n_1495)
);

INVx1_ASAP7_75t_SL g1496 ( 
.A(n_1487),
.Y(n_1496)
);

AOI21xp33_ASAP7_75t_L g1497 ( 
.A1(n_1496),
.A2(n_1492),
.B(n_1490),
.Y(n_1497)
);

OAI211xp5_ASAP7_75t_L g1498 ( 
.A1(n_1495),
.A2(n_1189),
.B(n_1204),
.C(n_1421),
.Y(n_1498)
);

NAND4xp25_ASAP7_75t_SL g1499 ( 
.A(n_1493),
.B(n_1432),
.C(n_1430),
.D(n_1316),
.Y(n_1499)
);

NOR2x1_ASAP7_75t_L g1500 ( 
.A(n_1494),
.B(n_1308),
.Y(n_1500)
);

AOI221xp5_ASAP7_75t_SL g1501 ( 
.A1(n_1491),
.A2(n_1301),
.B1(n_1379),
.B2(n_1277),
.C(n_1250),
.Y(n_1501)
);

NAND3xp33_ASAP7_75t_L g1502 ( 
.A(n_1492),
.B(n_1237),
.C(n_1250),
.Y(n_1502)
);

NOR2x1_ASAP7_75t_L g1503 ( 
.A(n_1499),
.B(n_1268),
.Y(n_1503)
);

BUFx2_ASAP7_75t_L g1504 ( 
.A(n_1500),
.Y(n_1504)
);

AOI22xp5_ASAP7_75t_L g1505 ( 
.A1(n_1497),
.A2(n_1341),
.B1(n_1385),
.B2(n_1377),
.Y(n_1505)
);

AOI221x1_ASAP7_75t_L g1506 ( 
.A1(n_1502),
.A2(n_1313),
.B1(n_1250),
.B2(n_1236),
.C(n_1219),
.Y(n_1506)
);

OAI22xp5_ASAP7_75t_L g1507 ( 
.A1(n_1498),
.A2(n_1365),
.B1(n_1385),
.B2(n_1377),
.Y(n_1507)
);

NOR2xp33_ASAP7_75t_L g1508 ( 
.A(n_1497),
.B(n_1377),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1501),
.B(n_1329),
.Y(n_1509)
);

AOI21xp5_ASAP7_75t_L g1510 ( 
.A1(n_1497),
.A2(n_1345),
.B(n_1292),
.Y(n_1510)
);

OAI21xp5_ASAP7_75t_L g1511 ( 
.A1(n_1497),
.A2(n_1345),
.B(n_1347),
.Y(n_1511)
);

INVx1_ASAP7_75t_SL g1512 ( 
.A(n_1497),
.Y(n_1512)
);

OAI211xp5_ASAP7_75t_SL g1513 ( 
.A1(n_1512),
.A2(n_133),
.B(n_134),
.C(n_135),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1504),
.Y(n_1514)
);

NAND4xp25_ASAP7_75t_L g1515 ( 
.A(n_1508),
.B(n_1385),
.C(n_1364),
.D(n_1358),
.Y(n_1515)
);

CKINVDCx5p33_ASAP7_75t_R g1516 ( 
.A(n_1505),
.Y(n_1516)
);

OAI211xp5_ASAP7_75t_SL g1517 ( 
.A1(n_1510),
.A2(n_137),
.B(n_141),
.C(n_143),
.Y(n_1517)
);

NAND3xp33_ASAP7_75t_L g1518 ( 
.A(n_1506),
.B(n_1219),
.C(n_1187),
.Y(n_1518)
);

NOR2xp33_ASAP7_75t_SL g1519 ( 
.A(n_1503),
.B(n_1276),
.Y(n_1519)
);

OR5x1_ASAP7_75t_L g1520 ( 
.A(n_1517),
.B(n_1509),
.C(n_1511),
.D(n_1507),
.E(n_151),
.Y(n_1520)
);

HB1xp67_ASAP7_75t_L g1521 ( 
.A(n_1516),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1515),
.Y(n_1522)
);

AND5x1_ASAP7_75t_L g1523 ( 
.A(n_1519),
.B(n_147),
.C(n_149),
.D(n_152),
.E(n_154),
.Y(n_1523)
);

NAND3xp33_ASAP7_75t_SL g1524 ( 
.A(n_1518),
.B(n_156),
.C(n_158),
.Y(n_1524)
);

AND4x1_ASAP7_75t_L g1525 ( 
.A(n_1513),
.B(n_159),
.C(n_160),
.D(n_162),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1514),
.Y(n_1526)
);

NOR2xp33_ASAP7_75t_L g1527 ( 
.A(n_1526),
.B(n_1521),
.Y(n_1527)
);

BUFx2_ASAP7_75t_L g1528 ( 
.A(n_1522),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1525),
.Y(n_1529)
);

INVx1_ASAP7_75t_SL g1530 ( 
.A(n_1520),
.Y(n_1530)
);

AOI21xp5_ASAP7_75t_L g1531 ( 
.A1(n_1527),
.A2(n_1524),
.B(n_1523),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1528),
.Y(n_1532)
);

OAI21x1_ASAP7_75t_L g1533 ( 
.A1(n_1529),
.A2(n_1355),
.B(n_1354),
.Y(n_1533)
);

AOI22xp5_ASAP7_75t_L g1534 ( 
.A1(n_1530),
.A2(n_1354),
.B1(n_1331),
.B2(n_1334),
.Y(n_1534)
);

AOI21xp5_ASAP7_75t_L g1535 ( 
.A1(n_1531),
.A2(n_1253),
.B(n_180),
.Y(n_1535)
);

OAI21x1_ASAP7_75t_SL g1536 ( 
.A1(n_1532),
.A2(n_181),
.B(n_184),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1536),
.Y(n_1537)
);

OAI22xp5_ASAP7_75t_L g1538 ( 
.A1(n_1537),
.A2(n_1535),
.B1(n_1534),
.B2(n_1533),
.Y(n_1538)
);

INVxp67_ASAP7_75t_L g1539 ( 
.A(n_1538),
.Y(n_1539)
);

OAI222xp33_ASAP7_75t_L g1540 ( 
.A1(n_1539),
.A2(n_1309),
.B1(n_185),
.B2(n_188),
.C1(n_191),
.C2(n_193),
.Y(n_1540)
);

AOI322xp5_ASAP7_75t_L g1541 ( 
.A1(n_1539),
.A2(n_1309),
.A3(n_194),
.B1(n_195),
.B2(n_199),
.C1(n_203),
.C2(n_204),
.Y(n_1541)
);

OAI221xp5_ASAP7_75t_R g1542 ( 
.A1(n_1540),
.A2(n_209),
.B1(n_211),
.B2(n_213),
.C(n_214),
.Y(n_1542)
);

AOI211xp5_ASAP7_75t_L g1543 ( 
.A1(n_1542),
.A2(n_1541),
.B(n_218),
.C(n_221),
.Y(n_1543)
);


endmodule