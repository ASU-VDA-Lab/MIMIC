module fake_netlist_5_860_n_1746 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_173, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_134, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1746);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_173;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_134;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1746;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_1723;
wire n_955;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1097;
wire n_1036;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_677;
wire n_293;
wire n_244;
wire n_1333;
wire n_1121;
wire n_433;
wire n_368;
wire n_314;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_259;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_968;
wire n_315;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1735;
wire n_1697;
wire n_1575;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_1722;
wire n_661;
wire n_849;
wire n_584;
wire n_336;
wire n_681;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_1683;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVx1_ASAP7_75t_SL g175 ( 
.A(n_132),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_98),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_174),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_68),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_75),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_101),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_49),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_38),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_87),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_48),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_0),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_33),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_48),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_37),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_115),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_19),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_12),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_73),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_92),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_163),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_100),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_126),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_15),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_81),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_14),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_162),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_24),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_120),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_102),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_62),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_88),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_35),
.Y(n_206)
);

BUFx10_ASAP7_75t_L g207 ( 
.A(n_122),
.Y(n_207)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_89),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_145),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_42),
.Y(n_210)
);

BUFx5_ASAP7_75t_L g211 ( 
.A(n_15),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_94),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_61),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_56),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_134),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_67),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_109),
.Y(n_217)
);

CKINVDCx14_ASAP7_75t_R g218 ( 
.A(n_123),
.Y(n_218)
);

BUFx10_ASAP7_75t_L g219 ( 
.A(n_152),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_6),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_125),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_170),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_24),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_76),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_129),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_18),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_168),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_66),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_71),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_164),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_91),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_36),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_58),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g234 ( 
.A(n_135),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_90),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_70),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_140),
.Y(n_237)
);

BUFx10_ASAP7_75t_L g238 ( 
.A(n_148),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_138),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_111),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_21),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_18),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_166),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_52),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_173),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_82),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_16),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_104),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_36),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_0),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_2),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_8),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_149),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_59),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_121),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_22),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_40),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_25),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_150),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_2),
.Y(n_260)
);

INVx2_ASAP7_75t_SL g261 ( 
.A(n_12),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_155),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_165),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_7),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_14),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_63),
.Y(n_266)
);

INVx2_ASAP7_75t_SL g267 ( 
.A(n_133),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_6),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_99),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_108),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_5),
.Y(n_271)
);

INVx1_ASAP7_75t_SL g272 ( 
.A(n_17),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_128),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_43),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_143),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_49),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_131),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_77),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_31),
.Y(n_279)
);

BUFx10_ASAP7_75t_L g280 ( 
.A(n_97),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_19),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_80),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_172),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_112),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_118),
.Y(n_285)
);

BUFx10_ASAP7_75t_L g286 ( 
.A(n_5),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_8),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_38),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_10),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_146),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_57),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_110),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_139),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_41),
.Y(n_294)
);

BUFx2_ASAP7_75t_L g295 ( 
.A(n_46),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_64),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_10),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_96),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_16),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_157),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_167),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_144),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_147),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_119),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_106),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_124),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_60),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_142),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_33),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_43),
.Y(n_310)
);

BUFx10_ASAP7_75t_L g311 ( 
.A(n_39),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_11),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_93),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_39),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_159),
.Y(n_315)
);

BUFx5_ASAP7_75t_L g316 ( 
.A(n_22),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_20),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_72),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_78),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_160),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_44),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_1),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_53),
.Y(n_323)
);

BUFx10_ASAP7_75t_L g324 ( 
.A(n_45),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_40),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_65),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_4),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_34),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_54),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_26),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_127),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_47),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_34),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_114),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_105),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_83),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_28),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_161),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_117),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_27),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_3),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_28),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_50),
.Y(n_343)
);

INVx2_ASAP7_75t_SL g344 ( 
.A(n_51),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_20),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_32),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_21),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_26),
.Y(n_348)
);

BUFx3_ASAP7_75t_L g349 ( 
.A(n_209),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_211),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_211),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_211),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_211),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_211),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_211),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_211),
.Y(n_356)
);

INVxp33_ASAP7_75t_SL g357 ( 
.A(n_190),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_316),
.Y(n_358)
);

BUFx3_ASAP7_75t_L g359 ( 
.A(n_209),
.Y(n_359)
);

CKINVDCx14_ASAP7_75t_R g360 ( 
.A(n_218),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_316),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_316),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_176),
.Y(n_363)
);

INVx1_ASAP7_75t_SL g364 ( 
.A(n_295),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_316),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_316),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_177),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_227),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_316),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_227),
.Y(n_370)
);

INVx3_ASAP7_75t_L g371 ( 
.A(n_182),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_316),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_182),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_182),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_182),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_179),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_230),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_230),
.Y(n_378)
);

HB1xp67_ASAP7_75t_L g379 ( 
.A(n_190),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_342),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_342),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_183),
.Y(n_382)
);

BUFx6f_ASAP7_75t_SL g383 ( 
.A(n_207),
.Y(n_383)
);

INVxp67_ASAP7_75t_SL g384 ( 
.A(n_203),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_342),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_200),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_342),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_187),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_187),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_282),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_202),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_205),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_327),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_210),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_210),
.Y(n_395)
);

INVxp67_ASAP7_75t_SL g396 ( 
.A(n_273),
.Y(n_396)
);

INVxp67_ASAP7_75t_SL g397 ( 
.A(n_300),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g398 ( 
.A(n_197),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_327),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_282),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_345),
.Y(n_401)
);

INVxp67_ASAP7_75t_SL g402 ( 
.A(n_285),
.Y(n_402)
);

INVxp67_ASAP7_75t_SL g403 ( 
.A(n_178),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_345),
.Y(n_404)
);

CKINVDCx16_ASAP7_75t_R g405 ( 
.A(n_222),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_184),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_348),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_188),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_347),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_213),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_199),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_197),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_214),
.Y(n_413)
);

INVxp67_ASAP7_75t_SL g414 ( 
.A(n_180),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_201),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_226),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_232),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_216),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_247),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_250),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_251),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_252),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_256),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_268),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_307),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_333),
.Y(n_426)
);

BUFx3_ASAP7_75t_L g427 ( 
.A(n_207),
.Y(n_427)
);

INVxp67_ASAP7_75t_SL g428 ( 
.A(n_189),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_341),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_307),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_261),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_261),
.Y(n_432)
);

INVxp67_ASAP7_75t_SL g433 ( 
.A(n_194),
.Y(n_433)
);

INVx3_ASAP7_75t_L g434 ( 
.A(n_217),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_204),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_361),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_361),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_373),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_350),
.Y(n_439)
);

HB1xp67_ASAP7_75t_L g440 ( 
.A(n_379),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_402),
.B(n_267),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_350),
.Y(n_442)
);

HB1xp67_ASAP7_75t_L g443 ( 
.A(n_398),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_403),
.B(n_414),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_428),
.B(n_267),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_351),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_373),
.Y(n_447)
);

INVxp67_ASAP7_75t_L g448 ( 
.A(n_412),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g449 ( 
.A(n_433),
.B(n_344),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_351),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_364),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_375),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_352),
.Y(n_453)
);

INVxp67_ASAP7_75t_SL g454 ( 
.A(n_371),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_375),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_368),
.Y(n_456)
);

INVxp67_ASAP7_75t_L g457 ( 
.A(n_349),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_370),
.Y(n_458)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_352),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_371),
.B(n_344),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_353),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_405),
.B(n_207),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_380),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_353),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_380),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_363),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_354),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_367),
.Y(n_468)
);

INVx3_ASAP7_75t_L g469 ( 
.A(n_354),
.Y(n_469)
);

INVxp67_ASAP7_75t_SL g470 ( 
.A(n_371),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_R g471 ( 
.A(n_360),
.B(n_221),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_355),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_374),
.B(n_192),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_381),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_355),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_356),
.Y(n_476)
);

BUFx3_ASAP7_75t_L g477 ( 
.A(n_374),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_356),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_381),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_435),
.B(n_192),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_385),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_358),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_385),
.B(n_193),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_387),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_358),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_362),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_387),
.B(n_193),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_362),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_365),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_365),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_366),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_366),
.Y(n_492)
);

NAND2xp33_ASAP7_75t_L g493 ( 
.A(n_434),
.B(n_304),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_369),
.Y(n_494)
);

INVx3_ASAP7_75t_L g495 ( 
.A(n_369),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_372),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_357),
.B(n_175),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_372),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_377),
.Y(n_499)
);

BUFx12f_ASAP7_75t_L g500 ( 
.A(n_376),
.Y(n_500)
);

INVx4_ASAP7_75t_L g501 ( 
.A(n_434),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_411),
.Y(n_502)
);

AND2x2_ASAP7_75t_SL g503 ( 
.A(n_434),
.B(n_217),
.Y(n_503)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_388),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_388),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_389),
.Y(n_506)
);

AND2x4_ASAP7_75t_L g507 ( 
.A(n_411),
.B(n_235),
.Y(n_507)
);

INVx4_ASAP7_75t_L g508 ( 
.A(n_349),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_389),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_359),
.B(n_195),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_393),
.Y(n_511)
);

HB1xp67_ASAP7_75t_L g512 ( 
.A(n_359),
.Y(n_512)
);

INVx3_ASAP7_75t_L g513 ( 
.A(n_393),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_488),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_497),
.B(n_382),
.Y(n_515)
);

CKINVDCx16_ASAP7_75t_R g516 ( 
.A(n_456),
.Y(n_516)
);

INVx3_ASAP7_75t_L g517 ( 
.A(n_459),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_437),
.Y(n_518)
);

BUFx2_ASAP7_75t_L g519 ( 
.A(n_451),
.Y(n_519)
);

INVx2_ASAP7_75t_SL g520 ( 
.A(n_451),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_445),
.B(n_384),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_437),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_437),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_497),
.B(n_386),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_448),
.A2(n_397),
.B1(n_396),
.B2(n_391),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_466),
.B(n_392),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_454),
.B(n_410),
.Y(n_527)
);

BUFx3_ASAP7_75t_L g528 ( 
.A(n_494),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_500),
.Y(n_529)
);

INVx4_ASAP7_75t_L g530 ( 
.A(n_459),
.Y(n_530)
);

OAI21xp33_ASAP7_75t_SL g531 ( 
.A1(n_441),
.A2(n_326),
.B(n_235),
.Y(n_531)
);

INVx3_ASAP7_75t_L g532 ( 
.A(n_459),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_437),
.Y(n_533)
);

INVx4_ASAP7_75t_SL g534 ( 
.A(n_459),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_477),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_494),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_475),
.Y(n_537)
);

INVx3_ASAP7_75t_L g538 ( 
.A(n_459),
.Y(n_538)
);

BUFx6f_ASAP7_75t_L g539 ( 
.A(n_459),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_444),
.B(n_413),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_459),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_454),
.B(n_418),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_466),
.B(n_427),
.Y(n_543)
);

INVx3_ASAP7_75t_L g544 ( 
.A(n_459),
.Y(n_544)
);

BUFx2_ASAP7_75t_L g545 ( 
.A(n_512),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_470),
.B(n_427),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_475),
.Y(n_547)
);

BUFx3_ASAP7_75t_L g548 ( 
.A(n_512),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_477),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_477),
.Y(n_550)
);

AOI22xp33_ASAP7_75t_L g551 ( 
.A1(n_445),
.A2(n_395),
.B1(n_394),
.B2(n_304),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_477),
.Y(n_552)
);

INVx2_ASAP7_75t_SL g553 ( 
.A(n_510),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_475),
.Y(n_554)
);

NAND3xp33_ASAP7_75t_L g555 ( 
.A(n_448),
.B(n_206),
.C(n_186),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_439),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_439),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_470),
.B(n_208),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_468),
.B(n_219),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_469),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_469),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_439),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_439),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_464),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_469),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_442),
.Y(n_566)
);

OAI22x1_ASAP7_75t_L g567 ( 
.A1(n_440),
.A2(n_443),
.B1(n_462),
.B2(n_340),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_R g568 ( 
.A(n_468),
.B(n_378),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_442),
.Y(n_569)
);

AOI22xp33_ASAP7_75t_L g570 ( 
.A1(n_445),
.A2(n_304),
.B1(n_420),
.B2(n_429),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_449),
.B(n_234),
.Y(n_571)
);

INVx3_ASAP7_75t_L g572 ( 
.A(n_464),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_442),
.Y(n_573)
);

NAND2xp33_ASAP7_75t_L g574 ( 
.A(n_449),
.B(n_304),
.Y(n_574)
);

INVx3_ASAP7_75t_L g575 ( 
.A(n_464),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_449),
.B(n_255),
.Y(n_576)
);

INVx2_ASAP7_75t_SL g577 ( 
.A(n_510),
.Y(n_577)
);

BUFx4f_ASAP7_75t_L g578 ( 
.A(n_503),
.Y(n_578)
);

INVx5_ASAP7_75t_L g579 ( 
.A(n_464),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_469),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_495),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_495),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_457),
.B(n_219),
.Y(n_583)
);

XNOR2xp5_ASAP7_75t_L g584 ( 
.A(n_456),
.B(n_390),
.Y(n_584)
);

INVxp67_ASAP7_75t_SL g585 ( 
.A(n_457),
.Y(n_585)
);

NAND3xp33_ASAP7_75t_L g586 ( 
.A(n_480),
.B(n_223),
.C(n_220),
.Y(n_586)
);

HB1xp67_ASAP7_75t_L g587 ( 
.A(n_440),
.Y(n_587)
);

BUFx3_ASAP7_75t_L g588 ( 
.A(n_508),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_442),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_495),
.Y(n_590)
);

OAI22xp33_ASAP7_75t_L g591 ( 
.A1(n_444),
.A2(n_272),
.B1(n_242),
.B2(n_343),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_508),
.B(n_383),
.Y(n_592)
);

AND2x4_ASAP7_75t_L g593 ( 
.A(n_508),
.B(n_406),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_471),
.B(n_219),
.Y(n_594)
);

NAND3xp33_ASAP7_75t_L g595 ( 
.A(n_480),
.B(n_249),
.C(n_241),
.Y(n_595)
);

BUFx6f_ASAP7_75t_L g596 ( 
.A(n_464),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_495),
.Y(n_597)
);

INVx3_ASAP7_75t_L g598 ( 
.A(n_464),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_508),
.B(n_399),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_495),
.Y(n_600)
);

BUFx6f_ASAP7_75t_L g601 ( 
.A(n_464),
.Y(n_601)
);

INVx3_ASAP7_75t_L g602 ( 
.A(n_464),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_508),
.B(n_277),
.Y(n_603)
);

BUFx10_ASAP7_75t_L g604 ( 
.A(n_503),
.Y(n_604)
);

BUFx4f_ASAP7_75t_L g605 ( 
.A(n_503),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_446),
.Y(n_606)
);

BUFx6f_ASAP7_75t_L g607 ( 
.A(n_476),
.Y(n_607)
);

BUFx6f_ASAP7_75t_L g608 ( 
.A(n_476),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_483),
.B(n_383),
.Y(n_609)
);

AND2x6_ASAP7_75t_L g610 ( 
.A(n_446),
.B(n_212),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_446),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_446),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_450),
.Y(n_613)
);

OR2x2_ASAP7_75t_L g614 ( 
.A(n_443),
.B(n_432),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_450),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_450),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_483),
.B(n_487),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_450),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_471),
.B(n_462),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_453),
.Y(n_620)
);

BUFx3_ASAP7_75t_L g621 ( 
.A(n_507),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_453),
.Y(n_622)
);

NAND2xp33_ASAP7_75t_L g623 ( 
.A(n_476),
.B(n_215),
.Y(n_623)
);

AOI21x1_ASAP7_75t_L g624 ( 
.A1(n_460),
.A2(n_229),
.B(n_225),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_453),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_501),
.B(n_302),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_453),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_461),
.Y(n_628)
);

AO22x2_ASAP7_75t_L g629 ( 
.A1(n_507),
.A2(n_269),
.B1(n_338),
.B2(n_278),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_461),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_461),
.Y(n_631)
);

NAND2xp33_ASAP7_75t_SL g632 ( 
.A(n_473),
.B(n_181),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_502),
.B(n_473),
.Y(n_633)
);

INVx3_ASAP7_75t_L g634 ( 
.A(n_476),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_500),
.B(n_238),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_487),
.B(n_383),
.Y(n_636)
);

CKINVDCx20_ASAP7_75t_R g637 ( 
.A(n_458),
.Y(n_637)
);

INVx5_ASAP7_75t_L g638 ( 
.A(n_476),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_461),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_467),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_467),
.Y(n_641)
);

OR2x6_ASAP7_75t_L g642 ( 
.A(n_500),
.B(n_431),
.Y(n_642)
);

NAND2xp33_ASAP7_75t_L g643 ( 
.A(n_476),
.B(n_233),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_467),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_500),
.B(n_238),
.Y(n_645)
);

INVx2_ASAP7_75t_SL g646 ( 
.A(n_460),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_467),
.Y(n_647)
);

XNOR2xp5_ASAP7_75t_L g648 ( 
.A(n_458),
.B(n_400),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_472),
.Y(n_649)
);

INVx2_ASAP7_75t_SL g650 ( 
.A(n_507),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_472),
.Y(n_651)
);

BUFx6f_ASAP7_75t_SL g652 ( 
.A(n_507),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_507),
.B(n_238),
.Y(n_653)
);

INVx3_ASAP7_75t_L g654 ( 
.A(n_476),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_472),
.Y(n_655)
);

INVx2_ASAP7_75t_SL g656 ( 
.A(n_507),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_472),
.Y(n_657)
);

OR2x6_ASAP7_75t_L g658 ( 
.A(n_502),
.B(n_431),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_438),
.B(n_399),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_501),
.B(n_224),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_478),
.Y(n_661)
);

INVx2_ASAP7_75t_SL g662 ( 
.A(n_501),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_659),
.Y(n_663)
);

AND2x4_ASAP7_75t_L g664 ( 
.A(n_548),
.B(n_406),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_R g665 ( 
.A(n_529),
.B(n_499),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_547),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_617),
.B(n_501),
.Y(n_667)
);

BUFx3_ASAP7_75t_L g668 ( 
.A(n_548),
.Y(n_668)
);

OR2x6_ASAP7_75t_L g669 ( 
.A(n_520),
.B(n_432),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_659),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_518),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_553),
.B(n_195),
.Y(n_672)
);

NOR3xp33_ASAP7_75t_L g673 ( 
.A(n_520),
.B(n_408),
.C(n_407),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_577),
.B(n_476),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_578),
.B(n_478),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_518),
.Y(n_676)
);

AOI221xp5_ASAP7_75t_L g677 ( 
.A1(n_591),
.A2(n_265),
.B1(n_314),
.B2(n_279),
.C(n_191),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_577),
.B(n_478),
.Y(n_678)
);

AND2x6_ASAP7_75t_L g679 ( 
.A(n_633),
.B(n_237),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_540),
.B(n_478),
.Y(n_680)
);

OAI22xp5_ASAP7_75t_L g681 ( 
.A1(n_578),
.A2(n_323),
.B1(n_303),
.B2(n_296),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_519),
.B(n_425),
.Y(n_682)
);

BUFx12f_ASAP7_75t_L g683 ( 
.A(n_519),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_SL g684 ( 
.A(n_529),
.B(n_181),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_SL g685 ( 
.A(n_587),
.B(n_185),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_578),
.B(n_482),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_522),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_522),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_646),
.B(n_482),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_605),
.B(n_604),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_621),
.Y(n_691)
);

AND2x4_ASAP7_75t_SL g692 ( 
.A(n_642),
.B(n_430),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_605),
.B(n_482),
.Y(n_693)
);

INVx3_ASAP7_75t_L g694 ( 
.A(n_621),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_547),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_528),
.Y(n_696)
);

BUFx6f_ASAP7_75t_L g697 ( 
.A(n_528),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_646),
.B(n_485),
.Y(n_698)
);

NOR2xp67_ASAP7_75t_L g699 ( 
.A(n_586),
.B(n_438),
.Y(n_699)
);

HB1xp67_ASAP7_75t_L g700 ( 
.A(n_545),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_662),
.B(n_485),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_514),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_554),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_662),
.B(n_486),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_604),
.B(n_486),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_650),
.B(n_486),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_523),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_521),
.B(n_286),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_527),
.B(n_196),
.Y(n_709)
);

HB1xp67_ASAP7_75t_L g710 ( 
.A(n_545),
.Y(n_710)
);

AOI22xp33_ASAP7_75t_L g711 ( 
.A1(n_629),
.A2(n_185),
.B1(n_191),
.B2(n_322),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_536),
.B(n_486),
.Y(n_712)
);

BUFx2_ASAP7_75t_L g713 ( 
.A(n_637),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_523),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_521),
.B(n_489),
.Y(n_715)
);

HB1xp67_ASAP7_75t_L g716 ( 
.A(n_614),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_650),
.B(n_489),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_533),
.Y(n_718)
);

AOI22xp5_ASAP7_75t_L g719 ( 
.A1(n_571),
.A2(n_290),
.B1(n_291),
.B2(n_292),
.Y(n_719)
);

NAND2xp33_ASAP7_75t_L g720 ( 
.A(n_576),
.B(n_626),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_537),
.B(n_489),
.Y(n_721)
);

INVx2_ASAP7_75t_SL g722 ( 
.A(n_614),
.Y(n_722)
);

NOR2xp67_ASAP7_75t_L g723 ( 
.A(n_595),
.B(n_447),
.Y(n_723)
);

INVx8_ASAP7_75t_L g724 ( 
.A(n_642),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_656),
.Y(n_725)
);

OAI22xp5_ASAP7_75t_L g726 ( 
.A1(n_542),
.A2(n_329),
.B1(n_283),
.B2(n_263),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_556),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_546),
.B(n_196),
.Y(n_728)
);

INVx4_ASAP7_75t_L g729 ( 
.A(n_588),
.Y(n_729)
);

NOR2x1p5_ASAP7_75t_L g730 ( 
.A(n_585),
.B(n_337),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_656),
.B(n_490),
.Y(n_731)
);

INVxp67_ASAP7_75t_SL g732 ( 
.A(n_539),
.Y(n_732)
);

OAI22xp33_ASAP7_75t_L g733 ( 
.A1(n_567),
.A2(n_322),
.B1(n_265),
.B2(n_314),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_515),
.B(n_198),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_593),
.B(n_490),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_599),
.Y(n_736)
);

INVx2_ASAP7_75t_SL g737 ( 
.A(n_558),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_554),
.B(n_490),
.Y(n_738)
);

NAND2xp33_ASAP7_75t_L g739 ( 
.A(n_603),
.B(n_228),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_535),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_599),
.B(n_491),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_597),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_597),
.B(n_491),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_600),
.B(n_491),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_535),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_524),
.B(n_198),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_600),
.B(n_492),
.Y(n_747)
);

NAND2xp33_ASAP7_75t_L g748 ( 
.A(n_660),
.B(n_560),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_658),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_561),
.B(n_492),
.Y(n_750)
);

AOI22xp5_ASAP7_75t_L g751 ( 
.A1(n_632),
.A2(n_239),
.B1(n_320),
.B2(n_319),
.Y(n_751)
);

INVx3_ASAP7_75t_L g752 ( 
.A(n_549),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_556),
.Y(n_753)
);

NOR2xp67_ASAP7_75t_L g754 ( 
.A(n_525),
.B(n_447),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_565),
.B(n_492),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_557),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_658),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_658),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_580),
.B(n_496),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_557),
.Y(n_760)
);

HB1xp67_ASAP7_75t_L g761 ( 
.A(n_658),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_562),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_581),
.B(n_496),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_582),
.B(n_496),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_590),
.B(n_498),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_562),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_568),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_609),
.B(n_498),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_570),
.B(n_498),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_636),
.B(n_574),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_531),
.B(n_243),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_637),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_543),
.B(n_286),
.Y(n_773)
);

OAI22xp5_ASAP7_75t_L g774 ( 
.A1(n_551),
.A2(n_334),
.B1(n_331),
.B2(n_318),
.Y(n_774)
);

OR2x6_ASAP7_75t_L g775 ( 
.A(n_642),
.B(n_407),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_574),
.B(n_436),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_549),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_550),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_550),
.B(n_253),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_R g780 ( 
.A(n_516),
.B(n_499),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_552),
.B(n_436),
.Y(n_781)
);

BUFx2_ASAP7_75t_L g782 ( 
.A(n_632),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_552),
.B(n_436),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_539),
.B(n_259),
.Y(n_784)
);

NAND2xp33_ASAP7_75t_L g785 ( 
.A(n_610),
.B(n_231),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_517),
.B(n_532),
.Y(n_786)
);

AOI22xp5_ASAP7_75t_L g787 ( 
.A1(n_619),
.A2(n_306),
.B1(n_240),
.B2(n_244),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_517),
.B(n_504),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_563),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_539),
.B(n_305),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_559),
.B(n_339),
.Y(n_791)
);

BUFx2_ASAP7_75t_L g792 ( 
.A(n_584),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_539),
.B(n_541),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_606),
.Y(n_794)
);

AND2x4_ASAP7_75t_SL g795 ( 
.A(n_642),
.B(n_280),
.Y(n_795)
);

AND2x4_ASAP7_75t_L g796 ( 
.A(n_653),
.B(n_408),
.Y(n_796)
);

AND2x2_ASAP7_75t_L g797 ( 
.A(n_526),
.B(n_311),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_563),
.Y(n_798)
);

INVx2_ASAP7_75t_SL g799 ( 
.A(n_583),
.Y(n_799)
);

NAND3xp33_ASAP7_75t_SL g800 ( 
.A(n_635),
.B(n_279),
.C(n_337),
.Y(n_800)
);

OR2x2_ASAP7_75t_L g801 ( 
.A(n_555),
.B(n_409),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_539),
.B(n_236),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_657),
.Y(n_803)
);

A2O1A1Ixp33_ASAP7_75t_L g804 ( 
.A1(n_592),
.A2(n_426),
.B(n_409),
.C(n_415),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_657),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_541),
.B(n_245),
.Y(n_806)
);

INVx2_ASAP7_75t_SL g807 ( 
.A(n_567),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_566),
.Y(n_808)
);

INVx8_ASAP7_75t_L g809 ( 
.A(n_652),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_594),
.B(n_339),
.Y(n_810)
);

BUFx3_ASAP7_75t_L g811 ( 
.A(n_610),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_566),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_569),
.Y(n_813)
);

AND2x4_ASAP7_75t_L g814 ( 
.A(n_645),
.B(n_415),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_L g815 ( 
.A(n_611),
.B(n_257),
.Y(n_815)
);

AOI22xp5_ASAP7_75t_L g816 ( 
.A1(n_652),
.A2(n_629),
.B1(n_610),
.B2(n_623),
.Y(n_816)
);

AOI22xp33_ASAP7_75t_L g817 ( 
.A1(n_629),
.A2(n_513),
.B1(n_504),
.B2(n_340),
.Y(n_817)
);

OR2x2_ASAP7_75t_L g818 ( 
.A(n_584),
.B(n_416),
.Y(n_818)
);

BUFx3_ASAP7_75t_L g819 ( 
.A(n_683),
.Y(n_819)
);

AOI22xp33_ASAP7_75t_L g820 ( 
.A1(n_679),
.A2(n_652),
.B1(n_610),
.B2(n_615),
.Y(n_820)
);

INVx5_ASAP7_75t_L g821 ( 
.A(n_809),
.Y(n_821)
);

BUFx2_ASAP7_75t_L g822 ( 
.A(n_700),
.Y(n_822)
);

AOI22xp5_ASAP7_75t_L g823 ( 
.A1(n_720),
.A2(n_610),
.B1(n_538),
.B2(n_654),
.Y(n_823)
);

NOR2x2_ASAP7_75t_L g824 ( 
.A(n_775),
.B(n_648),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_L g825 ( 
.A(n_737),
.B(n_648),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_666),
.Y(n_826)
);

AND2x4_ASAP7_75t_L g827 ( 
.A(n_668),
.B(n_416),
.Y(n_827)
);

OR2x6_ASAP7_75t_SL g828 ( 
.A(n_767),
.B(n_258),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_695),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_695),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_752),
.Y(n_831)
);

INVx2_ASAP7_75t_SL g832 ( 
.A(n_710),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_703),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_780),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_722),
.B(n_530),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_703),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_742),
.Y(n_837)
);

INVxp67_ASAP7_75t_L g838 ( 
.A(n_716),
.Y(n_838)
);

AOI22xp5_ASAP7_75t_L g839 ( 
.A1(n_679),
.A2(n_602),
.B1(n_538),
.B2(n_654),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_725),
.Y(n_840)
);

BUFx6f_ASAP7_75t_SL g841 ( 
.A(n_668),
.Y(n_841)
);

CKINVDCx20_ASAP7_75t_R g842 ( 
.A(n_780),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_702),
.Y(n_843)
);

INVx5_ASAP7_75t_L g844 ( 
.A(n_809),
.Y(n_844)
);

BUFx12f_ASAP7_75t_L g845 ( 
.A(n_772),
.Y(n_845)
);

BUFx6f_ASAP7_75t_L g846 ( 
.A(n_809),
.Y(n_846)
);

INVx2_ASAP7_75t_SL g847 ( 
.A(n_664),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_697),
.B(n_246),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_667),
.B(n_544),
.Y(n_849)
);

AOI22xp33_ASAP7_75t_L g850 ( 
.A1(n_679),
.A2(n_612),
.B1(n_616),
.B2(n_620),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_680),
.B(n_544),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_691),
.Y(n_852)
);

AND2x4_ASAP7_75t_L g853 ( 
.A(n_696),
.B(n_417),
.Y(n_853)
);

NAND2x1p5_ASAP7_75t_L g854 ( 
.A(n_694),
.B(n_544),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_665),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_R g856 ( 
.A(n_800),
.B(n_684),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_752),
.Y(n_857)
);

BUFx2_ASAP7_75t_L g858 ( 
.A(n_682),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_740),
.Y(n_859)
);

AOI22xp5_ASAP7_75t_L g860 ( 
.A1(n_679),
.A2(n_634),
.B1(n_564),
.B2(n_572),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_709),
.B(n_564),
.Y(n_861)
);

XOR2xp5_ASAP7_75t_L g862 ( 
.A(n_792),
.B(n_248),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_740),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_745),
.Y(n_864)
);

AOI22xp33_ASAP7_75t_L g865 ( 
.A1(n_679),
.A2(n_631),
.B1(n_625),
.B2(n_630),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_794),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_715),
.B(n_639),
.Y(n_867)
);

AND2x6_ASAP7_75t_SL g868 ( 
.A(n_734),
.B(n_417),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_736),
.B(n_641),
.Y(n_869)
);

INVxp67_ASAP7_75t_L g870 ( 
.A(n_708),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_678),
.B(n_647),
.Y(n_871)
);

AND2x4_ASAP7_75t_L g872 ( 
.A(n_749),
.B(n_419),
.Y(n_872)
);

NAND3xp33_ASAP7_75t_SL g873 ( 
.A(n_677),
.B(n_264),
.C(n_260),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_709),
.B(n_564),
.Y(n_874)
);

AOI22xp5_ASAP7_75t_L g875 ( 
.A1(n_690),
.A2(n_575),
.B1(n_598),
.B2(n_572),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_665),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_728),
.B(n_572),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_689),
.B(n_569),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_697),
.B(n_254),
.Y(n_879)
);

AND2x4_ASAP7_75t_L g880 ( 
.A(n_757),
.B(n_419),
.Y(n_880)
);

OAI22xp5_ASAP7_75t_SL g881 ( 
.A1(n_711),
.A2(n_309),
.B1(n_274),
.B2(n_271),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_698),
.B(n_573),
.Y(n_882)
);

AO22x1_ASAP7_75t_L g883 ( 
.A1(n_791),
.A2(n_330),
.B1(n_281),
.B2(n_276),
.Y(n_883)
);

BUFx2_ASAP7_75t_L g884 ( 
.A(n_713),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_728),
.B(n_575),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_803),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_672),
.B(n_575),
.Y(n_887)
);

AND2x4_ASAP7_75t_L g888 ( 
.A(n_758),
.B(n_420),
.Y(n_888)
);

AND2x4_ASAP7_75t_L g889 ( 
.A(n_663),
.B(n_421),
.Y(n_889)
);

INVx5_ASAP7_75t_L g890 ( 
.A(n_775),
.Y(n_890)
);

OR2x6_ASAP7_75t_L g891 ( 
.A(n_724),
.B(n_421),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_697),
.B(n_262),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_805),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_670),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_777),
.Y(n_895)
);

AND2x2_ASAP7_75t_SL g896 ( 
.A(n_711),
.B(n_623),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_672),
.B(n_598),
.Y(n_897)
);

NAND2xp33_ASAP7_75t_L g898 ( 
.A(n_770),
.B(n_541),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_664),
.B(n_311),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_L g900 ( 
.A(n_734),
.B(n_530),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_SL g901 ( 
.A(n_697),
.B(n_266),
.Y(n_901)
);

NOR3xp33_ASAP7_75t_SL g902 ( 
.A(n_733),
.B(n_310),
.C(n_287),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_778),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_745),
.Y(n_904)
);

AOI22xp5_ASAP7_75t_L g905 ( 
.A1(n_690),
.A2(n_746),
.B1(n_694),
.B2(n_723),
.Y(n_905)
);

INVx2_ASAP7_75t_SL g906 ( 
.A(n_669),
.Y(n_906)
);

BUFx4f_ASAP7_75t_SL g907 ( 
.A(n_782),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_L g908 ( 
.A(n_818),
.B(n_288),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_674),
.B(n_573),
.Y(n_909)
);

AND2x4_ASAP7_75t_L g910 ( 
.A(n_761),
.B(n_422),
.Y(n_910)
);

INVx3_ASAP7_75t_L g911 ( 
.A(n_729),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_789),
.Y(n_912)
);

AND2x6_ASAP7_75t_SL g913 ( 
.A(n_791),
.B(n_422),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_735),
.A2(n_608),
.B(n_541),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_768),
.B(n_589),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_808),
.Y(n_916)
);

AND2x4_ASAP7_75t_L g917 ( 
.A(n_775),
.B(n_814),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_671),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_L g919 ( 
.A(n_685),
.B(n_289),
.Y(n_919)
);

INVx2_ASAP7_75t_SL g920 ( 
.A(n_669),
.Y(n_920)
);

HB1xp67_ASAP7_75t_L g921 ( 
.A(n_669),
.Y(n_921)
);

INVx3_ASAP7_75t_L g922 ( 
.A(n_729),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_676),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_796),
.B(n_613),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_812),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_813),
.Y(n_926)
);

INVx2_ASAP7_75t_SL g927 ( 
.A(n_801),
.Y(n_927)
);

INVx2_ASAP7_75t_SL g928 ( 
.A(n_730),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_687),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_741),
.B(n_675),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_744),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_744),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_675),
.B(n_618),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_747),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_688),
.Y(n_935)
);

AND2x4_ASAP7_75t_L g936 ( 
.A(n_814),
.B(n_423),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_686),
.B(n_618),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_686),
.B(n_622),
.Y(n_938)
);

OAI21xp5_ASAP7_75t_L g939 ( 
.A1(n_693),
.A2(n_661),
.B(n_655),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_SL g940 ( 
.A(n_799),
.B(n_270),
.Y(n_940)
);

INVx2_ASAP7_75t_SL g941 ( 
.A(n_797),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_692),
.Y(n_942)
);

INVx8_ASAP7_75t_L g943 ( 
.A(n_724),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_SL g944 ( 
.A(n_810),
.B(n_275),
.Y(n_944)
);

BUFx3_ASAP7_75t_L g945 ( 
.A(n_724),
.Y(n_945)
);

AOI22xp5_ASAP7_75t_L g946 ( 
.A1(n_699),
.A2(n_643),
.B1(n_649),
.B2(n_644),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_747),
.Y(n_947)
);

OAI21xp5_ASAP7_75t_L g948 ( 
.A1(n_693),
.A2(n_651),
.B(n_649),
.Y(n_948)
);

BUFx3_ASAP7_75t_L g949 ( 
.A(n_773),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_L g950 ( 
.A(n_810),
.B(n_294),
.Y(n_950)
);

INVx3_ASAP7_75t_L g951 ( 
.A(n_811),
.Y(n_951)
);

NAND2x1p5_ASAP7_75t_L g952 ( 
.A(n_811),
.B(n_541),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_738),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_707),
.Y(n_954)
);

AOI22xp33_ASAP7_75t_L g955 ( 
.A1(n_771),
.A2(n_640),
.B1(n_628),
.B2(n_627),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_738),
.Y(n_956)
);

OR2x2_ASAP7_75t_L g957 ( 
.A(n_673),
.B(n_424),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_712),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_SL g959 ( 
.A(n_719),
.B(n_284),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_727),
.Y(n_960)
);

A2O1A1Ixp33_ASAP7_75t_L g961 ( 
.A1(n_815),
.A2(n_627),
.B(n_513),
.C(n_463),
.Y(n_961)
);

NOR2xp33_ASAP7_75t_L g962 ( 
.A(n_733),
.B(n_751),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_753),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_756),
.Y(n_964)
);

INVx3_ASAP7_75t_L g965 ( 
.A(n_760),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_705),
.B(n_596),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_762),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_766),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_795),
.Y(n_969)
);

AOI22xp5_ASAP7_75t_L g970 ( 
.A1(n_802),
.A2(n_293),
.B1(n_336),
.B2(n_315),
.Y(n_970)
);

INVx3_ASAP7_75t_L g971 ( 
.A(n_798),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_SL g972 ( 
.A(n_754),
.B(n_298),
.Y(n_972)
);

BUFx4f_ASAP7_75t_L g973 ( 
.A(n_795),
.Y(n_973)
);

BUFx3_ASAP7_75t_L g974 ( 
.A(n_787),
.Y(n_974)
);

OR2x6_ASAP7_75t_L g975 ( 
.A(n_771),
.B(n_424),
.Y(n_975)
);

INVxp67_ASAP7_75t_L g976 ( 
.A(n_815),
.Y(n_976)
);

BUFx2_ASAP7_75t_L g977 ( 
.A(n_804),
.Y(n_977)
);

NAND3xp33_ASAP7_75t_SL g978 ( 
.A(n_817),
.B(n_726),
.C(n_816),
.Y(n_978)
);

AOI22xp5_ASAP7_75t_L g979 ( 
.A1(n_802),
.A2(n_335),
.B1(n_301),
.B2(n_313),
.Y(n_979)
);

BUFx3_ASAP7_75t_L g980 ( 
.A(n_714),
.Y(n_980)
);

NOR2xp33_ASAP7_75t_L g981 ( 
.A(n_806),
.B(n_297),
.Y(n_981)
);

AND2x4_ASAP7_75t_L g982 ( 
.A(n_804),
.B(n_732),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_706),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_R g984 ( 
.A(n_739),
.B(n_624),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_701),
.B(n_601),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_704),
.B(n_601),
.Y(n_986)
);

BUFx6f_ASAP7_75t_L g987 ( 
.A(n_793),
.Y(n_987)
);

BUFx12f_ASAP7_75t_SL g988 ( 
.A(n_817),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_748),
.A2(n_608),
.B(n_607),
.Y(n_989)
);

BUFx2_ASAP7_75t_L g990 ( 
.A(n_884),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_859),
.Y(n_991)
);

BUFx4f_ASAP7_75t_L g992 ( 
.A(n_846),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_930),
.A2(n_898),
.B(n_900),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_976),
.B(n_743),
.Y(n_994)
);

BUFx2_ASAP7_75t_L g995 ( 
.A(n_822),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_SL g996 ( 
.A(n_927),
.B(n_806),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_950),
.B(n_838),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_863),
.Y(n_998)
);

OAI22xp5_ASAP7_75t_L g999 ( 
.A1(n_905),
.A2(n_731),
.B1(n_717),
.B2(n_786),
.Y(n_999)
);

BUFx3_ASAP7_75t_L g1000 ( 
.A(n_846),
.Y(n_1000)
);

OAI21xp33_ASAP7_75t_L g1001 ( 
.A1(n_908),
.A2(n_774),
.B(n_317),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_R g1002 ( 
.A(n_834),
.B(n_785),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_864),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_958),
.B(n_721),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_843),
.B(n_781),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_930),
.A2(n_717),
.B(n_769),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_826),
.Y(n_1007)
);

AOI22x1_ASAP7_75t_SL g1008 ( 
.A1(n_855),
.A2(n_312),
.B1(n_299),
.B2(n_346),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_849),
.A2(n_769),
.B(n_783),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_870),
.B(n_718),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_904),
.Y(n_1011)
);

INVx3_ASAP7_75t_SL g1012 ( 
.A(n_824),
.Y(n_1012)
);

A2O1A1Ixp33_ASAP7_75t_L g1013 ( 
.A1(n_981),
.A2(n_788),
.B(n_776),
.C(n_790),
.Y(n_1013)
);

O2A1O1Ixp33_ASAP7_75t_L g1014 ( 
.A1(n_978),
.A2(n_779),
.B(n_790),
.C(n_784),
.Y(n_1014)
);

AOI22xp5_ASAP7_75t_L g1015 ( 
.A1(n_941),
.A2(n_974),
.B1(n_825),
.B2(n_873),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_894),
.B(n_755),
.Y(n_1016)
);

CKINVDCx8_ASAP7_75t_R g1017 ( 
.A(n_868),
.Y(n_1017)
);

BUFx6f_ASAP7_75t_L g1018 ( 
.A(n_846),
.Y(n_1018)
);

INVx3_ASAP7_75t_SL g1019 ( 
.A(n_942),
.Y(n_1019)
);

HB1xp67_ASAP7_75t_L g1020 ( 
.A(n_832),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_829),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_845),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_842),
.Y(n_1023)
);

OR2x6_ASAP7_75t_SL g1024 ( 
.A(n_876),
.B(n_321),
.Y(n_1024)
);

OAI21x1_ASAP7_75t_L g1025 ( 
.A1(n_939),
.A2(n_764),
.B(n_763),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_830),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_833),
.Y(n_1027)
);

INVx1_ASAP7_75t_SL g1028 ( 
.A(n_858),
.Y(n_1028)
);

INVx3_ASAP7_75t_SL g1029 ( 
.A(n_969),
.Y(n_1029)
);

OAI22xp5_ASAP7_75t_SL g1030 ( 
.A1(n_881),
.A2(n_328),
.B1(n_325),
.B2(n_332),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_936),
.B(n_311),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_840),
.B(n_866),
.Y(n_1032)
);

O2A1O1Ixp33_ASAP7_75t_L g1033 ( 
.A1(n_977),
.A2(n_750),
.B(n_765),
.C(n_759),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_836),
.Y(n_1034)
);

OR2x2_ASAP7_75t_L g1035 ( 
.A(n_847),
.B(n_426),
.Y(n_1035)
);

AOI33xp33_ASAP7_75t_L g1036 ( 
.A1(n_889),
.A2(n_429),
.A3(n_404),
.B1(n_401),
.B2(n_455),
.B3(n_465),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_886),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_861),
.A2(n_793),
.B(n_607),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_912),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_SL g1040 ( 
.A(n_917),
.B(n_308),
.Y(n_1040)
);

BUFx2_ASAP7_75t_L g1041 ( 
.A(n_917),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_893),
.B(n_837),
.Y(n_1042)
);

NOR3xp33_ASAP7_75t_L g1043 ( 
.A(n_919),
.B(n_624),
.C(n_401),
.Y(n_1043)
);

AOI22xp5_ASAP7_75t_L g1044 ( 
.A1(n_896),
.A2(n_608),
.B1(n_607),
.B2(n_601),
.Y(n_1044)
);

INVxp67_ASAP7_75t_L g1045 ( 
.A(n_921),
.Y(n_1045)
);

OAI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_951),
.A2(n_608),
.B1(n_607),
.B2(n_601),
.Y(n_1046)
);

AOI22xp33_ASAP7_75t_L g1047 ( 
.A1(n_988),
.A2(n_324),
.B1(n_280),
.B2(n_513),
.Y(n_1047)
);

HB1xp67_ASAP7_75t_L g1048 ( 
.A(n_827),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_895),
.Y(n_1049)
);

BUFx3_ASAP7_75t_L g1050 ( 
.A(n_819),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_936),
.B(n_452),
.Y(n_1051)
);

AO22x1_ASAP7_75t_L g1052 ( 
.A1(n_890),
.A2(n_404),
.B1(n_324),
.B2(n_465),
.Y(n_1052)
);

A2O1A1Ixp33_ASAP7_75t_SL g1053 ( 
.A1(n_835),
.A2(n_479),
.B(n_452),
.C(n_455),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_874),
.A2(n_608),
.B(n_607),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_877),
.A2(n_493),
.B(n_579),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_983),
.B(n_479),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_885),
.A2(n_493),
.B(n_579),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_889),
.B(n_474),
.Y(n_1058)
);

NOR2xp33_ASAP7_75t_L g1059 ( 
.A(n_949),
.B(n_1),
.Y(n_1059)
);

A2O1A1Ixp33_ASAP7_75t_L g1060 ( 
.A1(n_902),
.A2(n_513),
.B(n_481),
.C(n_474),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_965),
.Y(n_1061)
);

BUFx6f_ASAP7_75t_L g1062 ( 
.A(n_943),
.Y(n_1062)
);

NOR2xp33_ASAP7_75t_L g1063 ( 
.A(n_868),
.B(n_3),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_899),
.B(n_513),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_841),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_SL g1066 ( 
.A(n_890),
.B(n_534),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_903),
.Y(n_1067)
);

OR2x2_ASAP7_75t_L g1068 ( 
.A(n_957),
.B(n_481),
.Y(n_1068)
);

AND2x2_ASAP7_75t_L g1069 ( 
.A(n_827),
.B(n_484),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_SL g1070 ( 
.A(n_890),
.B(n_534),
.Y(n_1070)
);

BUFx12f_ASAP7_75t_L g1071 ( 
.A(n_928),
.Y(n_1071)
);

INVx5_ASAP7_75t_L g1072 ( 
.A(n_951),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_841),
.Y(n_1073)
);

BUFx12f_ASAP7_75t_L g1074 ( 
.A(n_821),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_867),
.A2(n_638),
.B(n_534),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_L g1076 ( 
.A(n_907),
.B(n_4),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_911),
.B(n_922),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_L g1078 ( 
.A(n_913),
.B(n_7),
.Y(n_1078)
);

O2A1O1Ixp33_ASAP7_75t_L g1079 ( 
.A1(n_869),
.A2(n_484),
.B(n_505),
.C(n_509),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_SL g1080 ( 
.A(n_973),
.B(n_534),
.Y(n_1080)
);

A2O1A1Ixp33_ASAP7_75t_L g1081 ( 
.A1(n_953),
.A2(n_511),
.B(n_509),
.C(n_505),
.Y(n_1081)
);

O2A1O1Ixp33_ASAP7_75t_L g1082 ( 
.A1(n_869),
.A2(n_505),
.B(n_509),
.C(n_511),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_916),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_965),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_867),
.A2(n_638),
.B(n_511),
.Y(n_1085)
);

INVx3_ASAP7_75t_L g1086 ( 
.A(n_922),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_852),
.B(n_511),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_SL g1088 ( 
.A(n_973),
.B(n_506),
.Y(n_1088)
);

NOR2xp33_ASAP7_75t_L g1089 ( 
.A(n_913),
.B(n_9),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_851),
.A2(n_986),
.B(n_985),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_956),
.B(n_924),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_971),
.Y(n_1092)
);

OAI21xp33_ASAP7_75t_L g1093 ( 
.A1(n_856),
.A2(n_509),
.B(n_505),
.Y(n_1093)
);

BUFx6f_ASAP7_75t_SL g1094 ( 
.A(n_945),
.Y(n_1094)
);

AND2x2_ASAP7_75t_L g1095 ( 
.A(n_910),
.B(n_506),
.Y(n_1095)
);

BUFx4f_ASAP7_75t_L g1096 ( 
.A(n_943),
.Y(n_1096)
);

BUFx2_ASAP7_75t_L g1097 ( 
.A(n_910),
.Y(n_1097)
);

A2O1A1Ixp33_ASAP7_75t_L g1098 ( 
.A1(n_982),
.A2(n_506),
.B(n_11),
.C(n_13),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_971),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_925),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_831),
.Y(n_1101)
);

BUFx8_ASAP7_75t_L g1102 ( 
.A(n_906),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_926),
.Y(n_1103)
);

OAI22xp5_ASAP7_75t_L g1104 ( 
.A1(n_887),
.A2(n_506),
.B1(n_74),
.B2(n_79),
.Y(n_1104)
);

OR2x6_ASAP7_75t_SL g1105 ( 
.A(n_918),
.B(n_9),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_SL g1106 ( 
.A(n_920),
.B(n_506),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_857),
.Y(n_1107)
);

NOR2xp33_ASAP7_75t_L g1108 ( 
.A(n_862),
.B(n_13),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_931),
.B(n_506),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_985),
.A2(n_506),
.B(n_84),
.Y(n_1110)
);

NOR2xp67_ASAP7_75t_L g1111 ( 
.A(n_821),
.B(n_69),
.Y(n_1111)
);

OAI21x1_ASAP7_75t_L g1112 ( 
.A1(n_939),
.A2(n_85),
.B(n_169),
.Y(n_1112)
);

AOI22xp33_ASAP7_75t_L g1113 ( 
.A1(n_982),
.A2(n_17),
.B1(n_23),
.B2(n_25),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_932),
.B(n_23),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_853),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_923),
.Y(n_1116)
);

AND2x2_ASAP7_75t_L g1117 ( 
.A(n_853),
.B(n_27),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_934),
.B(n_29),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_929),
.Y(n_1119)
);

OAI22xp5_ASAP7_75t_L g1120 ( 
.A1(n_897),
.A2(n_95),
.B1(n_158),
.B2(n_156),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_986),
.A2(n_55),
.B(n_154),
.Y(n_1121)
);

NOR2xp33_ASAP7_75t_SL g1122 ( 
.A(n_844),
.B(n_171),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_947),
.B(n_29),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_960),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_871),
.B(n_30),
.Y(n_1125)
);

OAI21xp33_ASAP7_75t_L g1126 ( 
.A1(n_872),
.A2(n_30),
.B(n_31),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_SL g1127 ( 
.A(n_844),
.B(n_86),
.Y(n_1127)
);

INVx3_ASAP7_75t_L g1128 ( 
.A(n_854),
.Y(n_1128)
);

O2A1O1Ixp33_ASAP7_75t_L g1129 ( 
.A1(n_961),
.A2(n_32),
.B(n_35),
.C(n_37),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_915),
.A2(n_107),
.B(n_151),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_963),
.Y(n_1131)
);

INVx4_ASAP7_75t_L g1132 ( 
.A(n_844),
.Y(n_1132)
);

O2A1O1Ixp33_ASAP7_75t_L g1133 ( 
.A1(n_871),
.A2(n_41),
.B(n_42),
.C(n_44),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_878),
.B(n_45),
.Y(n_1134)
);

OAI21x1_ASAP7_75t_L g1135 ( 
.A1(n_948),
.A2(n_116),
.B(n_141),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_SL g1136 ( 
.A(n_987),
.B(n_113),
.Y(n_1136)
);

AOI21x1_ASAP7_75t_L g1137 ( 
.A1(n_993),
.A2(n_989),
.B(n_909),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_997),
.B(n_872),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_994),
.B(n_880),
.Y(n_1139)
);

BUFx3_ASAP7_75t_L g1140 ( 
.A(n_995),
.Y(n_1140)
);

INVx1_ASAP7_75t_SL g1141 ( 
.A(n_1028),
.Y(n_1141)
);

OAI21x1_ASAP7_75t_L g1142 ( 
.A1(n_1054),
.A2(n_948),
.B(n_914),
.Y(n_1142)
);

BUFx3_ASAP7_75t_L g1143 ( 
.A(n_990),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_1004),
.B(n_1091),
.Y(n_1144)
);

BUFx3_ASAP7_75t_L g1145 ( 
.A(n_1050),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_1039),
.Y(n_1146)
);

OAI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_1006),
.A2(n_933),
.B(n_937),
.Y(n_1147)
);

OAI22xp5_ASAP7_75t_L g1148 ( 
.A1(n_1015),
.A2(n_987),
.B1(n_850),
.B2(n_865),
.Y(n_1148)
);

NOR4xp25_ASAP7_75t_L g1149 ( 
.A(n_1133),
.B(n_944),
.C(n_959),
.D(n_972),
.Y(n_1149)
);

INVx1_ASAP7_75t_SL g1150 ( 
.A(n_1020),
.Y(n_1150)
);

AND2x2_ASAP7_75t_L g1151 ( 
.A(n_1048),
.B(n_888),
.Y(n_1151)
);

AOI22xp5_ASAP7_75t_L g1152 ( 
.A1(n_1126),
.A2(n_888),
.B1(n_975),
.B2(n_891),
.Y(n_1152)
);

AND2x2_ASAP7_75t_SL g1153 ( 
.A(n_1113),
.B(n_987),
.Y(n_1153)
);

CKINVDCx20_ASAP7_75t_R g1154 ( 
.A(n_1023),
.Y(n_1154)
);

NOR2xp67_ASAP7_75t_SL g1155 ( 
.A(n_1017),
.B(n_980),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1016),
.B(n_883),
.Y(n_1156)
);

NOR2xp33_ASAP7_75t_L g1157 ( 
.A(n_1020),
.B(n_1048),
.Y(n_1157)
);

BUFx2_ASAP7_75t_L g1158 ( 
.A(n_1041),
.Y(n_1158)
);

BUFx6f_ASAP7_75t_L g1159 ( 
.A(n_992),
.Y(n_1159)
);

AO21x2_ASAP7_75t_L g1160 ( 
.A1(n_1043),
.A2(n_984),
.B(n_823),
.Y(n_1160)
);

BUFx6f_ASAP7_75t_L g1161 ( 
.A(n_992),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1005),
.B(n_882),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1068),
.B(n_882),
.Y(n_1163)
);

AND2x2_ASAP7_75t_L g1164 ( 
.A(n_1031),
.B(n_975),
.Y(n_1164)
);

AO21x2_ASAP7_75t_L g1165 ( 
.A1(n_1043),
.A2(n_966),
.B(n_946),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1009),
.A2(n_966),
.B(n_938),
.Y(n_1166)
);

OR2x2_ASAP7_75t_L g1167 ( 
.A(n_1035),
.B(n_891),
.Y(n_1167)
);

OAI22xp5_ASAP7_75t_L g1168 ( 
.A1(n_1042),
.A2(n_1032),
.B1(n_1037),
.B2(n_1083),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_SL g1169 ( 
.A(n_1097),
.B(n_940),
.Y(n_1169)
);

OR2x6_ASAP7_75t_L g1170 ( 
.A(n_1074),
.B(n_943),
.Y(n_1170)
);

NOR2xp33_ASAP7_75t_L g1171 ( 
.A(n_1045),
.B(n_891),
.Y(n_1171)
);

OAI21xp5_ASAP7_75t_SL g1172 ( 
.A1(n_1113),
.A2(n_970),
.B(n_979),
.Y(n_1172)
);

OAI22xp5_ASAP7_75t_L g1173 ( 
.A1(n_1049),
.A2(n_952),
.B1(n_820),
.B2(n_854),
.Y(n_1173)
);

INVx3_ASAP7_75t_L g1174 ( 
.A(n_1072),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_1009),
.A2(n_879),
.B(n_848),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1069),
.B(n_975),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_1021),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_999),
.A2(n_1077),
.B(n_1038),
.Y(n_1178)
);

BUFx8_ASAP7_75t_L g1179 ( 
.A(n_1094),
.Y(n_1179)
);

AO31x2_ASAP7_75t_L g1180 ( 
.A1(n_1110),
.A2(n_964),
.A3(n_968),
.B(n_967),
.Y(n_1180)
);

OAI22xp5_ASAP7_75t_L g1181 ( 
.A1(n_1067),
.A2(n_952),
.B1(n_860),
.B2(n_839),
.Y(n_1181)
);

BUFx3_ASAP7_75t_L g1182 ( 
.A(n_1000),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1100),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1103),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1038),
.A2(n_901),
.B(n_892),
.Y(n_1185)
);

AND3x2_ASAP7_75t_L g1186 ( 
.A(n_1122),
.B(n_1078),
.C(n_1063),
.Y(n_1186)
);

OA22x2_ASAP7_75t_L g1187 ( 
.A1(n_1030),
.A2(n_875),
.B1(n_828),
.B2(n_935),
.Y(n_1187)
);

NAND3x1_ASAP7_75t_L g1188 ( 
.A(n_1108),
.B(n_46),
.C(n_47),
.Y(n_1188)
);

AOI22xp5_ASAP7_75t_L g1189 ( 
.A1(n_1001),
.A2(n_1089),
.B1(n_1059),
.B2(n_1115),
.Y(n_1189)
);

OAI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1014),
.A2(n_954),
.B(n_955),
.Y(n_1190)
);

NOR2xp33_ASAP7_75t_L g1191 ( 
.A(n_1045),
.B(n_50),
.Y(n_1191)
);

OAI22xp5_ASAP7_75t_L g1192 ( 
.A1(n_1072),
.A2(n_103),
.B1(n_130),
.B2(n_136),
.Y(n_1192)
);

OAI21x1_ASAP7_75t_L g1193 ( 
.A1(n_1025),
.A2(n_137),
.B(n_153),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_1072),
.A2(n_1055),
.B(n_1057),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1064),
.B(n_1125),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1058),
.B(n_1051),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1134),
.B(n_1010),
.Y(n_1197)
);

O2A1O1Ixp5_ASAP7_75t_SL g1198 ( 
.A1(n_996),
.A2(n_1106),
.B(n_1104),
.C(n_1136),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1124),
.B(n_1131),
.Y(n_1199)
);

CKINVDCx20_ASAP7_75t_R g1200 ( 
.A(n_1022),
.Y(n_1200)
);

A2O1A1Ixp33_ASAP7_75t_L g1201 ( 
.A1(n_1060),
.A2(n_1118),
.B(n_1114),
.C(n_1123),
.Y(n_1201)
);

INVx2_ASAP7_75t_SL g1202 ( 
.A(n_1102),
.Y(n_1202)
);

AOI221x1_ASAP7_75t_L g1203 ( 
.A1(n_1110),
.A2(n_1098),
.B1(n_1121),
.B2(n_1130),
.C(n_1055),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1057),
.A2(n_1033),
.B(n_1046),
.Y(n_1204)
);

OR2x2_ASAP7_75t_L g1205 ( 
.A(n_1012),
.B(n_1116),
.Y(n_1205)
);

A2O1A1Ixp33_ASAP7_75t_L g1206 ( 
.A1(n_1036),
.A2(n_1130),
.B(n_1129),
.C(n_1121),
.Y(n_1206)
);

INVx2_ASAP7_75t_SL g1207 ( 
.A(n_1102),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_SL g1208 ( 
.A(n_1002),
.B(n_1047),
.Y(n_1208)
);

BUFx10_ASAP7_75t_L g1209 ( 
.A(n_1094),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1047),
.B(n_1095),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1075),
.A2(n_1085),
.B(n_1088),
.Y(n_1211)
);

BUFx2_ASAP7_75t_L g1212 ( 
.A(n_1065),
.Y(n_1212)
);

BUFx2_ASAP7_75t_SL g1213 ( 
.A(n_1018),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1034),
.B(n_1027),
.Y(n_1214)
);

NAND3x1_ASAP7_75t_L g1215 ( 
.A(n_1076),
.B(n_1059),
.C(n_1117),
.Y(n_1215)
);

AOI22xp5_ASAP7_75t_L g1216 ( 
.A1(n_1040),
.A2(n_1007),
.B1(n_1026),
.B2(n_1119),
.Y(n_1216)
);

OAI21xp33_ASAP7_75t_L g1217 ( 
.A1(n_1133),
.A2(n_1129),
.B(n_1056),
.Y(n_1217)
);

BUFx10_ASAP7_75t_L g1218 ( 
.A(n_1073),
.Y(n_1218)
);

OA21x2_ASAP7_75t_L g1219 ( 
.A1(n_1085),
.A2(n_1135),
.B(n_1112),
.Y(n_1219)
);

BUFx8_ASAP7_75t_SL g1220 ( 
.A(n_1071),
.Y(n_1220)
);

AO21x2_ASAP7_75t_L g1221 ( 
.A1(n_1053),
.A2(n_1075),
.B(n_1079),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1061),
.B(n_1099),
.Y(n_1222)
);

AOI21x1_ASAP7_75t_L g1223 ( 
.A1(n_1109),
.A2(n_1087),
.B(n_1080),
.Y(n_1223)
);

NOR2xp33_ASAP7_75t_R g1224 ( 
.A(n_1096),
.B(n_1062),
.Y(n_1224)
);

OAI21x1_ASAP7_75t_L g1225 ( 
.A1(n_1082),
.A2(n_1079),
.B(n_1044),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_SL g1226 ( 
.A(n_1096),
.B(n_1084),
.Y(n_1226)
);

AO22x2_ASAP7_75t_L g1227 ( 
.A1(n_1120),
.A2(n_1127),
.B1(n_1092),
.B2(n_1107),
.Y(n_1227)
);

A2O1A1Ixp33_ASAP7_75t_L g1228 ( 
.A1(n_1093),
.A2(n_1101),
.B(n_998),
.C(n_1003),
.Y(n_1228)
);

AND2x2_ASAP7_75t_L g1229 ( 
.A(n_1105),
.B(n_1012),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1086),
.A2(n_1082),
.B(n_1066),
.Y(n_1230)
);

AO31x2_ASAP7_75t_L g1231 ( 
.A1(n_1081),
.A2(n_991),
.A3(n_1011),
.B(n_1132),
.Y(n_1231)
);

OAI21x1_ASAP7_75t_L g1232 ( 
.A1(n_1128),
.A2(n_1070),
.B(n_1111),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1128),
.A2(n_1052),
.B(n_1132),
.Y(n_1233)
);

OAI21x1_ASAP7_75t_L g1234 ( 
.A1(n_1019),
.A2(n_1029),
.B(n_1008),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1019),
.B(n_1029),
.Y(n_1235)
);

AO32x2_ASAP7_75t_L g1236 ( 
.A1(n_1024),
.A2(n_807),
.A3(n_999),
.B1(n_681),
.B2(n_881),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_997),
.B(n_540),
.Y(n_1237)
);

OAI21x1_ASAP7_75t_L g1238 ( 
.A1(n_1054),
.A2(n_1038),
.B(n_1025),
.Y(n_1238)
);

AOI21x1_ASAP7_75t_L g1239 ( 
.A1(n_993),
.A2(n_1038),
.B(n_1090),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_997),
.B(n_540),
.Y(n_1240)
);

INVx5_ASAP7_75t_L g1241 ( 
.A(n_1018),
.Y(n_1241)
);

AO21x2_ASAP7_75t_L g1242 ( 
.A1(n_993),
.A2(n_1090),
.B(n_1043),
.Y(n_1242)
);

AOI22xp5_ASAP7_75t_L g1243 ( 
.A1(n_997),
.A2(n_962),
.B1(n_950),
.B2(n_873),
.Y(n_1243)
);

NAND3xp33_ASAP7_75t_SL g1244 ( 
.A(n_1015),
.B(n_950),
.C(n_568),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_997),
.B(n_540),
.Y(n_1245)
);

AOI21x1_ASAP7_75t_L g1246 ( 
.A1(n_993),
.A2(n_1038),
.B(n_1090),
.Y(n_1246)
);

AND2x4_ASAP7_75t_L g1247 ( 
.A(n_1062),
.B(n_945),
.Y(n_1247)
);

A2O1A1Ixp33_ASAP7_75t_L g1248 ( 
.A1(n_1001),
.A2(n_950),
.B(n_962),
.C(n_734),
.Y(n_1248)
);

BUFx6f_ASAP7_75t_L g1249 ( 
.A(n_992),
.Y(n_1249)
);

AND2x2_ASAP7_75t_L g1250 ( 
.A(n_997),
.B(n_520),
.Y(n_1250)
);

INVx5_ASAP7_75t_L g1251 ( 
.A(n_1018),
.Y(n_1251)
);

NAND3x1_ASAP7_75t_L g1252 ( 
.A(n_1108),
.B(n_677),
.C(n_1063),
.Y(n_1252)
);

O2A1O1Ixp33_ASAP7_75t_L g1253 ( 
.A1(n_997),
.A2(n_950),
.B(n_962),
.C(n_976),
.Y(n_1253)
);

OAI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_993),
.A2(n_976),
.B(n_950),
.Y(n_1254)
);

OA21x2_ASAP7_75t_L g1255 ( 
.A1(n_993),
.A2(n_1090),
.B(n_1038),
.Y(n_1255)
);

CKINVDCx6p67_ASAP7_75t_R g1256 ( 
.A(n_1029),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1037),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1037),
.Y(n_1258)
);

AOI221x1_ASAP7_75t_L g1259 ( 
.A1(n_993),
.A2(n_962),
.B1(n_950),
.B2(n_1043),
.C(n_1110),
.Y(n_1259)
);

AOI21xp5_ASAP7_75t_SL g1260 ( 
.A1(n_1013),
.A2(n_690),
.B(n_900),
.Y(n_1260)
);

BUFx3_ASAP7_75t_L g1261 ( 
.A(n_995),
.Y(n_1261)
);

BUFx6f_ASAP7_75t_L g1262 ( 
.A(n_992),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_997),
.B(n_540),
.Y(n_1263)
);

BUFx2_ASAP7_75t_L g1264 ( 
.A(n_995),
.Y(n_1264)
);

AOI21xp33_ASAP7_75t_L g1265 ( 
.A1(n_1001),
.A2(n_950),
.B(n_962),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_997),
.B(n_540),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_997),
.B(n_540),
.Y(n_1267)
);

INVx2_ASAP7_75t_L g1268 ( 
.A(n_1039),
.Y(n_1268)
);

AOI221xp5_ASAP7_75t_SL g1269 ( 
.A1(n_1113),
.A2(n_962),
.B1(n_733),
.B2(n_1129),
.C(n_1126),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_997),
.B(n_540),
.Y(n_1270)
);

AOI211x1_ASAP7_75t_L g1271 ( 
.A1(n_1126),
.A2(n_733),
.B(n_873),
.C(n_978),
.Y(n_1271)
);

OAI22x1_ASAP7_75t_L g1272 ( 
.A1(n_1015),
.A2(n_962),
.B1(n_1078),
.B2(n_1063),
.Y(n_1272)
);

A2O1A1Ixp33_ASAP7_75t_L g1273 ( 
.A1(n_1001),
.A2(n_950),
.B(n_962),
.C(n_734),
.Y(n_1273)
);

AND2x4_ASAP7_75t_L g1274 ( 
.A(n_1062),
.B(n_945),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_997),
.B(n_540),
.Y(n_1275)
);

NAND3x1_ASAP7_75t_L g1276 ( 
.A(n_1108),
.B(n_677),
.C(n_1063),
.Y(n_1276)
);

OR2x2_ASAP7_75t_L g1277 ( 
.A(n_1138),
.B(n_1139),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1263),
.B(n_1266),
.Y(n_1278)
);

BUFx6f_ASAP7_75t_L g1279 ( 
.A(n_1159),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1267),
.B(n_1270),
.Y(n_1280)
);

AND2x2_ASAP7_75t_L g1281 ( 
.A(n_1250),
.B(n_1151),
.Y(n_1281)
);

NOR2x1_ASAP7_75t_R g1282 ( 
.A(n_1145),
.B(n_1143),
.Y(n_1282)
);

OAI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1248),
.A2(n_1273),
.B(n_1265),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1199),
.Y(n_1284)
);

A2O1A1Ixp33_ASAP7_75t_L g1285 ( 
.A1(n_1253),
.A2(n_1243),
.B(n_1172),
.C(n_1275),
.Y(n_1285)
);

AND2x2_ASAP7_75t_L g1286 ( 
.A(n_1164),
.B(n_1272),
.Y(n_1286)
);

OAI22xp5_ASAP7_75t_L g1287 ( 
.A1(n_1243),
.A2(n_1153),
.B1(n_1189),
.B2(n_1144),
.Y(n_1287)
);

BUFx6f_ASAP7_75t_L g1288 ( 
.A(n_1159),
.Y(n_1288)
);

CKINVDCx20_ASAP7_75t_R g1289 ( 
.A(n_1154),
.Y(n_1289)
);

OAI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1254),
.A2(n_1201),
.B(n_1259),
.Y(n_1290)
);

BUFx3_ASAP7_75t_L g1291 ( 
.A(n_1159),
.Y(n_1291)
);

BUFx2_ASAP7_75t_L g1292 ( 
.A(n_1140),
.Y(n_1292)
);

AO31x2_ASAP7_75t_L g1293 ( 
.A1(n_1203),
.A2(n_1204),
.A3(n_1211),
.B(n_1206),
.Y(n_1293)
);

AND2x4_ASAP7_75t_L g1294 ( 
.A(n_1247),
.B(n_1274),
.Y(n_1294)
);

AO32x2_ASAP7_75t_L g1295 ( 
.A1(n_1168),
.A2(n_1148),
.A3(n_1181),
.B1(n_1173),
.B2(n_1269),
.Y(n_1295)
);

AND2x2_ASAP7_75t_SL g1296 ( 
.A(n_1149),
.B(n_1269),
.Y(n_1296)
);

OA21x2_ASAP7_75t_L g1297 ( 
.A1(n_1225),
.A2(n_1238),
.B(n_1178),
.Y(n_1297)
);

AOI22x1_ASAP7_75t_L g1298 ( 
.A1(n_1227),
.A2(n_1233),
.B1(n_1175),
.B2(n_1185),
.Y(n_1298)
);

OR2x2_ASAP7_75t_L g1299 ( 
.A(n_1141),
.B(n_1176),
.Y(n_1299)
);

BUFx2_ASAP7_75t_SL g1300 ( 
.A(n_1161),
.Y(n_1300)
);

AOI22xp33_ASAP7_75t_L g1301 ( 
.A1(n_1244),
.A2(n_1217),
.B1(n_1208),
.B2(n_1186),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1184),
.Y(n_1302)
);

AOI22xp33_ASAP7_75t_L g1303 ( 
.A1(n_1217),
.A2(n_1187),
.B1(n_1189),
.B2(n_1197),
.Y(n_1303)
);

OAI22xp33_ASAP7_75t_L g1304 ( 
.A1(n_1172),
.A2(n_1152),
.B1(n_1163),
.B2(n_1196),
.Y(n_1304)
);

INVx3_ASAP7_75t_L g1305 ( 
.A(n_1161),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1257),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1258),
.Y(n_1307)
);

NAND3xp33_ASAP7_75t_L g1308 ( 
.A(n_1271),
.B(n_1156),
.C(n_1152),
.Y(n_1308)
);

OAI21x1_ASAP7_75t_L g1309 ( 
.A1(n_1142),
.A2(n_1137),
.B(n_1239),
.Y(n_1309)
);

OAI21xp5_ASAP7_75t_L g1310 ( 
.A1(n_1198),
.A2(n_1149),
.B(n_1195),
.Y(n_1310)
);

AOI22xp5_ASAP7_75t_L g1311 ( 
.A1(n_1252),
.A2(n_1276),
.B1(n_1215),
.B2(n_1229),
.Y(n_1311)
);

OAI21x1_ASAP7_75t_L g1312 ( 
.A1(n_1246),
.A2(n_1166),
.B(n_1193),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1214),
.Y(n_1313)
);

OA21x2_ASAP7_75t_L g1314 ( 
.A1(n_1147),
.A2(n_1190),
.B(n_1230),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1146),
.Y(n_1315)
);

OA21x2_ASAP7_75t_L g1316 ( 
.A1(n_1223),
.A2(n_1228),
.B(n_1210),
.Y(n_1316)
);

AOI22xp5_ASAP7_75t_L g1317 ( 
.A1(n_1169),
.A2(n_1155),
.B1(n_1171),
.B2(n_1188),
.Y(n_1317)
);

BUFx6f_ASAP7_75t_L g1318 ( 
.A(n_1161),
.Y(n_1318)
);

AOI22xp33_ASAP7_75t_L g1319 ( 
.A1(n_1191),
.A2(n_1162),
.B1(n_1268),
.B2(n_1177),
.Y(n_1319)
);

AOI21xp33_ASAP7_75t_L g1320 ( 
.A1(n_1227),
.A2(n_1160),
.B(n_1216),
.Y(n_1320)
);

INVx2_ASAP7_75t_L g1321 ( 
.A(n_1180),
.Y(n_1321)
);

OAI21x1_ASAP7_75t_L g1322 ( 
.A1(n_1232),
.A2(n_1219),
.B(n_1255),
.Y(n_1322)
);

AOI22xp33_ASAP7_75t_L g1323 ( 
.A1(n_1150),
.A2(n_1167),
.B1(n_1242),
.B2(n_1157),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1150),
.B(n_1158),
.Y(n_1324)
);

OAI21xp5_ASAP7_75t_L g1325 ( 
.A1(n_1205),
.A2(n_1226),
.B(n_1222),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1264),
.B(n_1261),
.Y(n_1326)
);

INVxp67_ASAP7_75t_SL g1327 ( 
.A(n_1249),
.Y(n_1327)
);

INVx4_ASAP7_75t_L g1328 ( 
.A(n_1249),
.Y(n_1328)
);

AOI22xp33_ASAP7_75t_L g1329 ( 
.A1(n_1160),
.A2(n_1192),
.B1(n_1165),
.B2(n_1236),
.Y(n_1329)
);

O2A1O1Ixp33_ASAP7_75t_L g1330 ( 
.A1(n_1202),
.A2(n_1207),
.B(n_1235),
.C(n_1221),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1231),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1231),
.Y(n_1332)
);

OAI221xp5_ASAP7_75t_L g1333 ( 
.A1(n_1170),
.A2(n_1212),
.B1(n_1182),
.B2(n_1249),
.C(n_1262),
.Y(n_1333)
);

OAI21xp5_ASAP7_75t_L g1334 ( 
.A1(n_1234),
.A2(n_1236),
.B(n_1251),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_1221),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_1220),
.Y(n_1336)
);

INVx1_ASAP7_75t_SL g1337 ( 
.A(n_1256),
.Y(n_1337)
);

CKINVDCx5p33_ASAP7_75t_R g1338 ( 
.A(n_1200),
.Y(n_1338)
);

INVxp67_ASAP7_75t_SL g1339 ( 
.A(n_1262),
.Y(n_1339)
);

OAI21x1_ASAP7_75t_L g1340 ( 
.A1(n_1224),
.A2(n_1170),
.B(n_1241),
.Y(n_1340)
);

AND2x4_ASAP7_75t_L g1341 ( 
.A(n_1170),
.B(n_1251),
.Y(n_1341)
);

A2O1A1Ixp33_ASAP7_75t_L g1342 ( 
.A1(n_1213),
.A2(n_1209),
.B(n_1179),
.C(n_1218),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1209),
.Y(n_1343)
);

AO21x2_ASAP7_75t_L g1344 ( 
.A1(n_1218),
.A2(n_1194),
.B(n_1204),
.Y(n_1344)
);

AOI22xp33_ASAP7_75t_L g1345 ( 
.A1(n_1265),
.A2(n_962),
.B1(n_1272),
.B2(n_1243),
.Y(n_1345)
);

OR2x2_ASAP7_75t_L g1346 ( 
.A(n_1138),
.B(n_1139),
.Y(n_1346)
);

NAND2xp33_ASAP7_75t_SL g1347 ( 
.A(n_1224),
.B(n_1113),
.Y(n_1347)
);

AOI22xp33_ASAP7_75t_L g1348 ( 
.A1(n_1265),
.A2(n_962),
.B1(n_1272),
.B2(n_1243),
.Y(n_1348)
);

AO21x2_ASAP7_75t_L g1349 ( 
.A1(n_1194),
.A2(n_1204),
.B(n_1211),
.Y(n_1349)
);

NOR2xp33_ASAP7_75t_L g1350 ( 
.A(n_1243),
.B(n_1237),
.Y(n_1350)
);

OAI21x1_ASAP7_75t_SL g1351 ( 
.A1(n_1233),
.A2(n_1129),
.B(n_1197),
.Y(n_1351)
);

CKINVDCx5p33_ASAP7_75t_R g1352 ( 
.A(n_1154),
.Y(n_1352)
);

AND2x4_ASAP7_75t_L g1353 ( 
.A(n_1247),
.B(n_1274),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1183),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_1183),
.Y(n_1355)
);

BUFx3_ASAP7_75t_L g1356 ( 
.A(n_1145),
.Y(n_1356)
);

OAI21xp5_ASAP7_75t_L g1357 ( 
.A1(n_1248),
.A2(n_1273),
.B(n_1265),
.Y(n_1357)
);

BUFx2_ASAP7_75t_L g1358 ( 
.A(n_1140),
.Y(n_1358)
);

AOI21xp5_ASAP7_75t_L g1359 ( 
.A1(n_1248),
.A2(n_1273),
.B(n_1260),
.Y(n_1359)
);

NOR2xp33_ASAP7_75t_L g1360 ( 
.A(n_1243),
.B(n_1237),
.Y(n_1360)
);

BUFx12f_ASAP7_75t_L g1361 ( 
.A(n_1179),
.Y(n_1361)
);

BUFx2_ASAP7_75t_L g1362 ( 
.A(n_1140),
.Y(n_1362)
);

AND2x4_ASAP7_75t_L g1363 ( 
.A(n_1247),
.B(n_1274),
.Y(n_1363)
);

NAND3xp33_ASAP7_75t_L g1364 ( 
.A(n_1243),
.B(n_1273),
.C(n_1248),
.Y(n_1364)
);

AO31x2_ASAP7_75t_L g1365 ( 
.A1(n_1203),
.A2(n_1259),
.A3(n_1204),
.B(n_1194),
.Y(n_1365)
);

BUFx4f_ASAP7_75t_SL g1366 ( 
.A(n_1179),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1250),
.B(n_1151),
.Y(n_1367)
);

AO31x2_ASAP7_75t_L g1368 ( 
.A1(n_1203),
.A2(n_1259),
.A3(n_1204),
.B(n_1194),
.Y(n_1368)
);

INVx3_ASAP7_75t_L g1369 ( 
.A(n_1174),
.Y(n_1369)
);

NAND3xp33_ASAP7_75t_L g1370 ( 
.A(n_1243),
.B(n_1273),
.C(n_1248),
.Y(n_1370)
);

AND2x4_ASAP7_75t_L g1371 ( 
.A(n_1247),
.B(n_1274),
.Y(n_1371)
);

OA21x2_ASAP7_75t_L g1372 ( 
.A1(n_1203),
.A2(n_1259),
.B(n_1204),
.Y(n_1372)
);

OAI22xp5_ASAP7_75t_L g1373 ( 
.A1(n_1243),
.A2(n_1237),
.B1(n_1245),
.B2(n_1240),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1237),
.B(n_1240),
.Y(n_1374)
);

INVx4_ASAP7_75t_L g1375 ( 
.A(n_1159),
.Y(n_1375)
);

BUFx2_ASAP7_75t_L g1376 ( 
.A(n_1140),
.Y(n_1376)
);

NAND2xp33_ASAP7_75t_SL g1377 ( 
.A(n_1224),
.B(n_1113),
.Y(n_1377)
);

NOR2xp33_ASAP7_75t_L g1378 ( 
.A(n_1243),
.B(n_1237),
.Y(n_1378)
);

INVx3_ASAP7_75t_L g1379 ( 
.A(n_1174),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1237),
.B(n_1240),
.Y(n_1380)
);

OA21x2_ASAP7_75t_L g1381 ( 
.A1(n_1203),
.A2(n_1259),
.B(n_1204),
.Y(n_1381)
);

O2A1O1Ixp33_ASAP7_75t_L g1382 ( 
.A1(n_1248),
.A2(n_1273),
.B(n_1265),
.C(n_1253),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1183),
.Y(n_1383)
);

OAI222xp33_ASAP7_75t_L g1384 ( 
.A1(n_1243),
.A2(n_1113),
.B1(n_733),
.B2(n_962),
.C1(n_1240),
.C2(n_1237),
.Y(n_1384)
);

NOR2xp67_ASAP7_75t_L g1385 ( 
.A(n_1343),
.B(n_1315),
.Y(n_1385)
);

OAI22xp5_ASAP7_75t_L g1386 ( 
.A1(n_1345),
.A2(n_1348),
.B1(n_1364),
.B2(n_1370),
.Y(n_1386)
);

INVx6_ASAP7_75t_L g1387 ( 
.A(n_1328),
.Y(n_1387)
);

OAI22xp5_ASAP7_75t_SL g1388 ( 
.A1(n_1311),
.A2(n_1301),
.B1(n_1360),
.B2(n_1378),
.Y(n_1388)
);

OR2x2_ASAP7_75t_L g1389 ( 
.A(n_1299),
.B(n_1277),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1373),
.B(n_1350),
.Y(n_1390)
);

OAI22xp5_ASAP7_75t_L g1391 ( 
.A1(n_1345),
.A2(n_1348),
.B1(n_1378),
.B2(n_1360),
.Y(n_1391)
);

OA21x2_ASAP7_75t_L g1392 ( 
.A1(n_1290),
.A2(n_1320),
.B(n_1359),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1350),
.B(n_1285),
.Y(n_1393)
);

CKINVDCx5p33_ASAP7_75t_R g1394 ( 
.A(n_1352),
.Y(n_1394)
);

CKINVDCx20_ASAP7_75t_R g1395 ( 
.A(n_1289),
.Y(n_1395)
);

OA22x2_ASAP7_75t_L g1396 ( 
.A1(n_1317),
.A2(n_1334),
.B1(n_1357),
.B2(n_1283),
.Y(n_1396)
);

OAI22xp5_ASAP7_75t_L g1397 ( 
.A1(n_1303),
.A2(n_1301),
.B1(n_1287),
.B2(n_1285),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1304),
.B(n_1346),
.Y(n_1398)
);

O2A1O1Ixp5_ASAP7_75t_L g1399 ( 
.A1(n_1384),
.A2(n_1310),
.B(n_1347),
.C(n_1377),
.Y(n_1399)
);

O2A1O1Ixp5_ASAP7_75t_L g1400 ( 
.A1(n_1384),
.A2(n_1347),
.B(n_1377),
.C(n_1304),
.Y(n_1400)
);

BUFx6f_ASAP7_75t_L g1401 ( 
.A(n_1356),
.Y(n_1401)
);

AOI221x1_ASAP7_75t_SL g1402 ( 
.A1(n_1278),
.A2(n_1380),
.B1(n_1280),
.B2(n_1374),
.C(n_1308),
.Y(n_1402)
);

O2A1O1Ixp33_ASAP7_75t_L g1403 ( 
.A1(n_1330),
.A2(n_1351),
.B(n_1303),
.C(n_1333),
.Y(n_1403)
);

OA22x2_ASAP7_75t_L g1404 ( 
.A1(n_1325),
.A2(n_1284),
.B1(n_1286),
.B2(n_1313),
.Y(n_1404)
);

AOI21xp5_ASAP7_75t_SL g1405 ( 
.A1(n_1342),
.A2(n_1330),
.B(n_1341),
.Y(n_1405)
);

AOI21xp5_ASAP7_75t_SL g1406 ( 
.A1(n_1342),
.A2(n_1327),
.B(n_1339),
.Y(n_1406)
);

AOI21xp5_ASAP7_75t_SL g1407 ( 
.A1(n_1282),
.A2(n_1314),
.B(n_1371),
.Y(n_1407)
);

AOI21xp5_ASAP7_75t_SL g1408 ( 
.A1(n_1294),
.A2(n_1353),
.B(n_1371),
.Y(n_1408)
);

O2A1O1Ixp33_ASAP7_75t_L g1409 ( 
.A1(n_1326),
.A2(n_1319),
.B(n_1306),
.C(n_1302),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1319),
.B(n_1307),
.Y(n_1410)
);

OAI22xp5_ASAP7_75t_L g1411 ( 
.A1(n_1296),
.A2(n_1329),
.B1(n_1323),
.B2(n_1355),
.Y(n_1411)
);

O2A1O1Ixp33_ASAP7_75t_L g1412 ( 
.A1(n_1305),
.A2(n_1329),
.B(n_1344),
.C(n_1383),
.Y(n_1412)
);

OAI22xp5_ASAP7_75t_L g1413 ( 
.A1(n_1296),
.A2(n_1323),
.B1(n_1354),
.B2(n_1383),
.Y(n_1413)
);

OA21x2_ASAP7_75t_L g1414 ( 
.A1(n_1309),
.A2(n_1322),
.B(n_1312),
.Y(n_1414)
);

O2A1O1Ixp5_ASAP7_75t_L g1415 ( 
.A1(n_1335),
.A2(n_1321),
.B(n_1332),
.C(n_1331),
.Y(n_1415)
);

AOI21xp5_ASAP7_75t_SL g1416 ( 
.A1(n_1363),
.A2(n_1344),
.B(n_1291),
.Y(n_1416)
);

BUFx3_ASAP7_75t_L g1417 ( 
.A(n_1292),
.Y(n_1417)
);

NOR2x1_ASAP7_75t_SL g1418 ( 
.A(n_1331),
.B(n_1349),
.Y(n_1418)
);

BUFx3_ASAP7_75t_L g1419 ( 
.A(n_1358),
.Y(n_1419)
);

O2A1O1Ixp33_ASAP7_75t_L g1420 ( 
.A1(n_1305),
.A2(n_1337),
.B(n_1362),
.C(n_1376),
.Y(n_1420)
);

AND2x4_ASAP7_75t_L g1421 ( 
.A(n_1340),
.B(n_1369),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1372),
.B(n_1381),
.Y(n_1422)
);

AOI221xp5_ASAP7_75t_L g1423 ( 
.A1(n_1295),
.A2(n_1375),
.B1(n_1300),
.B2(n_1379),
.C(n_1288),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1316),
.Y(n_1424)
);

OAI22xp5_ASAP7_75t_SL g1425 ( 
.A1(n_1366),
.A2(n_1289),
.B1(n_1361),
.B2(n_1338),
.Y(n_1425)
);

AND2x4_ASAP7_75t_L g1426 ( 
.A(n_1375),
.B(n_1279),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1316),
.B(n_1293),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1318),
.B(n_1293),
.Y(n_1428)
);

OAI22xp5_ASAP7_75t_L g1429 ( 
.A1(n_1318),
.A2(n_1298),
.B1(n_1295),
.B2(n_1336),
.Y(n_1429)
);

OAI22xp5_ASAP7_75t_SL g1430 ( 
.A1(n_1297),
.A2(n_1293),
.B1(n_1368),
.B2(n_1365),
.Y(n_1430)
);

OR2x2_ASAP7_75t_L g1431 ( 
.A(n_1293),
.B(n_1368),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1365),
.B(n_1368),
.Y(n_1432)
);

CKINVDCx9p33_ASAP7_75t_R g1433 ( 
.A(n_1292),
.Y(n_1433)
);

OAI22xp5_ASAP7_75t_L g1434 ( 
.A1(n_1345),
.A2(n_1113),
.B1(n_1153),
.B2(n_1243),
.Y(n_1434)
);

OAI22xp5_ASAP7_75t_L g1435 ( 
.A1(n_1345),
.A2(n_1113),
.B1(n_1153),
.B2(n_1243),
.Y(n_1435)
);

O2A1O1Ixp33_ASAP7_75t_L g1436 ( 
.A1(n_1384),
.A2(n_1273),
.B(n_1248),
.C(n_1253),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1373),
.B(n_1350),
.Y(n_1437)
);

OA21x2_ASAP7_75t_L g1438 ( 
.A1(n_1290),
.A2(n_1203),
.B(n_1259),
.Y(n_1438)
);

OR2x2_ASAP7_75t_L g1439 ( 
.A(n_1299),
.B(n_1277),
.Y(n_1439)
);

NOR2xp67_ASAP7_75t_L g1440 ( 
.A(n_1343),
.B(n_1235),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1281),
.B(n_1367),
.Y(n_1441)
);

OAI22xp5_ASAP7_75t_L g1442 ( 
.A1(n_1345),
.A2(n_1113),
.B1(n_1153),
.B2(n_1243),
.Y(n_1442)
);

OA21x2_ASAP7_75t_L g1443 ( 
.A1(n_1290),
.A2(n_1203),
.B(n_1259),
.Y(n_1443)
);

AOI221x1_ASAP7_75t_SL g1444 ( 
.A1(n_1373),
.A2(n_733),
.B1(n_1089),
.B2(n_1078),
.C(n_1063),
.Y(n_1444)
);

BUFx6f_ASAP7_75t_L g1445 ( 
.A(n_1356),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1281),
.B(n_1367),
.Y(n_1446)
);

BUFx2_ASAP7_75t_L g1447 ( 
.A(n_1324),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1281),
.B(n_1367),
.Y(n_1448)
);

OAI22xp5_ASAP7_75t_L g1449 ( 
.A1(n_1345),
.A2(n_1113),
.B1(n_1153),
.B2(n_1243),
.Y(n_1449)
);

O2A1O1Ixp33_ASAP7_75t_L g1450 ( 
.A1(n_1384),
.A2(n_1273),
.B(n_1248),
.C(n_1253),
.Y(n_1450)
);

AOI21xp5_ASAP7_75t_SL g1451 ( 
.A1(n_1382),
.A2(n_1273),
.B(n_1248),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1424),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1432),
.B(n_1431),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1415),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1438),
.B(n_1443),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1438),
.B(n_1443),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1390),
.B(n_1437),
.Y(n_1457)
);

CKINVDCx5p33_ASAP7_75t_R g1458 ( 
.A(n_1395),
.Y(n_1458)
);

OR2x2_ASAP7_75t_L g1459 ( 
.A(n_1427),
.B(n_1422),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1418),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1392),
.B(n_1428),
.Y(n_1461)
);

INVx1_ASAP7_75t_SL g1462 ( 
.A(n_1389),
.Y(n_1462)
);

NOR2xp33_ASAP7_75t_L g1463 ( 
.A(n_1388),
.B(n_1393),
.Y(n_1463)
);

OR2x2_ASAP7_75t_L g1464 ( 
.A(n_1430),
.B(n_1392),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1411),
.B(n_1413),
.Y(n_1465)
);

OR2x2_ASAP7_75t_L g1466 ( 
.A(n_1413),
.B(n_1411),
.Y(n_1466)
);

AO21x2_ASAP7_75t_L g1467 ( 
.A1(n_1451),
.A2(n_1391),
.B(n_1435),
.Y(n_1467)
);

OAI21xp5_ASAP7_75t_L g1468 ( 
.A1(n_1436),
.A2(n_1450),
.B(n_1400),
.Y(n_1468)
);

AO21x2_ASAP7_75t_L g1469 ( 
.A1(n_1391),
.A2(n_1434),
.B(n_1435),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1414),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1396),
.B(n_1404),
.Y(n_1471)
);

OR2x2_ASAP7_75t_L g1472 ( 
.A(n_1398),
.B(n_1439),
.Y(n_1472)
);

INVxp67_ASAP7_75t_L g1473 ( 
.A(n_1404),
.Y(n_1473)
);

AO21x2_ASAP7_75t_L g1474 ( 
.A1(n_1434),
.A2(n_1442),
.B(n_1449),
.Y(n_1474)
);

INVx3_ASAP7_75t_L g1475 ( 
.A(n_1421),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1398),
.B(n_1386),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1396),
.B(n_1429),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1399),
.B(n_1423),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1421),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1410),
.Y(n_1480)
);

HB1xp67_ASAP7_75t_L g1481 ( 
.A(n_1385),
.Y(n_1481)
);

AO21x2_ASAP7_75t_L g1482 ( 
.A1(n_1442),
.A2(n_1449),
.B(n_1412),
.Y(n_1482)
);

AO21x2_ASAP7_75t_L g1483 ( 
.A1(n_1397),
.A2(n_1403),
.B(n_1409),
.Y(n_1483)
);

AO21x2_ASAP7_75t_L g1484 ( 
.A1(n_1397),
.A2(n_1416),
.B(n_1405),
.Y(n_1484)
);

AOI22xp33_ASAP7_75t_L g1485 ( 
.A1(n_1444),
.A2(n_1447),
.B1(n_1448),
.B2(n_1446),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1407),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1402),
.Y(n_1487)
);

BUFx2_ASAP7_75t_L g1488 ( 
.A(n_1433),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1455),
.B(n_1441),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1480),
.B(n_1420),
.Y(n_1490)
);

AOI22xp33_ASAP7_75t_SL g1491 ( 
.A1(n_1467),
.A2(n_1417),
.B1(n_1419),
.B2(n_1425),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1480),
.B(n_1440),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1452),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1455),
.B(n_1456),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1452),
.Y(n_1495)
);

INVx2_ASAP7_75t_SL g1496 ( 
.A(n_1475),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1472),
.B(n_1406),
.Y(n_1497)
);

INVxp67_ASAP7_75t_L g1498 ( 
.A(n_1481),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1456),
.B(n_1445),
.Y(n_1499)
);

AOI22xp33_ASAP7_75t_L g1500 ( 
.A1(n_1467),
.A2(n_1469),
.B1(n_1474),
.B2(n_1463),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1461),
.B(n_1453),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1470),
.Y(n_1502)
);

AND2x4_ASAP7_75t_L g1503 ( 
.A(n_1479),
.B(n_1426),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1472),
.B(n_1401),
.Y(n_1504)
);

CKINVDCx6p67_ASAP7_75t_R g1505 ( 
.A(n_1488),
.Y(n_1505)
);

BUFx2_ASAP7_75t_L g1506 ( 
.A(n_1460),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1470),
.Y(n_1507)
);

AOI33xp33_ASAP7_75t_L g1508 ( 
.A1(n_1487),
.A2(n_1477),
.A3(n_1478),
.B1(n_1485),
.B2(n_1465),
.B3(n_1471),
.Y(n_1508)
);

OR2x2_ASAP7_75t_L g1509 ( 
.A(n_1459),
.B(n_1408),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1493),
.Y(n_1510)
);

AND2x2_ASAP7_75t_SL g1511 ( 
.A(n_1500),
.B(n_1465),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1501),
.B(n_1475),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1492),
.B(n_1462),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1493),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1501),
.B(n_1475),
.Y(n_1515)
);

AOI22xp33_ASAP7_75t_L g1516 ( 
.A1(n_1500),
.A2(n_1467),
.B1(n_1469),
.B2(n_1474),
.Y(n_1516)
);

AO21x2_ASAP7_75t_L g1517 ( 
.A1(n_1502),
.A2(n_1454),
.B(n_1460),
.Y(n_1517)
);

OR2x6_ASAP7_75t_L g1518 ( 
.A(n_1509),
.B(n_1486),
.Y(n_1518)
);

AOI22xp33_ASAP7_75t_L g1519 ( 
.A1(n_1491),
.A2(n_1467),
.B1(n_1469),
.B2(n_1474),
.Y(n_1519)
);

CKINVDCx8_ASAP7_75t_R g1520 ( 
.A(n_1503),
.Y(n_1520)
);

AOI22xp33_ASAP7_75t_L g1521 ( 
.A1(n_1491),
.A2(n_1469),
.B1(n_1474),
.B2(n_1482),
.Y(n_1521)
);

INVx1_ASAP7_75t_SL g1522 ( 
.A(n_1499),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1492),
.B(n_1462),
.Y(n_1523)
);

NOR2xp33_ASAP7_75t_R g1524 ( 
.A(n_1505),
.B(n_1458),
.Y(n_1524)
);

OR2x2_ASAP7_75t_L g1525 ( 
.A(n_1494),
.B(n_1464),
.Y(n_1525)
);

AND2x4_ASAP7_75t_L g1526 ( 
.A(n_1496),
.B(n_1475),
.Y(n_1526)
);

AOI221xp5_ASAP7_75t_SL g1527 ( 
.A1(n_1497),
.A2(n_1463),
.B1(n_1487),
.B2(n_1468),
.C(n_1477),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1493),
.Y(n_1528)
);

AOI22xp33_ASAP7_75t_SL g1529 ( 
.A1(n_1497),
.A2(n_1484),
.B1(n_1469),
.B2(n_1474),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1504),
.B(n_1472),
.Y(n_1530)
);

AOI21xp5_ASAP7_75t_L g1531 ( 
.A1(n_1490),
.A2(n_1484),
.B(n_1468),
.Y(n_1531)
);

INVx3_ASAP7_75t_L g1532 ( 
.A(n_1502),
.Y(n_1532)
);

OAI31xp33_ASAP7_75t_SL g1533 ( 
.A1(n_1508),
.A2(n_1477),
.A3(n_1465),
.B(n_1478),
.Y(n_1533)
);

NOR2x2_ASAP7_75t_L g1534 ( 
.A(n_1505),
.B(n_1486),
.Y(n_1534)
);

AOI22xp33_ASAP7_75t_L g1535 ( 
.A1(n_1509),
.A2(n_1482),
.B1(n_1483),
.B2(n_1484),
.Y(n_1535)
);

BUFx3_ASAP7_75t_L g1536 ( 
.A(n_1505),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1495),
.Y(n_1537)
);

AOI22xp33_ASAP7_75t_L g1538 ( 
.A1(n_1509),
.A2(n_1482),
.B1(n_1483),
.B2(n_1484),
.Y(n_1538)
);

OR2x2_ASAP7_75t_L g1539 ( 
.A(n_1494),
.B(n_1464),
.Y(n_1539)
);

OR2x2_ASAP7_75t_L g1540 ( 
.A(n_1494),
.B(n_1464),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1495),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1510),
.Y(n_1542)
);

OAI21xp5_ASAP7_75t_L g1543 ( 
.A1(n_1531),
.A2(n_1476),
.B(n_1478),
.Y(n_1543)
);

OR2x2_ASAP7_75t_L g1544 ( 
.A(n_1525),
.B(n_1494),
.Y(n_1544)
);

AND2x4_ASAP7_75t_SL g1545 ( 
.A(n_1518),
.B(n_1505),
.Y(n_1545)
);

OA21x2_ASAP7_75t_L g1546 ( 
.A1(n_1521),
.A2(n_1507),
.B(n_1506),
.Y(n_1546)
);

HB1xp67_ASAP7_75t_L g1547 ( 
.A(n_1510),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1514),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1530),
.B(n_1489),
.Y(n_1549)
);

OAI21xp5_ASAP7_75t_L g1550 ( 
.A1(n_1519),
.A2(n_1476),
.B(n_1471),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_SL g1551 ( 
.A(n_1533),
.B(n_1488),
.Y(n_1551)
);

HB1xp67_ASAP7_75t_L g1552 ( 
.A(n_1514),
.Y(n_1552)
);

INVx3_ASAP7_75t_L g1553 ( 
.A(n_1520),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1528),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1528),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1537),
.Y(n_1556)
);

INVxp67_ASAP7_75t_L g1557 ( 
.A(n_1513),
.Y(n_1557)
);

INVx4_ASAP7_75t_SL g1558 ( 
.A(n_1536),
.Y(n_1558)
);

INVxp67_ASAP7_75t_SL g1559 ( 
.A(n_1532),
.Y(n_1559)
);

BUFx6f_ASAP7_75t_L g1560 ( 
.A(n_1536),
.Y(n_1560)
);

BUFx2_ASAP7_75t_L g1561 ( 
.A(n_1534),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1517),
.Y(n_1562)
);

AND2x6_ASAP7_75t_SL g1563 ( 
.A(n_1523),
.B(n_1457),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1541),
.Y(n_1564)
);

HB1xp67_ASAP7_75t_L g1565 ( 
.A(n_1525),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1547),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1547),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1557),
.B(n_1543),
.Y(n_1568)
);

BUFx2_ASAP7_75t_L g1569 ( 
.A(n_1561),
.Y(n_1569)
);

AND2x4_ASAP7_75t_L g1570 ( 
.A(n_1558),
.B(n_1518),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1552),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1561),
.B(n_1518),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1562),
.Y(n_1573)
);

HB1xp67_ASAP7_75t_L g1574 ( 
.A(n_1565),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1562),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1552),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1561),
.B(n_1518),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1542),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1557),
.B(n_1527),
.Y(n_1579)
);

HB1xp67_ASAP7_75t_L g1580 ( 
.A(n_1565),
.Y(n_1580)
);

HB1xp67_ASAP7_75t_L g1581 ( 
.A(n_1551),
.Y(n_1581)
);

OR2x2_ASAP7_75t_L g1582 ( 
.A(n_1544),
.B(n_1539),
.Y(n_1582)
);

AOI211xp5_ASAP7_75t_L g1583 ( 
.A1(n_1543),
.A2(n_1533),
.B(n_1527),
.C(n_1487),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1542),
.Y(n_1584)
);

AOI221xp5_ASAP7_75t_SL g1585 ( 
.A1(n_1551),
.A2(n_1516),
.B1(n_1538),
.B2(n_1535),
.C(n_1473),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1553),
.B(n_1518),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1563),
.B(n_1548),
.Y(n_1587)
);

BUFx2_ASAP7_75t_L g1588 ( 
.A(n_1553),
.Y(n_1588)
);

INVx2_ASAP7_75t_L g1589 ( 
.A(n_1562),
.Y(n_1589)
);

CKINVDCx16_ASAP7_75t_R g1590 ( 
.A(n_1550),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1548),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1562),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1553),
.B(n_1512),
.Y(n_1593)
);

AND2x4_ASAP7_75t_L g1594 ( 
.A(n_1558),
.B(n_1536),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1554),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1554),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1563),
.B(n_1489),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1553),
.B(n_1558),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1558),
.B(n_1515),
.Y(n_1599)
);

AND2x4_ASAP7_75t_L g1600 ( 
.A(n_1558),
.B(n_1526),
.Y(n_1600)
);

INVx2_ASAP7_75t_SL g1601 ( 
.A(n_1545),
.Y(n_1601)
);

NAND4xp25_ASAP7_75t_L g1602 ( 
.A(n_1550),
.B(n_1529),
.C(n_1508),
.D(n_1457),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1558),
.B(n_1515),
.Y(n_1603)
);

NAND2x1_ASAP7_75t_SL g1604 ( 
.A(n_1546),
.B(n_1526),
.Y(n_1604)
);

HB1xp67_ASAP7_75t_L g1605 ( 
.A(n_1555),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_SL g1606 ( 
.A(n_1590),
.B(n_1524),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1605),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1605),
.Y(n_1608)
);

OR2x2_ASAP7_75t_L g1609 ( 
.A(n_1568),
.B(n_1549),
.Y(n_1609)
);

AOI32xp33_ASAP7_75t_L g1610 ( 
.A1(n_1583),
.A2(n_1545),
.A3(n_1471),
.B1(n_1488),
.B2(n_1522),
.Y(n_1610)
);

INVx3_ASAP7_75t_L g1611 ( 
.A(n_1570),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1583),
.B(n_1511),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1578),
.Y(n_1613)
);

OR2x2_ASAP7_75t_L g1614 ( 
.A(n_1568),
.B(n_1549),
.Y(n_1614)
);

OR2x2_ASAP7_75t_L g1615 ( 
.A(n_1569),
.B(n_1544),
.Y(n_1615)
);

OR2x6_ASAP7_75t_L g1616 ( 
.A(n_1569),
.B(n_1560),
.Y(n_1616)
);

HB1xp67_ASAP7_75t_L g1617 ( 
.A(n_1574),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1598),
.B(n_1560),
.Y(n_1618)
);

OAI22xp5_ASAP7_75t_L g1619 ( 
.A1(n_1590),
.A2(n_1511),
.B1(n_1466),
.B2(n_1520),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1578),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1584),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1588),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1584),
.Y(n_1623)
);

NOR5xp2_ASAP7_75t_L g1624 ( 
.A(n_1581),
.B(n_1498),
.C(n_1559),
.D(n_1564),
.E(n_1556),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1591),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1591),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1595),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1595),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1598),
.B(n_1560),
.Y(n_1629)
);

AND2x4_ASAP7_75t_L g1630 ( 
.A(n_1594),
.B(n_1545),
.Y(n_1630)
);

OR2x2_ASAP7_75t_L g1631 ( 
.A(n_1579),
.B(n_1540),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1579),
.B(n_1511),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1596),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1594),
.B(n_1599),
.Y(n_1634)
);

INVx2_ASAP7_75t_SL g1635 ( 
.A(n_1600),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1596),
.Y(n_1636)
);

HB1xp67_ASAP7_75t_L g1637 ( 
.A(n_1580),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1566),
.Y(n_1638)
);

OAI21xp33_ASAP7_75t_L g1639 ( 
.A1(n_1602),
.A2(n_1490),
.B(n_1466),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1585),
.B(n_1489),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1570),
.B(n_1545),
.Y(n_1641)
);

CKINVDCx16_ASAP7_75t_R g1642 ( 
.A(n_1616),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1617),
.Y(n_1643)
);

INVx1_ASAP7_75t_SL g1644 ( 
.A(n_1634),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1618),
.B(n_1588),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1617),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1616),
.Y(n_1647)
);

INVx2_ASAP7_75t_L g1648 ( 
.A(n_1616),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1639),
.B(n_1587),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1615),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1637),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1637),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1613),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1629),
.B(n_1594),
.Y(n_1654)
);

NAND3xp33_ASAP7_75t_L g1655 ( 
.A(n_1612),
.B(n_1585),
.C(n_1602),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1620),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1632),
.B(n_1587),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1635),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1635),
.B(n_1594),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1611),
.B(n_1601),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1621),
.Y(n_1661)
);

BUFx12f_ASAP7_75t_L g1662 ( 
.A(n_1630),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1623),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1622),
.Y(n_1664)
);

INVx1_ASAP7_75t_SL g1665 ( 
.A(n_1606),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1625),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1626),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1660),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1643),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1643),
.Y(n_1670)
);

O2A1O1Ixp33_ASAP7_75t_SL g1671 ( 
.A1(n_1655),
.A2(n_1606),
.B(n_1601),
.C(n_1622),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1646),
.B(n_1607),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1646),
.Y(n_1673)
);

OR2x2_ASAP7_75t_L g1674 ( 
.A(n_1650),
.B(n_1609),
.Y(n_1674)
);

AOI221xp5_ASAP7_75t_SL g1675 ( 
.A1(n_1649),
.A2(n_1619),
.B1(n_1640),
.B2(n_1577),
.C(n_1572),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1651),
.Y(n_1676)
);

INVxp67_ASAP7_75t_L g1677 ( 
.A(n_1645),
.Y(n_1677)
);

OAI32xp33_ASAP7_75t_L g1678 ( 
.A1(n_1642),
.A2(n_1611),
.A3(n_1631),
.B1(n_1608),
.B2(n_1624),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1654),
.B(n_1630),
.Y(n_1679)
);

OR2x2_ASAP7_75t_L g1680 ( 
.A(n_1650),
.B(n_1614),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1651),
.Y(n_1681)
);

AOI221x1_ASAP7_75t_L g1682 ( 
.A1(n_1652),
.A2(n_1638),
.B1(n_1611),
.B2(n_1566),
.C(n_1571),
.Y(n_1682)
);

AOI22xp5_ASAP7_75t_L g1683 ( 
.A1(n_1665),
.A2(n_1630),
.B1(n_1641),
.B2(n_1601),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1652),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1664),
.B(n_1657),
.Y(n_1685)
);

AOI22xp5_ASAP7_75t_L g1686 ( 
.A1(n_1662),
.A2(n_1641),
.B1(n_1577),
.B2(n_1572),
.Y(n_1686)
);

AOI31xp33_ASAP7_75t_L g1687 ( 
.A1(n_1644),
.A2(n_1458),
.A3(n_1394),
.B(n_1570),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1669),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1670),
.Y(n_1689)
);

INVx1_ASAP7_75t_SL g1690 ( 
.A(n_1679),
.Y(n_1690)
);

HB1xp67_ASAP7_75t_L g1691 ( 
.A(n_1677),
.Y(n_1691)
);

INVx2_ASAP7_75t_L g1692 ( 
.A(n_1668),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1673),
.Y(n_1693)
);

NOR2xp33_ASAP7_75t_L g1694 ( 
.A(n_1687),
.B(n_1662),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1683),
.B(n_1645),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1686),
.B(n_1654),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1676),
.Y(n_1697)
);

AOI22xp5_ASAP7_75t_L g1698 ( 
.A1(n_1675),
.A2(n_1642),
.B1(n_1659),
.B2(n_1660),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1681),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1674),
.B(n_1659),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1700),
.Y(n_1701)
);

AOI221xp5_ASAP7_75t_L g1702 ( 
.A1(n_1695),
.A2(n_1678),
.B1(n_1671),
.B2(n_1687),
.C(n_1685),
.Y(n_1702)
);

OAI221xp5_ASAP7_75t_SL g1703 ( 
.A1(n_1698),
.A2(n_1610),
.B1(n_1680),
.B2(n_1685),
.C(n_1672),
.Y(n_1703)
);

O2A1O1Ixp33_ASAP7_75t_L g1704 ( 
.A1(n_1691),
.A2(n_1672),
.B(n_1684),
.C(n_1648),
.Y(n_1704)
);

OAI221xp5_ASAP7_75t_L g1705 ( 
.A1(n_1694),
.A2(n_1648),
.B1(n_1647),
.B2(n_1664),
.C(n_1666),
.Y(n_1705)
);

NAND4xp75_ASAP7_75t_L g1706 ( 
.A(n_1694),
.B(n_1682),
.C(n_1647),
.D(n_1658),
.Y(n_1706)
);

AOI221xp5_ASAP7_75t_SL g1707 ( 
.A1(n_1690),
.A2(n_1658),
.B1(n_1667),
.B2(n_1663),
.C(n_1656),
.Y(n_1707)
);

INVx1_ASAP7_75t_SL g1708 ( 
.A(n_1700),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1692),
.Y(n_1709)
);

NAND4xp25_ASAP7_75t_SL g1710 ( 
.A(n_1696),
.B(n_1586),
.C(n_1667),
.D(n_1666),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_SL g1711 ( 
.A(n_1696),
.B(n_1570),
.Y(n_1711)
);

AOI22xp5_ASAP7_75t_L g1712 ( 
.A1(n_1702),
.A2(n_1692),
.B1(n_1697),
.B2(n_1693),
.Y(n_1712)
);

XNOR2x1_ASAP7_75t_L g1713 ( 
.A(n_1706),
.B(n_1688),
.Y(n_1713)
);

OAI21xp33_ASAP7_75t_SL g1714 ( 
.A1(n_1708),
.A2(n_1604),
.B(n_1689),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1701),
.B(n_1699),
.Y(n_1715)
);

OAI21xp33_ASAP7_75t_SL g1716 ( 
.A1(n_1711),
.A2(n_1604),
.B(n_1663),
.Y(n_1716)
);

OAI22xp5_ASAP7_75t_L g1717 ( 
.A1(n_1703),
.A2(n_1600),
.B1(n_1597),
.B2(n_1560),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1713),
.B(n_1709),
.Y(n_1718)
);

XOR2x2_ASAP7_75t_L g1719 ( 
.A(n_1717),
.B(n_1705),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1712),
.B(n_1707),
.Y(n_1720)
);

NOR2x1_ASAP7_75t_L g1721 ( 
.A(n_1715),
.B(n_1705),
.Y(n_1721)
);

OR2x2_ASAP7_75t_L g1722 ( 
.A(n_1714),
.B(n_1710),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1716),
.B(n_1704),
.Y(n_1723)
);

NOR2x1_ASAP7_75t_L g1724 ( 
.A(n_1713),
.B(n_1653),
.Y(n_1724)
);

NOR2xp67_ASAP7_75t_L g1725 ( 
.A(n_1722),
.B(n_1718),
.Y(n_1725)
);

O2A1O1Ixp5_ASAP7_75t_SL g1726 ( 
.A1(n_1723),
.A2(n_1661),
.B(n_1656),
.C(n_1653),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1720),
.B(n_1661),
.Y(n_1727)
);

AOI322xp5_ASAP7_75t_L g1728 ( 
.A1(n_1721),
.A2(n_1636),
.A3(n_1633),
.B1(n_1628),
.B2(n_1627),
.C1(n_1597),
.C2(n_1567),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1724),
.B(n_1593),
.Y(n_1729)
);

OR3x1_ASAP7_75t_L g1730 ( 
.A(n_1725),
.B(n_1719),
.C(n_1571),
.Y(n_1730)
);

NOR2xp33_ASAP7_75t_SL g1731 ( 
.A(n_1729),
.B(n_1560),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1727),
.Y(n_1732)
);

XNOR2x1_ASAP7_75t_L g1733 ( 
.A(n_1732),
.B(n_1726),
.Y(n_1733)
);

AOI22xp33_ASAP7_75t_L g1734 ( 
.A1(n_1733),
.A2(n_1731),
.B1(n_1730),
.B2(n_1560),
.Y(n_1734)
);

XNOR2xp5_ASAP7_75t_L g1735 ( 
.A(n_1734),
.B(n_1728),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1734),
.B(n_1593),
.Y(n_1736)
);

OAI22xp5_ASAP7_75t_L g1737 ( 
.A1(n_1735),
.A2(n_1736),
.B1(n_1567),
.B2(n_1576),
.Y(n_1737)
);

XNOR2xp5_ASAP7_75t_L g1738 ( 
.A(n_1735),
.B(n_1586),
.Y(n_1738)
);

OAI22xp5_ASAP7_75t_SL g1739 ( 
.A1(n_1738),
.A2(n_1576),
.B1(n_1600),
.B2(n_1560),
.Y(n_1739)
);

OAI22x1_ASAP7_75t_L g1740 ( 
.A1(n_1737),
.A2(n_1600),
.B1(n_1589),
.B2(n_1575),
.Y(n_1740)
);

AOI21x1_ASAP7_75t_L g1741 ( 
.A1(n_1740),
.A2(n_1575),
.B(n_1573),
.Y(n_1741)
);

OAI22xp5_ASAP7_75t_L g1742 ( 
.A1(n_1741),
.A2(n_1739),
.B1(n_1589),
.B2(n_1573),
.Y(n_1742)
);

OAI21xp5_ASAP7_75t_L g1743 ( 
.A1(n_1742),
.A2(n_1575),
.B(n_1573),
.Y(n_1743)
);

OR2x6_ASAP7_75t_L g1744 ( 
.A(n_1743),
.B(n_1387),
.Y(n_1744)
);

OAI22xp5_ASAP7_75t_L g1745 ( 
.A1(n_1744),
.A2(n_1592),
.B1(n_1589),
.B2(n_1582),
.Y(n_1745)
);

AOI211xp5_ASAP7_75t_L g1746 ( 
.A1(n_1745),
.A2(n_1592),
.B(n_1560),
.C(n_1603),
.Y(n_1746)
);


endmodule