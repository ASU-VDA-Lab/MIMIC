module fake_jpeg_31779_n_140 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_140);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_140;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_2),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_30),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_3),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

BUFx10_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_9),
.Y(n_46)
);

INVx6_ASAP7_75t_SL g47 ( 
.A(n_22),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_6),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_15),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

CKINVDCx14_ASAP7_75t_R g52 ( 
.A(n_4),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_16),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_54),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

BUFx16f_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

CKINVDCx6p67_ASAP7_75t_R g68 ( 
.A(n_57),
.Y(n_68)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_44),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_62),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

A2O1A1Ixp33_ASAP7_75t_L g63 ( 
.A1(n_57),
.A2(n_40),
.B(n_43),
.C(n_48),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_63),
.A2(n_51),
.B(n_47),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_58),
.B(n_42),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_50),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_52),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_70),
.B(n_73),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_60),
.B(n_52),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_72),
.B(n_74),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_53),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_44),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_69),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_77),
.B(n_79),
.Y(n_97)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_78),
.B(n_85),
.Y(n_95)
);

CKINVDCx14_ASAP7_75t_R g79 ( 
.A(n_68),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_80),
.B(n_2),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_49),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_81),
.B(n_88),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_71),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_82),
.B(n_83),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_45),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_67),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_84),
.B(n_86),
.Y(n_110)
);

INVx13_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_75),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_87),
.B(n_1),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_64),
.B(n_0),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_72),
.A2(n_46),
.B(n_41),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_89),
.A2(n_0),
.B(n_1),
.Y(n_93)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_90),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_93),
.B(n_94),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_81),
.Y(n_94)
);

OAI21xp33_ASAP7_75t_L g113 ( 
.A1(n_98),
.A2(n_8),
.B(n_10),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_99),
.B(n_105),
.Y(n_121)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_76),
.Y(n_100)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_100),
.Y(n_114)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_79),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_101),
.B(n_109),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_80),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_102),
.B(n_104),
.C(n_7),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_76),
.B(n_4),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_81),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_81),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_106),
.B(n_107),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_77),
.B(n_36),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_76),
.B(n_5),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_108),
.B(n_18),
.Y(n_122)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_81),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_112),
.B(n_115),
.Y(n_126)
);

NAND3xp33_ASAP7_75t_L g125 ( 
.A(n_113),
.B(n_120),
.C(n_122),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_110),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_103),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_116)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_116),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_97),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_117),
.B(n_118),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_97),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_96),
.B(n_14),
.Y(n_120)
);

AOI322xp5_ASAP7_75t_L g128 ( 
.A1(n_114),
.A2(n_104),
.A3(n_102),
.B1(n_95),
.B2(n_92),
.C1(n_27),
.C2(n_28),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_128),
.B(n_120),
.C(n_119),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_123),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_121),
.Y(n_130)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_130),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_125),
.B(n_111),
.Y(n_131)
);

NAND4xp25_ASAP7_75t_L g133 ( 
.A(n_131),
.B(n_132),
.C(n_125),
.D(n_126),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_133),
.A2(n_127),
.B(n_124),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_135),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_136),
.A2(n_134),
.B(n_23),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_137),
.B(n_21),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_25),
.C(n_26),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_29),
.Y(n_140)
);


endmodule