module fake_jpeg_8142_n_109 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_109);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_109;

wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_0),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_23),
.Y(n_38)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_25),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_12),
.A2(n_0),
.B(n_1),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_17),
.B(n_2),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_27),
.Y(n_34)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_28),
.B(n_29),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_11),
.B(n_2),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_27),
.A2(n_13),
.B1(n_15),
.B2(n_12),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_30),
.A2(n_31),
.B1(n_36),
.B2(n_10),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_27),
.A2(n_15),
.B1(n_12),
.B2(n_11),
.Y(n_31)
);

OAI22xp33_ASAP7_75t_L g32 ( 
.A1(n_24),
.A2(n_19),
.B1(n_16),
.B2(n_11),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_32),
.A2(n_15),
.B1(n_10),
.B2(n_25),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_25),
.A2(n_24),
.B1(n_16),
.B2(n_19),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_39),
.A2(n_17),
.B1(n_21),
.B2(n_20),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_37),
.B(n_29),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_40),
.B(n_46),
.Y(n_66)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_43),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_37),
.B(n_29),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_42),
.B(n_49),
.Y(n_58)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_28),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_SL g65 ( 
.A1(n_44),
.A2(n_50),
.B(n_52),
.Y(n_65)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_53),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_28),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_30),
.Y(n_47)
);

XOR2xp5_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_22),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_26),
.Y(n_48)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_38),
.B(n_18),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_28),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_51),
.A2(n_10),
.B1(n_21),
.B2(n_20),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_23),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx6_ASAP7_75t_SL g67 ( 
.A(n_54),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_30),
.Y(n_55)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_63),
.Y(n_73)
);

OA22x2_ASAP7_75t_L g61 ( 
.A1(n_47),
.A2(n_23),
.B1(n_22),
.B2(n_18),
.Y(n_61)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_54),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_68),
.Y(n_81)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_69),
.B(n_70),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_66),
.B(n_44),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_71),
.B(n_75),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_67),
.Y(n_72)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_72),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_56),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_70),
.B(n_44),
.C(n_46),
.Y(n_76)
);

XNOR2x1_ASAP7_75t_L g84 ( 
.A(n_76),
.B(n_80),
.Y(n_84)
);

NAND3xp33_ASAP7_75t_L g77 ( 
.A(n_59),
.B(n_40),
.C(n_6),
.Y(n_77)
);

NAND3xp33_ASAP7_75t_L g83 ( 
.A(n_77),
.B(n_6),
.C(n_7),
.Y(n_83)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

AO21x1_ASAP7_75t_L g87 ( 
.A1(n_78),
.A2(n_57),
.B(n_67),
.Y(n_87)
);

XOR2x2_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_51),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_83),
.B(n_86),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_79),
.A2(n_62),
.B1(n_61),
.B2(n_69),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_85),
.A2(n_88),
.B1(n_79),
.B2(n_73),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_81),
.Y(n_86)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_87),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_80),
.A2(n_62),
.B1(n_68),
.B2(n_63),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_84),
.B(n_76),
.C(n_71),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_92),
.B(n_94),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_93),
.B(n_95),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_84),
.B(n_65),
.C(n_74),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_89),
.B(n_74),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_91),
.A2(n_82),
.B1(n_61),
.B2(n_87),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_96),
.B(n_99),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_90),
.B(n_58),
.Y(n_99)
);

AOI31xp67_ASAP7_75t_L g100 ( 
.A1(n_98),
.A2(n_95),
.A3(n_61),
.B(n_83),
.Y(n_100)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_100),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_97),
.A2(n_52),
.B(n_7),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_101),
.B(n_103),
.C(n_3),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_97),
.A2(n_52),
.B(n_4),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_102),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_104),
.B(n_106),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_105),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_108),
.A2(n_3),
.B(n_4),
.Y(n_109)
);


endmodule