module fake_ariane_1032_n_3113 (n_295, n_356, n_556, n_170, n_190, n_698, n_695, n_160, n_64, n_180, n_730, n_119, n_124, n_386, n_307, n_516, n_589, n_332, n_581, n_294, n_646, n_197, n_640, n_463, n_830, n_176, n_691, n_34, n_404, n_172, n_678, n_651, n_347, n_423, n_183, n_469, n_479, n_726, n_603, n_373, n_299, n_836, n_541, n_499, n_789, n_788, n_12, n_850, n_771, n_564, n_133, n_610, n_66, n_205, n_752, n_341, n_71, n_109, n_245, n_421, n_96, n_549, n_522, n_319, n_49, n_591, n_760, n_20, n_690, n_416, n_283, n_50, n_187, n_525, n_806, n_367, n_713, n_649, n_598, n_345, n_374, n_318, n_817, n_103, n_244, n_643, n_679, n_226, n_781, n_220, n_261, n_682, n_36, n_663, n_370, n_706, n_189, n_717, n_819, n_72, n_286, n_443, n_586, n_57, n_686, n_605, n_776, n_424, n_528, n_584, n_387, n_406, n_826, n_117, n_139, n_524, n_85, n_130, n_349, n_391, n_634, n_466, n_756, n_346, n_214, n_764, n_348, n_552, n_2, n_462, n_607, n_670, n_32, n_410, n_379, n_445, n_515, n_807, n_138, n_162, n_765, n_264, n_737, n_137, n_122, n_198, n_232, n_52, n_441, n_568, n_385, n_637, n_73, n_327, n_77, n_766, n_372, n_377, n_15, n_396, n_802, n_631, n_23, n_399, n_554, n_520, n_87, n_714, n_279, n_702, n_207, n_790, n_363, n_720, n_354, n_41, n_813, n_140, n_725, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_633, n_154, n_338, n_142, n_285, n_473, n_186, n_801, n_202, n_145, n_193, n_733, n_761, n_818, n_500, n_665, n_59, n_336, n_731, n_754, n_779, n_315, n_594, n_311, n_239, n_402, n_35, n_272, n_54, n_829, n_8, n_668, n_339, n_738, n_758, n_833, n_672, n_487, n_740, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_648, n_784, n_269, n_597, n_816, n_75, n_158, n_69, n_259, n_835, n_95, n_808, n_446, n_553, n_143, n_753, n_566, n_814, n_578, n_701, n_625, n_152, n_405, n_557, n_120, n_169, n_106, n_173, n_242, n_645, n_309, n_320, n_115, n_331, n_559, n_401, n_485, n_267, n_495, n_504, n_647, n_483, n_335, n_435, n_350, n_291, n_822, n_344, n_381, n_795, n_426, n_433, n_481, n_600, n_721, n_840, n_398, n_62, n_210, n_200, n_529, n_502, n_166, n_253, n_561, n_770, n_218, n_821, n_79, n_839, n_3, n_271, n_465, n_486, n_507, n_759, n_247, n_569, n_567, n_825, n_732, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_787, n_31, n_547, n_420, n_562, n_518, n_439, n_604, n_614, n_677, n_222, n_478, n_703, n_748, n_786, n_510, n_831, n_256, n_326, n_681, n_778, n_227, n_48, n_188, n_323, n_550, n_635, n_707, n_330, n_400, n_689, n_694, n_11, n_129, n_126, n_282, n_328, n_368, n_590, n_699, n_727, n_277, n_248, n_301, n_467, n_432, n_545, n_536, n_644, n_293, n_823, n_620, n_228, n_325, n_276, n_93, n_688, n_636, n_427, n_108, n_587, n_497, n_693, n_303, n_671, n_442, n_777, n_168, n_81, n_1, n_206, n_352, n_538, n_576, n_843, n_511, n_611, n_238, n_365, n_429, n_455, n_654, n_588, n_638, n_136, n_334, n_192, n_729, n_661, n_488, n_775, n_667, n_300, n_533, n_505, n_14, n_163, n_88, n_141, n_846, n_390, n_498, n_104, n_501, n_438, n_314, n_684, n_16, n_440, n_627, n_273, n_305, n_539, n_312, n_233, n_56, n_60, n_728, n_388, n_333, n_449, n_612, n_413, n_392, n_376, n_512, n_715, n_579, n_844, n_459, n_685, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_623, n_838, n_237, n_780, n_175, n_711, n_453, n_734, n_74, n_491, n_810, n_19, n_40, n_181, n_723, n_616, n_617, n_658, n_630, n_705, n_570, n_53, n_260, n_362, n_543, n_310, n_709, n_236, n_601, n_683, n_565, n_281, n_24, n_7, n_628, n_809, n_461, n_209, n_262, n_490, n_743, n_17, n_225, n_235, n_660, n_464, n_735, n_575, n_546, n_297, n_662, n_641, n_503, n_700, n_290, n_527, n_46, n_741, n_747, n_772, n_84, n_847, n_371, n_845, n_199, n_107, n_639, n_217, n_452, n_673, n_676, n_178, n_42, n_551, n_308, n_708, n_417, n_201, n_70, n_572, n_343, n_10, n_414, n_571, n_680, n_287, n_302, n_380, n_6, n_582, n_94, n_284, n_4, n_448, n_593, n_755, n_710, n_249, n_534, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_609, n_278, n_851, n_255, n_560, n_450, n_257, n_842, n_148, n_652, n_451, n_613, n_745, n_475, n_135, n_409, n_171, n_519, n_384, n_468, n_853, n_61, n_526, n_716, n_102, n_742, n_182, n_696, n_674, n_482, n_316, n_196, n_125, n_798, n_769, n_820, n_43, n_577, n_407, n_774, n_13, n_27, n_254, n_596, n_476, n_460, n_219, n_832, n_55, n_535, n_231, n_366, n_744, n_762, n_656, n_555, n_234, n_492, n_574, n_848, n_804, n_280, n_215, n_252, n_629, n_664, n_161, n_454, n_298, n_532, n_68, n_415, n_794, n_763, n_78, n_63, n_655, n_99, n_540, n_216, n_544, n_692, n_5, n_599, n_768, n_514, n_418, n_537, n_223, n_403, n_25, n_750, n_834, n_83, n_389, n_800, n_657, n_513, n_837, n_288, n_179, n_812, n_395, n_621, n_195, n_606, n_213, n_110, n_304, n_659, n_67, n_509, n_583, n_724, n_306, n_666, n_313, n_92, n_430, n_626, n_493, n_722, n_203, n_378, n_436, n_150, n_98, n_757, n_375, n_113, n_114, n_33, n_324, n_585, n_669, n_785, n_827, n_619, n_337, n_437, n_111, n_21, n_274, n_622, n_697, n_472, n_296, n_265, n_746, n_208, n_456, n_156, n_292, n_793, n_852, n_174, n_275, n_100, n_704, n_132, n_147, n_204, n_751, n_615, n_521, n_51, n_496, n_739, n_76, n_342, n_26, n_246, n_517, n_530, n_0, n_792, n_824, n_428, n_159, n_358, n_105, n_580, n_608, n_30, n_494, n_719, n_131, n_263, n_434, n_360, n_563, n_229, n_394, n_250, n_773, n_165, n_144, n_317, n_101, n_243, n_803, n_134, n_329, n_718, n_185, n_340, n_749, n_289, n_9, n_112, n_45, n_542, n_548, n_815, n_523, n_268, n_266, n_470, n_457, n_164, n_157, n_632, n_184, n_177, n_477, n_364, n_258, n_650, n_782, n_425, n_431, n_811, n_508, n_624, n_118, n_121, n_791, n_618, n_411, n_484, n_712, n_849, n_353, n_22, n_736, n_767, n_241, n_29, n_357, n_412, n_687, n_447, n_191, n_382, n_797, n_489, n_80, n_480, n_211, n_642, n_97, n_408, n_828, n_595, n_322, n_251, n_506, n_602, n_799, n_558, n_592, n_116, n_397, n_841, n_471, n_351, n_39, n_393, n_474, n_653, n_359, n_155, n_573, n_796, n_805, n_127, n_531, n_783, n_675, n_3113);

input n_295;
input n_356;
input n_556;
input n_170;
input n_190;
input n_698;
input n_695;
input n_160;
input n_64;
input n_180;
input n_730;
input n_119;
input n_124;
input n_386;
input n_307;
input n_516;
input n_589;
input n_332;
input n_581;
input n_294;
input n_646;
input n_197;
input n_640;
input n_463;
input n_830;
input n_176;
input n_691;
input n_34;
input n_404;
input n_172;
input n_678;
input n_651;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_726;
input n_603;
input n_373;
input n_299;
input n_836;
input n_541;
input n_499;
input n_789;
input n_788;
input n_12;
input n_850;
input n_771;
input n_564;
input n_133;
input n_610;
input n_66;
input n_205;
input n_752;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_549;
input n_522;
input n_319;
input n_49;
input n_591;
input n_760;
input n_20;
input n_690;
input n_416;
input n_283;
input n_50;
input n_187;
input n_525;
input n_806;
input n_367;
input n_713;
input n_649;
input n_598;
input n_345;
input n_374;
input n_318;
input n_817;
input n_103;
input n_244;
input n_643;
input n_679;
input n_226;
input n_781;
input n_220;
input n_261;
input n_682;
input n_36;
input n_663;
input n_370;
input n_706;
input n_189;
input n_717;
input n_819;
input n_72;
input n_286;
input n_443;
input n_586;
input n_57;
input n_686;
input n_605;
input n_776;
input n_424;
input n_528;
input n_584;
input n_387;
input n_406;
input n_826;
input n_117;
input n_139;
input n_524;
input n_85;
input n_130;
input n_349;
input n_391;
input n_634;
input n_466;
input n_756;
input n_346;
input n_214;
input n_764;
input n_348;
input n_552;
input n_2;
input n_462;
input n_607;
input n_670;
input n_32;
input n_410;
input n_379;
input n_445;
input n_515;
input n_807;
input n_138;
input n_162;
input n_765;
input n_264;
input n_737;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_568;
input n_385;
input n_637;
input n_73;
input n_327;
input n_77;
input n_766;
input n_372;
input n_377;
input n_15;
input n_396;
input n_802;
input n_631;
input n_23;
input n_399;
input n_554;
input n_520;
input n_87;
input n_714;
input n_279;
input n_702;
input n_207;
input n_790;
input n_363;
input n_720;
input n_354;
input n_41;
input n_813;
input n_140;
input n_725;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_633;
input n_154;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_801;
input n_202;
input n_145;
input n_193;
input n_733;
input n_761;
input n_818;
input n_500;
input n_665;
input n_59;
input n_336;
input n_731;
input n_754;
input n_779;
input n_315;
input n_594;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_829;
input n_8;
input n_668;
input n_339;
input n_738;
input n_758;
input n_833;
input n_672;
input n_487;
input n_740;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_648;
input n_784;
input n_269;
input n_597;
input n_816;
input n_75;
input n_158;
input n_69;
input n_259;
input n_835;
input n_95;
input n_808;
input n_446;
input n_553;
input n_143;
input n_753;
input n_566;
input n_814;
input n_578;
input n_701;
input n_625;
input n_152;
input n_405;
input n_557;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_645;
input n_309;
input n_320;
input n_115;
input n_331;
input n_559;
input n_401;
input n_485;
input n_267;
input n_495;
input n_504;
input n_647;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_822;
input n_344;
input n_381;
input n_795;
input n_426;
input n_433;
input n_481;
input n_600;
input n_721;
input n_840;
input n_398;
input n_62;
input n_210;
input n_200;
input n_529;
input n_502;
input n_166;
input n_253;
input n_561;
input n_770;
input n_218;
input n_821;
input n_79;
input n_839;
input n_3;
input n_271;
input n_465;
input n_486;
input n_507;
input n_759;
input n_247;
input n_569;
input n_567;
input n_825;
input n_732;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_787;
input n_31;
input n_547;
input n_420;
input n_562;
input n_518;
input n_439;
input n_604;
input n_614;
input n_677;
input n_222;
input n_478;
input n_703;
input n_748;
input n_786;
input n_510;
input n_831;
input n_256;
input n_326;
input n_681;
input n_778;
input n_227;
input n_48;
input n_188;
input n_323;
input n_550;
input n_635;
input n_707;
input n_330;
input n_400;
input n_689;
input n_694;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_590;
input n_699;
input n_727;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_545;
input n_536;
input n_644;
input n_293;
input n_823;
input n_620;
input n_228;
input n_325;
input n_276;
input n_93;
input n_688;
input n_636;
input n_427;
input n_108;
input n_587;
input n_497;
input n_693;
input n_303;
input n_671;
input n_442;
input n_777;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_538;
input n_576;
input n_843;
input n_511;
input n_611;
input n_238;
input n_365;
input n_429;
input n_455;
input n_654;
input n_588;
input n_638;
input n_136;
input n_334;
input n_192;
input n_729;
input n_661;
input n_488;
input n_775;
input n_667;
input n_300;
input n_533;
input n_505;
input n_14;
input n_163;
input n_88;
input n_141;
input n_846;
input n_390;
input n_498;
input n_104;
input n_501;
input n_438;
input n_314;
input n_684;
input n_16;
input n_440;
input n_627;
input n_273;
input n_305;
input n_539;
input n_312;
input n_233;
input n_56;
input n_60;
input n_728;
input n_388;
input n_333;
input n_449;
input n_612;
input n_413;
input n_392;
input n_376;
input n_512;
input n_715;
input n_579;
input n_844;
input n_459;
input n_685;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_623;
input n_838;
input n_237;
input n_780;
input n_175;
input n_711;
input n_453;
input n_734;
input n_74;
input n_491;
input n_810;
input n_19;
input n_40;
input n_181;
input n_723;
input n_616;
input n_617;
input n_658;
input n_630;
input n_705;
input n_570;
input n_53;
input n_260;
input n_362;
input n_543;
input n_310;
input n_709;
input n_236;
input n_601;
input n_683;
input n_565;
input n_281;
input n_24;
input n_7;
input n_628;
input n_809;
input n_461;
input n_209;
input n_262;
input n_490;
input n_743;
input n_17;
input n_225;
input n_235;
input n_660;
input n_464;
input n_735;
input n_575;
input n_546;
input n_297;
input n_662;
input n_641;
input n_503;
input n_700;
input n_290;
input n_527;
input n_46;
input n_741;
input n_747;
input n_772;
input n_84;
input n_847;
input n_371;
input n_845;
input n_199;
input n_107;
input n_639;
input n_217;
input n_452;
input n_673;
input n_676;
input n_178;
input n_42;
input n_551;
input n_308;
input n_708;
input n_417;
input n_201;
input n_70;
input n_572;
input n_343;
input n_10;
input n_414;
input n_571;
input n_680;
input n_287;
input n_302;
input n_380;
input n_6;
input n_582;
input n_94;
input n_284;
input n_4;
input n_448;
input n_593;
input n_755;
input n_710;
input n_249;
input n_534;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_609;
input n_278;
input n_851;
input n_255;
input n_560;
input n_450;
input n_257;
input n_842;
input n_148;
input n_652;
input n_451;
input n_613;
input n_745;
input n_475;
input n_135;
input n_409;
input n_171;
input n_519;
input n_384;
input n_468;
input n_853;
input n_61;
input n_526;
input n_716;
input n_102;
input n_742;
input n_182;
input n_696;
input n_674;
input n_482;
input n_316;
input n_196;
input n_125;
input n_798;
input n_769;
input n_820;
input n_43;
input n_577;
input n_407;
input n_774;
input n_13;
input n_27;
input n_254;
input n_596;
input n_476;
input n_460;
input n_219;
input n_832;
input n_55;
input n_535;
input n_231;
input n_366;
input n_744;
input n_762;
input n_656;
input n_555;
input n_234;
input n_492;
input n_574;
input n_848;
input n_804;
input n_280;
input n_215;
input n_252;
input n_629;
input n_664;
input n_161;
input n_454;
input n_298;
input n_532;
input n_68;
input n_415;
input n_794;
input n_763;
input n_78;
input n_63;
input n_655;
input n_99;
input n_540;
input n_216;
input n_544;
input n_692;
input n_5;
input n_599;
input n_768;
input n_514;
input n_418;
input n_537;
input n_223;
input n_403;
input n_25;
input n_750;
input n_834;
input n_83;
input n_389;
input n_800;
input n_657;
input n_513;
input n_837;
input n_288;
input n_179;
input n_812;
input n_395;
input n_621;
input n_195;
input n_606;
input n_213;
input n_110;
input n_304;
input n_659;
input n_67;
input n_509;
input n_583;
input n_724;
input n_306;
input n_666;
input n_313;
input n_92;
input n_430;
input n_626;
input n_493;
input n_722;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_757;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_585;
input n_669;
input n_785;
input n_827;
input n_619;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_622;
input n_697;
input n_472;
input n_296;
input n_265;
input n_746;
input n_208;
input n_456;
input n_156;
input n_292;
input n_793;
input n_852;
input n_174;
input n_275;
input n_100;
input n_704;
input n_132;
input n_147;
input n_204;
input n_751;
input n_615;
input n_521;
input n_51;
input n_496;
input n_739;
input n_76;
input n_342;
input n_26;
input n_246;
input n_517;
input n_530;
input n_0;
input n_792;
input n_824;
input n_428;
input n_159;
input n_358;
input n_105;
input n_580;
input n_608;
input n_30;
input n_494;
input n_719;
input n_131;
input n_263;
input n_434;
input n_360;
input n_563;
input n_229;
input n_394;
input n_250;
input n_773;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_803;
input n_134;
input n_329;
input n_718;
input n_185;
input n_340;
input n_749;
input n_289;
input n_9;
input n_112;
input n_45;
input n_542;
input n_548;
input n_815;
input n_523;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_632;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_650;
input n_782;
input n_425;
input n_431;
input n_811;
input n_508;
input n_624;
input n_118;
input n_121;
input n_791;
input n_618;
input n_411;
input n_484;
input n_712;
input n_849;
input n_353;
input n_22;
input n_736;
input n_767;
input n_241;
input n_29;
input n_357;
input n_412;
input n_687;
input n_447;
input n_191;
input n_382;
input n_797;
input n_489;
input n_80;
input n_480;
input n_211;
input n_642;
input n_97;
input n_408;
input n_828;
input n_595;
input n_322;
input n_251;
input n_506;
input n_602;
input n_799;
input n_558;
input n_592;
input n_116;
input n_397;
input n_841;
input n_471;
input n_351;
input n_39;
input n_393;
input n_474;
input n_653;
input n_359;
input n_155;
input n_573;
input n_796;
input n_805;
input n_127;
input n_531;
input n_783;
input n_675;

output n_3113;

wire n_2752;
wire n_913;
wire n_1681;
wire n_2163;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_2484;
wire n_2866;
wire n_1174;
wire n_2346;
wire n_1469;
wire n_1353;
wire n_3056;
wire n_2679;
wire n_1355;
wire n_2131;
wire n_2559;
wire n_2500;
wire n_2509;
wire n_1383;
wire n_2182;
wire n_2135;
wire n_2334;
wire n_2680;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_2993;
wire n_1916;
wire n_2879;
wire n_1713;
wire n_1436;
wire n_2407;
wire n_2818;
wire n_1109;
wire n_1430;
wire n_2537;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_1238;
wire n_2694;
wire n_2011;
wire n_2729;
wire n_1515;
wire n_1837;
wire n_924;
wire n_2013;
wire n_2786;
wire n_1566;
wire n_2837;
wire n_2006;
wire n_952;
wire n_864;
wire n_2446;
wire n_1096;
wire n_1379;
wire n_2436;
wire n_2376;
wire n_2367;
wire n_2671;
wire n_2790;
wire n_1706;
wire n_2207;
wire n_2461;
wire n_2702;
wire n_2731;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_1503;
wire n_2238;
wire n_2529;
wire n_2374;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_2380;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_2646;
wire n_1298;
wire n_2653;
wire n_1745;
wire n_2873;
wire n_1366;
wire n_2084;
wire n_2278;
wire n_1088;
wire n_1424;
wire n_2976;
wire n_1835;
wire n_1457;
wire n_2482;
wire n_1682;
wire n_2750;
wire n_1836;
wire n_870;
wire n_2547;
wire n_1453;
wire n_945;
wire n_958;
wire n_2554;
wire n_2248;
wire n_3063;
wire n_1985;
wire n_2288;
wire n_2621;
wire n_2908;
wire n_3081;
wire n_995;
wire n_2579;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_2960;
wire n_903;
wire n_871;
wire n_2323;
wire n_1073;
wire n_2844;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_1761;
wire n_1062;
wire n_1690;
wire n_2221;
wire n_2807;
wire n_1283;
wire n_2317;
wire n_2838;
wire n_1974;
wire n_2906;
wire n_1736;
wire n_1018;
wire n_2342;
wire n_2200;
wire n_2781;
wire n_2442;
wire n_2735;
wire n_953;
wire n_1364;
wire n_2390;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_2709;
wire n_2634;
wire n_2322;
wire n_2746;
wire n_1107;
wire n_2832;
wire n_1688;
wire n_989;
wire n_2370;
wire n_1944;
wire n_2233;
wire n_2663;
wire n_2914;
wire n_1988;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_1428;
wire n_1284;
wire n_2878;
wire n_1241;
wire n_1514;
wire n_2539;
wire n_1528;
wire n_901;
wire n_2782;
wire n_2078;
wire n_1145;
wire n_971;
wire n_2359;
wire n_2201;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_1207;
wire n_1404;
wire n_868;
wire n_2232;
wire n_1847;
wire n_2458;
wire n_2779;
wire n_2950;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_2227;
wire n_2301;
wire n_1539;
wire n_2859;
wire n_2847;
wire n_884;
wire n_1851;
wire n_2162;
wire n_3015;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_2988;
wire n_1636;
wire n_1900;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_1977;
wire n_2650;
wire n_863;
wire n_1254;
wire n_929;
wire n_2433;
wire n_1703;
wire n_899;
wire n_2332;
wire n_2391;
wire n_3073;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_2571;
wire n_2427;
wire n_2885;
wire n_2098;
wire n_2616;
wire n_1751;
wire n_2874;
wire n_3003;
wire n_3049;
wire n_2867;
wire n_1917;
wire n_2456;
wire n_2769;
wire n_1924;
wire n_1560;
wire n_1654;
wire n_2341;
wire n_2899;
wire n_1548;
wire n_3066;
wire n_1811;
wire n_2045;
wire n_3013;
wire n_2575;
wire n_2722;
wire n_1396;
wire n_1230;
wire n_1840;
wire n_2739;
wire n_1597;
wire n_2942;
wire n_1771;
wire n_2902;
wire n_1544;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2685;
wire n_2094;
wire n_2512;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_2382;
wire n_2956;
wire n_2043;
wire n_2349;
wire n_1918;
wire n_2788;
wire n_1021;
wire n_1443;
wire n_3089;
wire n_2595;
wire n_1465;
wire n_2686;
wire n_3084;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_2727;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_1121;
wire n_1416;
wire n_2909;
wire n_1461;
wire n_2717;
wire n_3012;
wire n_1391;
wire n_2981;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_2527;
wire n_1112;
wire n_1159;
wire n_1216;
wire n_2759;
wire n_1245;
wire n_2743;
wire n_1669;
wire n_2969;
wire n_1675;
wire n_2466;
wire n_2038;
wire n_2263;
wire n_2800;
wire n_2568;
wire n_2116;
wire n_2271;
wire n_2145;
wire n_2326;
wire n_1838;
wire n_1594;
wire n_1935;
wire n_2806;
wire n_1716;
wire n_1872;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_1108;
wire n_1590;
wire n_1351;
wire n_2216;
wire n_1274;
wire n_2426;
wire n_1819;
wire n_3095;
wire n_947;
wire n_2134;
wire n_1260;
wire n_930;
wire n_1179;
wire n_2703;
wire n_1442;
wire n_2926;
wire n_2620;
wire n_1833;
wire n_1691;
wire n_916;
wire n_1386;
wire n_2810;
wire n_912;
wire n_1884;
wire n_1555;
wire n_1842;
wire n_2499;
wire n_2549;
wire n_1253;
wire n_1661;
wire n_1468;
wire n_2791;
wire n_2683;
wire n_1656;
wire n_1382;
wire n_3093;
wire n_2970;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_2855;
wire n_2166;
wire n_2848;
wire n_1692;
wire n_2611;
wire n_1562;
wire n_2748;
wire n_2185;
wire n_3029;
wire n_2398;
wire n_1376;
wire n_1292;
wire n_1178;
wire n_2015;
wire n_1972;
wire n_2925;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_2952;
wire n_2415;
wire n_2693;
wire n_2877;
wire n_2922;
wire n_3000;
wire n_2871;
wire n_2930;
wire n_2745;
wire n_2087;
wire n_931;
wire n_1491;
wire n_2628;
wire n_967;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_1357;
wire n_1079;
wire n_1787;
wire n_2462;
wire n_1389;
wire n_2155;
wire n_2659;
wire n_1139;
wire n_2836;
wire n_2439;
wire n_2864;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_2172;
wire n_2601;
wire n_892;
wire n_1880;
wire n_959;
wire n_2365;
wire n_2257;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_2219;
wire n_1855;
wire n_2100;
wire n_2333;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_2435;
wire n_1226;
wire n_2224;
wire n_944;
wire n_1932;
wire n_1780;
wire n_2825;
wire n_2888;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_2167;
wire n_2293;
wire n_2753;
wire n_1340;
wire n_2668;
wire n_1240;
wire n_2921;
wire n_3046;
wire n_1087;
wire n_2701;
wire n_2400;
wire n_3021;
wire n_2388;
wire n_2273;
wire n_2712;
wire n_1433;
wire n_1911;
wire n_2567;
wire n_2557;
wire n_2695;
wire n_2898;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_2755;
wire n_1071;
wire n_2598;
wire n_976;
wire n_909;
wire n_1392;
wire n_1832;
wire n_2795;
wire n_2682;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_2762;
wire n_964;
wire n_1627;
wire n_2220;
wire n_2954;
wire n_3014;
wire n_2294;
wire n_2274;
wire n_2895;
wire n_2903;
wire n_974;
wire n_1731;
wire n_1147;
wire n_2829;
wire n_2378;
wire n_2467;
wire n_2768;
wire n_965;
wire n_1914;
wire n_2253;
wire n_934;
wire n_2213;
wire n_1447;
wire n_2363;
wire n_1220;
wire n_2019;
wire n_2728;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_3010;
wire n_2160;
wire n_1992;
wire n_2924;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_3052;
wire n_2507;
wire n_2142;
wire n_1633;
wire n_2625;
wire n_2896;
wire n_1913;
wire n_2069;
wire n_2495;
wire n_1058;
wire n_2328;
wire n_2434;
wire n_1042;
wire n_1234;
wire n_2311;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_2287;
wire n_2223;
wire n_3082;
wire n_1279;
wire n_2473;
wire n_2144;
wire n_2511;
wire n_1029;
wire n_2649;
wire n_1247;
wire n_2438;
wire n_1568;
wire n_2919;
wire n_1483;
wire n_3108;
wire n_1363;
wire n_2681;
wire n_1111;
wire n_970;
wire n_1689;
wire n_2535;
wire n_1255;
wire n_2632;
wire n_1646;
wire n_3031;
wire n_2262;
wire n_2565;
wire n_1237;
wire n_927;
wire n_1095;
wire n_2980;
wire n_1728;
wire n_2335;
wire n_3078;
wire n_2120;
wire n_2631;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_2860;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_3087;
wire n_2697;
wire n_1387;
wire n_1263;
wire n_1817;
wire n_2404;
wire n_2168;
wire n_2757;
wire n_2312;
wire n_2677;
wire n_1826;
wire n_2834;
wire n_2483;
wire n_1951;
wire n_2490;
wire n_1032;
wire n_1217;
wire n_2558;
wire n_1496;
wire n_2996;
wire n_1592;
wire n_2812;
wire n_2662;
wire n_1259;
wire n_2801;
wire n_1177;
wire n_3104;
wire n_3074;
wire n_2655;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_2718;
wire n_926;
wire n_1943;
wire n_2687;
wire n_2296;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_2765;
wire n_1163;
wire n_2640;
wire n_3054;
wire n_2811;
wire n_3019;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2146;
wire n_2983;
wire n_1868;
wire n_1501;
wire n_2241;
wire n_2373;
wire n_1173;
wire n_2350;
wire n_1068;
wire n_1198;
wire n_2531;
wire n_1570;
wire n_2099;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2617;
wire n_2481;
wire n_2129;
wire n_855;
wire n_2327;
wire n_1365;
wire n_2476;
wire n_2814;
wire n_2059;
wire n_2437;
wire n_2636;
wire n_1439;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_2841;
wire n_1611;
wire n_2122;
wire n_2975;
wire n_2399;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_2055;
wire n_2998;
wire n_2027;
wire n_2932;
wire n_1423;
wire n_2117;
wire n_1609;
wire n_1053;
wire n_2822;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_1906;
wire n_1899;
wire n_3039;
wire n_2195;
wire n_2194;
wire n_2937;
wire n_1467;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_3057;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_3007;
wire n_2267;
wire n_1105;
wire n_3022;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_874;
wire n_2286;
wire n_2023;
wire n_1278;
wire n_983;
wire n_3036;
wire n_2783;
wire n_2599;
wire n_1726;
wire n_2075;
wire n_2523;
wire n_1945;
wire n_1015;
wire n_2496;
wire n_1377;
wire n_1162;
wire n_1614;
wire n_2031;
wire n_2418;
wire n_2118;
wire n_1740;
wire n_1602;
wire n_2853;
wire n_1098;
wire n_3009;
wire n_1490;
wire n_2338;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_3025;
wire n_3051;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_2802;
wire n_3035;
wire n_887;
wire n_2057;
wire n_2218;
wire n_1122;
wire n_1408;
wire n_1205;
wire n_2593;
wire n_1693;
wire n_2125;
wire n_2716;
wire n_1132;
wire n_1156;
wire n_2741;
wire n_2184;
wire n_2714;
wire n_1823;
wire n_2944;
wire n_2861;
wire n_2780;
wire n_3023;
wire n_1120;
wire n_1202;
wire n_2254;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_2618;
wire n_1402;
wire n_957;
wire n_1242;
wire n_2774;
wire n_2707;
wire n_2754;
wire n_2849;
wire n_1607;
wire n_1489;
wire n_2799;
wire n_1218;
wire n_2756;
wire n_2217;
wire n_2226;
wire n_1586;
wire n_861;
wire n_2962;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_2763;
wire n_2256;
wire n_1189;
wire n_1089;
wire n_1859;
wire n_2660;
wire n_1502;
wire n_3044;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_2732;
wire n_1883;
wire n_2516;
wire n_2776;
wire n_2555;
wire n_1969;
wire n_2708;
wire n_3070;
wire n_1005;
wire n_2379;
wire n_1294;
wire n_2661;
wire n_1667;
wire n_888;
wire n_2894;
wire n_2300;
wire n_2949;
wire n_1649;
wire n_2452;
wire n_1677;
wire n_2470;
wire n_1927;
wire n_1297;
wire n_2827;
wire n_1708;
wire n_3085;
wire n_1222;
wire n_2284;
wire n_3005;
wire n_1844;
wire n_2283;
wire n_2526;
wire n_1957;
wire n_1953;
wire n_2643;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_1919;
wire n_2994;
wire n_2508;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_2594;
wire n_2266;
wire n_2449;
wire n_890;
wire n_1898;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_2742;
wire n_1797;
wire n_2366;
wire n_2493;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_1895;
wire n_2821;
wire n_2690;
wire n_3090;
wire n_2474;
wire n_2623;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_1331;
wire n_1890;
wire n_2904;
wire n_3064;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_2946;
wire n_1734;
wire n_1860;
wire n_3065;
wire n_3016;
wire n_2460;
wire n_2840;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_2448;
wire n_2211;
wire n_2292;
wire n_2480;
wire n_951;
wire n_3024;
wire n_2772;
wire n_862;
wire n_1700;
wire n_2637;
wire n_1332;
wire n_2306;
wire n_1854;
wire n_1747;
wire n_2071;
wire n_2424;
wire n_1206;
wire n_1729;
wire n_1508;
wire n_2414;
wire n_2082;
wire n_2893;
wire n_2959;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_2389;
wire n_1309;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_2978;
wire n_1342;
wire n_2737;
wire n_1867;
wire n_1394;
wire n_2916;
wire n_2576;
wire n_2958;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_2696;
wire n_2140;
wire n_1748;
wire n_873;
wire n_1301;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_2468;
wire n_1400;
wire n_2035;
wire n_2614;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_2581;
wire n_1783;
wire n_2494;
wire n_1538;
wire n_2831;
wire n_2457;
wire n_2128;
wire n_3069;
wire n_2992;
wire n_1037;
wire n_1329;
wire n_1993;
wire n_1545;
wire n_2629;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_2540;
wire n_1605;
wire n_1078;
wire n_3060;
wire n_2486;
wire n_1897;
wire n_2984;
wire n_2520;
wire n_2137;
wire n_1161;
wire n_2489;
wire n_3097;
wire n_876;
wire n_1191;
wire n_2492;
wire n_2939;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_2337;
wire n_2265;
wire n_2900;
wire n_2026;
wire n_2912;
wire n_1786;
wire n_2627;
wire n_1327;
wire n_1475;
wire n_1804;
wire n_2106;
wire n_1406;
wire n_1405;
wire n_2684;
wire n_2726;
wire n_2622;
wire n_2272;
wire n_1757;
wire n_3102;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_1632;
wire n_1769;
wire n_1929;
wire n_1950;
wire n_2264;
wire n_2691;
wire n_2032;
wire n_2090;
wire n_2929;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_1526;
wire n_2991;
wire n_1305;
wire n_1596;
wire n_2348;
wire n_2785;
wire n_1281;
wire n_2574;
wire n_2364;
wire n_1997;
wire n_2656;
wire n_1873;
wire n_1137;
wire n_1258;
wire n_1733;
wire n_1856;
wire n_1476;
wire n_1524;
wire n_2016;
wire n_2723;
wire n_2667;
wire n_2725;
wire n_2928;
wire n_1118;
wire n_943;
wire n_2905;
wire n_2884;
wire n_2850;
wire n_1874;
wire n_1293;
wire n_961;
wire n_1046;
wire n_1807;
wire n_1123;
wire n_1657;
wire n_878;
wire n_2857;
wire n_1784;
wire n_3110;
wire n_1321;
wire n_3050;
wire n_2307;
wire n_1488;
wire n_985;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_2730;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_1561;
wire n_2720;
wire n_2412;
wire n_3107;
wire n_1352;
wire n_2405;
wire n_2815;
wire n_1824;
wire n_2700;
wire n_2606;
wire n_1492;
wire n_2383;
wire n_2764;
wire n_1441;
wire n_1822;
wire n_1616;
wire n_2633;
wire n_2416;
wire n_2386;
wire n_2907;
wire n_1971;
wire n_2945;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_2353;
wire n_2528;
wire n_1778;
wire n_1776;
wire n_2936;
wire n_1154;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_2325;
wire n_1130;
wire n_1450;
wire n_2022;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_1505;
wire n_2408;
wire n_2698;
wire n_2986;
wire n_2320;
wire n_3017;
wire n_979;
wire n_2329;
wire n_2570;
wire n_1642;
wire n_2417;
wire n_2789;
wire n_2525;
wire n_1815;
wire n_2813;
wire n_897;
wire n_2546;
wire n_949;
wire n_2454;
wire n_1493;
wire n_2890;
wire n_2911;
wire n_891;
wire n_885;
wire n_1659;
wire n_2354;
wire n_1864;
wire n_2760;
wire n_3086;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_2368;
wire n_1151;
wire n_960;
wire n_2352;
wire n_2502;
wire n_1256;
wire n_2170;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_2377;
wire n_1577;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_2652;
wire n_1133;
wire n_3067;
wire n_883;
wire n_1852;
wire n_1286;
wire n_2612;
wire n_1685;
wire n_2410;
wire n_2314;
wire n_2477;
wire n_2279;
wire n_2222;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2133;
wire n_2203;
wire n_2943;
wire n_1426;
wire n_2250;
wire n_2497;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_2001;
wire n_1047;
wire n_2506;
wire n_1472;
wire n_2413;
wire n_1593;
wire n_2610;
wire n_1050;
wire n_2626;
wire n_2158;
wire n_2578;
wire n_2607;
wire n_2285;
wire n_2892;
wire n_1288;
wire n_1201;
wire n_2796;
wire n_858;
wire n_2804;
wire n_1185;
wire n_2605;
wire n_2475;
wire n_2173;
wire n_2715;
wire n_1035;
wire n_1143;
wire n_2665;
wire n_2070;
wire n_2136;
wire n_2771;
wire n_1090;
wire n_2403;
wire n_2947;
wire n_1367;
wire n_2044;
wire n_928;
wire n_1153;
wire n_1103;
wire n_2619;
wire n_1565;
wire n_1192;
wire n_894;
wire n_3098;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_2854;
wire n_3055;
wire n_1291;
wire n_2020;
wire n_2310;
wire n_1045;
wire n_1160;
wire n_2968;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_2711;
wire n_1881;
wire n_2635;
wire n_2999;
wire n_988;
wire n_914;
wire n_1116;
wire n_3043;
wire n_1958;
wire n_2747;
wire n_3027;
wire n_1511;
wire n_2177;
wire n_2713;
wire n_1422;
wire n_2766;
wire n_1965;
wire n_1197;
wire n_3011;
wire n_2820;
wire n_2613;
wire n_1165;
wire n_2934;
wire n_1641;
wire n_2845;
wire n_1517;
wire n_2036;
wire n_2647;
wire n_2003;
wire n_2533;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_2343;
wire n_3096;
wire n_2419;
wire n_1049;
wire n_2330;
wire n_2826;
wire n_869;
wire n_1398;
wire n_1921;
wire n_2777;
wire n_2450;
wire n_2411;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_2309;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_2431;
wire n_1773;
wire n_1440;
wire n_2666;
wire n_1370;
wire n_1603;
wire n_2401;
wire n_2935;
wire n_889;
wire n_1066;
wire n_1549;
wire n_2588;
wire n_2863;
wire n_2331;
wire n_935;
wire n_2886;
wire n_2478;
wire n_911;
wire n_2658;
wire n_2608;
wire n_2920;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_1534;
wire n_1948;
wire n_3006;
wire n_2767;
wire n_1290;
wire n_1959;
wire n_2396;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_2692;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_1194;
wire n_2862;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_2553;
wire n_2645;
wire n_907;
wire n_2749;
wire n_1454;
wire n_2592;
wire n_2459;
wire n_962;
wire n_941;
wire n_1210;
wire n_1622;
wire n_1135;
wire n_2566;
wire n_2751;
wire n_3101;
wire n_918;
wire n_1968;
wire n_1885;
wire n_2842;
wire n_2833;
wire n_2196;
wire n_1038;
wire n_2371;
wire n_1978;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_3008;
wire n_1695;
wire n_2560;
wire n_1164;
wire n_2313;
wire n_3077;
wire n_1193;
wire n_3048;
wire n_1345;
wire n_3037;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_3062;
wire n_1774;
wire n_2963;
wire n_2609;
wire n_2561;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_1158;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_1749;
wire n_872;
wire n_1653;
wire n_2882;
wire n_2303;
wire n_2669;
wire n_1157;
wire n_1584;
wire n_1664;
wire n_1739;
wire n_2642;
wire n_1814;
wire n_2154;
wire n_2441;
wire n_2236;
wire n_1789;
wire n_1986;
wire n_2174;
wire n_2688;
wire n_2624;
wire n_2054;
wire n_1857;
wire n_2315;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_2938;
wire n_1612;
wire n_2498;
wire n_2638;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_2803;
wire n_1756;
wire n_2887;
wire n_1606;
wire n_2189;
wire n_2648;
wire n_1587;
wire n_2093;
wire n_2340;
wire n_2018;
wire n_2672;
wire n_1772;
wire n_2444;
wire n_2602;
wire n_1014;
wire n_2204;
wire n_2931;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_1311;
wire n_2977;
wire n_3106;
wire n_2199;
wire n_2881;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_875;
wire n_1617;
wire n_2455;
wire n_2600;
wire n_3092;
wire n_2231;
wire n_2828;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_2305;
wire n_880;
wire n_2114;
wire n_2927;
wire n_1175;
wire n_2289;
wire n_2530;
wire n_2299;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_1621;
wire n_1485;
wire n_1028;
wire n_2883;
wire n_1221;
wire n_1785;
wire n_1262;
wire n_1942;
wire n_2180;
wire n_2951;
wire n_1579;
wire n_2809;
wire n_2181;
wire n_2014;
wire n_975;
wire n_2974;
wire n_1645;
wire n_923;
wire n_1381;
wire n_1124;
wire n_2870;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_2889;
wire n_2276;
wire n_1805;
wire n_2282;
wire n_981;
wire n_2910;
wire n_2141;
wire n_1758;
wire n_1110;
wire n_2503;
wire n_2270;
wire n_2443;
wire n_1407;
wire n_2465;
wire n_1204;
wire n_2865;
wire n_1554;
wire n_994;
wire n_2428;
wire n_2972;
wire n_2586;
wire n_2989;
wire n_1360;
wire n_973;
wire n_2858;
wire n_972;
wire n_2251;
wire n_2923;
wire n_3076;
wire n_2843;
wire n_856;
wire n_3100;
wire n_2572;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_1679;
wire n_2872;
wire n_2126;
wire n_3109;
wire n_1952;
wire n_2425;
wire n_2394;
wire n_1858;
wire n_1678;
wire n_2589;
wire n_1482;
wire n_1361;
wire n_2356;
wire n_1601;
wire n_1057;
wire n_2487;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_2534;
wire n_2488;
wire n_1509;
wire n_2941;
wire n_1411;
wire n_1359;
wire n_3079;
wire n_1721;
wire n_2564;
wire n_2591;
wire n_1445;
wire n_1317;
wire n_3034;
wire n_2050;
wire n_2197;
wire n_2550;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_2385;
wire n_2387;
wire n_1008;
wire n_3091;
wire n_1024;
wire n_2291;
wire n_2816;
wire n_1980;
wire n_2518;
wire n_987;
wire n_936;
wire n_2510;
wire n_1620;
wire n_2501;
wire n_2542;
wire n_3105;
wire n_1385;
wire n_1525;
wire n_2793;
wire n_1998;
wire n_2165;
wire n_2675;
wire n_2604;
wire n_1775;
wire n_908;
wire n_2639;
wire n_1036;
wire n_2169;
wire n_2985;
wire n_2603;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_2630;
wire n_2794;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2901;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_2773;
wire n_2817;
wire n_1926;
wire n_2402;
wire n_1458;
wire n_1630;
wire n_3047;
wire n_1720;
wire n_2409;
wire n_2966;
wire n_2176;
wire n_1412;
wire n_3059;
wire n_1738;
wire n_1550;
wire n_1358;
wire n_1200;
wire n_2808;
wire n_2453;
wire n_2344;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_940;
wire n_2392;
wire n_1537;
wire n_2138;
wire n_3040;
wire n_2065;
wire n_2543;
wire n_2321;
wire n_1077;
wire n_2597;
wire n_956;
wire n_1930;
wire n_1809;
wire n_2787;
wire n_1904;
wire n_1843;
wire n_2000;
wire n_2805;
wire n_1268;
wire n_2676;
wire n_2758;
wire n_2395;
wire n_917;
wire n_2868;
wire n_1271;
wire n_2096;
wire n_2440;
wire n_2556;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_2770;
wire n_1170;
wire n_2724;
wire n_2258;
wire n_1261;
wire n_2471;
wire n_857;
wire n_898;
wire n_3042;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_2584;
wire n_2375;
wire n_1462;
wire n_2012;
wire n_1937;
wire n_2967;
wire n_1064;
wire n_900;
wire n_1446;
wire n_1282;
wire n_3004;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_3111;
wire n_2212;
wire n_1813;
wire n_2268;
wire n_2997;
wire n_1452;
wire n_2835;
wire n_1573;
wire n_2734;
wire n_2569;
wire n_2252;
wire n_2111;
wire n_2420;
wire n_2948;
wire n_3099;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_2897;
wire n_1322;
wire n_2583;
wire n_2918;
wire n_2987;
wire n_1473;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_2651;
wire n_2445;
wire n_2733;
wire n_1770;
wire n_1003;
wire n_2469;
wire n_1125;
wire n_2103;
wire n_2358;
wire n_1710;
wire n_1865;
wire n_2522;
wire n_2641;
wire n_2463;
wire n_1344;
wire n_2355;
wire n_1390;
wire n_2580;
wire n_2699;
wire n_1792;
wire n_2062;
wire n_3068;
wire n_1141;
wire n_1629;
wire n_1640;
wire n_1094;
wire n_2973;
wire n_1459;
wire n_2153;
wire n_2324;
wire n_1510;
wire n_3002;
wire n_2710;
wire n_2505;
wire n_2139;
wire n_1099;
wire n_1754;
wire n_3038;
wire n_2397;
wire n_2521;
wire n_1727;
wire n_2740;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_2721;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_2615;
wire n_2775;
wire n_1212;
wire n_1619;
wire n_2351;
wire n_2260;
wire n_1660;
wire n_1315;
wire n_1902;
wire n_997;
wire n_2206;
wire n_2784;
wire n_2541;
wire n_1643;
wire n_1320;
wire n_3001;
wire n_1113;
wire n_2347;
wire n_1152;
wire n_2657;
wire n_2990;
wire n_2538;
wire n_2034;
wire n_1845;
wire n_2447;
wire n_1934;
wire n_2101;
wire n_2577;
wire n_921;
wire n_2362;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_1533;
wire n_1806;
wire n_2372;
wire n_2552;
wire n_1409;
wire n_1588;
wire n_1148;
wire n_1684;
wire n_1673;
wire n_2422;
wire n_2704;
wire n_1334;
wire n_2290;
wire n_2933;
wire n_2856;
wire n_2088;
wire n_1275;
wire n_3103;
wire n_3018;
wire n_904;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_3028;
wire n_1875;
wire n_1059;
wire n_2429;
wire n_2736;
wire n_2108;
wire n_1039;
wire n_2246;
wire n_1150;
wire n_977;
wire n_2339;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2532;
wire n_2191;
wire n_2971;
wire n_1497;
wire n_1866;
wire n_2472;
wire n_2705;
wire n_2664;
wire n_2056;
wire n_2852;
wire n_1136;
wire n_2515;
wire n_1782;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_2519;
wire n_950;
wire n_1017;
wire n_1915;
wire n_2360;
wire n_1393;
wire n_2240;
wire n_1369;
wire n_2846;
wire n_1781;
wire n_2917;
wire n_2544;
wire n_2085;
wire n_2432;
wire n_3032;
wire n_1686;
wire n_1964;
wire n_881;
wire n_1477;
wire n_1019;
wire n_1777;
wire n_2188;
wire n_1982;
wire n_2097;
wire n_2430;
wire n_2504;
wire n_910;
wire n_939;
wire n_1410;
wire n_2297;
wire n_3094;
wire n_3020;
wire n_2964;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_1223;
wire n_2545;
wire n_1768;
wire n_2513;
wire n_2193;
wire n_2369;
wire n_1199;
wire n_2957;
wire n_865;
wire n_1273;
wire n_1983;
wire n_2982;
wire n_1041;
wire n_2451;
wire n_2115;
wire n_2913;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_3061;
wire n_2587;
wire n_1347;
wire n_2839;
wire n_860;
wire n_3072;
wire n_1043;
wire n_2961;
wire n_2869;
wire n_1923;
wire n_2955;
wire n_2670;
wire n_1764;
wire n_2674;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_3026;
wire n_2644;
wire n_902;
wire n_1031;
wire n_2979;
wire n_1723;
wire n_1638;
wire n_3071;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_1946;
wire n_2148;
wire n_933;
wire n_1779;
wire n_2562;
wire n_954;
wire n_2051;
wire n_3112;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_2673;
wire n_1591;
wire n_2585;
wire n_2995;
wire n_1229;
wire n_1683;
wire n_2582;
wire n_2548;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_2381;
wire n_2744;
wire n_1967;
wire n_2384;
wire n_2678;
wire n_2179;
wire n_1280;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_1091;
wire n_2052;
wire n_2485;
wire n_1063;
wire n_991;
wire n_2183;
wire n_2205;
wire n_2275;
wire n_2563;
wire n_1724;
wire n_3088;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2761;
wire n_2357;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_2875;
wire n_1639;
wire n_2209;
wire n_2421;
wire n_1302;
wire n_1000;
wire n_1581;
wire n_1928;
wire n_946;
wire n_2047;
wire n_3058;
wire n_2792;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_2596;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_2269;
wire n_2081;
wire n_937;
wire n_1474;
wire n_2536;
wire n_2524;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_1794;
wire n_1375;
wire n_3053;
wire n_1232;
wire n_1211;
wire n_1368;
wire n_996;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_2891;
wire n_2318;
wire n_1827;
wire n_866;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_2361;
wire n_1115;
wire n_2229;
wire n_2819;
wire n_2880;
wire n_3030;
wire n_3075;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_2551;
wire n_1102;
wire n_2255;
wire n_1252;
wire n_1129;
wire n_2239;
wire n_3045;
wire n_1464;
wire n_1296;
wire n_2798;
wire n_2316;
wire n_2464;
wire n_1010;
wire n_2830;
wire n_882;
wire n_2706;
wire n_2304;
wire n_1249;
wire n_1871;
wire n_2514;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_2573;
wire n_2940;
wire n_2336;
wire n_1662;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_2915;
wire n_3083;
wire n_2654;
wire n_2491;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_2517;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_2259;
wire n_2095;
wire n_2719;
wire n_2965;
wire n_2738;
wire n_1820;
wire n_2590;
wire n_2876;
wire n_2797;
wire n_1251;
wire n_1989;
wire n_3041;
wire n_1421;
wire n_2208;
wire n_2423;
wire n_2689;
wire n_2778;
wire n_1762;
wire n_1233;
wire n_3080;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_3033;
wire n_1704;
wire n_893;
wire n_1582;
wire n_2479;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2824;
wire n_2037;
wire n_2953;
wire n_1308;
wire n_2851;
wire n_2823;
wire n_2345;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;

BUFx10_ASAP7_75t_L g854 ( 
.A(n_114),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_838),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_771),
.Y(n_856)
);

BUFx3_ASAP7_75t_L g857 ( 
.A(n_793),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_741),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_770),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_416),
.Y(n_860)
);

CKINVDCx20_ASAP7_75t_R g861 ( 
.A(n_779),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_719),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_748),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_84),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_412),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_728),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_390),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_760),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_738),
.Y(n_869)
);

BUFx3_ASAP7_75t_L g870 ( 
.A(n_824),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_807),
.Y(n_871)
);

BUFx3_ASAP7_75t_L g872 ( 
.A(n_638),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_58),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_849),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_590),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_789),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_821),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_544),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_734),
.Y(n_879)
);

HB1xp67_ASAP7_75t_L g880 ( 
.A(n_784),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_753),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_814),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_66),
.Y(n_883)
);

CKINVDCx20_ASAP7_75t_R g884 ( 
.A(n_668),
.Y(n_884)
);

BUFx3_ASAP7_75t_L g885 ( 
.A(n_763),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_722),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_5),
.Y(n_887)
);

CKINVDCx16_ASAP7_75t_R g888 ( 
.A(n_840),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_112),
.Y(n_889)
);

CKINVDCx20_ASAP7_75t_R g890 ( 
.A(n_711),
.Y(n_890)
);

BUFx3_ASAP7_75t_L g891 ( 
.A(n_820),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_718),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_841),
.Y(n_893)
);

INVx1_ASAP7_75t_SL g894 ( 
.A(n_9),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_184),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_777),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_612),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_743),
.Y(n_898)
);

BUFx6f_ASAP7_75t_L g899 ( 
.A(n_727),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_529),
.Y(n_900)
);

CKINVDCx20_ASAP7_75t_R g901 ( 
.A(n_195),
.Y(n_901)
);

CKINVDCx20_ASAP7_75t_R g902 ( 
.A(n_822),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_714),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_8),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_752),
.Y(n_905)
);

INVx2_ASAP7_75t_SL g906 ( 
.A(n_436),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_766),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_79),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_724),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_817),
.Y(n_910)
);

CKINVDCx20_ASAP7_75t_R g911 ( 
.A(n_680),
.Y(n_911)
);

BUFx3_ASAP7_75t_L g912 ( 
.A(n_832),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_572),
.Y(n_913)
);

INVx1_ASAP7_75t_SL g914 ( 
.A(n_826),
.Y(n_914)
);

BUFx3_ASAP7_75t_L g915 ( 
.A(n_445),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_705),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_835),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_617),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_358),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_536),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_759),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_531),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_778),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_422),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_675),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_136),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_322),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_844),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_622),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_512),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_553),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_169),
.Y(n_932)
);

INVx2_ASAP7_75t_SL g933 ( 
.A(n_651),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_803),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_781),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_740),
.Y(n_936)
);

BUFx10_ASAP7_75t_L g937 ( 
.A(n_746),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_754),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_570),
.Y(n_939)
);

CKINVDCx20_ASAP7_75t_R g940 ( 
.A(n_510),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_403),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_634),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_307),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_6),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_222),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_692),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_439),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_209),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_852),
.Y(n_949)
);

BUFx3_ASAP7_75t_L g950 ( 
.A(n_448),
.Y(n_950)
);

BUFx6f_ASAP7_75t_L g951 ( 
.A(n_555),
.Y(n_951)
);

BUFx10_ASAP7_75t_L g952 ( 
.A(n_102),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_702),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_244),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_496),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_324),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_580),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_561),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_810),
.Y(n_959)
);

CKINVDCx20_ASAP7_75t_R g960 ( 
.A(n_73),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_359),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_142),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_159),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_75),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_809),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_710),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_842),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_562),
.Y(n_968)
);

CKINVDCx20_ASAP7_75t_R g969 ( 
.A(n_441),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_816),
.Y(n_970)
);

BUFx3_ASAP7_75t_L g971 ( 
.A(n_457),
.Y(n_971)
);

INVxp67_ASAP7_75t_L g972 ( 
.A(n_767),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_466),
.Y(n_973)
);

INVx1_ASAP7_75t_SL g974 ( 
.A(n_792),
.Y(n_974)
);

BUFx6f_ASAP7_75t_L g975 ( 
.A(n_410),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_729),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_733),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_774),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_443),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_368),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_118),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_258),
.Y(n_982)
);

INVxp67_ASAP7_75t_SL g983 ( 
.A(n_96),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_519),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_742),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_415),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_5),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_794),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_843),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_269),
.Y(n_990)
);

BUFx10_ASAP7_75t_L g991 ( 
.A(n_137),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_281),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_2),
.Y(n_993)
);

HB1xp67_ASAP7_75t_L g994 ( 
.A(n_833),
.Y(n_994)
);

BUFx6f_ASAP7_75t_L g995 ( 
.A(n_611),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_630),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_586),
.Y(n_997)
);

BUFx10_ASAP7_75t_L g998 ( 
.A(n_178),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_776),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_310),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_449),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_805),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_115),
.Y(n_1003)
);

INVxp67_ASAP7_75t_L g1004 ( 
.A(n_761),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_747),
.Y(n_1005)
);

BUFx10_ASAP7_75t_L g1006 ( 
.A(n_147),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_515),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_315),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_138),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_400),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_352),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_431),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_785),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_737),
.Y(n_1014)
);

INVx1_ASAP7_75t_SL g1015 ( 
.A(n_279),
.Y(n_1015)
);

CKINVDCx16_ASAP7_75t_R g1016 ( 
.A(n_542),
.Y(n_1016)
);

BUFx6f_ASAP7_75t_L g1017 ( 
.A(n_802),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_797),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_433),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_142),
.Y(n_1020)
);

CKINVDCx20_ASAP7_75t_R g1021 ( 
.A(n_735),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_254),
.Y(n_1022)
);

INVxp67_ASAP7_75t_L g1023 ( 
.A(n_69),
.Y(n_1023)
);

BUFx6f_ASAP7_75t_L g1024 ( 
.A(n_801),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_661),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_581),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_381),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_234),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_319),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_489),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_819),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_749),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_839),
.Y(n_1033)
);

INVx1_ASAP7_75t_SL g1034 ( 
.A(n_588),
.Y(n_1034)
);

CKINVDCx20_ASAP7_75t_R g1035 ( 
.A(n_731),
.Y(n_1035)
);

CKINVDCx20_ASAP7_75t_R g1036 ( 
.A(n_273),
.Y(n_1036)
);

BUFx8_ASAP7_75t_SL g1037 ( 
.A(n_757),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_782),
.Y(n_1038)
);

CKINVDCx16_ASAP7_75t_R g1039 ( 
.A(n_606),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_800),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_847),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_302),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_582),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_357),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_811),
.Y(n_1045)
);

INVx4_ASAP7_75t_R g1046 ( 
.A(n_709),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_545),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_330),
.Y(n_1048)
);

INVx2_ASAP7_75t_SL g1049 ( 
.A(n_707),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_730),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_627),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_106),
.Y(n_1052)
);

CKINVDCx20_ASAP7_75t_R g1053 ( 
.A(n_351),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_769),
.Y(n_1054)
);

BUFx3_ASAP7_75t_L g1055 ( 
.A(n_723),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_736),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_134),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_755),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_823),
.Y(n_1059)
);

INVx3_ASAP7_75t_L g1060 ( 
.A(n_463),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_318),
.Y(n_1061)
);

HB1xp67_ASAP7_75t_L g1062 ( 
.A(n_775),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_726),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_488),
.Y(n_1064)
);

BUFx6f_ASAP7_75t_L g1065 ( 
.A(n_265),
.Y(n_1065)
);

CKINVDCx20_ASAP7_75t_R g1066 ( 
.A(n_177),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_699),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_657),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_323),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_0),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_136),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_125),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_831),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_713),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_164),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_732),
.Y(n_1076)
);

INVx1_ASAP7_75t_SL g1077 ( 
.A(n_813),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_397),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_768),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_666),
.Y(n_1080)
);

INVxp67_ASAP7_75t_SL g1081 ( 
.A(n_28),
.Y(n_1081)
);

CKINVDCx20_ASAP7_75t_R g1082 ( 
.A(n_329),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_806),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_574),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_708),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_716),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_830),
.Y(n_1087)
);

CKINVDCx20_ASAP7_75t_R g1088 ( 
.A(n_313),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_244),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_790),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_787),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_762),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_603),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_609),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_773),
.Y(n_1095)
);

INVxp67_ASAP7_75t_L g1096 ( 
.A(n_656),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_804),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_788),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_148),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_796),
.Y(n_1100)
);

CKINVDCx16_ASAP7_75t_R g1101 ( 
.A(n_270),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_256),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_783),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_258),
.Y(n_1104)
);

CKINVDCx20_ASAP7_75t_R g1105 ( 
.A(n_366),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_201),
.Y(n_1106)
);

BUFx6f_ASAP7_75t_L g1107 ( 
.A(n_815),
.Y(n_1107)
);

CKINVDCx20_ASAP7_75t_R g1108 ( 
.A(n_290),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_751),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_450),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_848),
.Y(n_1111)
);

INVx1_ASAP7_75t_SL g1112 ( 
.A(n_237),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_61),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_420),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_795),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_720),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_332),
.Y(n_1117)
);

BUFx2_ASAP7_75t_L g1118 ( 
.A(n_712),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_82),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_389),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_624),
.Y(n_1121)
);

INVx2_ASAP7_75t_SL g1122 ( 
.A(n_53),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_739),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_827),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_429),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_681),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_780),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_121),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_828),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_589),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_461),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_725),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_272),
.Y(n_1133)
);

CKINVDCx20_ASAP7_75t_R g1134 ( 
.A(n_745),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_791),
.Y(n_1135)
);

BUFx6f_ASAP7_75t_L g1136 ( 
.A(n_344),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_340),
.Y(n_1137)
);

INVx1_ASAP7_75t_SL g1138 ( 
.A(n_834),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_535),
.Y(n_1139)
);

BUFx3_ASAP7_75t_L g1140 ( 
.A(n_756),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_837),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_179),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_251),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_547),
.Y(n_1144)
);

INVx4_ASAP7_75t_R g1145 ( 
.A(n_36),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_808),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_345),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_195),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_518),
.Y(n_1149)
);

BUFx10_ASAP7_75t_L g1150 ( 
.A(n_374),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_419),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_786),
.Y(n_1152)
);

CKINVDCx20_ASAP7_75t_R g1153 ( 
.A(n_706),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_211),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_799),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_331),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_721),
.Y(n_1157)
);

CKINVDCx20_ASAP7_75t_R g1158 ( 
.A(n_70),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_593),
.Y(n_1159)
);

CKINVDCx20_ASAP7_75t_R g1160 ( 
.A(n_266),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_818),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_626),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_587),
.Y(n_1163)
);

CKINVDCx14_ASAP7_75t_R g1164 ( 
.A(n_303),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_812),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_432),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_522),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_685),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_764),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_369),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_356),
.Y(n_1171)
);

CKINVDCx20_ASAP7_75t_R g1172 ( 
.A(n_194),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_407),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_528),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_92),
.Y(n_1175)
);

INVxp67_ASAP7_75t_L g1176 ( 
.A(n_176),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_81),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_772),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_78),
.Y(n_1179)
);

BUFx10_ASAP7_75t_L g1180 ( 
.A(n_453),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_546),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_229),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_308),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_836),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_825),
.Y(n_1185)
);

BUFx10_ASAP7_75t_L g1186 ( 
.A(n_744),
.Y(n_1186)
);

CKINVDCx16_ASAP7_75t_R g1187 ( 
.A(n_758),
.Y(n_1187)
);

CKINVDCx20_ASAP7_75t_R g1188 ( 
.A(n_637),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_639),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_376),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_159),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_186),
.Y(n_1192)
);

INVx2_ASAP7_75t_L g1193 ( 
.A(n_798),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_765),
.Y(n_1194)
);

HB1xp67_ASAP7_75t_L g1195 ( 
.A(n_750),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_120),
.Y(n_1196)
);

CKINVDCx20_ASAP7_75t_R g1197 ( 
.A(n_261),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_715),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_435),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_216),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_717),
.Y(n_1201)
);

INVx2_ASAP7_75t_L g1202 ( 
.A(n_526),
.Y(n_1202)
);

INVxp67_ASAP7_75t_L g1203 ( 
.A(n_386),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_549),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_829),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_191),
.Y(n_1206)
);

CKINVDCx20_ASAP7_75t_R g1207 ( 
.A(n_615),
.Y(n_1207)
);

INVxp67_ASAP7_75t_SL g1208 ( 
.A(n_1065),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_895),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_1065),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_944),
.Y(n_1211)
);

INVxp33_ASAP7_75t_L g1212 ( 
.A(n_987),
.Y(n_1212)
);

INVxp33_ASAP7_75t_SL g1213 ( 
.A(n_864),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_982),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1003),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1009),
.Y(n_1216)
);

BUFx6f_ASAP7_75t_L g1217 ( 
.A(n_1065),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1020),
.Y(n_1218)
);

INVx2_ASAP7_75t_L g1219 ( 
.A(n_1022),
.Y(n_1219)
);

CKINVDCx16_ASAP7_75t_R g1220 ( 
.A(n_1101),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1028),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_1037),
.Y(n_1222)
);

CKINVDCx20_ASAP7_75t_R g1223 ( 
.A(n_861),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1057),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1072),
.Y(n_1225)
);

CKINVDCx16_ASAP7_75t_R g1226 ( 
.A(n_888),
.Y(n_1226)
);

INVxp67_ASAP7_75t_SL g1227 ( 
.A(n_1089),
.Y(n_1227)
);

INVxp67_ASAP7_75t_SL g1228 ( 
.A(n_1099),
.Y(n_1228)
);

INVx2_ASAP7_75t_L g1229 ( 
.A(n_1104),
.Y(n_1229)
);

INVxp67_ASAP7_75t_SL g1230 ( 
.A(n_1133),
.Y(n_1230)
);

CKINVDCx20_ASAP7_75t_R g1231 ( 
.A(n_884),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1142),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1148),
.Y(n_1233)
);

HB1xp67_ASAP7_75t_L g1234 ( 
.A(n_873),
.Y(n_1234)
);

CKINVDCx20_ASAP7_75t_R g1235 ( 
.A(n_890),
.Y(n_1235)
);

INVxp67_ASAP7_75t_SL g1236 ( 
.A(n_1196),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_880),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_994),
.Y(n_1238)
);

NOR2xp33_ASAP7_75t_L g1239 ( 
.A(n_1118),
.B(n_1),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_902),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1062),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1195),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1122),
.Y(n_1243)
);

CKINVDCx20_ASAP7_75t_R g1244 ( 
.A(n_911),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_937),
.Y(n_1245)
);

CKINVDCx14_ASAP7_75t_R g1246 ( 
.A(n_1164),
.Y(n_1246)
);

BUFx5_ASAP7_75t_L g1247 ( 
.A(n_856),
.Y(n_1247)
);

BUFx3_ASAP7_75t_L g1248 ( 
.A(n_937),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1150),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1150),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1180),
.Y(n_1251)
);

CKINVDCx16_ASAP7_75t_R g1252 ( 
.A(n_1016),
.Y(n_1252)
);

INVxp33_ASAP7_75t_L g1253 ( 
.A(n_854),
.Y(n_1253)
);

BUFx2_ASAP7_75t_L g1254 ( 
.A(n_883),
.Y(n_1254)
);

INVxp33_ASAP7_75t_L g1255 ( 
.A(n_854),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1180),
.Y(n_1256)
);

INVxp67_ASAP7_75t_L g1257 ( 
.A(n_952),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1186),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_940),
.Y(n_1259)
);

INVxp67_ASAP7_75t_SL g1260 ( 
.A(n_1023),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1186),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_952),
.Y(n_1262)
);

CKINVDCx5p33_ASAP7_75t_R g1263 ( 
.A(n_969),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_991),
.Y(n_1264)
);

CKINVDCx5p33_ASAP7_75t_R g1265 ( 
.A(n_1021),
.Y(n_1265)
);

BUFx3_ASAP7_75t_L g1266 ( 
.A(n_857),
.Y(n_1266)
);

INVxp33_ASAP7_75t_SL g1267 ( 
.A(n_887),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_991),
.Y(n_1268)
);

OA21x2_ASAP7_75t_L g1269 ( 
.A1(n_1208),
.A2(n_863),
.B(n_862),
.Y(n_1269)
);

HB1xp67_ASAP7_75t_L g1270 ( 
.A(n_1220),
.Y(n_1270)
);

INVx3_ASAP7_75t_L g1271 ( 
.A(n_1266),
.Y(n_1271)
);

BUFx12f_ASAP7_75t_L g1272 ( 
.A(n_1222),
.Y(n_1272)
);

BUFx3_ASAP7_75t_L g1273 ( 
.A(n_1248),
.Y(n_1273)
);

CKINVDCx16_ASAP7_75t_R g1274 ( 
.A(n_1226),
.Y(n_1274)
);

BUFx6f_ASAP7_75t_L g1275 ( 
.A(n_1217),
.Y(n_1275)
);

INVx5_ASAP7_75t_L g1276 ( 
.A(n_1217),
.Y(n_1276)
);

AND2x2_ASAP7_75t_SL g1277 ( 
.A(n_1239),
.B(n_1039),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_1210),
.Y(n_1278)
);

AND2x4_ASAP7_75t_L g1279 ( 
.A(n_1245),
.B(n_1176),
.Y(n_1279)
);

INVx4_ASAP7_75t_L g1280 ( 
.A(n_1254),
.Y(n_1280)
);

OA21x2_ASAP7_75t_L g1281 ( 
.A1(n_1227),
.A2(n_874),
.B(n_868),
.Y(n_1281)
);

OAI22xp5_ASAP7_75t_L g1282 ( 
.A1(n_1252),
.A2(n_901),
.B1(n_1036),
.B2(n_960),
.Y(n_1282)
);

OA21x2_ASAP7_75t_L g1283 ( 
.A1(n_1228),
.A2(n_879),
.B(n_875),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1209),
.Y(n_1284)
);

INVx5_ASAP7_75t_L g1285 ( 
.A(n_1219),
.Y(n_1285)
);

BUFx6f_ASAP7_75t_L g1286 ( 
.A(n_1229),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1211),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1246),
.B(n_1187),
.Y(n_1288)
);

INVx3_ASAP7_75t_L g1289 ( 
.A(n_1214),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1215),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1216),
.Y(n_1291)
);

BUFx3_ASAP7_75t_L g1292 ( 
.A(n_1247),
.Y(n_1292)
);

INVx3_ASAP7_75t_L g1293 ( 
.A(n_1218),
.Y(n_1293)
);

BUFx6f_ASAP7_75t_L g1294 ( 
.A(n_1221),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1249),
.B(n_882),
.Y(n_1295)
);

INVx4_ASAP7_75t_L g1296 ( 
.A(n_1247),
.Y(n_1296)
);

BUFx6f_ASAP7_75t_L g1297 ( 
.A(n_1224),
.Y(n_1297)
);

OA21x2_ASAP7_75t_L g1298 ( 
.A1(n_1230),
.A2(n_903),
.B(n_898),
.Y(n_1298)
);

AND2x4_ASAP7_75t_L g1299 ( 
.A(n_1250),
.B(n_983),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1225),
.Y(n_1300)
);

AND2x2_ASAP7_75t_L g1301 ( 
.A(n_1212),
.B(n_998),
.Y(n_1301)
);

BUFx6f_ASAP7_75t_L g1302 ( 
.A(n_1232),
.Y(n_1302)
);

BUFx6f_ASAP7_75t_L g1303 ( 
.A(n_1233),
.Y(n_1303)
);

INVx2_ASAP7_75t_L g1304 ( 
.A(n_1247),
.Y(n_1304)
);

BUFx12f_ASAP7_75t_L g1305 ( 
.A(n_1240),
.Y(n_1305)
);

BUFx3_ASAP7_75t_L g1306 ( 
.A(n_1247),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1243),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1251),
.B(n_909),
.Y(n_1308)
);

HB1xp67_ASAP7_75t_L g1309 ( 
.A(n_1234),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1236),
.Y(n_1310)
);

INVx2_ASAP7_75t_L g1311 ( 
.A(n_1237),
.Y(n_1311)
);

OAI22xp5_ASAP7_75t_SL g1312 ( 
.A1(n_1223),
.A2(n_1158),
.B1(n_1160),
.B2(n_1066),
.Y(n_1312)
);

AOI22x1_ASAP7_75t_SL g1313 ( 
.A1(n_1231),
.A2(n_1197),
.B1(n_1172),
.B2(n_981),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1294),
.Y(n_1314)
);

BUFx2_ASAP7_75t_L g1315 ( 
.A(n_1270),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1297),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1302),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1301),
.B(n_1253),
.Y(n_1318)
);

INVx3_ASAP7_75t_L g1319 ( 
.A(n_1271),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_1278),
.Y(n_1320)
);

AND2x4_ASAP7_75t_L g1321 ( 
.A(n_1273),
.B(n_1257),
.Y(n_1321)
);

INVx2_ASAP7_75t_L g1322 ( 
.A(n_1286),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1284),
.Y(n_1323)
);

INVx2_ASAP7_75t_L g1324 ( 
.A(n_1303),
.Y(n_1324)
);

BUFx6f_ASAP7_75t_L g1325 ( 
.A(n_1303),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1287),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1290),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1291),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1307),
.Y(n_1329)
);

CKINVDCx16_ASAP7_75t_R g1330 ( 
.A(n_1274),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1304),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1300),
.Y(n_1332)
);

BUFx3_ASAP7_75t_L g1333 ( 
.A(n_1272),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1309),
.B(n_1255),
.Y(n_1334)
);

HB1xp67_ASAP7_75t_L g1335 ( 
.A(n_1282),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1280),
.B(n_1260),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1289),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_1293),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1292),
.B(n_1256),
.Y(n_1339)
);

XNOR2xp5_ASAP7_75t_L g1340 ( 
.A(n_1277),
.B(n_1259),
.Y(n_1340)
);

INVxp67_ASAP7_75t_L g1341 ( 
.A(n_1288),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1310),
.Y(n_1342)
);

HB1xp67_ASAP7_75t_L g1343 ( 
.A(n_1305),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1281),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1283),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1298),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1311),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1269),
.Y(n_1348)
);

BUFx6f_ASAP7_75t_L g1349 ( 
.A(n_1275),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_SL g1350 ( 
.A(n_1277),
.B(n_1213),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1306),
.B(n_1258),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1295),
.Y(n_1352)
);

BUFx6f_ASAP7_75t_L g1353 ( 
.A(n_1276),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1308),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1285),
.Y(n_1355)
);

INVx3_ASAP7_75t_L g1356 ( 
.A(n_1285),
.Y(n_1356)
);

INVx3_ASAP7_75t_L g1357 ( 
.A(n_1276),
.Y(n_1357)
);

AND2x4_ASAP7_75t_L g1358 ( 
.A(n_1279),
.B(n_1261),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1296),
.Y(n_1359)
);

INVxp67_ASAP7_75t_L g1360 ( 
.A(n_1312),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_1299),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1313),
.Y(n_1362)
);

BUFx6f_ASAP7_75t_L g1363 ( 
.A(n_1286),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_1278),
.Y(n_1364)
);

BUFx2_ASAP7_75t_L g1365 ( 
.A(n_1270),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1278),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1294),
.Y(n_1367)
);

INVxp67_ASAP7_75t_L g1368 ( 
.A(n_1301),
.Y(n_1368)
);

INVx3_ASAP7_75t_L g1369 ( 
.A(n_1271),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1278),
.Y(n_1370)
);

BUFx2_ASAP7_75t_L g1371 ( 
.A(n_1270),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_SL g1372 ( 
.A(n_1277),
.B(n_1267),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1292),
.B(n_1238),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1294),
.Y(n_1374)
);

INVx3_ASAP7_75t_L g1375 ( 
.A(n_1271),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1294),
.Y(n_1376)
);

CKINVDCx5p33_ASAP7_75t_R g1377 ( 
.A(n_1272),
.Y(n_1377)
);

NAND2x1_ASAP7_75t_L g1378 ( 
.A(n_1296),
.B(n_1046),
.Y(n_1378)
);

OAI22xp33_ASAP7_75t_L g1379 ( 
.A1(n_1350),
.A2(n_1263),
.B1(n_1265),
.B2(n_1112),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1347),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1318),
.B(n_1262),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_1329),
.Y(n_1382)
);

INVx2_ASAP7_75t_SL g1383 ( 
.A(n_1315),
.Y(n_1383)
);

AO22x2_ASAP7_75t_L g1384 ( 
.A1(n_1360),
.A2(n_1244),
.B1(n_1235),
.B2(n_1242),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_SL g1385 ( 
.A(n_1341),
.B(n_1053),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_1320),
.Y(n_1386)
);

NOR2xp33_ASAP7_75t_L g1387 ( 
.A(n_1368),
.B(n_1264),
.Y(n_1387)
);

BUFx4f_ASAP7_75t_L g1388 ( 
.A(n_1321),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1334),
.B(n_1268),
.Y(n_1389)
);

BUFx3_ASAP7_75t_L g1390 ( 
.A(n_1333),
.Y(n_1390)
);

INVx3_ASAP7_75t_L g1391 ( 
.A(n_1363),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1352),
.B(n_1241),
.Y(n_1392)
);

AO21x2_ASAP7_75t_L g1393 ( 
.A1(n_1344),
.A2(n_919),
.B(n_913),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1336),
.B(n_998),
.Y(n_1394)
);

OAI22xp5_ASAP7_75t_L g1395 ( 
.A1(n_1354),
.A2(n_1081),
.B1(n_1082),
.B2(n_1035),
.Y(n_1395)
);

INVx6_ASAP7_75t_L g1396 ( 
.A(n_1330),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1323),
.Y(n_1397)
);

AND2x2_ASAP7_75t_SL g1398 ( 
.A(n_1365),
.B(n_1371),
.Y(n_1398)
);

BUFx10_ASAP7_75t_L g1399 ( 
.A(n_1377),
.Y(n_1399)
);

NOR2xp33_ASAP7_75t_L g1400 ( 
.A(n_1372),
.B(n_1088),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1342),
.B(n_914),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1326),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1327),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1335),
.B(n_1006),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1358),
.B(n_1006),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1328),
.B(n_974),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1361),
.B(n_894),
.Y(n_1407)
);

NOR2xp33_ASAP7_75t_L g1408 ( 
.A(n_1339),
.B(n_1105),
.Y(n_1408)
);

INVx5_ASAP7_75t_L g1409 ( 
.A(n_1363),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1332),
.B(n_1034),
.Y(n_1410)
);

BUFx6f_ASAP7_75t_L g1411 ( 
.A(n_1325),
.Y(n_1411)
);

INVx4_ASAP7_75t_L g1412 ( 
.A(n_1353),
.Y(n_1412)
);

NAND2xp33_ASAP7_75t_L g1413 ( 
.A(n_1359),
.B(n_889),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_SL g1414 ( 
.A(n_1351),
.B(n_1108),
.Y(n_1414)
);

NOR2xp33_ASAP7_75t_L g1415 ( 
.A(n_1373),
.B(n_1134),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1364),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1366),
.Y(n_1417)
);

AND2x4_ASAP7_75t_L g1418 ( 
.A(n_1343),
.B(n_1153),
.Y(n_1418)
);

INVx4_ASAP7_75t_L g1419 ( 
.A(n_1353),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1370),
.Y(n_1420)
);

INVx6_ASAP7_75t_L g1421 ( 
.A(n_1349),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_SL g1422 ( 
.A(n_1325),
.B(n_1188),
.Y(n_1422)
);

INVxp67_ASAP7_75t_L g1423 ( 
.A(n_1319),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1337),
.B(n_1077),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1338),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1331),
.B(n_1138),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1324),
.B(n_1207),
.Y(n_1427)
);

NAND2xp33_ASAP7_75t_SL g1428 ( 
.A(n_1378),
.B(n_904),
.Y(n_1428)
);

BUFx6f_ASAP7_75t_L g1429 ( 
.A(n_1349),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1345),
.B(n_908),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1346),
.Y(n_1431)
);

BUFx3_ASAP7_75t_L g1432 ( 
.A(n_1369),
.Y(n_1432)
);

NAND2x1p5_ASAP7_75t_L g1433 ( 
.A(n_1375),
.B(n_1015),
.Y(n_1433)
);

INVx4_ASAP7_75t_L g1434 ( 
.A(n_1357),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1348),
.B(n_926),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1314),
.Y(n_1436)
);

OR2x2_ASAP7_75t_L g1437 ( 
.A(n_1340),
.B(n_932),
.Y(n_1437)
);

CKINVDCx5p33_ASAP7_75t_R g1438 ( 
.A(n_1322),
.Y(n_1438)
);

CKINVDCx11_ASAP7_75t_R g1439 ( 
.A(n_1362),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1316),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1317),
.Y(n_1441)
);

OAI22xp33_ASAP7_75t_L g1442 ( 
.A1(n_1367),
.A2(n_948),
.B1(n_954),
.B2(n_945),
.Y(n_1442)
);

INVx2_ASAP7_75t_L g1443 ( 
.A(n_1374),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1376),
.Y(n_1444)
);

INVx2_ASAP7_75t_L g1445 ( 
.A(n_1355),
.Y(n_1445)
);

INVx4_ASAP7_75t_L g1446 ( 
.A(n_1356),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1329),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1318),
.B(n_962),
.Y(n_1448)
);

OR2x6_ASAP7_75t_L g1449 ( 
.A(n_1333),
.B(n_906),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1329),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1318),
.B(n_963),
.Y(n_1451)
);

BUFx2_ASAP7_75t_L g1452 ( 
.A(n_1315),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1347),
.Y(n_1453)
);

INVx4_ASAP7_75t_SL g1454 ( 
.A(n_1333),
.Y(n_1454)
);

NOR2xp33_ASAP7_75t_L g1455 ( 
.A(n_1341),
.B(n_1191),
.Y(n_1455)
);

INVx3_ASAP7_75t_L g1456 ( 
.A(n_1363),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1329),
.Y(n_1457)
);

INVxp67_ASAP7_75t_SL g1458 ( 
.A(n_1319),
.Y(n_1458)
);

NOR2xp33_ASAP7_75t_L g1459 ( 
.A(n_1341),
.B(n_1192),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1347),
.Y(n_1460)
);

AOI22xp5_ASAP7_75t_L g1461 ( 
.A1(n_1350),
.A2(n_972),
.B1(n_1096),
.B2(n_1004),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1347),
.Y(n_1462)
);

OAI22xp33_ASAP7_75t_L g1463 ( 
.A1(n_1350),
.A2(n_990),
.B1(n_992),
.B2(n_964),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1347),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_SL g1465 ( 
.A(n_1341),
.B(n_1206),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1352),
.B(n_993),
.Y(n_1466)
);

OAI21xp33_ASAP7_75t_SL g1467 ( 
.A1(n_1352),
.A2(n_922),
.B(n_920),
.Y(n_1467)
);

BUFx3_ASAP7_75t_L g1468 ( 
.A(n_1333),
.Y(n_1468)
);

INVx5_ASAP7_75t_L g1469 ( 
.A(n_1330),
.Y(n_1469)
);

INVx1_ASAP7_75t_SL g1470 ( 
.A(n_1315),
.Y(n_1470)
);

OR2x6_ASAP7_75t_L g1471 ( 
.A(n_1333),
.B(n_933),
.Y(n_1471)
);

INVx1_ASAP7_75t_SL g1472 ( 
.A(n_1315),
.Y(n_1472)
);

AND2x2_ASAP7_75t_SL g1473 ( 
.A(n_1330),
.B(n_1145),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1329),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1347),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1347),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1329),
.Y(n_1477)
);

BUFx3_ASAP7_75t_L g1478 ( 
.A(n_1333),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1352),
.B(n_1052),
.Y(n_1479)
);

BUFx2_ASAP7_75t_L g1480 ( 
.A(n_1315),
.Y(n_1480)
);

BUFx10_ASAP7_75t_L g1481 ( 
.A(n_1377),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_SL g1482 ( 
.A(n_1341),
.B(n_1200),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1347),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1347),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1329),
.Y(n_1485)
);

INVx4_ASAP7_75t_L g1486 ( 
.A(n_1377),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1347),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1347),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1329),
.Y(n_1489)
);

AND2x4_ASAP7_75t_L g1490 ( 
.A(n_1333),
.B(n_1070),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1329),
.Y(n_1491)
);

AND2x2_ASAP7_75t_SL g1492 ( 
.A(n_1330),
.B(n_878),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_SL g1493 ( 
.A(n_1398),
.B(n_1071),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1408),
.B(n_1075),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_SL g1495 ( 
.A(n_1470),
.B(n_1102),
.Y(n_1495)
);

NOR2xp33_ASAP7_75t_L g1496 ( 
.A(n_1472),
.B(n_1106),
.Y(n_1496)
);

OR2x6_ASAP7_75t_L g1497 ( 
.A(n_1396),
.B(n_1049),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_SL g1498 ( 
.A(n_1383),
.B(n_1113),
.Y(n_1498)
);

CKINVDCx5p33_ASAP7_75t_R g1499 ( 
.A(n_1399),
.Y(n_1499)
);

AOI21xp5_ASAP7_75t_L g1500 ( 
.A1(n_1466),
.A2(n_1203),
.B(n_858),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1397),
.Y(n_1501)
);

INVx2_ASAP7_75t_SL g1502 ( 
.A(n_1388),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1415),
.B(n_1119),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1386),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1402),
.Y(n_1505)
);

NOR2xp33_ASAP7_75t_L g1506 ( 
.A(n_1452),
.B(n_1128),
.Y(n_1506)
);

INVx2_ASAP7_75t_SL g1507 ( 
.A(n_1469),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1403),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_SL g1509 ( 
.A(n_1480),
.B(n_1143),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1380),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1453),
.Y(n_1511)
);

AOI22xp5_ASAP7_75t_L g1512 ( 
.A1(n_1455),
.A2(n_928),
.B1(n_929),
.B2(n_924),
.Y(n_1512)
);

NOR2xp33_ASAP7_75t_L g1513 ( 
.A(n_1400),
.B(n_1154),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1460),
.Y(n_1514)
);

NOR2xp33_ASAP7_75t_L g1515 ( 
.A(n_1385),
.B(n_1175),
.Y(n_1515)
);

OAI22xp5_ASAP7_75t_L g1516 ( 
.A1(n_1479),
.A2(n_1179),
.B1(n_1182),
.B2(n_1177),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1462),
.Y(n_1517)
);

AOI22xp5_ASAP7_75t_L g1518 ( 
.A1(n_1459),
.A2(n_934),
.B1(n_939),
.B2(n_930),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_SL g1519 ( 
.A(n_1463),
.B(n_855),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1394),
.B(n_1201),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_SL g1521 ( 
.A(n_1379),
.B(n_859),
.Y(n_1521)
);

O2A1O1Ixp33_ASAP7_75t_L g1522 ( 
.A1(n_1392),
.A2(n_942),
.B(n_946),
.C(n_943),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1401),
.B(n_1174),
.Y(n_1523)
);

NAND2xp33_ASAP7_75t_L g1524 ( 
.A(n_1428),
.B(n_860),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1389),
.B(n_1181),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1464),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1382),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1447),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1450),
.Y(n_1529)
);

A2O1A1Ixp33_ASAP7_75t_L g1530 ( 
.A1(n_1467),
.A2(n_956),
.B(n_959),
.C(n_957),
.Y(n_1530)
);

BUFx4f_ASAP7_75t_L g1531 ( 
.A(n_1429),
.Y(n_1531)
);

INVx8_ASAP7_75t_L g1532 ( 
.A(n_1469),
.Y(n_1532)
);

XNOR2xp5_ASAP7_75t_L g1533 ( 
.A(n_1473),
.B(n_865),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1407),
.B(n_0),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1475),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1381),
.B(n_1),
.Y(n_1536)
);

BUFx2_ASAP7_75t_L g1537 ( 
.A(n_1390),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1457),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1448),
.B(n_1198),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1451),
.B(n_966),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1474),
.Y(n_1541)
);

INVx3_ASAP7_75t_L g1542 ( 
.A(n_1468),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1476),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1477),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1406),
.B(n_977),
.Y(n_1545)
);

AOI22xp33_ASAP7_75t_L g1546 ( 
.A1(n_1395),
.A2(n_872),
.B1(n_891),
.B2(n_870),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_SL g1547 ( 
.A(n_1411),
.B(n_1410),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1387),
.B(n_980),
.Y(n_1548)
);

OR2x2_ASAP7_75t_L g1549 ( 
.A(n_1437),
.B(n_2),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_SL g1550 ( 
.A(n_1411),
.B(n_866),
.Y(n_1550)
);

HB1xp67_ASAP7_75t_L g1551 ( 
.A(n_1478),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_SL g1552 ( 
.A(n_1424),
.B(n_867),
.Y(n_1552)
);

AND2x2_ASAP7_75t_SL g1553 ( 
.A(n_1492),
.B(n_1090),
.Y(n_1553)
);

CKINVDCx5p33_ASAP7_75t_R g1554 ( 
.A(n_1481),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1404),
.B(n_1185),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1483),
.B(n_986),
.Y(n_1556)
);

NOR2xp33_ASAP7_75t_L g1557 ( 
.A(n_1414),
.B(n_988),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1484),
.B(n_999),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1487),
.B(n_1005),
.Y(n_1559)
);

XOR2x2_ASAP7_75t_L g1560 ( 
.A(n_1422),
.B(n_4),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1488),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1485),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1489),
.B(n_1007),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_SL g1564 ( 
.A(n_1461),
.B(n_869),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1491),
.B(n_1013),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_SL g1566 ( 
.A(n_1486),
.B(n_871),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1458),
.B(n_1025),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_SL g1568 ( 
.A(n_1434),
.B(n_876),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_SL g1569 ( 
.A(n_1446),
.B(n_877),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1405),
.B(n_3),
.Y(n_1570)
);

AOI21xp5_ASAP7_75t_L g1571 ( 
.A1(n_1430),
.A2(n_892),
.B(n_886),
.Y(n_1571)
);

HB1xp67_ASAP7_75t_L g1572 ( 
.A(n_1454),
.Y(n_1572)
);

INVxp67_ASAP7_75t_L g1573 ( 
.A(n_1427),
.Y(n_1573)
);

CKINVDCx5p33_ASAP7_75t_R g1574 ( 
.A(n_1438),
.Y(n_1574)
);

NAND2xp33_ASAP7_75t_L g1575 ( 
.A(n_1465),
.B(n_893),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1416),
.B(n_1178),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1417),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1420),
.Y(n_1578)
);

INVx8_ASAP7_75t_L g1579 ( 
.A(n_1409),
.Y(n_1579)
);

NOR2xp33_ASAP7_75t_L g1580 ( 
.A(n_1482),
.B(n_1030),
.Y(n_1580)
);

NOR3xp33_ASAP7_75t_L g1581 ( 
.A(n_1442),
.B(n_1032),
.C(n_1031),
.Y(n_1581)
);

AOI22xp5_ASAP7_75t_L g1582 ( 
.A1(n_1413),
.A2(n_1043),
.B1(n_1050),
.B2(n_1040),
.Y(n_1582)
);

AOI22xp5_ASAP7_75t_L g1583 ( 
.A1(n_1435),
.A2(n_1078),
.B1(n_1087),
.B2(n_1063),
.Y(n_1583)
);

AND2x6_ASAP7_75t_L g1584 ( 
.A(n_1431),
.B(n_1060),
.Y(n_1584)
);

NOR2xp33_ASAP7_75t_L g1585 ( 
.A(n_1423),
.B(n_1091),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1425),
.Y(n_1586)
);

BUFx3_ASAP7_75t_L g1587 ( 
.A(n_1409),
.Y(n_1587)
);

NOR2xp33_ASAP7_75t_L g1588 ( 
.A(n_1445),
.B(n_1093),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_SL g1589 ( 
.A(n_1432),
.B(n_896),
.Y(n_1589)
);

NOR2xp33_ASAP7_75t_L g1590 ( 
.A(n_1418),
.B(n_1094),
.Y(n_1590)
);

AND2x6_ASAP7_75t_SL g1591 ( 
.A(n_1490),
.B(n_1116),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1441),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_SL g1593 ( 
.A(n_1433),
.B(n_897),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1436),
.Y(n_1594)
);

OAI22xp5_ASAP7_75t_L g1595 ( 
.A1(n_1426),
.A2(n_1124),
.B1(n_1146),
.B2(n_1141),
.Y(n_1595)
);

NOR2xp33_ASAP7_75t_L g1596 ( 
.A(n_1440),
.B(n_1155),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_SL g1597 ( 
.A(n_1429),
.B(n_900),
.Y(n_1597)
);

AOI22xp5_ASAP7_75t_L g1598 ( 
.A1(n_1444),
.A2(n_1159),
.B1(n_1166),
.B2(n_1157),
.Y(n_1598)
);

NOR2xp33_ASAP7_75t_L g1599 ( 
.A(n_1443),
.B(n_1170),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1391),
.B(n_905),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1456),
.B(n_907),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1393),
.Y(n_1602)
);

INVx2_ASAP7_75t_L g1603 ( 
.A(n_1421),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1412),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1419),
.B(n_910),
.Y(n_1605)
);

AOI21xp5_ASAP7_75t_L g1606 ( 
.A1(n_1449),
.A2(n_917),
.B(n_916),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1384),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1471),
.B(n_918),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_SL g1609 ( 
.A(n_1449),
.B(n_921),
.Y(n_1609)
);

CKINVDCx20_ASAP7_75t_R g1610 ( 
.A(n_1439),
.Y(n_1610)
);

NOR2xp33_ASAP7_75t_L g1611 ( 
.A(n_1471),
.B(n_923),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_1386),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1408),
.B(n_925),
.Y(n_1613)
);

AOI22xp33_ASAP7_75t_L g1614 ( 
.A1(n_1395),
.A2(n_885),
.B1(n_915),
.B2(n_912),
.Y(n_1614)
);

NOR2x1p5_ASAP7_75t_L g1615 ( 
.A(n_1486),
.B(n_1060),
.Y(n_1615)
);

NOR2xp67_ASAP7_75t_L g1616 ( 
.A(n_1469),
.B(n_927),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1408),
.B(n_931),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1397),
.Y(n_1618)
);

AOI22xp33_ASAP7_75t_L g1619 ( 
.A1(n_1395),
.A2(n_950),
.B1(n_1140),
.B2(n_1055),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1408),
.B(n_935),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1408),
.B(n_936),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_SL g1622 ( 
.A(n_1398),
.B(n_938),
.Y(n_1622)
);

NOR2xp33_ASAP7_75t_L g1623 ( 
.A(n_1470),
.B(n_941),
.Y(n_1623)
);

NOR2x1p5_ASAP7_75t_L g1624 ( 
.A(n_1486),
.B(n_971),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1397),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1386),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1408),
.B(n_947),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1386),
.Y(n_1628)
);

AOI21xp5_ASAP7_75t_L g1629 ( 
.A1(n_1466),
.A2(n_953),
.B(n_949),
.Y(n_1629)
);

AOI22xp5_ASAP7_75t_L g1630 ( 
.A1(n_1408),
.A2(n_955),
.B1(n_961),
.B2(n_958),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1386),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1397),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1408),
.B(n_965),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1408),
.B(n_967),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1386),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1397),
.Y(n_1636)
);

INVx2_ASAP7_75t_SL g1637 ( 
.A(n_1388),
.Y(n_1637)
);

NOR2xp33_ASAP7_75t_L g1638 ( 
.A(n_1470),
.B(n_970),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1408),
.B(n_973),
.Y(n_1639)
);

INVx1_ASAP7_75t_SL g1640 ( 
.A(n_1470),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1397),
.Y(n_1641)
);

INVx1_ASAP7_75t_SL g1642 ( 
.A(n_1470),
.Y(n_1642)
);

CKINVDCx5p33_ASAP7_75t_R g1643 ( 
.A(n_1399),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1386),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1386),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_SL g1646 ( 
.A(n_1398),
.B(n_976),
.Y(n_1646)
);

NAND3xp33_ASAP7_75t_L g1647 ( 
.A(n_1455),
.B(n_979),
.C(n_978),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1408),
.B(n_985),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1397),
.Y(n_1649)
);

NAND2xp33_ASAP7_75t_L g1650 ( 
.A(n_1397),
.B(n_989),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1408),
.B(n_996),
.Y(n_1651)
);

AOI22xp33_ASAP7_75t_L g1652 ( 
.A1(n_1553),
.A2(n_968),
.B1(n_984),
.B2(n_881),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1640),
.B(n_3),
.Y(n_1653)
);

AOI22xp5_ASAP7_75t_L g1654 ( 
.A1(n_1513),
.A2(n_1000),
.B1(n_1001),
.B2(n_997),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1578),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1586),
.Y(n_1656)
);

INVx2_ASAP7_75t_SL g1657 ( 
.A(n_1579),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_SL g1658 ( 
.A(n_1574),
.B(n_1194),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_SL g1659 ( 
.A(n_1642),
.B(n_1199),
.Y(n_1659)
);

O2A1O1Ixp33_ASAP7_75t_L g1660 ( 
.A1(n_1548),
.A2(n_1033),
.B(n_1038),
.C(n_1018),
.Y(n_1660)
);

HB1xp67_ASAP7_75t_L g1661 ( 
.A(n_1537),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1573),
.B(n_4),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1501),
.Y(n_1663)
);

OR2x4_ASAP7_75t_L g1664 ( 
.A(n_1506),
.B(n_6),
.Y(n_1664)
);

AND2x4_ASAP7_75t_L g1665 ( 
.A(n_1502),
.B(n_1056),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1505),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_SL g1667 ( 
.A(n_1531),
.B(n_1168),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1496),
.B(n_7),
.Y(n_1668)
);

INVx5_ASAP7_75t_L g1669 ( 
.A(n_1532),
.Y(n_1669)
);

BUFx4f_ASAP7_75t_L g1670 ( 
.A(n_1579),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1508),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1618),
.Y(n_1672)
);

BUFx12f_ASAP7_75t_L g1673 ( 
.A(n_1499),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_SL g1674 ( 
.A(n_1637),
.B(n_1169),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1534),
.B(n_7),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1536),
.B(n_8),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1494),
.B(n_9),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_SL g1678 ( 
.A(n_1623),
.B(n_1183),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1638),
.B(n_10),
.Y(n_1679)
);

BUFx8_ASAP7_75t_SL g1680 ( 
.A(n_1610),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1577),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_SL g1682 ( 
.A(n_1542),
.B(n_1184),
.Y(n_1682)
);

NAND2x1p5_ASAP7_75t_L g1683 ( 
.A(n_1587),
.B(n_899),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1503),
.B(n_10),
.Y(n_1684)
);

NAND2x1p5_ASAP7_75t_L g1685 ( 
.A(n_1507),
.B(n_899),
.Y(n_1685)
);

NAND2x1p5_ASAP7_75t_L g1686 ( 
.A(n_1603),
.B(n_899),
.Y(n_1686)
);

NOR2xp33_ASAP7_75t_L g1687 ( 
.A(n_1493),
.B(n_1002),
.Y(n_1687)
);

HB1xp67_ASAP7_75t_L g1688 ( 
.A(n_1551),
.Y(n_1688)
);

INVx3_ASAP7_75t_L g1689 ( 
.A(n_1532),
.Y(n_1689)
);

NAND3xp33_ASAP7_75t_SL g1690 ( 
.A(n_1512),
.B(n_1045),
.C(n_1019),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1625),
.Y(n_1691)
);

NAND2xp33_ASAP7_75t_L g1692 ( 
.A(n_1554),
.B(n_1643),
.Y(n_1692)
);

INVx2_ASAP7_75t_SL g1693 ( 
.A(n_1572),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1570),
.B(n_11),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1632),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1525),
.B(n_1636),
.Y(n_1696)
);

INVx5_ASAP7_75t_L g1697 ( 
.A(n_1497),
.Y(n_1697)
);

INVx5_ASAP7_75t_L g1698 ( 
.A(n_1497),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1641),
.Y(n_1699)
);

INVx2_ASAP7_75t_L g1700 ( 
.A(n_1504),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1649),
.B(n_11),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1510),
.Y(n_1702)
);

AND3x1_ASAP7_75t_L g1703 ( 
.A(n_1611),
.B(n_1069),
.C(n_1059),
.Y(n_1703)
);

INVx3_ASAP7_75t_L g1704 ( 
.A(n_1604),
.Y(n_1704)
);

O2A1O1Ixp33_ASAP7_75t_L g1705 ( 
.A1(n_1530),
.A2(n_1127),
.B(n_1139),
.C(n_1123),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1520),
.B(n_12),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1555),
.B(n_12),
.Y(n_1707)
);

HB1xp67_ASAP7_75t_L g1708 ( 
.A(n_1549),
.Y(n_1708)
);

AND2x4_ASAP7_75t_L g1709 ( 
.A(n_1615),
.B(n_1624),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1511),
.B(n_13),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1590),
.B(n_13),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1527),
.Y(n_1712)
);

INVx4_ASAP7_75t_L g1713 ( 
.A(n_1591),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1514),
.B(n_14),
.Y(n_1714)
);

CKINVDCx5p33_ASAP7_75t_R g1715 ( 
.A(n_1533),
.Y(n_1715)
);

INVx3_ASAP7_75t_L g1716 ( 
.A(n_1592),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1517),
.B(n_14),
.Y(n_1717)
);

AOI22xp33_ASAP7_75t_L g1718 ( 
.A1(n_1557),
.A2(n_1167),
.B1(n_1193),
.B2(n_1165),
.Y(n_1718)
);

AOI22xp5_ASAP7_75t_L g1719 ( 
.A1(n_1581),
.A2(n_1010),
.B1(n_1011),
.B2(n_1008),
.Y(n_1719)
);

AOI22xp33_ASAP7_75t_L g1720 ( 
.A1(n_1607),
.A2(n_1202),
.B1(n_975),
.B2(n_995),
.Y(n_1720)
);

AOI22xp5_ASAP7_75t_L g1721 ( 
.A1(n_1515),
.A2(n_1014),
.B1(n_1026),
.B2(n_1012),
.Y(n_1721)
);

INVx3_ASAP7_75t_L g1722 ( 
.A(n_1528),
.Y(n_1722)
);

INVx2_ASAP7_75t_L g1723 ( 
.A(n_1529),
.Y(n_1723)
);

AOI22xp5_ASAP7_75t_L g1724 ( 
.A1(n_1518),
.A2(n_1029),
.B1(n_1041),
.B2(n_1027),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1526),
.Y(n_1725)
);

AOI22xp33_ASAP7_75t_L g1726 ( 
.A1(n_1546),
.A2(n_975),
.B1(n_995),
.B2(n_951),
.Y(n_1726)
);

AOI22xp5_ASAP7_75t_L g1727 ( 
.A1(n_1580),
.A2(n_1044),
.B1(n_1047),
.B2(n_1042),
.Y(n_1727)
);

OAI22xp5_ASAP7_75t_L g1728 ( 
.A1(n_1613),
.A2(n_1162),
.B1(n_1073),
.B2(n_1086),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1535),
.Y(n_1729)
);

NOR2xp33_ASAP7_75t_R g1730 ( 
.A(n_1650),
.B(n_1048),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1538),
.Y(n_1731)
);

INVx1_ASAP7_75t_SL g1732 ( 
.A(n_1509),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1543),
.Y(n_1733)
);

NOR2x1p5_ASAP7_75t_L g1734 ( 
.A(n_1608),
.B(n_1051),
.Y(n_1734)
);

OR2x6_ASAP7_75t_L g1735 ( 
.A(n_1609),
.B(n_951),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1561),
.B(n_15),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1541),
.Y(n_1737)
);

INVx2_ASAP7_75t_SL g1738 ( 
.A(n_1594),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1544),
.Y(n_1739)
);

NOR2xp33_ASAP7_75t_SL g1740 ( 
.A(n_1616),
.B(n_1190),
.Y(n_1740)
);

INVx2_ASAP7_75t_L g1741 ( 
.A(n_1562),
.Y(n_1741)
);

BUFx2_ASAP7_75t_SL g1742 ( 
.A(n_1560),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_SL g1743 ( 
.A(n_1617),
.B(n_1204),
.Y(n_1743)
);

BUFx2_ASAP7_75t_L g1744 ( 
.A(n_1584),
.Y(n_1744)
);

CKINVDCx20_ASAP7_75t_R g1745 ( 
.A(n_1622),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1612),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1620),
.B(n_15),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1621),
.B(n_16),
.Y(n_1748)
);

INVx3_ASAP7_75t_L g1749 ( 
.A(n_1626),
.Y(n_1749)
);

OAI22xp5_ASAP7_75t_SL g1750 ( 
.A1(n_1614),
.A2(n_1058),
.B1(n_1100),
.B2(n_1080),
.Y(n_1750)
);

INVx3_ASAP7_75t_SL g1751 ( 
.A(n_1495),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1628),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1627),
.B(n_16),
.Y(n_1753)
);

INVx2_ASAP7_75t_L g1754 ( 
.A(n_1631),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_SL g1755 ( 
.A(n_1633),
.B(n_1144),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1634),
.B(n_17),
.Y(n_1756)
);

BUFx2_ASAP7_75t_L g1757 ( 
.A(n_1584),
.Y(n_1757)
);

HB1xp67_ASAP7_75t_L g1758 ( 
.A(n_1635),
.Y(n_1758)
);

CKINVDCx11_ASAP7_75t_R g1759 ( 
.A(n_1644),
.Y(n_1759)
);

AND2x4_ASAP7_75t_SL g1760 ( 
.A(n_1645),
.B(n_1582),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1539),
.B(n_17),
.Y(n_1761)
);

INVxp67_ASAP7_75t_L g1762 ( 
.A(n_1585),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_SL g1763 ( 
.A(n_1639),
.B(n_1149),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1563),
.Y(n_1764)
);

HB1xp67_ASAP7_75t_L g1765 ( 
.A(n_1547),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1648),
.B(n_18),
.Y(n_1766)
);

INVx3_ASAP7_75t_L g1767 ( 
.A(n_1584),
.Y(n_1767)
);

CKINVDCx5p33_ASAP7_75t_R g1768 ( 
.A(n_1646),
.Y(n_1768)
);

AOI22xp33_ASAP7_75t_L g1769 ( 
.A1(n_1619),
.A2(n_975),
.B1(n_995),
.B2(n_951),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1762),
.B(n_1651),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1656),
.Y(n_1771)
);

INVx2_ASAP7_75t_L g1772 ( 
.A(n_1681),
.Y(n_1772)
);

NAND2x1p5_ASAP7_75t_L g1773 ( 
.A(n_1670),
.B(n_1593),
.Y(n_1773)
);

OR2x2_ASAP7_75t_L g1774 ( 
.A(n_1708),
.B(n_1661),
.Y(n_1774)
);

AND2x4_ASAP7_75t_L g1775 ( 
.A(n_1669),
.B(n_1498),
.Y(n_1775)
);

AND2x4_ASAP7_75t_L g1776 ( 
.A(n_1669),
.B(n_1589),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1663),
.Y(n_1777)
);

INVx2_ASAP7_75t_L g1778 ( 
.A(n_1655),
.Y(n_1778)
);

INVx2_ASAP7_75t_L g1779 ( 
.A(n_1700),
.Y(n_1779)
);

BUFx6f_ASAP7_75t_L g1780 ( 
.A(n_1759),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_SL g1781 ( 
.A(n_1697),
.B(n_1647),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1696),
.B(n_1523),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1666),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1671),
.Y(n_1784)
);

INVx2_ASAP7_75t_L g1785 ( 
.A(n_1712),
.Y(n_1785)
);

INVx4_ASAP7_75t_L g1786 ( 
.A(n_1673),
.Y(n_1786)
);

BUFx4f_ASAP7_75t_L g1787 ( 
.A(n_1751),
.Y(n_1787)
);

INVx2_ASAP7_75t_L g1788 ( 
.A(n_1723),
.Y(n_1788)
);

AND2x4_ASAP7_75t_L g1789 ( 
.A(n_1697),
.B(n_1597),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1672),
.Y(n_1790)
);

INVx2_ASAP7_75t_L g1791 ( 
.A(n_1731),
.Y(n_1791)
);

AND2x2_ASAP7_75t_L g1792 ( 
.A(n_1653),
.B(n_1540),
.Y(n_1792)
);

INVx4_ASAP7_75t_L g1793 ( 
.A(n_1698),
.Y(n_1793)
);

NOR2xp33_ASAP7_75t_L g1794 ( 
.A(n_1732),
.B(n_1630),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1691),
.Y(n_1795)
);

BUFx6f_ASAP7_75t_L g1796 ( 
.A(n_1657),
.Y(n_1796)
);

BUFx3_ASAP7_75t_L g1797 ( 
.A(n_1689),
.Y(n_1797)
);

CKINVDCx5p33_ASAP7_75t_R g1798 ( 
.A(n_1680),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1764),
.B(n_1545),
.Y(n_1799)
);

AND2x6_ASAP7_75t_SL g1800 ( 
.A(n_1709),
.B(n_1735),
.Y(n_1800)
);

BUFx2_ASAP7_75t_L g1801 ( 
.A(n_1688),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1761),
.B(n_1596),
.Y(n_1802)
);

BUFx2_ASAP7_75t_SL g1803 ( 
.A(n_1698),
.Y(n_1803)
);

CKINVDCx5p33_ASAP7_75t_R g1804 ( 
.A(n_1715),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1695),
.Y(n_1805)
);

BUFx6f_ASAP7_75t_L g1806 ( 
.A(n_1693),
.Y(n_1806)
);

OR2x2_ASAP7_75t_L g1807 ( 
.A(n_1738),
.B(n_1556),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1699),
.Y(n_1808)
);

INVx2_ASAP7_75t_L g1809 ( 
.A(n_1737),
.Y(n_1809)
);

A2O1A1Ixp33_ASAP7_75t_L g1810 ( 
.A1(n_1677),
.A2(n_1522),
.B(n_1583),
.C(n_1500),
.Y(n_1810)
);

INVx1_ASAP7_75t_SL g1811 ( 
.A(n_1745),
.Y(n_1811)
);

INVx2_ASAP7_75t_L g1812 ( 
.A(n_1741),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1702),
.B(n_1725),
.Y(n_1813)
);

BUFx4f_ASAP7_75t_L g1814 ( 
.A(n_1735),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1729),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1733),
.B(n_1588),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1711),
.B(n_1599),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1758),
.Y(n_1818)
);

BUFx6f_ASAP7_75t_L g1819 ( 
.A(n_1683),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1707),
.B(n_1516),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_L g1821 ( 
.A(n_1679),
.B(n_1558),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_SL g1822 ( 
.A(n_1703),
.B(n_1567),
.Y(n_1822)
);

INVx1_ASAP7_75t_SL g1823 ( 
.A(n_1768),
.Y(n_1823)
);

BUFx3_ASAP7_75t_L g1824 ( 
.A(n_1704),
.Y(n_1824)
);

NOR2xp33_ASAP7_75t_L g1825 ( 
.A(n_1678),
.B(n_1564),
.Y(n_1825)
);

BUFx6f_ASAP7_75t_L g1826 ( 
.A(n_1716),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1739),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_L g1828 ( 
.A(n_1668),
.B(n_1559),
.Y(n_1828)
);

OR2x2_ASAP7_75t_L g1829 ( 
.A(n_1742),
.B(n_1576),
.Y(n_1829)
);

BUFx6f_ASAP7_75t_L g1830 ( 
.A(n_1722),
.Y(n_1830)
);

OAI21xp33_ASAP7_75t_L g1831 ( 
.A1(n_1684),
.A2(n_1519),
.B(n_1575),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1706),
.B(n_1598),
.Y(n_1832)
);

OR2x2_ASAP7_75t_L g1833 ( 
.A(n_1676),
.B(n_1565),
.Y(n_1833)
);

INVx2_ASAP7_75t_SL g1834 ( 
.A(n_1734),
.Y(n_1834)
);

NAND2x1p5_ASAP7_75t_L g1835 ( 
.A(n_1744),
.B(n_1566),
.Y(n_1835)
);

INVx2_ASAP7_75t_L g1836 ( 
.A(n_1754),
.Y(n_1836)
);

NOR2xp67_ASAP7_75t_L g1837 ( 
.A(n_1749),
.B(n_1605),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1746),
.Y(n_1838)
);

INVxp67_ASAP7_75t_L g1839 ( 
.A(n_1662),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1752),
.Y(n_1840)
);

OAI22xp33_ASAP7_75t_L g1841 ( 
.A1(n_1664),
.A2(n_1521),
.B1(n_1595),
.B2(n_1600),
.Y(n_1841)
);

INVxp67_ASAP7_75t_L g1842 ( 
.A(n_1765),
.Y(n_1842)
);

INVx5_ASAP7_75t_L g1843 ( 
.A(n_1713),
.Y(n_1843)
);

INVx2_ASAP7_75t_L g1844 ( 
.A(n_1701),
.Y(n_1844)
);

INVx3_ASAP7_75t_L g1845 ( 
.A(n_1685),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1675),
.B(n_1584),
.Y(n_1846)
);

OR2x2_ASAP7_75t_L g1847 ( 
.A(n_1710),
.B(n_1601),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1694),
.B(n_1606),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_SL g1849 ( 
.A(n_1730),
.B(n_1552),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1652),
.B(n_1568),
.Y(n_1850)
);

HB1xp67_ASAP7_75t_L g1851 ( 
.A(n_1757),
.Y(n_1851)
);

NAND2x1p5_ASAP7_75t_L g1852 ( 
.A(n_1767),
.B(n_1569),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_L g1853 ( 
.A(n_1727),
.B(n_1550),
.Y(n_1853)
);

INVx2_ASAP7_75t_L g1854 ( 
.A(n_1714),
.Y(n_1854)
);

INVx2_ASAP7_75t_L g1855 ( 
.A(n_1717),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1760),
.B(n_1629),
.Y(n_1856)
);

OR2x2_ASAP7_75t_L g1857 ( 
.A(n_1736),
.B(n_1602),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_L g1858 ( 
.A(n_1687),
.B(n_1571),
.Y(n_1858)
);

CKINVDCx8_ASAP7_75t_R g1859 ( 
.A(n_1665),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_SL g1860 ( 
.A(n_1747),
.B(n_1163),
.Y(n_1860)
);

AOI22xp33_ASAP7_75t_L g1861 ( 
.A1(n_1718),
.A2(n_1524),
.B1(n_1024),
.B2(n_1107),
.Y(n_1861)
);

CKINVDCx5p33_ASAP7_75t_R g1862 ( 
.A(n_1658),
.Y(n_1862)
);

BUFx12f_ASAP7_75t_L g1863 ( 
.A(n_1686),
.Y(n_1863)
);

OAI22xp5_ASAP7_75t_L g1864 ( 
.A1(n_1748),
.A2(n_1061),
.B1(n_1064),
.B2(n_1054),
.Y(n_1864)
);

BUFx5_ASAP7_75t_L g1865 ( 
.A(n_1740),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_SL g1866 ( 
.A(n_1753),
.B(n_1205),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1654),
.B(n_18),
.Y(n_1867)
);

BUFx3_ASAP7_75t_L g1868 ( 
.A(n_1756),
.Y(n_1868)
);

INVx2_ASAP7_75t_L g1869 ( 
.A(n_1766),
.Y(n_1869)
);

AND3x1_ASAP7_75t_SL g1870 ( 
.A(n_1692),
.B(n_19),
.C(n_20),
.Y(n_1870)
);

INVx2_ASAP7_75t_SL g1871 ( 
.A(n_1667),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1721),
.B(n_1719),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1705),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_SL g1874 ( 
.A(n_1750),
.B(n_1067),
.Y(n_1874)
);

NOR2xp33_ASAP7_75t_L g1875 ( 
.A(n_1659),
.B(n_1068),
.Y(n_1875)
);

CKINVDCx5p33_ASAP7_75t_R g1876 ( 
.A(n_1674),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1724),
.B(n_19),
.Y(n_1877)
);

CKINVDCx5p33_ASAP7_75t_R g1878 ( 
.A(n_1682),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_L g1879 ( 
.A(n_1728),
.B(n_20),
.Y(n_1879)
);

NAND2x1_ASAP7_75t_L g1880 ( 
.A(n_1720),
.B(n_1017),
.Y(n_1880)
);

BUFx12f_ASAP7_75t_L g1881 ( 
.A(n_1690),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1743),
.B(n_21),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1660),
.Y(n_1883)
);

AOI22xp5_ASAP7_75t_L g1884 ( 
.A1(n_1755),
.A2(n_1763),
.B1(n_1769),
.B2(n_1726),
.Y(n_1884)
);

INVx2_ASAP7_75t_L g1885 ( 
.A(n_1656),
.Y(n_1885)
);

BUFx12f_ASAP7_75t_L g1886 ( 
.A(n_1759),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1656),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1656),
.Y(n_1888)
);

INVx2_ASAP7_75t_L g1889 ( 
.A(n_1656),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_L g1890 ( 
.A(n_1762),
.B(n_21),
.Y(n_1890)
);

INVx2_ASAP7_75t_SL g1891 ( 
.A(n_1670),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_L g1892 ( 
.A(n_1762),
.B(n_22),
.Y(n_1892)
);

BUFx6f_ASAP7_75t_L g1893 ( 
.A(n_1670),
.Y(n_1893)
);

AOI22xp5_ASAP7_75t_L g1894 ( 
.A1(n_1762),
.A2(n_1076),
.B1(n_1079),
.B2(n_1074),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_L g1895 ( 
.A(n_1762),
.B(n_22),
.Y(n_1895)
);

INVxp67_ASAP7_75t_SL g1896 ( 
.A(n_1688),
.Y(n_1896)
);

NOR2xp67_ASAP7_75t_L g1897 ( 
.A(n_1697),
.B(n_282),
.Y(n_1897)
);

BUFx3_ASAP7_75t_L g1898 ( 
.A(n_1893),
.Y(n_1898)
);

OAI21x1_ASAP7_75t_L g1899 ( 
.A1(n_1873),
.A2(n_284),
.B(n_283),
.Y(n_1899)
);

AND2x2_ASAP7_75t_L g1900 ( 
.A(n_1792),
.B(n_23),
.Y(n_1900)
);

INVx2_ASAP7_75t_L g1901 ( 
.A(n_1772),
.Y(n_1901)
);

NOR2xp67_ASAP7_75t_L g1902 ( 
.A(n_1793),
.B(n_285),
.Y(n_1902)
);

OA22x2_ASAP7_75t_L g1903 ( 
.A1(n_1802),
.A2(n_1084),
.B1(n_1085),
.B2(n_1083),
.Y(n_1903)
);

BUFx10_ASAP7_75t_L g1904 ( 
.A(n_1798),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1782),
.B(n_23),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1817),
.B(n_24),
.Y(n_1906)
);

AOI21xp5_ASAP7_75t_L g1907 ( 
.A1(n_1858),
.A2(n_1024),
.B(n_1017),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1799),
.B(n_24),
.Y(n_1908)
);

OAI21x1_ASAP7_75t_L g1909 ( 
.A1(n_1856),
.A2(n_1883),
.B(n_1857),
.Y(n_1909)
);

AOI21xp5_ASAP7_75t_L g1910 ( 
.A1(n_1831),
.A2(n_1024),
.B(n_1017),
.Y(n_1910)
);

OAI21x1_ASAP7_75t_L g1911 ( 
.A1(n_1813),
.A2(n_287),
.B(n_286),
.Y(n_1911)
);

AOI21x1_ASAP7_75t_L g1912 ( 
.A1(n_1822),
.A2(n_1136),
.B(n_1107),
.Y(n_1912)
);

AOI21xp5_ASAP7_75t_L g1913 ( 
.A1(n_1810),
.A2(n_1136),
.B(n_1107),
.Y(n_1913)
);

NAND2x1p5_ASAP7_75t_L g1914 ( 
.A(n_1787),
.B(n_1136),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1771),
.Y(n_1915)
);

AOI21xp5_ASAP7_75t_L g1916 ( 
.A1(n_1820),
.A2(n_1095),
.B(n_1092),
.Y(n_1916)
);

OAI21x1_ASAP7_75t_L g1917 ( 
.A1(n_1777),
.A2(n_289),
.B(n_288),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1887),
.Y(n_1918)
);

BUFx2_ASAP7_75t_SL g1919 ( 
.A(n_1893),
.Y(n_1919)
);

NOR2x1_ASAP7_75t_L g1920 ( 
.A(n_1868),
.B(n_1097),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1888),
.Y(n_1921)
);

OAI21x1_ASAP7_75t_L g1922 ( 
.A1(n_1783),
.A2(n_1790),
.B(n_1784),
.Y(n_1922)
);

OAI21x1_ASAP7_75t_L g1923 ( 
.A1(n_1795),
.A2(n_292),
.B(n_291),
.Y(n_1923)
);

AOI21xp5_ASAP7_75t_L g1924 ( 
.A1(n_1872),
.A2(n_1103),
.B(n_1098),
.Y(n_1924)
);

AND2x2_ASAP7_75t_L g1925 ( 
.A(n_1794),
.B(n_25),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1816),
.B(n_25),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_SL g1927 ( 
.A(n_1865),
.B(n_1109),
.Y(n_1927)
);

OAI21x1_ASAP7_75t_L g1928 ( 
.A1(n_1805),
.A2(n_294),
.B(n_293),
.Y(n_1928)
);

BUFx2_ASAP7_75t_L g1929 ( 
.A(n_1801),
.Y(n_1929)
);

INVx5_ASAP7_75t_L g1930 ( 
.A(n_1800),
.Y(n_1930)
);

AND2x2_ASAP7_75t_L g1931 ( 
.A(n_1896),
.B(n_26),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_L g1932 ( 
.A(n_1770),
.B(n_26),
.Y(n_1932)
);

NOR2xp33_ASAP7_75t_L g1933 ( 
.A(n_1804),
.B(n_27),
.Y(n_1933)
);

AOI21xp5_ASAP7_75t_L g1934 ( 
.A1(n_1821),
.A2(n_1111),
.B(n_1110),
.Y(n_1934)
);

AND2x2_ASAP7_75t_L g1935 ( 
.A(n_1774),
.B(n_27),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1808),
.Y(n_1936)
);

OAI21x1_ASAP7_75t_L g1937 ( 
.A1(n_1815),
.A2(n_296),
.B(n_295),
.Y(n_1937)
);

A2O1A1Ixp33_ASAP7_75t_L g1938 ( 
.A1(n_1832),
.A2(n_1115),
.B(n_1117),
.C(n_1114),
.Y(n_1938)
);

HB1xp67_ASAP7_75t_L g1939 ( 
.A(n_1851),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_L g1940 ( 
.A(n_1828),
.B(n_28),
.Y(n_1940)
);

AND2x2_ASAP7_75t_L g1941 ( 
.A(n_1811),
.B(n_29),
.Y(n_1941)
);

OAI21x1_ASAP7_75t_L g1942 ( 
.A1(n_1869),
.A2(n_298),
.B(n_297),
.Y(n_1942)
);

AO31x2_ASAP7_75t_L g1943 ( 
.A1(n_1844),
.A2(n_300),
.A3(n_301),
.B(n_299),
.Y(n_1943)
);

AO31x2_ASAP7_75t_L g1944 ( 
.A1(n_1854),
.A2(n_305),
.A3(n_306),
.B(n_304),
.Y(n_1944)
);

INVx2_ASAP7_75t_L g1945 ( 
.A(n_1885),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_SL g1946 ( 
.A(n_1865),
.B(n_1120),
.Y(n_1946)
);

INVx5_ASAP7_75t_L g1947 ( 
.A(n_1886),
.Y(n_1947)
);

OAI21x1_ASAP7_75t_L g1948 ( 
.A1(n_1852),
.A2(n_311),
.B(n_309),
.Y(n_1948)
);

AO31x2_ASAP7_75t_L g1949 ( 
.A1(n_1855),
.A2(n_314),
.A3(n_316),
.B(n_312),
.Y(n_1949)
);

OAI21xp5_ASAP7_75t_L g1950 ( 
.A1(n_1839),
.A2(n_1125),
.B(n_1121),
.Y(n_1950)
);

AOI21xp5_ASAP7_75t_L g1951 ( 
.A1(n_1848),
.A2(n_1129),
.B(n_1126),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1827),
.Y(n_1952)
);

OAI21xp5_ASAP7_75t_L g1953 ( 
.A1(n_1879),
.A2(n_1131),
.B(n_1130),
.Y(n_1953)
);

INVx3_ASAP7_75t_L g1954 ( 
.A(n_1863),
.Y(n_1954)
);

OAI21x1_ASAP7_75t_L g1955 ( 
.A1(n_1838),
.A2(n_320),
.B(n_317),
.Y(n_1955)
);

BUFx3_ASAP7_75t_L g1956 ( 
.A(n_1806),
.Y(n_1956)
);

OAI21x1_ASAP7_75t_L g1957 ( 
.A1(n_1840),
.A2(n_1846),
.B(n_1835),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_L g1958 ( 
.A(n_1807),
.B(n_29),
.Y(n_1958)
);

INVx1_ASAP7_75t_SL g1959 ( 
.A(n_1823),
.Y(n_1959)
);

NOR2x1_ASAP7_75t_SL g1960 ( 
.A(n_1803),
.B(n_30),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_L g1961 ( 
.A(n_1865),
.B(n_30),
.Y(n_1961)
);

AOI221xp5_ASAP7_75t_SL g1962 ( 
.A1(n_1841),
.A2(n_1867),
.B1(n_1877),
.B2(n_1895),
.C(n_1892),
.Y(n_1962)
);

INVx4_ASAP7_75t_L g1963 ( 
.A(n_1780),
.Y(n_1963)
);

INVx2_ASAP7_75t_L g1964 ( 
.A(n_1889),
.Y(n_1964)
);

OAI21xp5_ASAP7_75t_L g1965 ( 
.A1(n_1847),
.A2(n_1135),
.B(n_1132),
.Y(n_1965)
);

AOI21xp5_ASAP7_75t_L g1966 ( 
.A1(n_1860),
.A2(n_1147),
.B(n_1137),
.Y(n_1966)
);

INVx2_ASAP7_75t_L g1967 ( 
.A(n_1778),
.Y(n_1967)
);

OAI21x1_ASAP7_75t_SL g1968 ( 
.A1(n_1882),
.A2(n_31),
.B(n_32),
.Y(n_1968)
);

NOR2xp33_ASAP7_75t_L g1969 ( 
.A(n_1862),
.B(n_31),
.Y(n_1969)
);

OAI21x1_ASAP7_75t_L g1970 ( 
.A1(n_1779),
.A2(n_325),
.B(n_321),
.Y(n_1970)
);

OAI21xp5_ASAP7_75t_L g1971 ( 
.A1(n_1833),
.A2(n_1152),
.B(n_1151),
.Y(n_1971)
);

OAI21x1_ASAP7_75t_L g1972 ( 
.A1(n_1785),
.A2(n_327),
.B(n_326),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_L g1973 ( 
.A(n_1818),
.B(n_32),
.Y(n_1973)
);

AND2x4_ASAP7_75t_L g1974 ( 
.A(n_1891),
.B(n_33),
.Y(n_1974)
);

AO31x2_ASAP7_75t_L g1975 ( 
.A1(n_1788),
.A2(n_333),
.A3(n_334),
.B(n_328),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_L g1976 ( 
.A(n_1829),
.B(n_33),
.Y(n_1976)
);

NAND2xp5_ASAP7_75t_L g1977 ( 
.A(n_1842),
.B(n_34),
.Y(n_1977)
);

AO31x2_ASAP7_75t_L g1978 ( 
.A1(n_1791),
.A2(n_336),
.A3(n_337),
.B(n_335),
.Y(n_1978)
);

INVx3_ASAP7_75t_L g1979 ( 
.A(n_1898),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_L g1980 ( 
.A(n_1929),
.B(n_1824),
.Y(n_1980)
);

INVx3_ASAP7_75t_L g1981 ( 
.A(n_1956),
.Y(n_1981)
);

HB1xp67_ASAP7_75t_L g1982 ( 
.A(n_1939),
.Y(n_1982)
);

AND2x6_ASAP7_75t_L g1983 ( 
.A(n_1961),
.B(n_1819),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1936),
.Y(n_1984)
);

AND2x4_ASAP7_75t_L g1985 ( 
.A(n_1930),
.B(n_1780),
.Y(n_1985)
);

OAI22xp33_ASAP7_75t_L g1986 ( 
.A1(n_1925),
.A2(n_1814),
.B1(n_1850),
.B2(n_1853),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1922),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1952),
.Y(n_1988)
);

AND2x2_ASAP7_75t_L g1989 ( 
.A(n_1900),
.B(n_1935),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_L g1990 ( 
.A(n_1931),
.B(n_1890),
.Y(n_1990)
);

OAI22xp5_ASAP7_75t_SL g1991 ( 
.A1(n_1947),
.A2(n_1878),
.B1(n_1876),
.B2(n_1881),
.Y(n_1991)
);

OR2x6_ASAP7_75t_L g1992 ( 
.A(n_1919),
.B(n_1786),
.Y(n_1992)
);

AOI21xp5_ASAP7_75t_L g1993 ( 
.A1(n_1913),
.A2(n_1866),
.B(n_1825),
.Y(n_1993)
);

OAI22xp5_ASAP7_75t_L g1994 ( 
.A1(n_1932),
.A2(n_1894),
.B1(n_1884),
.B2(n_1871),
.Y(n_1994)
);

AOI21xp5_ASAP7_75t_L g1995 ( 
.A1(n_1910),
.A2(n_1861),
.B(n_1849),
.Y(n_1995)
);

AND2x2_ASAP7_75t_L g1996 ( 
.A(n_1941),
.B(n_1806),
.Y(n_1996)
);

INVx2_ASAP7_75t_L g1997 ( 
.A(n_1901),
.Y(n_1997)
);

O2A1O1Ixp33_ASAP7_75t_L g1998 ( 
.A1(n_1965),
.A2(n_1874),
.B(n_1864),
.C(n_1781),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_L g1999 ( 
.A(n_1905),
.B(n_1826),
.Y(n_1999)
);

CKINVDCx20_ASAP7_75t_R g2000 ( 
.A(n_1947),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_L g2001 ( 
.A(n_1962),
.B(n_1826),
.Y(n_2001)
);

INVxp67_ASAP7_75t_L g2002 ( 
.A(n_1906),
.Y(n_2002)
);

BUFx6f_ASAP7_75t_L g2003 ( 
.A(n_1954),
.Y(n_2003)
);

AOI22xp33_ASAP7_75t_L g2004 ( 
.A1(n_1903),
.A2(n_1836),
.B1(n_1809),
.B2(n_1812),
.Y(n_2004)
);

BUFx2_ASAP7_75t_L g2005 ( 
.A(n_1957),
.Y(n_2005)
);

BUFx3_ASAP7_75t_L g2006 ( 
.A(n_1904),
.Y(n_2006)
);

OAI22xp5_ASAP7_75t_L g2007 ( 
.A1(n_1971),
.A2(n_1773),
.B1(n_1837),
.B2(n_1875),
.Y(n_2007)
);

BUFx2_ASAP7_75t_L g2008 ( 
.A(n_1959),
.Y(n_2008)
);

OA21x2_ASAP7_75t_L g2009 ( 
.A1(n_1909),
.A2(n_1907),
.B(n_1899),
.Y(n_2009)
);

BUFx12f_ASAP7_75t_L g2010 ( 
.A(n_1963),
.Y(n_2010)
);

CKINVDCx16_ASAP7_75t_R g2011 ( 
.A(n_1969),
.Y(n_2011)
);

HB1xp67_ASAP7_75t_L g2012 ( 
.A(n_1915),
.Y(n_2012)
);

OR2x2_ASAP7_75t_L g2013 ( 
.A(n_1918),
.B(n_1830),
.Y(n_2013)
);

CKINVDCx16_ASAP7_75t_R g2014 ( 
.A(n_1933),
.Y(n_2014)
);

BUFx6f_ASAP7_75t_L g2015 ( 
.A(n_1930),
.Y(n_2015)
);

INVx2_ASAP7_75t_L g2016 ( 
.A(n_1945),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_L g2017 ( 
.A(n_1908),
.B(n_1921),
.Y(n_2017)
);

BUFx3_ASAP7_75t_L g2018 ( 
.A(n_1914),
.Y(n_2018)
);

AOI21xp5_ASAP7_75t_L g2019 ( 
.A1(n_1951),
.A2(n_1880),
.B(n_1776),
.Y(n_2019)
);

AOI21xp5_ASAP7_75t_L g2020 ( 
.A1(n_1924),
.A2(n_1897),
.B(n_1775),
.Y(n_2020)
);

CKINVDCx5p33_ASAP7_75t_R g2021 ( 
.A(n_1974),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1964),
.Y(n_2022)
);

AND2x2_ASAP7_75t_L g2023 ( 
.A(n_1976),
.B(n_1830),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_L g2024 ( 
.A(n_1926),
.B(n_1789),
.Y(n_2024)
);

INVx2_ASAP7_75t_L g2025 ( 
.A(n_1967),
.Y(n_2025)
);

BUFx4f_ASAP7_75t_L g2026 ( 
.A(n_1960),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1973),
.Y(n_2027)
);

INVx2_ASAP7_75t_L g2028 ( 
.A(n_1997),
.Y(n_2028)
);

BUFx12f_ASAP7_75t_L g2029 ( 
.A(n_2015),
.Y(n_2029)
);

OAI22xp5_ASAP7_75t_L g2030 ( 
.A1(n_2014),
.A2(n_1938),
.B1(n_1940),
.B2(n_1977),
.Y(n_2030)
);

AND2x4_ASAP7_75t_L g2031 ( 
.A(n_2008),
.B(n_1843),
.Y(n_2031)
);

AND2x2_ASAP7_75t_L g2032 ( 
.A(n_1989),
.B(n_1982),
.Y(n_2032)
);

INVxp67_ASAP7_75t_L g2033 ( 
.A(n_1980),
.Y(n_2033)
);

OR2x6_ASAP7_75t_SL g2034 ( 
.A(n_2021),
.B(n_1958),
.Y(n_2034)
);

OAI211xp5_ASAP7_75t_L g2035 ( 
.A1(n_2001),
.A2(n_1953),
.B(n_1950),
.C(n_1916),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_L g2036 ( 
.A(n_2012),
.B(n_1920),
.Y(n_2036)
);

BUFx6f_ASAP7_75t_L g2037 ( 
.A(n_1992),
.Y(n_2037)
);

OR2x2_ASAP7_75t_L g2038 ( 
.A(n_1984),
.B(n_1834),
.Y(n_2038)
);

AND2x4_ASAP7_75t_L g2039 ( 
.A(n_1981),
.B(n_1843),
.Y(n_2039)
);

NAND2xp5_ASAP7_75t_L g2040 ( 
.A(n_2017),
.B(n_2027),
.Y(n_2040)
);

AOI21xp5_ASAP7_75t_SL g2041 ( 
.A1(n_1993),
.A2(n_1946),
.B(n_1927),
.Y(n_2041)
);

AND2x2_ASAP7_75t_L g2042 ( 
.A(n_1996),
.B(n_1796),
.Y(n_2042)
);

O2A1O1Ixp33_ASAP7_75t_L g2043 ( 
.A1(n_1994),
.A2(n_1968),
.B(n_1934),
.C(n_1966),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_L g2044 ( 
.A(n_1988),
.B(n_34),
.Y(n_2044)
);

OA21x2_ASAP7_75t_L g2045 ( 
.A1(n_2005),
.A2(n_1911),
.B(n_1917),
.Y(n_2045)
);

A2O1A1Ixp33_ASAP7_75t_SL g2046 ( 
.A1(n_1979),
.A2(n_1870),
.B(n_1845),
.C(n_1797),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_L g2047 ( 
.A(n_2002),
.B(n_35),
.Y(n_2047)
);

AOI21xp5_ASAP7_75t_L g2048 ( 
.A1(n_2009),
.A2(n_1955),
.B(n_1928),
.Y(n_2048)
);

A2O1A1Ixp33_ASAP7_75t_SL g2049 ( 
.A1(n_1998),
.A2(n_1796),
.B(n_37),
.C(n_35),
.Y(n_2049)
);

OR2x2_ASAP7_75t_L g2050 ( 
.A(n_1990),
.B(n_1943),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_2022),
.Y(n_2051)
);

A2O1A1Ixp33_ASAP7_75t_L g2052 ( 
.A1(n_2020),
.A2(n_1902),
.B(n_1948),
.C(n_1937),
.Y(n_2052)
);

HB1xp67_ASAP7_75t_L g2053 ( 
.A(n_1987),
.Y(n_2053)
);

BUFx6f_ASAP7_75t_L g2054 ( 
.A(n_1992),
.Y(n_2054)
);

A2O1A1Ixp33_ASAP7_75t_L g2055 ( 
.A1(n_2007),
.A2(n_1923),
.B(n_1942),
.C(n_1970),
.Y(n_2055)
);

A2O1A1Ixp33_ASAP7_75t_SL g2056 ( 
.A1(n_1999),
.A2(n_38),
.B(n_36),
.C(n_37),
.Y(n_2056)
);

INVx2_ASAP7_75t_L g2057 ( 
.A(n_2016),
.Y(n_2057)
);

O2A1O1Ixp33_ASAP7_75t_L g2058 ( 
.A1(n_1986),
.A2(n_1859),
.B(n_40),
.C(n_38),
.Y(n_2058)
);

HB1xp67_ASAP7_75t_L g2059 ( 
.A(n_2013),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_2025),
.Y(n_2060)
);

NOR2xp67_ASAP7_75t_L g2061 ( 
.A(n_2015),
.B(n_1912),
.Y(n_2061)
);

OAI22xp5_ASAP7_75t_L g2062 ( 
.A1(n_2011),
.A2(n_1819),
.B1(n_1161),
.B2(n_1171),
.Y(n_2062)
);

AND2x4_ASAP7_75t_L g2063 ( 
.A(n_1985),
.B(n_1943),
.Y(n_2063)
);

AND2x2_ASAP7_75t_L g2064 ( 
.A(n_2023),
.B(n_1949),
.Y(n_2064)
);

OR2x2_ASAP7_75t_L g2065 ( 
.A(n_2024),
.B(n_1944),
.Y(n_2065)
);

NAND2x1p5_ASAP7_75t_L g2066 ( 
.A(n_2018),
.B(n_1972),
.Y(n_2066)
);

OAI21xp5_ASAP7_75t_L g2067 ( 
.A1(n_1995),
.A2(n_1173),
.B(n_1156),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_1983),
.Y(n_2068)
);

NAND2xp5_ASAP7_75t_L g2069 ( 
.A(n_1983),
.B(n_39),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_1983),
.Y(n_2070)
);

HB1xp67_ASAP7_75t_L g2071 ( 
.A(n_2003),
.Y(n_2071)
);

A2O1A1Ixp33_ASAP7_75t_SL g2072 ( 
.A1(n_2004),
.A2(n_41),
.B(n_39),
.C(n_40),
.Y(n_2072)
);

AOI21xp5_ASAP7_75t_L g2073 ( 
.A1(n_2019),
.A2(n_1949),
.B(n_1944),
.Y(n_2073)
);

NAND2xp5_ASAP7_75t_L g2074 ( 
.A(n_2003),
.B(n_41),
.Y(n_2074)
);

A2O1A1Ixp33_ASAP7_75t_SL g2075 ( 
.A1(n_2026),
.A2(n_44),
.B(n_42),
.C(n_43),
.Y(n_2075)
);

OAI21xp33_ASAP7_75t_L g2076 ( 
.A1(n_2006),
.A2(n_1189),
.B(n_42),
.Y(n_2076)
);

NAND2xp5_ASAP7_75t_L g2077 ( 
.A(n_2000),
.B(n_43),
.Y(n_2077)
);

AND2x4_ASAP7_75t_L g2078 ( 
.A(n_2010),
.B(n_1975),
.Y(n_2078)
);

AND2x4_ASAP7_75t_L g2079 ( 
.A(n_1991),
.B(n_1975),
.Y(n_2079)
);

NAND2xp5_ASAP7_75t_L g2080 ( 
.A(n_2032),
.B(n_44),
.Y(n_2080)
);

INVx2_ASAP7_75t_L g2081 ( 
.A(n_2028),
.Y(n_2081)
);

INVx2_ASAP7_75t_SL g2082 ( 
.A(n_2071),
.Y(n_2082)
);

AOI21xp5_ASAP7_75t_SL g2083 ( 
.A1(n_2052),
.A2(n_1978),
.B(n_47),
.Y(n_2083)
);

BUFx3_ASAP7_75t_L g2084 ( 
.A(n_2029),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_2051),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_2040),
.Y(n_2086)
);

OAI21x1_ASAP7_75t_L g2087 ( 
.A1(n_2073),
.A2(n_1978),
.B(n_45),
.Y(n_2087)
);

INVx2_ASAP7_75t_L g2088 ( 
.A(n_2057),
.Y(n_2088)
);

INVx2_ASAP7_75t_L g2089 ( 
.A(n_2060),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_2059),
.Y(n_2090)
);

NAND2xp5_ASAP7_75t_L g2091 ( 
.A(n_2033),
.B(n_45),
.Y(n_2091)
);

AND2x2_ASAP7_75t_L g2092 ( 
.A(n_2034),
.B(n_46),
.Y(n_2092)
);

INVx2_ASAP7_75t_L g2093 ( 
.A(n_2050),
.Y(n_2093)
);

INVx2_ASAP7_75t_L g2094 ( 
.A(n_2065),
.Y(n_2094)
);

AND2x2_ASAP7_75t_L g2095 ( 
.A(n_2042),
.B(n_46),
.Y(n_2095)
);

OAI22xp5_ASAP7_75t_L g2096 ( 
.A1(n_2030),
.A2(n_49),
.B1(n_47),
.B2(n_48),
.Y(n_2096)
);

AND2x2_ASAP7_75t_L g2097 ( 
.A(n_2031),
.B(n_48),
.Y(n_2097)
);

HB1xp67_ASAP7_75t_L g2098 ( 
.A(n_2053),
.Y(n_2098)
);

AND2x2_ASAP7_75t_L g2099 ( 
.A(n_2064),
.B(n_49),
.Y(n_2099)
);

OAI22xp5_ASAP7_75t_L g2100 ( 
.A1(n_2069),
.A2(n_52),
.B1(n_50),
.B2(n_51),
.Y(n_2100)
);

INVx2_ASAP7_75t_L g2101 ( 
.A(n_2038),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_2044),
.Y(n_2102)
);

INVx4_ASAP7_75t_L g2103 ( 
.A(n_2037),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_2036),
.Y(n_2104)
);

OAI21x1_ASAP7_75t_L g2105 ( 
.A1(n_2048),
.A2(n_50),
.B(n_51),
.Y(n_2105)
);

AOI22xp33_ASAP7_75t_L g2106 ( 
.A1(n_2067),
.A2(n_54),
.B1(n_52),
.B2(n_53),
.Y(n_2106)
);

INVx2_ASAP7_75t_L g2107 ( 
.A(n_2068),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_2070),
.Y(n_2108)
);

AOI22xp33_ASAP7_75t_L g2109 ( 
.A1(n_2063),
.A2(n_56),
.B1(n_54),
.B2(n_55),
.Y(n_2109)
);

HB1xp67_ASAP7_75t_L g2110 ( 
.A(n_2045),
.Y(n_2110)
);

OAI21x1_ASAP7_75t_L g2111 ( 
.A1(n_2066),
.A2(n_55),
.B(n_56),
.Y(n_2111)
);

INVx1_ASAP7_75t_L g2112 ( 
.A(n_2047),
.Y(n_2112)
);

OAI21x1_ASAP7_75t_L g2113 ( 
.A1(n_2061),
.A2(n_57),
.B(n_58),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_2078),
.Y(n_2114)
);

HB1xp67_ASAP7_75t_L g2115 ( 
.A(n_2079),
.Y(n_2115)
);

HB1xp67_ASAP7_75t_L g2116 ( 
.A(n_2037),
.Y(n_2116)
);

BUFx4f_ASAP7_75t_SL g2117 ( 
.A(n_2054),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_2074),
.Y(n_2118)
);

AND2x4_ASAP7_75t_L g2119 ( 
.A(n_2054),
.B(n_57),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_2055),
.Y(n_2120)
);

CKINVDCx20_ASAP7_75t_R g2121 ( 
.A(n_2062),
.Y(n_2121)
);

AND2x2_ASAP7_75t_L g2122 ( 
.A(n_2039),
.B(n_59),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_2077),
.Y(n_2123)
);

CKINVDCx20_ASAP7_75t_R g2124 ( 
.A(n_2041),
.Y(n_2124)
);

AND2x4_ASAP7_75t_L g2125 ( 
.A(n_2046),
.B(n_59),
.Y(n_2125)
);

INVx2_ASAP7_75t_L g2126 ( 
.A(n_2072),
.Y(n_2126)
);

INVx2_ASAP7_75t_L g2127 ( 
.A(n_2056),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_2058),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_2043),
.Y(n_2129)
);

AND2x4_ASAP7_75t_L g2130 ( 
.A(n_2076),
.B(n_60),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_2035),
.Y(n_2131)
);

AOI21x1_ASAP7_75t_L g2132 ( 
.A1(n_2049),
.A2(n_60),
.B(n_61),
.Y(n_2132)
);

INVx2_ASAP7_75t_L g2133 ( 
.A(n_2075),
.Y(n_2133)
);

INVx2_ASAP7_75t_L g2134 ( 
.A(n_2028),
.Y(n_2134)
);

BUFx6f_ASAP7_75t_L g2135 ( 
.A(n_2037),
.Y(n_2135)
);

OAI21x1_ASAP7_75t_L g2136 ( 
.A1(n_2073),
.A2(n_62),
.B(n_63),
.Y(n_2136)
);

OAI21x1_ASAP7_75t_L g2137 ( 
.A1(n_2073),
.A2(n_62),
.B(n_63),
.Y(n_2137)
);

NOR2xp33_ASAP7_75t_L g2138 ( 
.A(n_2034),
.B(n_64),
.Y(n_2138)
);

AND2x2_ASAP7_75t_L g2139 ( 
.A(n_2032),
.B(n_64),
.Y(n_2139)
);

INVx2_ASAP7_75t_L g2140 ( 
.A(n_2028),
.Y(n_2140)
);

INVx2_ASAP7_75t_L g2141 ( 
.A(n_2028),
.Y(n_2141)
);

AND2x2_ASAP7_75t_L g2142 ( 
.A(n_2032),
.B(n_65),
.Y(n_2142)
);

INVx4_ASAP7_75t_SL g2143 ( 
.A(n_2029),
.Y(n_2143)
);

AND2x2_ASAP7_75t_L g2144 ( 
.A(n_2032),
.B(n_65),
.Y(n_2144)
);

OAI21xp5_ASAP7_75t_L g2145 ( 
.A1(n_2067),
.A2(n_66),
.B(n_67),
.Y(n_2145)
);

OAI21x1_ASAP7_75t_L g2146 ( 
.A1(n_2073),
.A2(n_67),
.B(n_68),
.Y(n_2146)
);

BUFx2_ASAP7_75t_L g2147 ( 
.A(n_2032),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_2051),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_2051),
.Y(n_2149)
);

INVx3_ASAP7_75t_SL g2150 ( 
.A(n_2031),
.Y(n_2150)
);

INVx2_ASAP7_75t_L g2151 ( 
.A(n_2028),
.Y(n_2151)
);

BUFx3_ASAP7_75t_L g2152 ( 
.A(n_2029),
.Y(n_2152)
);

INVx2_ASAP7_75t_L g2153 ( 
.A(n_2028),
.Y(n_2153)
);

NAND2x1p5_ASAP7_75t_L g2154 ( 
.A(n_2037),
.B(n_68),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_2051),
.Y(n_2155)
);

CKINVDCx20_ASAP7_75t_R g2156 ( 
.A(n_2071),
.Y(n_2156)
);

INVx2_ASAP7_75t_L g2157 ( 
.A(n_2094),
.Y(n_2157)
);

AND2x4_ASAP7_75t_L g2158 ( 
.A(n_2082),
.B(n_69),
.Y(n_2158)
);

BUFx2_ASAP7_75t_L g2159 ( 
.A(n_2147),
.Y(n_2159)
);

BUFx3_ASAP7_75t_L g2160 ( 
.A(n_2156),
.Y(n_2160)
);

OAI22xp5_ASAP7_75t_L g2161 ( 
.A1(n_2131),
.A2(n_72),
.B1(n_70),
.B2(n_71),
.Y(n_2161)
);

AND2x2_ASAP7_75t_L g2162 ( 
.A(n_2147),
.B(n_71),
.Y(n_2162)
);

NAND2xp5_ASAP7_75t_L g2163 ( 
.A(n_2102),
.B(n_72),
.Y(n_2163)
);

AND2x2_ASAP7_75t_L g2164 ( 
.A(n_2150),
.B(n_2090),
.Y(n_2164)
);

AOI22xp33_ASAP7_75t_SL g2165 ( 
.A1(n_2120),
.A2(n_75),
.B1(n_73),
.B2(n_74),
.Y(n_2165)
);

INVx2_ASAP7_75t_L g2166 ( 
.A(n_2093),
.Y(n_2166)
);

INVx2_ASAP7_75t_L g2167 ( 
.A(n_2107),
.Y(n_2167)
);

HB1xp67_ASAP7_75t_L g2168 ( 
.A(n_2098),
.Y(n_2168)
);

AND2x2_ASAP7_75t_L g2169 ( 
.A(n_2101),
.B(n_74),
.Y(n_2169)
);

AND2x2_ASAP7_75t_L g2170 ( 
.A(n_2104),
.B(n_76),
.Y(n_2170)
);

BUFx2_ASAP7_75t_L g2171 ( 
.A(n_2108),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_2085),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_2148),
.Y(n_2173)
);

INVx2_ASAP7_75t_L g2174 ( 
.A(n_2089),
.Y(n_2174)
);

INVx2_ASAP7_75t_SL g2175 ( 
.A(n_2117),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_2149),
.Y(n_2176)
);

AND2x2_ASAP7_75t_L g2177 ( 
.A(n_2115),
.B(n_76),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_2155),
.Y(n_2178)
);

AND2x2_ASAP7_75t_L g2179 ( 
.A(n_2123),
.B(n_77),
.Y(n_2179)
);

AOI22xp33_ASAP7_75t_L g2180 ( 
.A1(n_2128),
.A2(n_2129),
.B1(n_2130),
.B2(n_2126),
.Y(n_2180)
);

AOI22xp33_ASAP7_75t_SL g2181 ( 
.A1(n_2099),
.A2(n_79),
.B1(n_77),
.B2(n_78),
.Y(n_2181)
);

HB1xp67_ASAP7_75t_L g2182 ( 
.A(n_2110),
.Y(n_2182)
);

BUFx3_ASAP7_75t_L g2183 ( 
.A(n_2084),
.Y(n_2183)
);

NOR2x1_ASAP7_75t_L g2184 ( 
.A(n_2112),
.B(n_80),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_2086),
.Y(n_2185)
);

AND2x2_ASAP7_75t_L g2186 ( 
.A(n_2139),
.B(n_80),
.Y(n_2186)
);

NAND2xp5_ASAP7_75t_L g2187 ( 
.A(n_2118),
.B(n_81),
.Y(n_2187)
);

OR2x2_ASAP7_75t_L g2188 ( 
.A(n_2080),
.B(n_82),
.Y(n_2188)
);

AND2x4_ASAP7_75t_L g2189 ( 
.A(n_2116),
.B(n_83),
.Y(n_2189)
);

AND2x2_ASAP7_75t_L g2190 ( 
.A(n_2142),
.B(n_2144),
.Y(n_2190)
);

AND2x2_ASAP7_75t_L g2191 ( 
.A(n_2092),
.B(n_83),
.Y(n_2191)
);

AND2x4_ASAP7_75t_SL g2192 ( 
.A(n_2103),
.B(n_84),
.Y(n_2192)
);

AND2x4_ASAP7_75t_L g2193 ( 
.A(n_2114),
.B(n_85),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_2081),
.Y(n_2194)
);

CKINVDCx11_ASAP7_75t_R g2195 ( 
.A(n_2143),
.Y(n_2195)
);

AND2x2_ASAP7_75t_L g2196 ( 
.A(n_2152),
.B(n_85),
.Y(n_2196)
);

AND2x2_ASAP7_75t_L g2197 ( 
.A(n_2143),
.B(n_86),
.Y(n_2197)
);

NAND2xp5_ASAP7_75t_L g2198 ( 
.A(n_2091),
.B(n_86),
.Y(n_2198)
);

INVx1_ASAP7_75t_SL g2199 ( 
.A(n_2135),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_2088),
.Y(n_2200)
);

AND2x2_ASAP7_75t_L g2201 ( 
.A(n_2095),
.B(n_87),
.Y(n_2201)
);

AND2x2_ASAP7_75t_L g2202 ( 
.A(n_2138),
.B(n_87),
.Y(n_2202)
);

INVx1_ASAP7_75t_L g2203 ( 
.A(n_2134),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_2140),
.Y(n_2204)
);

INVx2_ASAP7_75t_L g2205 ( 
.A(n_2141),
.Y(n_2205)
);

INVx2_ASAP7_75t_L g2206 ( 
.A(n_2151),
.Y(n_2206)
);

INVx2_ASAP7_75t_L g2207 ( 
.A(n_2153),
.Y(n_2207)
);

INVx1_ASAP7_75t_L g2208 ( 
.A(n_2136),
.Y(n_2208)
);

AND2x2_ASAP7_75t_L g2209 ( 
.A(n_2097),
.B(n_88),
.Y(n_2209)
);

AND2x2_ASAP7_75t_L g2210 ( 
.A(n_2135),
.B(n_88),
.Y(n_2210)
);

BUFx12f_ASAP7_75t_L g2211 ( 
.A(n_2119),
.Y(n_2211)
);

AND2x4_ASAP7_75t_L g2212 ( 
.A(n_2122),
.B(n_89),
.Y(n_2212)
);

OR2x2_ASAP7_75t_L g2213 ( 
.A(n_2137),
.B(n_89),
.Y(n_2213)
);

AND2x2_ASAP7_75t_L g2214 ( 
.A(n_2124),
.B(n_2125),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_2146),
.Y(n_2215)
);

AOI22xp33_ASAP7_75t_L g2216 ( 
.A1(n_2133),
.A2(n_92),
.B1(n_90),
.B2(n_91),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_2087),
.Y(n_2217)
);

INVx2_ASAP7_75t_L g2218 ( 
.A(n_2105),
.Y(n_2218)
);

OR2x2_ASAP7_75t_L g2219 ( 
.A(n_2127),
.B(n_90),
.Y(n_2219)
);

AND2x2_ASAP7_75t_L g2220 ( 
.A(n_2111),
.B(n_91),
.Y(n_2220)
);

AND2x2_ASAP7_75t_L g2221 ( 
.A(n_2154),
.B(n_93),
.Y(n_2221)
);

AOI22xp33_ASAP7_75t_L g2222 ( 
.A1(n_2096),
.A2(n_95),
.B1(n_93),
.B2(n_94),
.Y(n_2222)
);

NAND2xp5_ASAP7_75t_L g2223 ( 
.A(n_2100),
.B(n_94),
.Y(n_2223)
);

NAND2xp5_ASAP7_75t_L g2224 ( 
.A(n_2083),
.B(n_2109),
.Y(n_2224)
);

HB1xp67_ASAP7_75t_L g2225 ( 
.A(n_2113),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_2132),
.Y(n_2226)
);

NAND2xp5_ASAP7_75t_L g2227 ( 
.A(n_2145),
.B(n_95),
.Y(n_2227)
);

OR2x2_ASAP7_75t_L g2228 ( 
.A(n_2106),
.B(n_96),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_2121),
.Y(n_2229)
);

BUFx2_ASAP7_75t_L g2230 ( 
.A(n_2110),
.Y(n_2230)
);

INVx2_ASAP7_75t_L g2231 ( 
.A(n_2094),
.Y(n_2231)
);

BUFx2_ASAP7_75t_L g2232 ( 
.A(n_2110),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_2098),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_2098),
.Y(n_2234)
);

INVx2_ASAP7_75t_L g2235 ( 
.A(n_2094),
.Y(n_2235)
);

AOI22xp5_ASAP7_75t_L g2236 ( 
.A1(n_2131),
.A2(n_99),
.B1(n_97),
.B2(n_98),
.Y(n_2236)
);

AND2x2_ASAP7_75t_L g2237 ( 
.A(n_2147),
.B(n_97),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_2098),
.Y(n_2238)
);

INVx2_ASAP7_75t_L g2239 ( 
.A(n_2094),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_2098),
.Y(n_2240)
);

HB1xp67_ASAP7_75t_L g2241 ( 
.A(n_2098),
.Y(n_2241)
);

INVx2_ASAP7_75t_L g2242 ( 
.A(n_2094),
.Y(n_2242)
);

NAND2xp5_ASAP7_75t_L g2243 ( 
.A(n_2102),
.B(n_98),
.Y(n_2243)
);

NAND2xp5_ASAP7_75t_L g2244 ( 
.A(n_2102),
.B(n_99),
.Y(n_2244)
);

BUFx3_ASAP7_75t_L g2245 ( 
.A(n_2156),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_2098),
.Y(n_2246)
);

AND2x2_ASAP7_75t_L g2247 ( 
.A(n_2147),
.B(n_100),
.Y(n_2247)
);

AND2x2_ASAP7_75t_L g2248 ( 
.A(n_2147),
.B(n_100),
.Y(n_2248)
);

INVx1_ASAP7_75t_L g2249 ( 
.A(n_2098),
.Y(n_2249)
);

BUFx3_ASAP7_75t_L g2250 ( 
.A(n_2156),
.Y(n_2250)
);

AND2x4_ASAP7_75t_L g2251 ( 
.A(n_2082),
.B(n_101),
.Y(n_2251)
);

AND2x2_ASAP7_75t_L g2252 ( 
.A(n_2147),
.B(n_101),
.Y(n_2252)
);

INVx2_ASAP7_75t_L g2253 ( 
.A(n_2094),
.Y(n_2253)
);

BUFx12f_ASAP7_75t_L g2254 ( 
.A(n_2119),
.Y(n_2254)
);

BUFx2_ASAP7_75t_L g2255 ( 
.A(n_2160),
.Y(n_2255)
);

OR2x2_ASAP7_75t_L g2256 ( 
.A(n_2159),
.B(n_102),
.Y(n_2256)
);

OR2x2_ASAP7_75t_L g2257 ( 
.A(n_2168),
.B(n_103),
.Y(n_2257)
);

AND2x2_ASAP7_75t_L g2258 ( 
.A(n_2164),
.B(n_2190),
.Y(n_2258)
);

BUFx3_ASAP7_75t_L g2259 ( 
.A(n_2245),
.Y(n_2259)
);

AND2x2_ASAP7_75t_L g2260 ( 
.A(n_2241),
.B(n_103),
.Y(n_2260)
);

OR2x2_ASAP7_75t_L g2261 ( 
.A(n_2233),
.B(n_2234),
.Y(n_2261)
);

INVx2_ASAP7_75t_L g2262 ( 
.A(n_2167),
.Y(n_2262)
);

AND2x2_ASAP7_75t_L g2263 ( 
.A(n_2238),
.B(n_104),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_2185),
.Y(n_2264)
);

AND2x2_ASAP7_75t_L g2265 ( 
.A(n_2240),
.B(n_104),
.Y(n_2265)
);

INVx2_ASAP7_75t_L g2266 ( 
.A(n_2174),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_2172),
.Y(n_2267)
);

NOR2xp33_ASAP7_75t_L g2268 ( 
.A(n_2195),
.B(n_105),
.Y(n_2268)
);

BUFx6f_ASAP7_75t_L g2269 ( 
.A(n_2183),
.Y(n_2269)
);

OAI22xp5_ASAP7_75t_L g2270 ( 
.A1(n_2224),
.A2(n_107),
.B1(n_105),
.B2(n_106),
.Y(n_2270)
);

INVx1_ASAP7_75t_L g2271 ( 
.A(n_2173),
.Y(n_2271)
);

OR2x2_ASAP7_75t_L g2272 ( 
.A(n_2246),
.B(n_2249),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_2176),
.Y(n_2273)
);

INVx2_ASAP7_75t_L g2274 ( 
.A(n_2218),
.Y(n_2274)
);

INVx1_ASAP7_75t_L g2275 ( 
.A(n_2178),
.Y(n_2275)
);

INVx2_ASAP7_75t_L g2276 ( 
.A(n_2225),
.Y(n_2276)
);

NOR2xp33_ASAP7_75t_L g2277 ( 
.A(n_2250),
.B(n_107),
.Y(n_2277)
);

INVx1_ASAP7_75t_L g2278 ( 
.A(n_2171),
.Y(n_2278)
);

NAND2xp5_ASAP7_75t_L g2279 ( 
.A(n_2162),
.B(n_108),
.Y(n_2279)
);

INVx2_ASAP7_75t_L g2280 ( 
.A(n_2205),
.Y(n_2280)
);

BUFx2_ASAP7_75t_L g2281 ( 
.A(n_2158),
.Y(n_2281)
);

INVx1_ASAP7_75t_L g2282 ( 
.A(n_2208),
.Y(n_2282)
);

AND2x2_ASAP7_75t_L g2283 ( 
.A(n_2237),
.B(n_108),
.Y(n_2283)
);

INVx2_ASAP7_75t_L g2284 ( 
.A(n_2206),
.Y(n_2284)
);

INVx2_ASAP7_75t_L g2285 ( 
.A(n_2207),
.Y(n_2285)
);

INVx2_ASAP7_75t_SL g2286 ( 
.A(n_2175),
.Y(n_2286)
);

AND2x2_ASAP7_75t_L g2287 ( 
.A(n_2247),
.B(n_109),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_2215),
.Y(n_2288)
);

INVx3_ASAP7_75t_L g2289 ( 
.A(n_2189),
.Y(n_2289)
);

INVx2_ASAP7_75t_L g2290 ( 
.A(n_2157),
.Y(n_2290)
);

AND2x4_ASAP7_75t_L g2291 ( 
.A(n_2248),
.B(n_109),
.Y(n_2291)
);

INVx2_ASAP7_75t_SL g2292 ( 
.A(n_2252),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_2217),
.Y(n_2293)
);

INVx1_ASAP7_75t_L g2294 ( 
.A(n_2182),
.Y(n_2294)
);

AND2x2_ASAP7_75t_L g2295 ( 
.A(n_2230),
.B(n_2232),
.Y(n_2295)
);

INVx1_ASAP7_75t_L g2296 ( 
.A(n_2230),
.Y(n_2296)
);

INVx2_ASAP7_75t_L g2297 ( 
.A(n_2166),
.Y(n_2297)
);

AOI33xp33_ASAP7_75t_L g2298 ( 
.A1(n_2180),
.A2(n_112),
.A3(n_114),
.B1(n_110),
.B2(n_111),
.B3(n_113),
.Y(n_2298)
);

OR2x2_ASAP7_75t_L g2299 ( 
.A(n_2232),
.B(n_110),
.Y(n_2299)
);

AO31x2_ASAP7_75t_L g2300 ( 
.A1(n_2226),
.A2(n_121),
.A3(n_129),
.B(n_111),
.Y(n_2300)
);

NAND2xp5_ASAP7_75t_L g2301 ( 
.A(n_2170),
.B(n_113),
.Y(n_2301)
);

AND2x2_ASAP7_75t_L g2302 ( 
.A(n_2199),
.B(n_115),
.Y(n_2302)
);

HB1xp67_ASAP7_75t_L g2303 ( 
.A(n_2219),
.Y(n_2303)
);

INVx2_ASAP7_75t_L g2304 ( 
.A(n_2231),
.Y(n_2304)
);

AND2x2_ASAP7_75t_L g2305 ( 
.A(n_2214),
.B(n_116),
.Y(n_2305)
);

AND2x2_ASAP7_75t_L g2306 ( 
.A(n_2251),
.B(n_116),
.Y(n_2306)
);

INVx3_ASAP7_75t_L g2307 ( 
.A(n_2211),
.Y(n_2307)
);

INVx1_ASAP7_75t_L g2308 ( 
.A(n_2194),
.Y(n_2308)
);

AND2x2_ASAP7_75t_L g2309 ( 
.A(n_2191),
.B(n_117),
.Y(n_2309)
);

BUFx2_ASAP7_75t_L g2310 ( 
.A(n_2177),
.Y(n_2310)
);

OR2x2_ASAP7_75t_L g2311 ( 
.A(n_2235),
.B(n_117),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_2200),
.Y(n_2312)
);

AND2x2_ASAP7_75t_L g2313 ( 
.A(n_2186),
.B(n_2202),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_2203),
.Y(n_2314)
);

INVx1_ASAP7_75t_L g2315 ( 
.A(n_2204),
.Y(n_2315)
);

AND2x2_ASAP7_75t_L g2316 ( 
.A(n_2179),
.B(n_118),
.Y(n_2316)
);

INVx2_ASAP7_75t_L g2317 ( 
.A(n_2239),
.Y(n_2317)
);

AND2x2_ASAP7_75t_L g2318 ( 
.A(n_2229),
.B(n_119),
.Y(n_2318)
);

HB1xp67_ASAP7_75t_L g2319 ( 
.A(n_2187),
.Y(n_2319)
);

AND2x2_ASAP7_75t_L g2320 ( 
.A(n_2209),
.B(n_119),
.Y(n_2320)
);

INVx3_ASAP7_75t_L g2321 ( 
.A(n_2254),
.Y(n_2321)
);

INVx2_ASAP7_75t_L g2322 ( 
.A(n_2242),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_2163),
.Y(n_2323)
);

NOR2xp33_ASAP7_75t_R g2324 ( 
.A(n_2197),
.B(n_120),
.Y(n_2324)
);

AND2x2_ASAP7_75t_L g2325 ( 
.A(n_2201),
.B(n_122),
.Y(n_2325)
);

AND2x2_ASAP7_75t_L g2326 ( 
.A(n_2212),
.B(n_122),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_2243),
.Y(n_2327)
);

INVx1_ASAP7_75t_L g2328 ( 
.A(n_2244),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_2253),
.Y(n_2329)
);

INVx1_ASAP7_75t_L g2330 ( 
.A(n_2169),
.Y(n_2330)
);

AND2x2_ASAP7_75t_L g2331 ( 
.A(n_2196),
.B(n_123),
.Y(n_2331)
);

BUFx3_ASAP7_75t_L g2332 ( 
.A(n_2192),
.Y(n_2332)
);

INVx2_ASAP7_75t_L g2333 ( 
.A(n_2193),
.Y(n_2333)
);

INVxp67_ASAP7_75t_L g2334 ( 
.A(n_2184),
.Y(n_2334)
);

INVx1_ASAP7_75t_L g2335 ( 
.A(n_2213),
.Y(n_2335)
);

BUFx6f_ASAP7_75t_L g2336 ( 
.A(n_2210),
.Y(n_2336)
);

AND2x2_ASAP7_75t_L g2337 ( 
.A(n_2188),
.B(n_123),
.Y(n_2337)
);

INVx1_ASAP7_75t_L g2338 ( 
.A(n_2198),
.Y(n_2338)
);

AND2x2_ASAP7_75t_L g2339 ( 
.A(n_2221),
.B(n_124),
.Y(n_2339)
);

HB1xp67_ASAP7_75t_L g2340 ( 
.A(n_2220),
.Y(n_2340)
);

AND2x2_ASAP7_75t_L g2341 ( 
.A(n_2223),
.B(n_124),
.Y(n_2341)
);

BUFx2_ASAP7_75t_L g2342 ( 
.A(n_2227),
.Y(n_2342)
);

OR2x2_ASAP7_75t_L g2343 ( 
.A(n_2228),
.B(n_125),
.Y(n_2343)
);

AND2x2_ASAP7_75t_L g2344 ( 
.A(n_2181),
.B(n_126),
.Y(n_2344)
);

HB1xp67_ASAP7_75t_L g2345 ( 
.A(n_2161),
.Y(n_2345)
);

INVx4_ASAP7_75t_L g2346 ( 
.A(n_2236),
.Y(n_2346)
);

NOR2x1_ASAP7_75t_SL g2347 ( 
.A(n_2165),
.B(n_126),
.Y(n_2347)
);

AND2x2_ASAP7_75t_L g2348 ( 
.A(n_2216),
.B(n_127),
.Y(n_2348)
);

AND2x2_ASAP7_75t_L g2349 ( 
.A(n_2222),
.B(n_127),
.Y(n_2349)
);

INVx2_ASAP7_75t_L g2350 ( 
.A(n_2167),
.Y(n_2350)
);

AND2x2_ASAP7_75t_L g2351 ( 
.A(n_2159),
.B(n_128),
.Y(n_2351)
);

INVx3_ASAP7_75t_L g2352 ( 
.A(n_2160),
.Y(n_2352)
);

INVxp67_ASAP7_75t_L g2353 ( 
.A(n_2168),
.Y(n_2353)
);

INVx2_ASAP7_75t_L g2354 ( 
.A(n_2167),
.Y(n_2354)
);

OR2x2_ASAP7_75t_L g2355 ( 
.A(n_2159),
.B(n_128),
.Y(n_2355)
);

AND2x4_ASAP7_75t_L g2356 ( 
.A(n_2160),
.B(n_129),
.Y(n_2356)
);

INVx2_ASAP7_75t_L g2357 ( 
.A(n_2167),
.Y(n_2357)
);

INVx1_ASAP7_75t_L g2358 ( 
.A(n_2185),
.Y(n_2358)
);

INVx2_ASAP7_75t_SL g2359 ( 
.A(n_2160),
.Y(n_2359)
);

INVx2_ASAP7_75t_L g2360 ( 
.A(n_2167),
.Y(n_2360)
);

OA21x2_ASAP7_75t_L g2361 ( 
.A1(n_2230),
.A2(n_130),
.B(n_131),
.Y(n_2361)
);

AND2x2_ASAP7_75t_L g2362 ( 
.A(n_2159),
.B(n_130),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_2185),
.Y(n_2363)
);

INVx1_ASAP7_75t_L g2364 ( 
.A(n_2185),
.Y(n_2364)
);

INVx2_ASAP7_75t_L g2365 ( 
.A(n_2167),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_2185),
.Y(n_2366)
);

INVx2_ASAP7_75t_L g2367 ( 
.A(n_2167),
.Y(n_2367)
);

AND2x2_ASAP7_75t_L g2368 ( 
.A(n_2159),
.B(n_131),
.Y(n_2368)
);

NAND2xp5_ASAP7_75t_L g2369 ( 
.A(n_2168),
.B(n_132),
.Y(n_2369)
);

AND2x4_ASAP7_75t_L g2370 ( 
.A(n_2160),
.B(n_132),
.Y(n_2370)
);

AND2x2_ASAP7_75t_L g2371 ( 
.A(n_2159),
.B(n_133),
.Y(n_2371)
);

OAI221xp5_ASAP7_75t_L g2372 ( 
.A1(n_2180),
.A2(n_135),
.B1(n_133),
.B2(n_134),
.C(n_137),
.Y(n_2372)
);

AND2x2_ASAP7_75t_L g2373 ( 
.A(n_2159),
.B(n_135),
.Y(n_2373)
);

BUFx3_ASAP7_75t_L g2374 ( 
.A(n_2160),
.Y(n_2374)
);

INVx1_ASAP7_75t_L g2375 ( 
.A(n_2267),
.Y(n_2375)
);

AND2x4_ASAP7_75t_SL g2376 ( 
.A(n_2269),
.B(n_138),
.Y(n_2376)
);

BUFx3_ASAP7_75t_L g2377 ( 
.A(n_2269),
.Y(n_2377)
);

HB1xp67_ASAP7_75t_L g2378 ( 
.A(n_2361),
.Y(n_2378)
);

INVx1_ASAP7_75t_L g2379 ( 
.A(n_2271),
.Y(n_2379)
);

AND2x2_ASAP7_75t_L g2380 ( 
.A(n_2258),
.B(n_139),
.Y(n_2380)
);

AND2x2_ASAP7_75t_L g2381 ( 
.A(n_2310),
.B(n_2340),
.Y(n_2381)
);

INVx2_ASAP7_75t_L g2382 ( 
.A(n_2274),
.Y(n_2382)
);

NOR2xp67_ASAP7_75t_L g2383 ( 
.A(n_2334),
.B(n_139),
.Y(n_2383)
);

AND2x2_ASAP7_75t_L g2384 ( 
.A(n_2342),
.B(n_140),
.Y(n_2384)
);

INVx2_ASAP7_75t_L g2385 ( 
.A(n_2290),
.Y(n_2385)
);

INVx1_ASAP7_75t_SL g2386 ( 
.A(n_2324),
.Y(n_2386)
);

INVx1_ASAP7_75t_L g2387 ( 
.A(n_2273),
.Y(n_2387)
);

OR2x2_ASAP7_75t_L g2388 ( 
.A(n_2261),
.B(n_140),
.Y(n_2388)
);

AND2x2_ASAP7_75t_L g2389 ( 
.A(n_2313),
.B(n_141),
.Y(n_2389)
);

INVx1_ASAP7_75t_L g2390 ( 
.A(n_2275),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_2264),
.Y(n_2391)
);

HB1xp67_ASAP7_75t_L g2392 ( 
.A(n_2353),
.Y(n_2392)
);

INVx1_ASAP7_75t_L g2393 ( 
.A(n_2358),
.Y(n_2393)
);

AND2x4_ASAP7_75t_L g2394 ( 
.A(n_2255),
.B(n_141),
.Y(n_2394)
);

NAND2xp5_ASAP7_75t_L g2395 ( 
.A(n_2319),
.B(n_143),
.Y(n_2395)
);

INVx1_ASAP7_75t_L g2396 ( 
.A(n_2363),
.Y(n_2396)
);

NAND2xp5_ASAP7_75t_L g2397 ( 
.A(n_2303),
.B(n_143),
.Y(n_2397)
);

AND2x2_ASAP7_75t_L g2398 ( 
.A(n_2292),
.B(n_144),
.Y(n_2398)
);

AND2x2_ASAP7_75t_L g2399 ( 
.A(n_2281),
.B(n_144),
.Y(n_2399)
);

AND2x2_ASAP7_75t_L g2400 ( 
.A(n_2289),
.B(n_145),
.Y(n_2400)
);

INVx1_ASAP7_75t_L g2401 ( 
.A(n_2364),
.Y(n_2401)
);

AND2x2_ASAP7_75t_L g2402 ( 
.A(n_2278),
.B(n_145),
.Y(n_2402)
);

HB1xp67_ASAP7_75t_L g2403 ( 
.A(n_2276),
.Y(n_2403)
);

NAND2xp5_ASAP7_75t_L g2404 ( 
.A(n_2323),
.B(n_146),
.Y(n_2404)
);

INVx1_ASAP7_75t_SL g2405 ( 
.A(n_2259),
.Y(n_2405)
);

INVx1_ASAP7_75t_L g2406 ( 
.A(n_2366),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_2272),
.Y(n_2407)
);

INVx1_ASAP7_75t_L g2408 ( 
.A(n_2293),
.Y(n_2408)
);

AND2x2_ASAP7_75t_L g2409 ( 
.A(n_2263),
.B(n_146),
.Y(n_2409)
);

NOR2x1_ASAP7_75t_L g2410 ( 
.A(n_2374),
.B(n_2299),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_2282),
.Y(n_2411)
);

AND2x4_ASAP7_75t_L g2412 ( 
.A(n_2335),
.B(n_147),
.Y(n_2412)
);

INVx1_ASAP7_75t_L g2413 ( 
.A(n_2288),
.Y(n_2413)
);

HB1xp67_ASAP7_75t_L g2414 ( 
.A(n_2294),
.Y(n_2414)
);

AND2x2_ASAP7_75t_L g2415 ( 
.A(n_2265),
.B(n_148),
.Y(n_2415)
);

AND2x4_ASAP7_75t_L g2416 ( 
.A(n_2286),
.B(n_149),
.Y(n_2416)
);

AND2x2_ASAP7_75t_SL g2417 ( 
.A(n_2346),
.B(n_149),
.Y(n_2417)
);

INVx2_ASAP7_75t_L g2418 ( 
.A(n_2297),
.Y(n_2418)
);

INVx1_ASAP7_75t_L g2419 ( 
.A(n_2308),
.Y(n_2419)
);

AND2x2_ASAP7_75t_L g2420 ( 
.A(n_2295),
.B(n_150),
.Y(n_2420)
);

INVx2_ASAP7_75t_L g2421 ( 
.A(n_2304),
.Y(n_2421)
);

INVx1_ASAP7_75t_L g2422 ( 
.A(n_2312),
.Y(n_2422)
);

AND2x2_ASAP7_75t_L g2423 ( 
.A(n_2338),
.B(n_150),
.Y(n_2423)
);

AND2x2_ASAP7_75t_L g2424 ( 
.A(n_2345),
.B(n_151),
.Y(n_2424)
);

NAND2xp5_ASAP7_75t_L g2425 ( 
.A(n_2327),
.B(n_151),
.Y(n_2425)
);

AND2x2_ASAP7_75t_L g2426 ( 
.A(n_2296),
.B(n_152),
.Y(n_2426)
);

INVx1_ASAP7_75t_L g2427 ( 
.A(n_2314),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_2315),
.Y(n_2428)
);

OR2x2_ASAP7_75t_L g2429 ( 
.A(n_2328),
.B(n_152),
.Y(n_2429)
);

AND2x2_ASAP7_75t_L g2430 ( 
.A(n_2351),
.B(n_153),
.Y(n_2430)
);

HB1xp67_ASAP7_75t_L g2431 ( 
.A(n_2300),
.Y(n_2431)
);

AND2x2_ASAP7_75t_L g2432 ( 
.A(n_2362),
.B(n_153),
.Y(n_2432)
);

INVx1_ASAP7_75t_L g2433 ( 
.A(n_2300),
.Y(n_2433)
);

INVx1_ASAP7_75t_SL g2434 ( 
.A(n_2332),
.Y(n_2434)
);

BUFx2_ASAP7_75t_L g2435 ( 
.A(n_2352),
.Y(n_2435)
);

OR2x2_ASAP7_75t_L g2436 ( 
.A(n_2257),
.B(n_154),
.Y(n_2436)
);

OR2x2_ASAP7_75t_L g2437 ( 
.A(n_2256),
.B(n_154),
.Y(n_2437)
);

HB1xp67_ASAP7_75t_L g2438 ( 
.A(n_2355),
.Y(n_2438)
);

INVx1_ASAP7_75t_SL g2439 ( 
.A(n_2291),
.Y(n_2439)
);

AOI22xp33_ASAP7_75t_L g2440 ( 
.A1(n_2343),
.A2(n_157),
.B1(n_155),
.B2(n_156),
.Y(n_2440)
);

BUFx2_ASAP7_75t_SL g2441 ( 
.A(n_2359),
.Y(n_2441)
);

INVx1_ASAP7_75t_L g2442 ( 
.A(n_2311),
.Y(n_2442)
);

INVx2_ASAP7_75t_L g2443 ( 
.A(n_2317),
.Y(n_2443)
);

INVx2_ASAP7_75t_L g2444 ( 
.A(n_2322),
.Y(n_2444)
);

NAND2xp5_ASAP7_75t_L g2445 ( 
.A(n_2260),
.B(n_155),
.Y(n_2445)
);

AND2x2_ASAP7_75t_L g2446 ( 
.A(n_2368),
.B(n_2371),
.Y(n_2446)
);

INVx1_ASAP7_75t_L g2447 ( 
.A(n_2369),
.Y(n_2447)
);

INVx1_ASAP7_75t_L g2448 ( 
.A(n_2330),
.Y(n_2448)
);

INVx1_ASAP7_75t_L g2449 ( 
.A(n_2373),
.Y(n_2449)
);

INVx1_ASAP7_75t_L g2450 ( 
.A(n_2329),
.Y(n_2450)
);

AND2x4_ASAP7_75t_SL g2451 ( 
.A(n_2307),
.B(n_156),
.Y(n_2451)
);

INVxp67_ASAP7_75t_L g2452 ( 
.A(n_2268),
.Y(n_2452)
);

NAND2xp5_ASAP7_75t_L g2453 ( 
.A(n_2341),
.B(n_157),
.Y(n_2453)
);

INVx1_ASAP7_75t_L g2454 ( 
.A(n_2262),
.Y(n_2454)
);

AND2x2_ASAP7_75t_L g2455 ( 
.A(n_2321),
.B(n_158),
.Y(n_2455)
);

AND2x2_ASAP7_75t_L g2456 ( 
.A(n_2318),
.B(n_158),
.Y(n_2456)
);

OR2x2_ASAP7_75t_L g2457 ( 
.A(n_2333),
.B(n_160),
.Y(n_2457)
);

OR2x2_ASAP7_75t_L g2458 ( 
.A(n_2279),
.B(n_160),
.Y(n_2458)
);

AND2x2_ASAP7_75t_L g2459 ( 
.A(n_2283),
.B(n_161),
.Y(n_2459)
);

INVx1_ASAP7_75t_L g2460 ( 
.A(n_2266),
.Y(n_2460)
);

AND2x2_ASAP7_75t_L g2461 ( 
.A(n_2287),
.B(n_161),
.Y(n_2461)
);

INVx2_ASAP7_75t_L g2462 ( 
.A(n_2280),
.Y(n_2462)
);

AND2x2_ASAP7_75t_L g2463 ( 
.A(n_2302),
.B(n_162),
.Y(n_2463)
);

NOR2xp33_ASAP7_75t_L g2464 ( 
.A(n_2336),
.B(n_2277),
.Y(n_2464)
);

INVx1_ASAP7_75t_L g2465 ( 
.A(n_2350),
.Y(n_2465)
);

NAND2xp5_ASAP7_75t_L g2466 ( 
.A(n_2337),
.B(n_162),
.Y(n_2466)
);

OR2x2_ASAP7_75t_SL g2467 ( 
.A(n_2336),
.B(n_163),
.Y(n_2467)
);

AND2x2_ASAP7_75t_L g2468 ( 
.A(n_2305),
.B(n_163),
.Y(n_2468)
);

AND2x2_ASAP7_75t_L g2469 ( 
.A(n_2309),
.B(n_164),
.Y(n_2469)
);

OR2x2_ASAP7_75t_L g2470 ( 
.A(n_2354),
.B(n_165),
.Y(n_2470)
);

AND2x4_ASAP7_75t_L g2471 ( 
.A(n_2356),
.B(n_165),
.Y(n_2471)
);

NAND2xp5_ASAP7_75t_SL g2472 ( 
.A(n_2370),
.B(n_166),
.Y(n_2472)
);

AND2x2_ASAP7_75t_L g2473 ( 
.A(n_2325),
.B(n_166),
.Y(n_2473)
);

AND2x2_ASAP7_75t_L g2474 ( 
.A(n_2306),
.B(n_167),
.Y(n_2474)
);

INVx1_ASAP7_75t_L g2475 ( 
.A(n_2357),
.Y(n_2475)
);

AND2x2_ASAP7_75t_L g2476 ( 
.A(n_2320),
.B(n_167),
.Y(n_2476)
);

AND2x2_ASAP7_75t_L g2477 ( 
.A(n_2331),
.B(n_168),
.Y(n_2477)
);

INVx1_ASAP7_75t_SL g2478 ( 
.A(n_2339),
.Y(n_2478)
);

CKINVDCx6p67_ASAP7_75t_R g2479 ( 
.A(n_2326),
.Y(n_2479)
);

INVx2_ASAP7_75t_SL g2480 ( 
.A(n_2316),
.Y(n_2480)
);

OR2x2_ASAP7_75t_L g2481 ( 
.A(n_2360),
.B(n_168),
.Y(n_2481)
);

INVx1_ASAP7_75t_L g2482 ( 
.A(n_2365),
.Y(n_2482)
);

INVx2_ASAP7_75t_L g2483 ( 
.A(n_2284),
.Y(n_2483)
);

INVx4_ASAP7_75t_L g2484 ( 
.A(n_2344),
.Y(n_2484)
);

INVx3_ASAP7_75t_L g2485 ( 
.A(n_2367),
.Y(n_2485)
);

AND2x4_ASAP7_75t_SL g2486 ( 
.A(n_2349),
.B(n_169),
.Y(n_2486)
);

AND2x2_ASAP7_75t_L g2487 ( 
.A(n_2301),
.B(n_170),
.Y(n_2487)
);

INVx2_ASAP7_75t_L g2488 ( 
.A(n_2285),
.Y(n_2488)
);

INVx1_ASAP7_75t_L g2489 ( 
.A(n_2270),
.Y(n_2489)
);

INVxp67_ASAP7_75t_SL g2490 ( 
.A(n_2347),
.Y(n_2490)
);

NOR2x1p5_ASAP7_75t_L g2491 ( 
.A(n_2348),
.B(n_170),
.Y(n_2491)
);

INVx3_ASAP7_75t_L g2492 ( 
.A(n_2298),
.Y(n_2492)
);

INVx1_ASAP7_75t_L g2493 ( 
.A(n_2372),
.Y(n_2493)
);

INVx2_ASAP7_75t_L g2494 ( 
.A(n_2361),
.Y(n_2494)
);

AND2x2_ASAP7_75t_L g2495 ( 
.A(n_2258),
.B(n_171),
.Y(n_2495)
);

AND2x2_ASAP7_75t_L g2496 ( 
.A(n_2258),
.B(n_171),
.Y(n_2496)
);

OR2x2_ASAP7_75t_L g2497 ( 
.A(n_2261),
.B(n_172),
.Y(n_2497)
);

NOR2x1_ASAP7_75t_SL g2498 ( 
.A(n_2299),
.B(n_172),
.Y(n_2498)
);

AND2x2_ASAP7_75t_L g2499 ( 
.A(n_2258),
.B(n_173),
.Y(n_2499)
);

AND2x4_ASAP7_75t_L g2500 ( 
.A(n_2258),
.B(n_173),
.Y(n_2500)
);

INVxp67_ASAP7_75t_SL g2501 ( 
.A(n_2334),
.Y(n_2501)
);

INVx2_ASAP7_75t_L g2502 ( 
.A(n_2361),
.Y(n_2502)
);

INVx1_ASAP7_75t_L g2503 ( 
.A(n_2267),
.Y(n_2503)
);

OR2x2_ASAP7_75t_L g2504 ( 
.A(n_2261),
.B(n_174),
.Y(n_2504)
);

BUFx2_ASAP7_75t_L g2505 ( 
.A(n_2255),
.Y(n_2505)
);

AND2x4_ASAP7_75t_L g2506 ( 
.A(n_2258),
.B(n_174),
.Y(n_2506)
);

INVx3_ASAP7_75t_L g2507 ( 
.A(n_2269),
.Y(n_2507)
);

INVx1_ASAP7_75t_L g2508 ( 
.A(n_2267),
.Y(n_2508)
);

AND2x2_ASAP7_75t_L g2509 ( 
.A(n_2258),
.B(n_175),
.Y(n_2509)
);

INVx1_ASAP7_75t_L g2510 ( 
.A(n_2267),
.Y(n_2510)
);

NAND2x1_ASAP7_75t_L g2511 ( 
.A(n_2295),
.B(n_175),
.Y(n_2511)
);

INVx1_ASAP7_75t_L g2512 ( 
.A(n_2267),
.Y(n_2512)
);

AND2x2_ASAP7_75t_L g2513 ( 
.A(n_2258),
.B(n_176),
.Y(n_2513)
);

INVx2_ASAP7_75t_L g2514 ( 
.A(n_2361),
.Y(n_2514)
);

NAND2xp5_ASAP7_75t_SL g2515 ( 
.A(n_2255),
.B(n_177),
.Y(n_2515)
);

AND2x2_ASAP7_75t_L g2516 ( 
.A(n_2258),
.B(n_178),
.Y(n_2516)
);

HB1xp67_ASAP7_75t_L g2517 ( 
.A(n_2361),
.Y(n_2517)
);

NAND2xp5_ASAP7_75t_L g2518 ( 
.A(n_2319),
.B(n_179),
.Y(n_2518)
);

AND2x2_ASAP7_75t_L g2519 ( 
.A(n_2258),
.B(n_180),
.Y(n_2519)
);

NAND2xp5_ASAP7_75t_L g2520 ( 
.A(n_2319),
.B(n_180),
.Y(n_2520)
);

AND2x4_ASAP7_75t_L g2521 ( 
.A(n_2258),
.B(n_181),
.Y(n_2521)
);

NAND2xp5_ASAP7_75t_L g2522 ( 
.A(n_2319),
.B(n_181),
.Y(n_2522)
);

HB1xp67_ASAP7_75t_L g2523 ( 
.A(n_2361),
.Y(n_2523)
);

AND2x2_ASAP7_75t_L g2524 ( 
.A(n_2258),
.B(n_182),
.Y(n_2524)
);

INVx3_ASAP7_75t_L g2525 ( 
.A(n_2269),
.Y(n_2525)
);

OR2x2_ASAP7_75t_L g2526 ( 
.A(n_2261),
.B(n_182),
.Y(n_2526)
);

INVx2_ASAP7_75t_L g2527 ( 
.A(n_2361),
.Y(n_2527)
);

AND2x2_ASAP7_75t_L g2528 ( 
.A(n_2258),
.B(n_183),
.Y(n_2528)
);

INVx1_ASAP7_75t_L g2529 ( 
.A(n_2267),
.Y(n_2529)
);

INVxp67_ASAP7_75t_L g2530 ( 
.A(n_2303),
.Y(n_2530)
);

NAND2xp5_ASAP7_75t_L g2531 ( 
.A(n_2319),
.B(n_183),
.Y(n_2531)
);

HB1xp67_ASAP7_75t_L g2532 ( 
.A(n_2361),
.Y(n_2532)
);

BUFx6f_ASAP7_75t_L g2533 ( 
.A(n_2269),
.Y(n_2533)
);

INVx1_ASAP7_75t_L g2534 ( 
.A(n_2267),
.Y(n_2534)
);

INVx4_ASAP7_75t_L g2535 ( 
.A(n_2269),
.Y(n_2535)
);

INVx2_ASAP7_75t_L g2536 ( 
.A(n_2361),
.Y(n_2536)
);

INVx1_ASAP7_75t_L g2537 ( 
.A(n_2267),
.Y(n_2537)
);

INVx2_ASAP7_75t_L g2538 ( 
.A(n_2361),
.Y(n_2538)
);

INVx2_ASAP7_75t_L g2539 ( 
.A(n_2361),
.Y(n_2539)
);

AND2x2_ASAP7_75t_L g2540 ( 
.A(n_2258),
.B(n_184),
.Y(n_2540)
);

NOR2xp67_ASAP7_75t_L g2541 ( 
.A(n_2334),
.B(n_185),
.Y(n_2541)
);

INVx1_ASAP7_75t_SL g2542 ( 
.A(n_2324),
.Y(n_2542)
);

AND2x2_ASAP7_75t_L g2543 ( 
.A(n_2258),
.B(n_185),
.Y(n_2543)
);

INVx2_ASAP7_75t_L g2544 ( 
.A(n_2361),
.Y(n_2544)
);

AND2x4_ASAP7_75t_L g2545 ( 
.A(n_2505),
.B(n_186),
.Y(n_2545)
);

INVx1_ASAP7_75t_L g2546 ( 
.A(n_2431),
.Y(n_2546)
);

INVx1_ASAP7_75t_L g2547 ( 
.A(n_2375),
.Y(n_2547)
);

INVx2_ASAP7_75t_L g2548 ( 
.A(n_2467),
.Y(n_2548)
);

OA211x2_ASAP7_75t_L g2549 ( 
.A1(n_2511),
.A2(n_2530),
.B(n_2452),
.C(n_2515),
.Y(n_2549)
);

AO21x1_ASAP7_75t_SL g2550 ( 
.A1(n_2392),
.A2(n_187),
.B(n_188),
.Y(n_2550)
);

BUFx2_ASAP7_75t_L g2551 ( 
.A(n_2435),
.Y(n_2551)
);

INVx1_ASAP7_75t_L g2552 ( 
.A(n_2379),
.Y(n_2552)
);

BUFx2_ASAP7_75t_L g2553 ( 
.A(n_2535),
.Y(n_2553)
);

NAND2xp5_ASAP7_75t_L g2554 ( 
.A(n_2378),
.B(n_187),
.Y(n_2554)
);

OAI21xp5_ASAP7_75t_SL g2555 ( 
.A1(n_2410),
.A2(n_188),
.B(n_189),
.Y(n_2555)
);

INVx1_ASAP7_75t_L g2556 ( 
.A(n_2387),
.Y(n_2556)
);

OR2x2_ASAP7_75t_L g2557 ( 
.A(n_2407),
.B(n_189),
.Y(n_2557)
);

INVx2_ASAP7_75t_L g2558 ( 
.A(n_2467),
.Y(n_2558)
);

INVx3_ASAP7_75t_L g2559 ( 
.A(n_2533),
.Y(n_2559)
);

AOI21xp5_ASAP7_75t_L g2560 ( 
.A1(n_2490),
.A2(n_190),
.B(n_191),
.Y(n_2560)
);

OAI31xp33_ASAP7_75t_L g2561 ( 
.A1(n_2517),
.A2(n_193),
.A3(n_190),
.B(n_192),
.Y(n_2561)
);

AND2x2_ASAP7_75t_L g2562 ( 
.A(n_2381),
.B(n_192),
.Y(n_2562)
);

INVx1_ASAP7_75t_L g2563 ( 
.A(n_2390),
.Y(n_2563)
);

AND2x2_ASAP7_75t_L g2564 ( 
.A(n_2441),
.B(n_193),
.Y(n_2564)
);

INVx3_ASAP7_75t_L g2565 ( 
.A(n_2533),
.Y(n_2565)
);

INVx2_ASAP7_75t_SL g2566 ( 
.A(n_2377),
.Y(n_2566)
);

NAND2xp5_ASAP7_75t_L g2567 ( 
.A(n_2523),
.B(n_194),
.Y(n_2567)
);

NAND4xp25_ASAP7_75t_L g2568 ( 
.A(n_2405),
.B(n_2434),
.C(n_2492),
.D(n_2489),
.Y(n_2568)
);

INVx1_ASAP7_75t_L g2569 ( 
.A(n_2391),
.Y(n_2569)
);

AND2x2_ASAP7_75t_L g2570 ( 
.A(n_2446),
.B(n_196),
.Y(n_2570)
);

NAND3xp33_ASAP7_75t_L g2571 ( 
.A(n_2532),
.B(n_196),
.C(n_197),
.Y(n_2571)
);

INVx2_ASAP7_75t_L g2572 ( 
.A(n_2480),
.Y(n_2572)
);

INVx2_ASAP7_75t_L g2573 ( 
.A(n_2478),
.Y(n_2573)
);

AOI221xp5_ASAP7_75t_L g2574 ( 
.A1(n_2494),
.A2(n_199),
.B1(n_197),
.B2(n_198),
.C(n_200),
.Y(n_2574)
);

AND2x2_ASAP7_75t_L g2575 ( 
.A(n_2438),
.B(n_198),
.Y(n_2575)
);

BUFx2_ASAP7_75t_L g2576 ( 
.A(n_2501),
.Y(n_2576)
);

INVx1_ASAP7_75t_L g2577 ( 
.A(n_2393),
.Y(n_2577)
);

AOI22xp33_ASAP7_75t_L g2578 ( 
.A1(n_2502),
.A2(n_201),
.B1(n_199),
.B2(n_200),
.Y(n_2578)
);

INVx1_ASAP7_75t_L g2579 ( 
.A(n_2396),
.Y(n_2579)
);

INVx1_ASAP7_75t_L g2580 ( 
.A(n_2401),
.Y(n_2580)
);

AOI211xp5_ASAP7_75t_L g2581 ( 
.A1(n_2514),
.A2(n_204),
.B(n_202),
.C(n_203),
.Y(n_2581)
);

INVx2_ASAP7_75t_L g2582 ( 
.A(n_2470),
.Y(n_2582)
);

NAND2xp5_ASAP7_75t_L g2583 ( 
.A(n_2527),
.B(n_202),
.Y(n_2583)
);

AND2x2_ASAP7_75t_L g2584 ( 
.A(n_2479),
.B(n_203),
.Y(n_2584)
);

AND2x2_ASAP7_75t_L g2585 ( 
.A(n_2449),
.B(n_204),
.Y(n_2585)
);

AOI222xp33_ASAP7_75t_L g2586 ( 
.A1(n_2536),
.A2(n_229),
.B1(n_213),
.B2(n_237),
.C1(n_221),
.C2(n_205),
.Y(n_2586)
);

AND2x2_ASAP7_75t_L g2587 ( 
.A(n_2389),
.B(n_205),
.Y(n_2587)
);

AOI22xp33_ASAP7_75t_L g2588 ( 
.A1(n_2538),
.A2(n_208),
.B1(n_206),
.B2(n_207),
.Y(n_2588)
);

INVx2_ASAP7_75t_SL g2589 ( 
.A(n_2507),
.Y(n_2589)
);

HB1xp67_ASAP7_75t_L g2590 ( 
.A(n_2539),
.Y(n_2590)
);

INVx1_ASAP7_75t_L g2591 ( 
.A(n_2406),
.Y(n_2591)
);

BUFx3_ASAP7_75t_L g2592 ( 
.A(n_2471),
.Y(n_2592)
);

AND2x2_ASAP7_75t_L g2593 ( 
.A(n_2380),
.B(n_206),
.Y(n_2593)
);

INVx1_ASAP7_75t_L g2594 ( 
.A(n_2503),
.Y(n_2594)
);

HB1xp67_ASAP7_75t_L g2595 ( 
.A(n_2544),
.Y(n_2595)
);

INVx2_ASAP7_75t_L g2596 ( 
.A(n_2481),
.Y(n_2596)
);

OR2x2_ASAP7_75t_L g2597 ( 
.A(n_2448),
.B(n_207),
.Y(n_2597)
);

AOI22xp33_ASAP7_75t_L g2598 ( 
.A1(n_2433),
.A2(n_210),
.B1(n_208),
.B2(n_209),
.Y(n_2598)
);

INVx2_ASAP7_75t_SL g2599 ( 
.A(n_2525),
.Y(n_2599)
);

INVx2_ASAP7_75t_L g2600 ( 
.A(n_2498),
.Y(n_2600)
);

AOI221xp5_ASAP7_75t_L g2601 ( 
.A1(n_2493),
.A2(n_212),
.B1(n_210),
.B2(n_211),
.C(n_213),
.Y(n_2601)
);

OAI22xp5_ASAP7_75t_L g2602 ( 
.A1(n_2388),
.A2(n_215),
.B1(n_212),
.B2(n_214),
.Y(n_2602)
);

AND2x2_ASAP7_75t_L g2603 ( 
.A(n_2495),
.B(n_214),
.Y(n_2603)
);

AO21x2_ASAP7_75t_L g2604 ( 
.A1(n_2395),
.A2(n_215),
.B(n_216),
.Y(n_2604)
);

INVx2_ASAP7_75t_L g2605 ( 
.A(n_2457),
.Y(n_2605)
);

AND2x2_ASAP7_75t_L g2606 ( 
.A(n_2496),
.B(n_217),
.Y(n_2606)
);

BUFx3_ASAP7_75t_L g2607 ( 
.A(n_2451),
.Y(n_2607)
);

INVx2_ASAP7_75t_L g2608 ( 
.A(n_2497),
.Y(n_2608)
);

INVx1_ASAP7_75t_L g2609 ( 
.A(n_2508),
.Y(n_2609)
);

AOI22xp33_ASAP7_75t_SL g2610 ( 
.A1(n_2484),
.A2(n_219),
.B1(n_217),
.B2(n_218),
.Y(n_2610)
);

INVx2_ASAP7_75t_L g2611 ( 
.A(n_2504),
.Y(n_2611)
);

INVx2_ASAP7_75t_L g2612 ( 
.A(n_2526),
.Y(n_2612)
);

OAI31xp33_ASAP7_75t_L g2613 ( 
.A1(n_2491),
.A2(n_220),
.A3(n_218),
.B(n_219),
.Y(n_2613)
);

AND2x2_ASAP7_75t_L g2614 ( 
.A(n_2499),
.B(n_220),
.Y(n_2614)
);

INVx1_ASAP7_75t_L g2615 ( 
.A(n_2510),
.Y(n_2615)
);

AND2x2_ASAP7_75t_L g2616 ( 
.A(n_2509),
.B(n_2513),
.Y(n_2616)
);

INVxp67_ASAP7_75t_L g2617 ( 
.A(n_2464),
.Y(n_2617)
);

BUFx2_ASAP7_75t_L g2618 ( 
.A(n_2414),
.Y(n_2618)
);

OAI221xp5_ASAP7_75t_L g2619 ( 
.A1(n_2383),
.A2(n_223),
.B1(n_221),
.B2(n_222),
.C(n_224),
.Y(n_2619)
);

INVx1_ASAP7_75t_L g2620 ( 
.A(n_2512),
.Y(n_2620)
);

INVx2_ASAP7_75t_L g2621 ( 
.A(n_2485),
.Y(n_2621)
);

INVx2_ASAP7_75t_L g2622 ( 
.A(n_2442),
.Y(n_2622)
);

INVxp67_ASAP7_75t_SL g2623 ( 
.A(n_2541),
.Y(n_2623)
);

INVx1_ASAP7_75t_L g2624 ( 
.A(n_2529),
.Y(n_2624)
);

NAND2xp5_ASAP7_75t_SL g2625 ( 
.A(n_2439),
.B(n_2447),
.Y(n_2625)
);

OAI22xp5_ASAP7_75t_L g2626 ( 
.A1(n_2417),
.A2(n_225),
.B1(n_223),
.B2(n_224),
.Y(n_2626)
);

BUFx2_ASAP7_75t_L g2627 ( 
.A(n_2403),
.Y(n_2627)
);

INVx1_ASAP7_75t_L g2628 ( 
.A(n_2534),
.Y(n_2628)
);

AOI222xp33_ASAP7_75t_L g2629 ( 
.A1(n_2424),
.A2(n_252),
.B1(n_234),
.B2(n_261),
.C1(n_243),
.C2(n_225),
.Y(n_2629)
);

BUFx3_ASAP7_75t_L g2630 ( 
.A(n_2394),
.Y(n_2630)
);

INVxp67_ASAP7_75t_L g2631 ( 
.A(n_2386),
.Y(n_2631)
);

AND2x2_ASAP7_75t_L g2632 ( 
.A(n_2516),
.B(n_226),
.Y(n_2632)
);

AOI22xp5_ASAP7_75t_L g2633 ( 
.A1(n_2542),
.A2(n_228),
.B1(n_226),
.B2(n_227),
.Y(n_2633)
);

INVx1_ASAP7_75t_L g2634 ( 
.A(n_2537),
.Y(n_2634)
);

OAI211xp5_ASAP7_75t_SL g2635 ( 
.A1(n_2472),
.A2(n_2445),
.B(n_2404),
.C(n_2425),
.Y(n_2635)
);

AOI322xp5_ASAP7_75t_L g2636 ( 
.A1(n_2440),
.A2(n_233),
.A3(n_232),
.B1(n_230),
.B2(n_227),
.C1(n_228),
.C2(n_231),
.Y(n_2636)
);

OAI221xp5_ASAP7_75t_L g2637 ( 
.A1(n_2450),
.A2(n_232),
.B1(n_230),
.B2(n_231),
.C(n_233),
.Y(n_2637)
);

OAI21xp5_ASAP7_75t_L g2638 ( 
.A1(n_2384),
.A2(n_235),
.B(n_236),
.Y(n_2638)
);

INVx1_ASAP7_75t_L g2639 ( 
.A(n_2419),
.Y(n_2639)
);

AO21x2_ASAP7_75t_L g2640 ( 
.A1(n_2518),
.A2(n_235),
.B(n_236),
.Y(n_2640)
);

INVx1_ASAP7_75t_L g2641 ( 
.A(n_2422),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_2427),
.Y(n_2642)
);

INVx2_ASAP7_75t_L g2643 ( 
.A(n_2385),
.Y(n_2643)
);

INVxp67_ASAP7_75t_SL g2644 ( 
.A(n_2429),
.Y(n_2644)
);

INVx2_ASAP7_75t_L g2645 ( 
.A(n_2418),
.Y(n_2645)
);

INVx1_ASAP7_75t_L g2646 ( 
.A(n_2428),
.Y(n_2646)
);

INVx1_ASAP7_75t_L g2647 ( 
.A(n_2408),
.Y(n_2647)
);

INVx1_ASAP7_75t_L g2648 ( 
.A(n_2411),
.Y(n_2648)
);

INVx1_ASAP7_75t_SL g2649 ( 
.A(n_2376),
.Y(n_2649)
);

NOR2xp67_ASAP7_75t_L g2650 ( 
.A(n_2437),
.B(n_238),
.Y(n_2650)
);

INVx1_ASAP7_75t_L g2651 ( 
.A(n_2413),
.Y(n_2651)
);

NAND3xp33_ASAP7_75t_L g2652 ( 
.A(n_2520),
.B(n_238),
.C(n_239),
.Y(n_2652)
);

AOI221xp5_ASAP7_75t_L g2653 ( 
.A1(n_2397),
.A2(n_241),
.B1(n_239),
.B2(n_240),
.C(n_242),
.Y(n_2653)
);

AND2x2_ASAP7_75t_L g2654 ( 
.A(n_2519),
.B(n_240),
.Y(n_2654)
);

INVx2_ASAP7_75t_L g2655 ( 
.A(n_2421),
.Y(n_2655)
);

AOI22xp33_ASAP7_75t_SL g2656 ( 
.A1(n_2486),
.A2(n_243),
.B1(n_241),
.B2(n_242),
.Y(n_2656)
);

NAND4xp25_ASAP7_75t_L g2657 ( 
.A(n_2420),
.B(n_247),
.C(n_245),
.D(n_246),
.Y(n_2657)
);

AND2x2_ASAP7_75t_L g2658 ( 
.A(n_2524),
.B(n_245),
.Y(n_2658)
);

OAI22xp5_ASAP7_75t_L g2659 ( 
.A1(n_2522),
.A2(n_248),
.B1(n_246),
.B2(n_247),
.Y(n_2659)
);

BUFx2_ASAP7_75t_L g2660 ( 
.A(n_2500),
.Y(n_2660)
);

INVx1_ASAP7_75t_L g2661 ( 
.A(n_2531),
.Y(n_2661)
);

NAND2xp5_ASAP7_75t_L g2662 ( 
.A(n_2423),
.B(n_248),
.Y(n_2662)
);

AND2x2_ASAP7_75t_SL g2663 ( 
.A(n_2528),
.B(n_249),
.Y(n_2663)
);

AND2x2_ASAP7_75t_L g2664 ( 
.A(n_2540),
.B(n_249),
.Y(n_2664)
);

INVx2_ASAP7_75t_L g2665 ( 
.A(n_2443),
.Y(n_2665)
);

INVx2_ASAP7_75t_L g2666 ( 
.A(n_2444),
.Y(n_2666)
);

AND4x1_ASAP7_75t_L g2667 ( 
.A(n_2543),
.B(n_252),
.C(n_250),
.D(n_251),
.Y(n_2667)
);

AND2x2_ASAP7_75t_L g2668 ( 
.A(n_2553),
.B(n_2426),
.Y(n_2668)
);

INVx1_ASAP7_75t_SL g2669 ( 
.A(n_2663),
.Y(n_2669)
);

AND2x2_ASAP7_75t_L g2670 ( 
.A(n_2616),
.B(n_2402),
.Y(n_2670)
);

INVx1_ASAP7_75t_L g2671 ( 
.A(n_2546),
.Y(n_2671)
);

AND2x2_ASAP7_75t_L g2672 ( 
.A(n_2566),
.B(n_2506),
.Y(n_2672)
);

OR2x2_ASAP7_75t_L g2673 ( 
.A(n_2576),
.B(n_2436),
.Y(n_2673)
);

NAND2x1p5_ASAP7_75t_L g2674 ( 
.A(n_2545),
.B(n_2416),
.Y(n_2674)
);

INVx1_ASAP7_75t_L g2675 ( 
.A(n_2575),
.Y(n_2675)
);

HB1xp67_ASAP7_75t_L g2676 ( 
.A(n_2631),
.Y(n_2676)
);

AND2x2_ASAP7_75t_L g2677 ( 
.A(n_2551),
.B(n_2521),
.Y(n_2677)
);

HB1xp67_ASAP7_75t_L g2678 ( 
.A(n_2590),
.Y(n_2678)
);

OR2x2_ASAP7_75t_L g2679 ( 
.A(n_2627),
.B(n_2458),
.Y(n_2679)
);

OR2x2_ASAP7_75t_L g2680 ( 
.A(n_2573),
.B(n_2466),
.Y(n_2680)
);

NOR2x1_ASAP7_75t_L g2681 ( 
.A(n_2555),
.B(n_2399),
.Y(n_2681)
);

INVx2_ASAP7_75t_L g2682 ( 
.A(n_2660),
.Y(n_2682)
);

NAND2xp5_ASAP7_75t_L g2683 ( 
.A(n_2644),
.B(n_2487),
.Y(n_2683)
);

INVx1_ASAP7_75t_L g2684 ( 
.A(n_2622),
.Y(n_2684)
);

INVxp67_ASAP7_75t_L g2685 ( 
.A(n_2550),
.Y(n_2685)
);

INVx1_ASAP7_75t_SL g2686 ( 
.A(n_2607),
.Y(n_2686)
);

INVx2_ASAP7_75t_L g2687 ( 
.A(n_2548),
.Y(n_2687)
);

AND2x4_ASAP7_75t_L g2688 ( 
.A(n_2630),
.B(n_2455),
.Y(n_2688)
);

INVx1_ASAP7_75t_L g2689 ( 
.A(n_2547),
.Y(n_2689)
);

NOR2xp33_ASAP7_75t_L g2690 ( 
.A(n_2635),
.B(n_2453),
.Y(n_2690)
);

INVx1_ASAP7_75t_L g2691 ( 
.A(n_2552),
.Y(n_2691)
);

NAND2xp5_ASAP7_75t_L g2692 ( 
.A(n_2608),
.B(n_2459),
.Y(n_2692)
);

INVx2_ASAP7_75t_L g2693 ( 
.A(n_2558),
.Y(n_2693)
);

AND2x2_ASAP7_75t_L g2694 ( 
.A(n_2559),
.B(n_2398),
.Y(n_2694)
);

NAND2xp5_ASAP7_75t_R g2695 ( 
.A(n_2589),
.B(n_2599),
.Y(n_2695)
);

AND2x2_ASAP7_75t_L g2696 ( 
.A(n_2565),
.B(n_2430),
.Y(n_2696)
);

OR2x2_ASAP7_75t_L g2697 ( 
.A(n_2568),
.B(n_2432),
.Y(n_2697)
);

INVx2_ASAP7_75t_L g2698 ( 
.A(n_2592),
.Y(n_2698)
);

AND2x2_ASAP7_75t_L g2699 ( 
.A(n_2562),
.B(n_2456),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_2556),
.Y(n_2700)
);

INVx2_ASAP7_75t_L g2701 ( 
.A(n_2545),
.Y(n_2701)
);

INVx1_ASAP7_75t_L g2702 ( 
.A(n_2563),
.Y(n_2702)
);

OR2x2_ASAP7_75t_L g2703 ( 
.A(n_2661),
.B(n_2409),
.Y(n_2703)
);

AND2x2_ASAP7_75t_L g2704 ( 
.A(n_2572),
.B(n_2468),
.Y(n_2704)
);

NAND2xp5_ASAP7_75t_L g2705 ( 
.A(n_2611),
.B(n_2461),
.Y(n_2705)
);

BUFx2_ASAP7_75t_L g2706 ( 
.A(n_2600),
.Y(n_2706)
);

AND2x2_ASAP7_75t_L g2707 ( 
.A(n_2584),
.B(n_2400),
.Y(n_2707)
);

NAND2xp5_ASAP7_75t_L g2708 ( 
.A(n_2612),
.B(n_2415),
.Y(n_2708)
);

OR2x2_ASAP7_75t_L g2709 ( 
.A(n_2618),
.B(n_2557),
.Y(n_2709)
);

OR2x2_ASAP7_75t_L g2710 ( 
.A(n_2583),
.B(n_2469),
.Y(n_2710)
);

INVx1_ASAP7_75t_SL g2711 ( 
.A(n_2649),
.Y(n_2711)
);

NAND2xp5_ASAP7_75t_L g2712 ( 
.A(n_2604),
.B(n_2473),
.Y(n_2712)
);

INVx1_ASAP7_75t_L g2713 ( 
.A(n_2569),
.Y(n_2713)
);

INVx1_ASAP7_75t_L g2714 ( 
.A(n_2577),
.Y(n_2714)
);

INVxp67_ASAP7_75t_SL g2715 ( 
.A(n_2617),
.Y(n_2715)
);

NAND2xp5_ASAP7_75t_L g2716 ( 
.A(n_2640),
.B(n_2476),
.Y(n_2716)
);

INVxp67_ASAP7_75t_L g2717 ( 
.A(n_2623),
.Y(n_2717)
);

INVxp33_ASAP7_75t_L g2718 ( 
.A(n_2650),
.Y(n_2718)
);

INVx2_ASAP7_75t_SL g2719 ( 
.A(n_2564),
.Y(n_2719)
);

AND2x2_ASAP7_75t_L g2720 ( 
.A(n_2570),
.B(n_2474),
.Y(n_2720)
);

INVx1_ASAP7_75t_L g2721 ( 
.A(n_2579),
.Y(n_2721)
);

AND2x2_ASAP7_75t_L g2722 ( 
.A(n_2585),
.B(n_2625),
.Y(n_2722)
);

HB1xp67_ASAP7_75t_L g2723 ( 
.A(n_2595),
.Y(n_2723)
);

INVx1_ASAP7_75t_L g2724 ( 
.A(n_2580),
.Y(n_2724)
);

NAND2xp5_ASAP7_75t_L g2725 ( 
.A(n_2554),
.B(n_2477),
.Y(n_2725)
);

OR2x2_ASAP7_75t_L g2726 ( 
.A(n_2567),
.B(n_2465),
.Y(n_2726)
);

AND2x2_ASAP7_75t_L g2727 ( 
.A(n_2621),
.B(n_2412),
.Y(n_2727)
);

NAND2xp5_ASAP7_75t_L g2728 ( 
.A(n_2676),
.B(n_2561),
.Y(n_2728)
);

AND2x2_ASAP7_75t_L g2729 ( 
.A(n_2670),
.B(n_2591),
.Y(n_2729)
);

INVx2_ASAP7_75t_L g2730 ( 
.A(n_2720),
.Y(n_2730)
);

HB1xp67_ASAP7_75t_L g2731 ( 
.A(n_2711),
.Y(n_2731)
);

AND2x2_ASAP7_75t_L g2732 ( 
.A(n_2685),
.B(n_2594),
.Y(n_2732)
);

OAI21xp5_ASAP7_75t_L g2733 ( 
.A1(n_2681),
.A2(n_2560),
.B(n_2571),
.Y(n_2733)
);

INVx2_ASAP7_75t_L g2734 ( 
.A(n_2699),
.Y(n_2734)
);

NAND4xp25_ASAP7_75t_L g2735 ( 
.A(n_2682),
.B(n_2549),
.C(n_2581),
.D(n_2657),
.Y(n_2735)
);

INVx1_ASAP7_75t_L g2736 ( 
.A(n_2678),
.Y(n_2736)
);

OR2x2_ASAP7_75t_L g2737 ( 
.A(n_2715),
.B(n_2597),
.Y(n_2737)
);

INVx1_ASAP7_75t_L g2738 ( 
.A(n_2723),
.Y(n_2738)
);

INVx1_ASAP7_75t_L g2739 ( 
.A(n_2703),
.Y(n_2739)
);

AND2x2_ASAP7_75t_L g2740 ( 
.A(n_2686),
.B(n_2668),
.Y(n_2740)
);

AND2x2_ASAP7_75t_L g2741 ( 
.A(n_2677),
.B(n_2696),
.Y(n_2741)
);

OR2x2_ASAP7_75t_L g2742 ( 
.A(n_2673),
.B(n_2609),
.Y(n_2742)
);

INVx2_ASAP7_75t_L g2743 ( 
.A(n_2674),
.Y(n_2743)
);

HB1xp67_ASAP7_75t_L g2744 ( 
.A(n_2717),
.Y(n_2744)
);

NAND2xp5_ASAP7_75t_L g2745 ( 
.A(n_2690),
.B(n_2610),
.Y(n_2745)
);

BUFx2_ASAP7_75t_L g2746 ( 
.A(n_2688),
.Y(n_2746)
);

OR2x2_ASAP7_75t_L g2747 ( 
.A(n_2683),
.B(n_2615),
.Y(n_2747)
);

AND2x2_ASAP7_75t_L g2748 ( 
.A(n_2672),
.B(n_2620),
.Y(n_2748)
);

INVx1_ASAP7_75t_L g2749 ( 
.A(n_2671),
.Y(n_2749)
);

INVx1_ASAP7_75t_L g2750 ( 
.A(n_2684),
.Y(n_2750)
);

INVx1_ASAP7_75t_L g2751 ( 
.A(n_2689),
.Y(n_2751)
);

INVx1_ASAP7_75t_L g2752 ( 
.A(n_2691),
.Y(n_2752)
);

NOR2xp33_ASAP7_75t_L g2753 ( 
.A(n_2710),
.B(n_2667),
.Y(n_2753)
);

INVx1_ASAP7_75t_L g2754 ( 
.A(n_2700),
.Y(n_2754)
);

INVx1_ASAP7_75t_L g2755 ( 
.A(n_2702),
.Y(n_2755)
);

INVx2_ASAP7_75t_L g2756 ( 
.A(n_2688),
.Y(n_2756)
);

INVx2_ASAP7_75t_L g2757 ( 
.A(n_2707),
.Y(n_2757)
);

INVx1_ASAP7_75t_L g2758 ( 
.A(n_2713),
.Y(n_2758)
);

AND2x2_ASAP7_75t_L g2759 ( 
.A(n_2694),
.B(n_2624),
.Y(n_2759)
);

OR2x2_ASAP7_75t_L g2760 ( 
.A(n_2731),
.B(n_2679),
.Y(n_2760)
);

INVx2_ASAP7_75t_L g2761 ( 
.A(n_2740),
.Y(n_2761)
);

AND2x2_ASAP7_75t_L g2762 ( 
.A(n_2746),
.B(n_2698),
.Y(n_2762)
);

NAND2xp5_ASAP7_75t_L g2763 ( 
.A(n_2729),
.B(n_2675),
.Y(n_2763)
);

NAND2xp5_ASAP7_75t_L g2764 ( 
.A(n_2759),
.B(n_2719),
.Y(n_2764)
);

AND2x2_ASAP7_75t_L g2765 ( 
.A(n_2741),
.B(n_2704),
.Y(n_2765)
);

AND2x2_ASAP7_75t_L g2766 ( 
.A(n_2730),
.B(n_2722),
.Y(n_2766)
);

INVx1_ASAP7_75t_L g2767 ( 
.A(n_2744),
.Y(n_2767)
);

NAND4xp25_ASAP7_75t_L g2768 ( 
.A(n_2756),
.B(n_2706),
.C(n_2709),
.D(n_2697),
.Y(n_2768)
);

AND2x2_ASAP7_75t_L g2769 ( 
.A(n_2734),
.B(n_2757),
.Y(n_2769)
);

INVx2_ASAP7_75t_L g2770 ( 
.A(n_2737),
.Y(n_2770)
);

NAND2xp5_ASAP7_75t_L g2771 ( 
.A(n_2753),
.B(n_2669),
.Y(n_2771)
);

NOR3xp33_ASAP7_75t_L g2772 ( 
.A(n_2728),
.B(n_2716),
.C(n_2712),
.Y(n_2772)
);

INVx1_ASAP7_75t_L g2773 ( 
.A(n_2736),
.Y(n_2773)
);

OR2x2_ASAP7_75t_L g2774 ( 
.A(n_2742),
.B(n_2680),
.Y(n_2774)
);

NAND2xp5_ASAP7_75t_L g2775 ( 
.A(n_2748),
.B(n_2708),
.Y(n_2775)
);

INVx1_ASAP7_75t_L g2776 ( 
.A(n_2738),
.Y(n_2776)
);

NAND2xp5_ASAP7_75t_L g2777 ( 
.A(n_2745),
.B(n_2692),
.Y(n_2777)
);

HB1xp67_ASAP7_75t_L g2778 ( 
.A(n_2732),
.Y(n_2778)
);

HB1xp67_ASAP7_75t_L g2779 ( 
.A(n_2743),
.Y(n_2779)
);

INVx1_ASAP7_75t_L g2780 ( 
.A(n_2760),
.Y(n_2780)
);

NAND2xp5_ASAP7_75t_L g2781 ( 
.A(n_2765),
.B(n_2761),
.Y(n_2781)
);

OR2x2_ASAP7_75t_L g2782 ( 
.A(n_2774),
.B(n_2739),
.Y(n_2782)
);

OR2x2_ASAP7_75t_L g2783 ( 
.A(n_2770),
.B(n_2747),
.Y(n_2783)
);

INVx4_ASAP7_75t_L g2784 ( 
.A(n_2762),
.Y(n_2784)
);

NAND2xp5_ASAP7_75t_L g2785 ( 
.A(n_2778),
.B(n_2766),
.Y(n_2785)
);

INVx2_ASAP7_75t_L g2786 ( 
.A(n_2769),
.Y(n_2786)
);

INVx1_ASAP7_75t_L g2787 ( 
.A(n_2779),
.Y(n_2787)
);

OR2x2_ASAP7_75t_L g2788 ( 
.A(n_2763),
.B(n_2735),
.Y(n_2788)
);

INVx2_ASAP7_75t_SL g2789 ( 
.A(n_2764),
.Y(n_2789)
);

INVx1_ASAP7_75t_L g2790 ( 
.A(n_2785),
.Y(n_2790)
);

INVx1_ASAP7_75t_L g2791 ( 
.A(n_2782),
.Y(n_2791)
);

INVx3_ASAP7_75t_L g2792 ( 
.A(n_2784),
.Y(n_2792)
);

INVx2_ASAP7_75t_L g2793 ( 
.A(n_2783),
.Y(n_2793)
);

AOI322xp5_ASAP7_75t_L g2794 ( 
.A1(n_2787),
.A2(n_2772),
.A3(n_2777),
.B1(n_2771),
.B2(n_2767),
.C1(n_2775),
.C2(n_2750),
.Y(n_2794)
);

INVx1_ASAP7_75t_L g2795 ( 
.A(n_2781),
.Y(n_2795)
);

XNOR2x1_ASAP7_75t_L g2796 ( 
.A(n_2788),
.B(n_2733),
.Y(n_2796)
);

NAND2xp5_ASAP7_75t_L g2797 ( 
.A(n_2786),
.B(n_2725),
.Y(n_2797)
);

A2O1A1Ixp33_ASAP7_75t_L g2798 ( 
.A1(n_2780),
.A2(n_2718),
.B(n_2638),
.C(n_2652),
.Y(n_2798)
);

NAND2x1_ASAP7_75t_L g2799 ( 
.A(n_2792),
.B(n_2789),
.Y(n_2799)
);

NAND2xp5_ASAP7_75t_L g2800 ( 
.A(n_2793),
.B(n_2701),
.Y(n_2800)
);

INVx1_ASAP7_75t_L g2801 ( 
.A(n_2791),
.Y(n_2801)
);

INVx1_ASAP7_75t_L g2802 ( 
.A(n_2797),
.Y(n_2802)
);

AND2x2_ASAP7_75t_L g2803 ( 
.A(n_2795),
.B(n_2727),
.Y(n_2803)
);

NAND2xp5_ASAP7_75t_SL g2804 ( 
.A(n_2794),
.B(n_2798),
.Y(n_2804)
);

INVx1_ASAP7_75t_L g2805 ( 
.A(n_2790),
.Y(n_2805)
);

NAND2xp5_ASAP7_75t_L g2806 ( 
.A(n_2796),
.B(n_2705),
.Y(n_2806)
);

INVx1_ASAP7_75t_SL g2807 ( 
.A(n_2796),
.Y(n_2807)
);

NAND2xp5_ASAP7_75t_L g2808 ( 
.A(n_2793),
.B(n_2749),
.Y(n_2808)
);

NAND2xp5_ASAP7_75t_L g2809 ( 
.A(n_2793),
.B(n_2752),
.Y(n_2809)
);

INVx2_ASAP7_75t_L g2810 ( 
.A(n_2793),
.Y(n_2810)
);

AND2x2_ASAP7_75t_L g2811 ( 
.A(n_2792),
.B(n_2773),
.Y(n_2811)
);

NAND2xp5_ASAP7_75t_L g2812 ( 
.A(n_2793),
.B(n_2754),
.Y(n_2812)
);

INVx1_ASAP7_75t_L g2813 ( 
.A(n_2793),
.Y(n_2813)
);

NOR2xp33_ASAP7_75t_L g2814 ( 
.A(n_2796),
.B(n_2768),
.Y(n_2814)
);

INVx1_ASAP7_75t_L g2815 ( 
.A(n_2793),
.Y(n_2815)
);

NAND2x1_ASAP7_75t_L g2816 ( 
.A(n_2792),
.B(n_2751),
.Y(n_2816)
);

NOR3xp33_ASAP7_75t_SL g2817 ( 
.A(n_2804),
.B(n_2776),
.C(n_2751),
.Y(n_2817)
);

AOI22xp5_ASAP7_75t_L g2818 ( 
.A1(n_2807),
.A2(n_2693),
.B1(n_2687),
.B2(n_2726),
.Y(n_2818)
);

INVx2_ASAP7_75t_L g2819 ( 
.A(n_2803),
.Y(n_2819)
);

INVx1_ASAP7_75t_L g2820 ( 
.A(n_2810),
.Y(n_2820)
);

NOR3xp33_ASAP7_75t_SL g2821 ( 
.A(n_2814),
.B(n_2758),
.C(n_2755),
.Y(n_2821)
);

OR2x2_ASAP7_75t_L g2822 ( 
.A(n_2806),
.B(n_2714),
.Y(n_2822)
);

NAND2xp5_ASAP7_75t_SL g2823 ( 
.A(n_2813),
.B(n_2721),
.Y(n_2823)
);

XOR2x2_ASAP7_75t_L g2824 ( 
.A(n_2800),
.B(n_2626),
.Y(n_2824)
);

BUFx3_ASAP7_75t_L g2825 ( 
.A(n_2799),
.Y(n_2825)
);

NAND3xp33_ASAP7_75t_L g2826 ( 
.A(n_2815),
.B(n_2601),
.C(n_2586),
.Y(n_2826)
);

XNOR2xp5_ASAP7_75t_L g2827 ( 
.A(n_2811),
.B(n_2633),
.Y(n_2827)
);

NAND2xp5_ASAP7_75t_L g2828 ( 
.A(n_2802),
.B(n_2724),
.Y(n_2828)
);

NAND2xp5_ASAP7_75t_L g2829 ( 
.A(n_2805),
.B(n_2587),
.Y(n_2829)
);

NOR2xp33_ASAP7_75t_L g2830 ( 
.A(n_2816),
.B(n_2808),
.Y(n_2830)
);

CKINVDCx20_ASAP7_75t_L g2831 ( 
.A(n_2812),
.Y(n_2831)
);

INVx1_ASAP7_75t_L g2832 ( 
.A(n_2809),
.Y(n_2832)
);

INVx1_ASAP7_75t_L g2833 ( 
.A(n_2801),
.Y(n_2833)
);

AND3x2_ASAP7_75t_L g2834 ( 
.A(n_2814),
.B(n_2603),
.C(n_2593),
.Y(n_2834)
);

AND2x2_ASAP7_75t_L g2835 ( 
.A(n_2803),
.B(n_2628),
.Y(n_2835)
);

AND2x4_ASAP7_75t_L g2836 ( 
.A(n_2810),
.B(n_2634),
.Y(n_2836)
);

INVx1_ASAP7_75t_L g2837 ( 
.A(n_2829),
.Y(n_2837)
);

OAI21xp33_ASAP7_75t_L g2838 ( 
.A1(n_2817),
.A2(n_2821),
.B(n_2825),
.Y(n_2838)
);

NAND2xp5_ASAP7_75t_L g2839 ( 
.A(n_2834),
.B(n_2639),
.Y(n_2839)
);

NOR2x1_ASAP7_75t_L g2840 ( 
.A(n_2819),
.B(n_2662),
.Y(n_2840)
);

OAI321xp33_ASAP7_75t_L g2841 ( 
.A1(n_2818),
.A2(n_2574),
.A3(n_2619),
.B1(n_2637),
.B2(n_2588),
.C(n_2578),
.Y(n_2841)
);

AND3x1_ASAP7_75t_L g2842 ( 
.A(n_2830),
.B(n_2832),
.C(n_2820),
.Y(n_2842)
);

NOR2xp33_ASAP7_75t_L g2843 ( 
.A(n_2827),
.B(n_2606),
.Y(n_2843)
);

OR2x2_ASAP7_75t_L g2844 ( 
.A(n_2822),
.B(n_2641),
.Y(n_2844)
);

AOI21xp33_ASAP7_75t_L g2845 ( 
.A1(n_2833),
.A2(n_2659),
.B(n_2629),
.Y(n_2845)
);

INVx1_ASAP7_75t_L g2846 ( 
.A(n_2835),
.Y(n_2846)
);

NOR3xp33_ASAP7_75t_L g2847 ( 
.A(n_2823),
.B(n_2828),
.C(n_2826),
.Y(n_2847)
);

NAND2xp5_ASAP7_75t_L g2848 ( 
.A(n_2836),
.B(n_2642),
.Y(n_2848)
);

NOR3xp33_ASAP7_75t_L g2849 ( 
.A(n_2831),
.B(n_2653),
.C(n_2602),
.Y(n_2849)
);

CKINVDCx5p33_ASAP7_75t_R g2850 ( 
.A(n_2824),
.Y(n_2850)
);

NAND4xp25_ASAP7_75t_L g2851 ( 
.A(n_2836),
.B(n_2636),
.C(n_2656),
.D(n_2613),
.Y(n_2851)
);

NOR3xp33_ASAP7_75t_L g2852 ( 
.A(n_2830),
.B(n_2632),
.C(n_2614),
.Y(n_2852)
);

AOI22xp5_ASAP7_75t_L g2853 ( 
.A1(n_2820),
.A2(n_2664),
.B1(n_2654),
.B2(n_2658),
.Y(n_2853)
);

NOR3x1_ASAP7_75t_SL g2854 ( 
.A(n_2831),
.B(n_2695),
.C(n_2463),
.Y(n_2854)
);

AOI21xp5_ASAP7_75t_L g2855 ( 
.A1(n_2829),
.A2(n_2647),
.B(n_2646),
.Y(n_2855)
);

AOI211xp5_ASAP7_75t_L g2856 ( 
.A1(n_2830),
.A2(n_2648),
.B(n_2651),
.C(n_2605),
.Y(n_2856)
);

NOR3xp33_ASAP7_75t_L g2857 ( 
.A(n_2830),
.B(n_2596),
.C(n_2582),
.Y(n_2857)
);

AOI221xp5_ASAP7_75t_L g2858 ( 
.A1(n_2845),
.A2(n_2598),
.B1(n_2655),
.B2(n_2645),
.C(n_2643),
.Y(n_2858)
);

NAND4xp25_ASAP7_75t_SL g2859 ( 
.A(n_2856),
.B(n_2666),
.C(n_2665),
.D(n_2454),
.Y(n_2859)
);

NAND3xp33_ASAP7_75t_SL g2860 ( 
.A(n_2850),
.B(n_2382),
.C(n_2460),
.Y(n_2860)
);

NAND2xp5_ASAP7_75t_SL g2861 ( 
.A(n_2843),
.B(n_2475),
.Y(n_2861)
);

INVx1_ASAP7_75t_L g2862 ( 
.A(n_2840),
.Y(n_2862)
);

INVx2_ASAP7_75t_L g2863 ( 
.A(n_2844),
.Y(n_2863)
);

NOR3xp33_ASAP7_75t_L g2864 ( 
.A(n_2838),
.B(n_2482),
.C(n_2462),
.Y(n_2864)
);

NAND3xp33_ASAP7_75t_L g2865 ( 
.A(n_2847),
.B(n_2488),
.C(n_2483),
.Y(n_2865)
);

INVx1_ASAP7_75t_L g2866 ( 
.A(n_2853),
.Y(n_2866)
);

NOR2xp33_ASAP7_75t_L g2867 ( 
.A(n_2851),
.B(n_250),
.Y(n_2867)
);

AOI211xp5_ASAP7_75t_L g2868 ( 
.A1(n_2839),
.A2(n_255),
.B(n_253),
.C(n_254),
.Y(n_2868)
);

INVx1_ASAP7_75t_L g2869 ( 
.A(n_2842),
.Y(n_2869)
);

AOI221xp5_ASAP7_75t_L g2870 ( 
.A1(n_2852),
.A2(n_256),
.B1(n_253),
.B2(n_255),
.C(n_257),
.Y(n_2870)
);

NAND2xp5_ASAP7_75t_L g2871 ( 
.A(n_2846),
.B(n_257),
.Y(n_2871)
);

AOI221xp5_ASAP7_75t_L g2872 ( 
.A1(n_2849),
.A2(n_262),
.B1(n_259),
.B2(n_260),
.C(n_263),
.Y(n_2872)
);

NOR2xp33_ASAP7_75t_L g2873 ( 
.A(n_2837),
.B(n_259),
.Y(n_2873)
);

NAND2xp5_ASAP7_75t_L g2874 ( 
.A(n_2857),
.B(n_2855),
.Y(n_2874)
);

NAND4xp75_ASAP7_75t_L g2875 ( 
.A(n_2848),
.B(n_2854),
.C(n_2841),
.D(n_263),
.Y(n_2875)
);

INVxp33_ASAP7_75t_SL g2876 ( 
.A(n_2850),
.Y(n_2876)
);

NOR2xp33_ASAP7_75t_L g2877 ( 
.A(n_2853),
.B(n_260),
.Y(n_2877)
);

NAND4xp25_ASAP7_75t_L g2878 ( 
.A(n_2847),
.B(n_265),
.C(n_262),
.D(n_264),
.Y(n_2878)
);

INVxp33_ASAP7_75t_L g2879 ( 
.A(n_2843),
.Y(n_2879)
);

OR2x2_ASAP7_75t_L g2880 ( 
.A(n_2846),
.B(n_264),
.Y(n_2880)
);

NAND2xp5_ASAP7_75t_L g2881 ( 
.A(n_2850),
.B(n_266),
.Y(n_2881)
);

NAND2xp5_ASAP7_75t_SL g2882 ( 
.A(n_2850),
.B(n_267),
.Y(n_2882)
);

NOR4xp75_ASAP7_75t_L g2883 ( 
.A(n_2838),
.B(n_269),
.C(n_267),
.D(n_268),
.Y(n_2883)
);

O2A1O1Ixp33_ASAP7_75t_L g2884 ( 
.A1(n_2838),
.A2(n_271),
.B(n_268),
.C(n_270),
.Y(n_2884)
);

O2A1O1Ixp33_ASAP7_75t_L g2885 ( 
.A1(n_2838),
.A2(n_273),
.B(n_271),
.C(n_272),
.Y(n_2885)
);

OAI211xp5_ASAP7_75t_SL g2886 ( 
.A1(n_2838),
.A2(n_276),
.B(n_274),
.C(n_275),
.Y(n_2886)
);

AOI22xp5_ASAP7_75t_L g2887 ( 
.A1(n_2852),
.A2(n_276),
.B1(n_274),
.B2(n_275),
.Y(n_2887)
);

AOI221xp5_ASAP7_75t_L g2888 ( 
.A1(n_2845),
.A2(n_279),
.B1(n_277),
.B2(n_278),
.C(n_280),
.Y(n_2888)
);

NAND5xp2_ASAP7_75t_L g2889 ( 
.A(n_2847),
.B(n_280),
.C(n_278),
.D(n_281),
.E(n_277),
.Y(n_2889)
);

NAND4xp75_ASAP7_75t_L g2890 ( 
.A(n_2842),
.B(n_341),
.C(n_338),
.D(n_339),
.Y(n_2890)
);

AOI211xp5_ASAP7_75t_L g2891 ( 
.A1(n_2847),
.A2(n_346),
.B(n_342),
.C(n_343),
.Y(n_2891)
);

INVx1_ASAP7_75t_L g2892 ( 
.A(n_2850),
.Y(n_2892)
);

NOR3xp33_ASAP7_75t_L g2893 ( 
.A(n_2850),
.B(n_347),
.C(n_348),
.Y(n_2893)
);

AND4x1_ASAP7_75t_L g2894 ( 
.A(n_2838),
.B(n_353),
.C(n_349),
.D(n_350),
.Y(n_2894)
);

NAND2xp5_ASAP7_75t_L g2895 ( 
.A(n_2876),
.B(n_354),
.Y(n_2895)
);

INVx2_ASAP7_75t_SL g2896 ( 
.A(n_2880),
.Y(n_2896)
);

INVx1_ASAP7_75t_L g2897 ( 
.A(n_2881),
.Y(n_2897)
);

HB1xp67_ASAP7_75t_L g2898 ( 
.A(n_2883),
.Y(n_2898)
);

INVx8_ASAP7_75t_L g2899 ( 
.A(n_2892),
.Y(n_2899)
);

NAND2xp5_ASAP7_75t_L g2900 ( 
.A(n_2862),
.B(n_355),
.Y(n_2900)
);

AOI21xp5_ASAP7_75t_L g2901 ( 
.A1(n_2874),
.A2(n_360),
.B(n_361),
.Y(n_2901)
);

AND2x2_ASAP7_75t_L g2902 ( 
.A(n_2863),
.B(n_362),
.Y(n_2902)
);

AND2x2_ASAP7_75t_L g2903 ( 
.A(n_2869),
.B(n_363),
.Y(n_2903)
);

AND2x2_ASAP7_75t_L g2904 ( 
.A(n_2879),
.B(n_364),
.Y(n_2904)
);

AOI21xp33_ASAP7_75t_L g2905 ( 
.A1(n_2877),
.A2(n_2873),
.B(n_2882),
.Y(n_2905)
);

NOR2x1_ASAP7_75t_L g2906 ( 
.A(n_2875),
.B(n_365),
.Y(n_2906)
);

AND3x4_ASAP7_75t_L g2907 ( 
.A(n_2864),
.B(n_367),
.C(n_370),
.Y(n_2907)
);

INVxp67_ASAP7_75t_SL g2908 ( 
.A(n_2871),
.Y(n_2908)
);

NAND2xp5_ASAP7_75t_L g2909 ( 
.A(n_2868),
.B(n_371),
.Y(n_2909)
);

INVx1_ASAP7_75t_L g2910 ( 
.A(n_2889),
.Y(n_2910)
);

INVx1_ASAP7_75t_L g2911 ( 
.A(n_2878),
.Y(n_2911)
);

INVx1_ASAP7_75t_L g2912 ( 
.A(n_2866),
.Y(n_2912)
);

OAI22xp5_ASAP7_75t_L g2913 ( 
.A1(n_2887),
.A2(n_375),
.B1(n_372),
.B2(n_373),
.Y(n_2913)
);

NAND2xp5_ASAP7_75t_L g2914 ( 
.A(n_2890),
.B(n_377),
.Y(n_2914)
);

AOI22xp5_ASAP7_75t_L g2915 ( 
.A1(n_2867),
.A2(n_380),
.B1(n_378),
.B2(n_379),
.Y(n_2915)
);

INVxp67_ASAP7_75t_SL g2916 ( 
.A(n_2884),
.Y(n_2916)
);

NOR2x1p5_ASAP7_75t_L g2917 ( 
.A(n_2860),
.B(n_382),
.Y(n_2917)
);

AOI22xp33_ASAP7_75t_SL g2918 ( 
.A1(n_2865),
.A2(n_2894),
.B1(n_2859),
.B2(n_2886),
.Y(n_2918)
);

NAND2xp5_ASAP7_75t_L g2919 ( 
.A(n_2872),
.B(n_2888),
.Y(n_2919)
);

INVx1_ASAP7_75t_L g2920 ( 
.A(n_2861),
.Y(n_2920)
);

NAND2xp5_ASAP7_75t_L g2921 ( 
.A(n_2891),
.B(n_383),
.Y(n_2921)
);

OR2x2_ASAP7_75t_L g2922 ( 
.A(n_2893),
.B(n_384),
.Y(n_2922)
);

INVx1_ASAP7_75t_L g2923 ( 
.A(n_2885),
.Y(n_2923)
);

CKINVDCx14_ASAP7_75t_R g2924 ( 
.A(n_2870),
.Y(n_2924)
);

XNOR2x1_ASAP7_75t_L g2925 ( 
.A(n_2858),
.B(n_385),
.Y(n_2925)
);

INVx1_ASAP7_75t_L g2926 ( 
.A(n_2881),
.Y(n_2926)
);

OR2x2_ASAP7_75t_L g2927 ( 
.A(n_2889),
.B(n_387),
.Y(n_2927)
);

NOR2x1_ASAP7_75t_L g2928 ( 
.A(n_2875),
.B(n_388),
.Y(n_2928)
);

NAND2xp5_ASAP7_75t_L g2929 ( 
.A(n_2876),
.B(n_391),
.Y(n_2929)
);

NOR2x1_ASAP7_75t_L g2930 ( 
.A(n_2875),
.B(n_392),
.Y(n_2930)
);

AND2x4_ASAP7_75t_L g2931 ( 
.A(n_2892),
.B(n_393),
.Y(n_2931)
);

INVx1_ASAP7_75t_L g2932 ( 
.A(n_2881),
.Y(n_2932)
);

INVx2_ASAP7_75t_L g2933 ( 
.A(n_2927),
.Y(n_2933)
);

AND2x2_ASAP7_75t_L g2934 ( 
.A(n_2916),
.B(n_2898),
.Y(n_2934)
);

NAND4xp75_ASAP7_75t_L g2935 ( 
.A(n_2906),
.B(n_396),
.C(n_394),
.D(n_395),
.Y(n_2935)
);

INVx1_ASAP7_75t_L g2936 ( 
.A(n_2910),
.Y(n_2936)
);

NAND2xp5_ASAP7_75t_L g2937 ( 
.A(n_2896),
.B(n_398),
.Y(n_2937)
);

NOR3xp33_ASAP7_75t_L g2938 ( 
.A(n_2895),
.B(n_399),
.C(n_401),
.Y(n_2938)
);

NOR2x1_ASAP7_75t_L g2939 ( 
.A(n_2920),
.B(n_402),
.Y(n_2939)
);

NOR3x2_ASAP7_75t_L g2940 ( 
.A(n_2899),
.B(n_2922),
.C(n_2928),
.Y(n_2940)
);

NOR2x1_ASAP7_75t_L g2941 ( 
.A(n_2930),
.B(n_404),
.Y(n_2941)
);

AND4x2_ASAP7_75t_L g2942 ( 
.A(n_2899),
.B(n_418),
.C(n_430),
.D(n_405),
.Y(n_2942)
);

INVx1_ASAP7_75t_L g2943 ( 
.A(n_2912),
.Y(n_2943)
);

AOI22xp5_ASAP7_75t_L g2944 ( 
.A1(n_2908),
.A2(n_409),
.B1(n_406),
.B2(n_408),
.Y(n_2944)
);

NOR3xp33_ASAP7_75t_L g2945 ( 
.A(n_2929),
.B(n_2926),
.C(n_2897),
.Y(n_2945)
);

NAND3xp33_ASAP7_75t_L g2946 ( 
.A(n_2901),
.B(n_411),
.C(n_413),
.Y(n_2946)
);

NAND2xp5_ASAP7_75t_L g2947 ( 
.A(n_2931),
.B(n_414),
.Y(n_2947)
);

NAND2xp5_ASAP7_75t_SL g2948 ( 
.A(n_2918),
.B(n_421),
.Y(n_2948)
);

AND2x2_ASAP7_75t_L g2949 ( 
.A(n_2923),
.B(n_417),
.Y(n_2949)
);

NOR3x2_ASAP7_75t_L g2950 ( 
.A(n_2924),
.B(n_423),
.C(n_424),
.Y(n_2950)
);

NOR2xp33_ASAP7_75t_L g2951 ( 
.A(n_2932),
.B(n_425),
.Y(n_2951)
);

OAI221xp5_ASAP7_75t_L g2952 ( 
.A1(n_2911),
.A2(n_428),
.B1(n_426),
.B2(n_427),
.C(n_434),
.Y(n_2952)
);

NOR2x1_ASAP7_75t_L g2953 ( 
.A(n_2900),
.B(n_437),
.Y(n_2953)
);

NOR3xp33_ASAP7_75t_L g2954 ( 
.A(n_2904),
.B(n_438),
.C(n_440),
.Y(n_2954)
);

NAND4xp75_ASAP7_75t_L g2955 ( 
.A(n_2903),
.B(n_446),
.C(n_442),
.D(n_444),
.Y(n_2955)
);

NAND4xp25_ASAP7_75t_L g2956 ( 
.A(n_2905),
.B(n_460),
.C(n_471),
.D(n_447),
.Y(n_2956)
);

NAND3xp33_ASAP7_75t_L g2957 ( 
.A(n_2915),
.B(n_451),
.C(n_452),
.Y(n_2957)
);

AND2x2_ASAP7_75t_L g2958 ( 
.A(n_2917),
.B(n_2902),
.Y(n_2958)
);

NOR3xp33_ASAP7_75t_L g2959 ( 
.A(n_2914),
.B(n_454),
.C(n_455),
.Y(n_2959)
);

NOR3xp33_ASAP7_75t_L g2960 ( 
.A(n_2909),
.B(n_456),
.C(n_458),
.Y(n_2960)
);

NAND4xp75_ASAP7_75t_L g2961 ( 
.A(n_2919),
.B(n_464),
.C(n_459),
.D(n_462),
.Y(n_2961)
);

NOR2x1_ASAP7_75t_L g2962 ( 
.A(n_2907),
.B(n_465),
.Y(n_2962)
);

NOR2x1_ASAP7_75t_L g2963 ( 
.A(n_2921),
.B(n_2925),
.Y(n_2963)
);

INVx1_ASAP7_75t_L g2964 ( 
.A(n_2913),
.Y(n_2964)
);

INVx1_ASAP7_75t_L g2965 ( 
.A(n_2898),
.Y(n_2965)
);

NAND3x2_ASAP7_75t_L g2966 ( 
.A(n_2920),
.B(n_467),
.C(n_468),
.Y(n_2966)
);

HB1xp67_ASAP7_75t_L g2967 ( 
.A(n_2898),
.Y(n_2967)
);

INVx1_ASAP7_75t_L g2968 ( 
.A(n_2898),
.Y(n_2968)
);

AOI21xp5_ASAP7_75t_L g2969 ( 
.A1(n_2899),
.A2(n_469),
.B(n_470),
.Y(n_2969)
);

NAND4xp75_ASAP7_75t_L g2970 ( 
.A(n_2906),
.B(n_474),
.C(n_472),
.D(n_473),
.Y(n_2970)
);

NAND4xp75_ASAP7_75t_L g2971 ( 
.A(n_2906),
.B(n_477),
.C(n_475),
.D(n_476),
.Y(n_2971)
);

NOR4xp75_ASAP7_75t_L g2972 ( 
.A(n_2919),
.B(n_480),
.C(n_478),
.D(n_479),
.Y(n_2972)
);

INVx1_ASAP7_75t_L g2973 ( 
.A(n_2898),
.Y(n_2973)
);

AOI22xp5_ASAP7_75t_L g2974 ( 
.A1(n_2916),
.A2(n_483),
.B1(n_481),
.B2(n_482),
.Y(n_2974)
);

NOR2x1_ASAP7_75t_L g2975 ( 
.A(n_2920),
.B(n_484),
.Y(n_2975)
);

NAND2xp5_ASAP7_75t_L g2976 ( 
.A(n_2898),
.B(n_485),
.Y(n_2976)
);

INVx1_ASAP7_75t_L g2977 ( 
.A(n_2898),
.Y(n_2977)
);

NOR2xp67_ASAP7_75t_SL g2978 ( 
.A(n_2912),
.B(n_486),
.Y(n_2978)
);

AND2x4_ASAP7_75t_L g2979 ( 
.A(n_2934),
.B(n_487),
.Y(n_2979)
);

XNOR2x1_ASAP7_75t_L g2980 ( 
.A(n_2963),
.B(n_490),
.Y(n_2980)
);

AND2x2_ASAP7_75t_SL g2981 ( 
.A(n_2943),
.B(n_491),
.Y(n_2981)
);

OA21x2_ASAP7_75t_L g2982 ( 
.A1(n_2965),
.A2(n_846),
.B(n_845),
.Y(n_2982)
);

CKINVDCx20_ASAP7_75t_R g2983 ( 
.A(n_2967),
.Y(n_2983)
);

NOR3x1_ASAP7_75t_L g2984 ( 
.A(n_2968),
.B(n_492),
.C(n_493),
.Y(n_2984)
);

AOI21xp33_ASAP7_75t_L g2985 ( 
.A1(n_2933),
.A2(n_494),
.B(n_495),
.Y(n_2985)
);

OR2x2_ASAP7_75t_L g2986 ( 
.A(n_2973),
.B(n_497),
.Y(n_2986)
);

NOR2xp33_ASAP7_75t_L g2987 ( 
.A(n_2977),
.B(n_498),
.Y(n_2987)
);

NAND2xp5_ASAP7_75t_L g2988 ( 
.A(n_2958),
.B(n_499),
.Y(n_2988)
);

INVx1_ASAP7_75t_L g2989 ( 
.A(n_2937),
.Y(n_2989)
);

INVx1_ASAP7_75t_L g2990 ( 
.A(n_2949),
.Y(n_2990)
);

AND4x1_ASAP7_75t_L g2991 ( 
.A(n_2945),
.B(n_502),
.C(n_500),
.D(n_501),
.Y(n_2991)
);

NAND5xp2_ASAP7_75t_L g2992 ( 
.A(n_2936),
.B(n_505),
.C(n_503),
.D(n_504),
.E(n_506),
.Y(n_2992)
);

OAI22x1_ASAP7_75t_L g2993 ( 
.A1(n_2941),
.A2(n_509),
.B1(n_507),
.B2(n_508),
.Y(n_2993)
);

INVx2_ASAP7_75t_L g2994 ( 
.A(n_2935),
.Y(n_2994)
);

CKINVDCx5p33_ASAP7_75t_R g2995 ( 
.A(n_2976),
.Y(n_2995)
);

NAND2x1p5_ASAP7_75t_L g2996 ( 
.A(n_2978),
.B(n_511),
.Y(n_2996)
);

AOI22xp5_ASAP7_75t_SL g2997 ( 
.A1(n_2947),
.A2(n_516),
.B1(n_513),
.B2(n_514),
.Y(n_2997)
);

AND2x4_ASAP7_75t_L g2998 ( 
.A(n_2948),
.B(n_517),
.Y(n_2998)
);

AND2x4_ASAP7_75t_L g2999 ( 
.A(n_2964),
.B(n_520),
.Y(n_2999)
);

NAND3x1_ASAP7_75t_L g3000 ( 
.A(n_2939),
.B(n_521),
.C(n_523),
.Y(n_3000)
);

INVx1_ASAP7_75t_L g3001 ( 
.A(n_2940),
.Y(n_3001)
);

NAND2xp5_ASAP7_75t_L g3002 ( 
.A(n_2959),
.B(n_524),
.Y(n_3002)
);

NOR2xp67_ASAP7_75t_L g3003 ( 
.A(n_2969),
.B(n_525),
.Y(n_3003)
);

INVx2_ASAP7_75t_L g3004 ( 
.A(n_2970),
.Y(n_3004)
);

AND2x4_ASAP7_75t_L g3005 ( 
.A(n_2962),
.B(n_527),
.Y(n_3005)
);

AND2x2_ASAP7_75t_L g3006 ( 
.A(n_2960),
.B(n_530),
.Y(n_3006)
);

NOR2x1p5_ASAP7_75t_L g3007 ( 
.A(n_2971),
.B(n_2946),
.Y(n_3007)
);

NOR3xp33_ASAP7_75t_L g3008 ( 
.A(n_2951),
.B(n_532),
.C(n_533),
.Y(n_3008)
);

NOR4xp75_ASAP7_75t_L g3009 ( 
.A(n_2961),
.B(n_538),
.C(n_534),
.D(n_537),
.Y(n_3009)
);

NAND3x1_ASAP7_75t_L g3010 ( 
.A(n_2975),
.B(n_539),
.C(n_540),
.Y(n_3010)
);

INVx1_ASAP7_75t_L g3011 ( 
.A(n_2953),
.Y(n_3011)
);

NOR4xp75_ASAP7_75t_SL g3012 ( 
.A(n_2966),
.B(n_548),
.C(n_541),
.D(n_543),
.Y(n_3012)
);

AOI21xp5_ASAP7_75t_L g3013 ( 
.A1(n_2957),
.A2(n_550),
.B(n_551),
.Y(n_3013)
);

NAND2x1_ASAP7_75t_L g3014 ( 
.A(n_2974),
.B(n_552),
.Y(n_3014)
);

NAND4xp75_ASAP7_75t_L g3015 ( 
.A(n_2944),
.B(n_557),
.C(n_554),
.D(n_556),
.Y(n_3015)
);

AND2x2_ASAP7_75t_SL g3016 ( 
.A(n_2938),
.B(n_558),
.Y(n_3016)
);

OAI22xp33_ASAP7_75t_L g3017 ( 
.A1(n_2983),
.A2(n_2956),
.B1(n_2952),
.B2(n_2950),
.Y(n_3017)
);

HB1xp67_ASAP7_75t_L g3018 ( 
.A(n_2982),
.Y(n_3018)
);

NAND2xp5_ASAP7_75t_SL g3019 ( 
.A(n_3012),
.B(n_2954),
.Y(n_3019)
);

AND3x1_ASAP7_75t_L g3020 ( 
.A(n_3001),
.B(n_3004),
.C(n_2994),
.Y(n_3020)
);

AOI21xp5_ASAP7_75t_L g3021 ( 
.A1(n_2988),
.A2(n_2942),
.B(n_2972),
.Y(n_3021)
);

NAND3xp33_ASAP7_75t_L g3022 ( 
.A(n_3011),
.B(n_2955),
.C(n_559),
.Y(n_3022)
);

NAND2xp5_ASAP7_75t_L g3023 ( 
.A(n_3005),
.B(n_2979),
.Y(n_3023)
);

CKINVDCx5p33_ASAP7_75t_R g3024 ( 
.A(n_2995),
.Y(n_3024)
);

XOR2xp5_ASAP7_75t_L g3025 ( 
.A(n_2980),
.B(n_560),
.Y(n_3025)
);

INVx1_ASAP7_75t_L g3026 ( 
.A(n_2981),
.Y(n_3026)
);

AOI22xp5_ASAP7_75t_L g3027 ( 
.A1(n_3003),
.A2(n_565),
.B1(n_563),
.B2(n_564),
.Y(n_3027)
);

NAND2xp5_ASAP7_75t_L g3028 ( 
.A(n_2987),
.B(n_566),
.Y(n_3028)
);

OAI222xp33_ASAP7_75t_L g3029 ( 
.A1(n_3014),
.A2(n_569),
.B1(n_573),
.B2(n_567),
.C1(n_568),
.C2(n_571),
.Y(n_3029)
);

OA22x2_ASAP7_75t_L g3030 ( 
.A1(n_2993),
.A2(n_577),
.B1(n_575),
.B2(n_576),
.Y(n_3030)
);

NAND3xp33_ASAP7_75t_L g3031 ( 
.A(n_2991),
.B(n_578),
.C(n_579),
.Y(n_3031)
);

OR2x2_ASAP7_75t_L g3032 ( 
.A(n_2986),
.B(n_583),
.Y(n_3032)
);

OAI22xp5_ASAP7_75t_L g3033 ( 
.A1(n_3007),
.A2(n_853),
.B1(n_591),
.B2(n_584),
.Y(n_3033)
);

OAI22xp5_ASAP7_75t_SL g3034 ( 
.A1(n_2996),
.A2(n_594),
.B1(n_585),
.B2(n_592),
.Y(n_3034)
);

INVx1_ASAP7_75t_L g3035 ( 
.A(n_2990),
.Y(n_3035)
);

NAND2xp5_ASAP7_75t_L g3036 ( 
.A(n_2984),
.B(n_595),
.Y(n_3036)
);

INVx1_ASAP7_75t_L g3037 ( 
.A(n_3000),
.Y(n_3037)
);

INVx2_ASAP7_75t_L g3038 ( 
.A(n_3010),
.Y(n_3038)
);

NOR2xp33_ASAP7_75t_L g3039 ( 
.A(n_2989),
.B(n_3002),
.Y(n_3039)
);

INVx1_ASAP7_75t_L g3040 ( 
.A(n_2999),
.Y(n_3040)
);

BUFx3_ASAP7_75t_L g3041 ( 
.A(n_2998),
.Y(n_3041)
);

NOR3xp33_ASAP7_75t_L g3042 ( 
.A(n_2985),
.B(n_3008),
.C(n_2992),
.Y(n_3042)
);

A2O1A1Ixp33_ASAP7_75t_SL g3043 ( 
.A1(n_3013),
.A2(n_598),
.B(n_596),
.C(n_597),
.Y(n_3043)
);

NAND2xp33_ASAP7_75t_R g3044 ( 
.A(n_3006),
.B(n_599),
.Y(n_3044)
);

INVx2_ASAP7_75t_L g3045 ( 
.A(n_3015),
.Y(n_3045)
);

INVx1_ASAP7_75t_L g3046 ( 
.A(n_3018),
.Y(n_3046)
);

OAI22xp33_ASAP7_75t_L g3047 ( 
.A1(n_3024),
.A2(n_3009),
.B1(n_3016),
.B2(n_2997),
.Y(n_3047)
);

NAND2xp5_ASAP7_75t_L g3048 ( 
.A(n_3026),
.B(n_3021),
.Y(n_3048)
);

AOI211x1_ASAP7_75t_L g3049 ( 
.A1(n_3017),
.A2(n_602),
.B(n_600),
.C(n_601),
.Y(n_3049)
);

OAI21xp33_ASAP7_75t_SL g3050 ( 
.A1(n_3019),
.A2(n_604),
.B(n_605),
.Y(n_3050)
);

INVx1_ASAP7_75t_L g3051 ( 
.A(n_3041),
.Y(n_3051)
);

NAND2xp5_ASAP7_75t_L g3052 ( 
.A(n_3025),
.B(n_3037),
.Y(n_3052)
);

AO22x2_ASAP7_75t_L g3053 ( 
.A1(n_3038),
.A2(n_610),
.B1(n_607),
.B2(n_608),
.Y(n_3053)
);

AOI22xp5_ASAP7_75t_L g3054 ( 
.A1(n_3020),
.A2(n_616),
.B1(n_613),
.B2(n_614),
.Y(n_3054)
);

AOI21xp33_ASAP7_75t_L g3055 ( 
.A1(n_3039),
.A2(n_851),
.B(n_618),
.Y(n_3055)
);

AND2x2_ASAP7_75t_L g3056 ( 
.A(n_3035),
.B(n_619),
.Y(n_3056)
);

INVx1_ASAP7_75t_L g3057 ( 
.A(n_3032),
.Y(n_3057)
);

BUFx2_ASAP7_75t_L g3058 ( 
.A(n_3030),
.Y(n_3058)
);

XOR2xp5_ASAP7_75t_L g3059 ( 
.A(n_3023),
.B(n_620),
.Y(n_3059)
);

INVx1_ASAP7_75t_L g3060 ( 
.A(n_3036),
.Y(n_3060)
);

INVxp33_ASAP7_75t_L g3061 ( 
.A(n_3034),
.Y(n_3061)
);

INVx2_ASAP7_75t_L g3062 ( 
.A(n_3040),
.Y(n_3062)
);

XNOR2xp5_ASAP7_75t_L g3063 ( 
.A(n_3042),
.B(n_621),
.Y(n_3063)
);

OAI22xp5_ASAP7_75t_L g3064 ( 
.A1(n_3022),
.A2(n_628),
.B1(n_623),
.B2(n_625),
.Y(n_3064)
);

INVx2_ASAP7_75t_L g3065 ( 
.A(n_3028),
.Y(n_3065)
);

NAND2xp5_ASAP7_75t_L g3066 ( 
.A(n_3027),
.B(n_629),
.Y(n_3066)
);

AND4x1_ASAP7_75t_L g3067 ( 
.A(n_3031),
.B(n_633),
.C(n_631),
.D(n_632),
.Y(n_3067)
);

NOR2xp33_ASAP7_75t_L g3068 ( 
.A(n_3046),
.B(n_3045),
.Y(n_3068)
);

AOI22xp33_ASAP7_75t_SL g3069 ( 
.A1(n_3058),
.A2(n_3033),
.B1(n_3044),
.B2(n_3043),
.Y(n_3069)
);

OAI22xp5_ASAP7_75t_L g3070 ( 
.A1(n_3048),
.A2(n_3029),
.B1(n_640),
.B2(n_635),
.Y(n_3070)
);

AOI22xp5_ASAP7_75t_L g3071 ( 
.A1(n_3052),
.A2(n_642),
.B1(n_636),
.B2(n_641),
.Y(n_3071)
);

NAND4xp75_ASAP7_75t_L g3072 ( 
.A(n_3051),
.B(n_645),
.C(n_643),
.D(n_644),
.Y(n_3072)
);

OAI22xp33_ASAP7_75t_L g3073 ( 
.A1(n_3061),
.A2(n_648),
.B1(n_646),
.B2(n_647),
.Y(n_3073)
);

NOR4xp75_ASAP7_75t_L g3074 ( 
.A(n_3064),
.B(n_652),
.C(n_649),
.D(n_650),
.Y(n_3074)
);

INVx1_ASAP7_75t_L g3075 ( 
.A(n_3057),
.Y(n_3075)
);

INVx1_ASAP7_75t_L g3076 ( 
.A(n_3065),
.Y(n_3076)
);

OR2x2_ASAP7_75t_L g3077 ( 
.A(n_3062),
.B(n_653),
.Y(n_3077)
);

NOR3xp33_ASAP7_75t_SL g3078 ( 
.A(n_3047),
.B(n_654),
.C(n_655),
.Y(n_3078)
);

OAI222xp33_ASAP7_75t_L g3079 ( 
.A1(n_3075),
.A2(n_3060),
.B1(n_3063),
.B2(n_3054),
.C1(n_3066),
.C2(n_3059),
.Y(n_3079)
);

NAND4xp25_ASAP7_75t_L g3080 ( 
.A(n_3068),
.B(n_3049),
.C(n_3056),
.D(n_3055),
.Y(n_3080)
);

AOI221x1_ASAP7_75t_L g3081 ( 
.A1(n_3076),
.A2(n_3070),
.B1(n_3053),
.B2(n_3069),
.C(n_3050),
.Y(n_3081)
);

NAND4xp75_ASAP7_75t_L g3082 ( 
.A(n_3078),
.B(n_3067),
.C(n_3053),
.D(n_660),
.Y(n_3082)
);

NOR4xp25_ASAP7_75t_SL g3083 ( 
.A(n_3074),
.B(n_662),
.C(n_658),
.D(n_659),
.Y(n_3083)
);

NAND3xp33_ASAP7_75t_SL g3084 ( 
.A(n_3077),
.B(n_663),
.C(n_664),
.Y(n_3084)
);

OA22x2_ASAP7_75t_L g3085 ( 
.A1(n_3071),
.A2(n_669),
.B1(n_665),
.B2(n_667),
.Y(n_3085)
);

INVx1_ASAP7_75t_L g3086 ( 
.A(n_3072),
.Y(n_3086)
);

NAND3xp33_ASAP7_75t_SL g3087 ( 
.A(n_3073),
.B(n_670),
.C(n_671),
.Y(n_3087)
);

INVxp67_ASAP7_75t_SL g3088 ( 
.A(n_3086),
.Y(n_3088)
);

OAI22xp5_ASAP7_75t_L g3089 ( 
.A1(n_3082),
.A2(n_674),
.B1(n_672),
.B2(n_673),
.Y(n_3089)
);

AO22x2_ASAP7_75t_SL g3090 ( 
.A1(n_3081),
.A2(n_678),
.B1(n_676),
.B2(n_677),
.Y(n_3090)
);

INVxp67_ASAP7_75t_SL g3091 ( 
.A(n_3080),
.Y(n_3091)
);

INVx1_ASAP7_75t_L g3092 ( 
.A(n_3084),
.Y(n_3092)
);

OAI21x1_ASAP7_75t_L g3093 ( 
.A1(n_3079),
.A2(n_679),
.B(n_682),
.Y(n_3093)
);

INVx1_ASAP7_75t_L g3094 ( 
.A(n_3085),
.Y(n_3094)
);

AOI322xp5_ASAP7_75t_L g3095 ( 
.A1(n_3088),
.A2(n_3087),
.A3(n_3083),
.B1(n_689),
.B2(n_686),
.C1(n_688),
.C2(n_683),
.Y(n_3095)
);

INVx1_ASAP7_75t_L g3096 ( 
.A(n_3091),
.Y(n_3096)
);

INVx1_ASAP7_75t_L g3097 ( 
.A(n_3090),
.Y(n_3097)
);

INVx2_ASAP7_75t_SL g3098 ( 
.A(n_3094),
.Y(n_3098)
);

INVx1_ASAP7_75t_L g3099 ( 
.A(n_3092),
.Y(n_3099)
);

OR2x2_ASAP7_75t_L g3100 ( 
.A(n_3093),
.B(n_3089),
.Y(n_3100)
);

OR2x6_ASAP7_75t_L g3101 ( 
.A(n_3092),
.B(n_684),
.Y(n_3101)
);

HB1xp67_ASAP7_75t_L g3102 ( 
.A(n_3096),
.Y(n_3102)
);

OAI22xp5_ASAP7_75t_SL g3103 ( 
.A1(n_3097),
.A2(n_691),
.B1(n_687),
.B2(n_690),
.Y(n_3103)
);

OAI22x1_ASAP7_75t_L g3104 ( 
.A1(n_3098),
.A2(n_850),
.B1(n_695),
.B2(n_693),
.Y(n_3104)
);

OAI22x1_ASAP7_75t_L g3105 ( 
.A1(n_3099),
.A2(n_697),
.B1(n_694),
.B2(n_696),
.Y(n_3105)
);

AOI21xp5_ASAP7_75t_L g3106 ( 
.A1(n_3100),
.A2(n_698),
.B(n_700),
.Y(n_3106)
);

INVxp33_ASAP7_75t_L g3107 ( 
.A(n_3102),
.Y(n_3107)
);

OAI221xp5_ASAP7_75t_L g3108 ( 
.A1(n_3106),
.A2(n_3095),
.B1(n_3101),
.B2(n_703),
.C(n_701),
.Y(n_3108)
);

CKINVDCx20_ASAP7_75t_R g3109 ( 
.A(n_3107),
.Y(n_3109)
);

INVx3_ASAP7_75t_L g3110 ( 
.A(n_3109),
.Y(n_3110)
);

NOR2xp33_ASAP7_75t_L g3111 ( 
.A(n_3110),
.B(n_3108),
.Y(n_3111)
);

AOI21xp5_ASAP7_75t_L g3112 ( 
.A1(n_3111),
.A2(n_3101),
.B(n_3104),
.Y(n_3112)
);

AOI211xp5_ASAP7_75t_L g3113 ( 
.A1(n_3112),
.A2(n_3103),
.B(n_3105),
.C(n_704),
.Y(n_3113)
);


endmodule