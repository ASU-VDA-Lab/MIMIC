module fake_jpeg_30008_n_120 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_120);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_120;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_5),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_24),
.Y(n_25)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g27 ( 
.A(n_15),
.B(n_0),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_27),
.B(n_30),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_13),
.B(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_15),
.B(n_1),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_16),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_16),
.B(n_1),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_34),
.B(n_36),
.Y(n_47)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx3_ASAP7_75t_SL g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx2_ASAP7_75t_SL g51 ( 
.A(n_37),
.Y(n_51)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_39),
.B(n_47),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_29),
.A2(n_19),
.B1(n_14),
.B2(n_12),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_46),
.A2(n_50),
.B1(n_23),
.B2(n_13),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_27),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_17),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_37),
.A2(n_18),
.B1(n_19),
.B2(n_14),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_51),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_61),
.Y(n_71)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_57),
.B(n_68),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_41),
.A2(n_25),
.B1(n_32),
.B2(n_26),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_58),
.A2(n_64),
.B1(n_70),
.B2(n_53),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_52),
.A2(n_38),
.B1(n_35),
.B2(n_19),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_12),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_45),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

AND2x2_ASAP7_75t_SL g62 ( 
.A(n_44),
.B(n_1),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_66),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_40),
.A2(n_22),
.B1(n_23),
.B2(n_17),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_65),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_43),
.B(n_2),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_67),
.Y(n_81)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_42),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_48),
.A2(n_2),
.B1(n_3),
.B2(n_6),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_80),
.Y(n_88)
);

O2A1O1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_61),
.A2(n_54),
.B(n_48),
.C(n_42),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_77),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_78),
.B(n_62),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_76),
.B(n_60),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_83),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_62),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_84),
.B(n_89),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_81),
.A2(n_70),
.B1(n_66),
.B2(n_53),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_85),
.A2(n_72),
.B1(n_66),
.B2(n_76),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_56),
.C(n_55),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_86),
.B(n_79),
.Y(n_96)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_82),
.B(n_78),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_90),
.B(n_92),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_86),
.B(n_75),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_88),
.B(n_71),
.Y(n_94)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_94),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_95),
.B(n_96),
.C(n_88),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_91),
.A2(n_72),
.B(n_88),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_99),
.A2(n_100),
.B(n_63),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g100 ( 
.A(n_96),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_93),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_101),
.A2(n_52),
.B1(n_41),
.B2(n_63),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_102),
.B(n_69),
.C(n_65),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_98),
.A2(n_95),
.B1(n_87),
.B2(n_74),
.Y(n_103)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_103),
.Y(n_108)
);

FAx1_ASAP7_75t_L g104 ( 
.A(n_97),
.B(n_77),
.CI(n_74),
.CON(n_104),
.SN(n_104)
);

XNOR2xp5_ASAP7_75t_SL g109 ( 
.A(n_104),
.B(n_100),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_105),
.B(n_107),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_106),
.B(n_2),
.Y(n_111)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_109),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_111),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_112),
.B(n_114),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_110),
.B(n_104),
.C(n_11),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_113),
.B(n_108),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_116),
.B(n_104),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_117),
.A2(n_109),
.B(n_115),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_3),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_3),
.Y(n_120)
);


endmodule