module fake_jpeg_84_n_216 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_216);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_216;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_38),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_20),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_15),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_52),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_11),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_13),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_49),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_0),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_30),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_28),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_31),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_12),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_15),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_7),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_35),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_79),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_54),
.B(n_0),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_80),
.B(n_81),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_77),
.B(n_1),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_83),
.Y(n_91)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_84),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_63),
.B(n_1),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_59),
.Y(n_92)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_86),
.B(n_57),
.Y(n_93)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_87),
.A2(n_65),
.B1(n_73),
.B2(n_57),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_82),
.B(n_55),
.C(n_76),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_88),
.B(n_93),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_85),
.B(n_55),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_97),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_92),
.B(n_81),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_94),
.A2(n_99),
.B1(n_87),
.B2(n_83),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_79),
.A2(n_76),
.B1(n_75),
.B2(n_65),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_96),
.A2(n_101),
.B1(n_87),
.B2(n_73),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_64),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_84),
.A2(n_75),
.B1(n_62),
.B2(n_71),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_79),
.A2(n_58),
.B1(n_60),
.B2(n_62),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_102),
.B(n_103),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_97),
.B(n_74),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_L g104 ( 
.A1(n_100),
.A2(n_101),
.B1(n_84),
.B2(n_86),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_104),
.A2(n_110),
.B1(n_91),
.B2(n_21),
.Y(n_122)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_100),
.Y(n_105)
);

HB1xp67_ASAP7_75t_L g132 ( 
.A(n_105),
.Y(n_132)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_100),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_98),
.B(n_74),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_107),
.B(n_116),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_108),
.Y(n_128)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_109),
.Y(n_133)
);

A2O1A1Ixp33_ASAP7_75t_L g111 ( 
.A1(n_90),
.A2(n_71),
.B(n_72),
.C(n_53),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_111),
.B(n_113),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_88),
.B(n_78),
.Y(n_113)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_89),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_115),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_68),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_95),
.Y(n_117)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_117),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_93),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_118),
.B(n_91),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_93),
.A2(n_69),
.B1(n_67),
.B2(n_60),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_119),
.Y(n_138)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_95),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_120),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_92),
.A2(n_66),
.B(n_61),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_121),
.B(n_111),
.Y(n_137)
);

INVxp33_ASAP7_75t_L g165 ( 
.A(n_122),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_121),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_124),
.B(n_126),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_125),
.B(n_131),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_115),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_113),
.B(n_2),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_127),
.B(n_129),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_112),
.B(n_2),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_112),
.B(n_114),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_114),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_134),
.A2(n_139),
.B1(n_14),
.B2(n_16),
.Y(n_155)
);

OR2x6_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_40),
.Y(n_136)
);

AO22x1_ASAP7_75t_L g167 ( 
.A1(n_136),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_137),
.B(n_14),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_104),
.A2(n_106),
.B1(n_105),
.B2(n_120),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_113),
.B(n_3),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_140),
.B(n_144),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_113),
.B(n_4),
.Y(n_144)
);

BUFx2_ASAP7_75t_L g145 ( 
.A(n_132),
.Y(n_145)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_145),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_141),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_146),
.B(n_150),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_130),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_147),
.A2(n_151),
.B1(n_155),
.B2(n_158),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_130),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_148),
.B(n_163),
.Y(n_173)
);

OAI32xp33_ASAP7_75t_L g149 ( 
.A1(n_137),
.A2(n_8),
.A3(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_149)
);

XOR2x2_ASAP7_75t_L g183 ( 
.A(n_149),
.B(n_17),
.Y(n_183)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_143),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_136),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_151)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_133),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_153),
.B(n_154),
.Y(n_178)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_141),
.Y(n_154)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_123),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_156),
.B(n_160),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_139),
.A2(n_34),
.B1(n_51),
.B2(n_48),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_123),
.Y(n_160)
);

NOR2x1_ASAP7_75t_SL g161 ( 
.A(n_136),
.B(n_32),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_161),
.B(n_162),
.Y(n_182)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_136),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_138),
.Y(n_163)
);

AO21x1_ASAP7_75t_L g170 ( 
.A1(n_164),
.A2(n_167),
.B(n_134),
.Y(n_170)
);

BUFx2_ASAP7_75t_L g166 ( 
.A(n_138),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_166),
.Y(n_181)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_136),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_169),
.A2(n_165),
.B1(n_167),
.B2(n_159),
.Y(n_186)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_170),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_168),
.B(n_135),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_171),
.B(n_172),
.C(n_176),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_152),
.B(n_128),
.C(n_142),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_164),
.B(n_128),
.C(n_37),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_166),
.A2(n_36),
.B(n_46),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_177),
.A2(n_183),
.B(n_184),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_162),
.A2(n_18),
.B(n_19),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_145),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_185),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_186),
.A2(n_24),
.B1(n_29),
.B2(n_42),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_172),
.A2(n_165),
.B1(n_155),
.B2(n_158),
.Y(n_187)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_187),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_171),
.B(n_174),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_189),
.B(n_176),
.Y(n_203)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_178),
.Y(n_192)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_192),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_173),
.A2(n_157),
.B1(n_19),
.B2(n_25),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_194),
.A2(n_196),
.B1(n_180),
.B2(n_183),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_179),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_195),
.B(n_173),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_197),
.B(n_199),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_193),
.A2(n_177),
.B(n_184),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_191),
.A2(n_182),
.B(n_170),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_200),
.A2(n_201),
.B1(n_202),
.B2(n_190),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_203),
.B(n_189),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_205),
.B(n_206),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_198),
.B(n_188),
.C(n_187),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_207),
.A2(n_194),
.B1(n_181),
.B2(n_175),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_209),
.B(n_204),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_210),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_211),
.B(n_206),
.Y(n_212)
);

NAND2xp33_ASAP7_75t_R g213 ( 
.A(n_212),
.B(n_208),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_213),
.A2(n_205),
.B(n_188),
.Y(n_214)
);

OAI21x1_ASAP7_75t_L g215 ( 
.A1(n_214),
.A2(n_209),
.B(n_44),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_215),
.B(n_43),
.Y(n_216)
);


endmodule