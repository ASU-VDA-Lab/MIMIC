module fake_jpeg_3157_n_73 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_73);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_73;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_51;
wire n_47;
wire n_40;
wire n_59;
wire n_71;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_31;
wire n_25;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;
wire n_70;
wire n_66;

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_20),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_16),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_26),
.Y(n_28)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_27),
.B(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_30),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_27),
.B(n_1),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_21),
.B(n_19),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_31),
.B(n_23),
.Y(n_34)
);

HB1xp67_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_31),
.B(n_24),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_1),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_34),
.B(n_25),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_31),
.A2(n_23),
.B1(n_25),
.B2(n_24),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_37),
.A2(n_22),
.B1(n_26),
.B2(n_3),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_22),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_40),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g41 ( 
.A1(n_38),
.A2(n_28),
.B(n_22),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_41),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_44),
.Y(n_46)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_45),
.B(n_3),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_35),
.C(n_36),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_48),
.B(n_4),
.C(n_9),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_2),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_51),
.B(n_52),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_SL g53 ( 
.A(n_50),
.B(n_41),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_54),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_SL g54 ( 
.A(n_52),
.B(n_46),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_49),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_55),
.B(n_59),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_47),
.A2(n_22),
.B1(n_5),
.B2(n_6),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_56),
.A2(n_58),
.B1(n_13),
.B2(n_14),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_47),
.A2(n_22),
.B1(n_5),
.B2(n_4),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_57),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_61)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_62),
.B(n_63),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_15),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g65 ( 
.A(n_64),
.B(n_17),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_65),
.B(n_60),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_68),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_65),
.A2(n_64),
.B(n_61),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_70),
.A2(n_69),
.B(n_67),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_71),
.B(n_66),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_72),
.B(n_18),
.Y(n_73)
);


endmodule