module fake_jpeg_1565_n_190 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_190);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_190;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_15),
.Y(n_46)
);

BUFx6f_ASAP7_75t_SL g47 ( 
.A(n_31),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_16),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_11),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_0),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_9),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_9),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_69),
.Y(n_74)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_46),
.B(n_1),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_71),
.B(n_48),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_1),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_72),
.B(n_2),
.Y(n_75)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_62),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_76),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_68),
.A2(n_62),
.B1(n_51),
.B2(n_60),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_77),
.A2(n_47),
.B1(n_58),
.B2(n_63),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g81 ( 
.A(n_71),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_83),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_65),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_49),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_84),
.B(n_85),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_70),
.B(n_50),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_82),
.A2(n_73),
.B1(n_67),
.B2(n_60),
.Y(n_87)
);

AO21x2_ASAP7_75t_L g119 ( 
.A1(n_87),
.A2(n_55),
.B(n_59),
.Y(n_119)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_89),
.Y(n_112)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

CKINVDCx14_ASAP7_75t_R g105 ( 
.A(n_90),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_100),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_80),
.A2(n_53),
.B1(n_70),
.B2(n_64),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g107 ( 
.A(n_93),
.Y(n_107)
);

XNOR2x1_ASAP7_75t_SL g94 ( 
.A(n_84),
.B(n_56),
.Y(n_94)
);

NOR2x1_ASAP7_75t_L g122 ( 
.A(n_94),
.B(n_4),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_96),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_78),
.Y(n_97)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_97),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_98),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_74),
.A2(n_86),
.B1(n_58),
.B2(n_53),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_74),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_101),
.B(n_102),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_76),
.Y(n_103)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_103),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_99),
.B(n_64),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_104),
.B(n_115),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_99),
.A2(n_53),
.B(n_54),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_110),
.B(n_119),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_88),
.B(n_2),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_113),
.B(n_114),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_92),
.B(n_3),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_102),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_87),
.B(n_64),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_116),
.B(n_117),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_101),
.B(n_55),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_119),
.A2(n_98),
.B1(n_97),
.B2(n_96),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_103),
.B(n_3),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_120),
.B(n_5),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_122),
.B(n_4),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_106),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_123),
.B(n_124),
.Y(n_146)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_112),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_126),
.A2(n_141),
.B1(n_119),
.B2(n_109),
.Y(n_148)
);

MAJx2_ASAP7_75t_L g127 ( 
.A(n_111),
.B(n_94),
.C(n_95),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_127),
.B(n_129),
.C(n_140),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_128),
.B(n_132),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_104),
.B(n_90),
.C(n_89),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_122),
.B(n_5),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_130),
.B(n_133),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_105),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_112),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_135),
.B(n_142),
.Y(n_149)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_108),
.Y(n_136)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_136),
.Y(n_144)
);

INVx1_ASAP7_75t_SL g137 ( 
.A(n_121),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_137),
.B(n_118),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_138),
.Y(n_145)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_117),
.Y(n_139)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_139),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_21),
.C(n_43),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_116),
.A2(n_20),
.B1(n_42),
.B2(n_39),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_6),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_131),
.A2(n_119),
.B1(n_109),
.B2(n_107),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_147),
.A2(n_134),
.B1(n_10),
.B2(n_11),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_148),
.A2(n_23),
.B1(n_35),
.B2(n_34),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_123),
.A2(n_118),
.B(n_19),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_151),
.B(n_12),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_152),
.B(n_155),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_127),
.B(n_18),
.C(n_38),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_153),
.B(n_157),
.C(n_13),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g155 ( 
.A(n_125),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_138),
.A2(n_126),
.B(n_129),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_156),
.A2(n_33),
.B(n_32),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_141),
.B(n_44),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_137),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_158),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_167)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_140),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_160),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_161),
.B(n_168),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_162),
.A2(n_167),
.B1(n_158),
.B2(n_150),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_163),
.B(n_157),
.Y(n_171)
);

OAI322xp33_ASAP7_75t_L g165 ( 
.A1(n_146),
.A2(n_29),
.A3(n_28),
.B1(n_27),
.B2(n_14),
.C1(n_15),
.C2(n_8),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_165),
.B(n_170),
.C(n_153),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_149),
.Y(n_168)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_169),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_171),
.B(n_172),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_166),
.B(n_143),
.C(n_145),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_174),
.A2(n_177),
.B1(n_156),
.B2(n_147),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g175 ( 
.A(n_163),
.B(n_143),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_175),
.A2(n_145),
.B1(n_166),
.B2(n_154),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_179),
.A2(n_181),
.B1(n_175),
.B2(n_178),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_173),
.A2(n_164),
.B(n_162),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_180),
.A2(n_159),
.B(n_176),
.Y(n_183)
);

OAI21xp33_ASAP7_75t_L g184 ( 
.A1(n_182),
.A2(n_183),
.B(n_179),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_184),
.B(n_144),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_185),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_186),
.B(n_170),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_187),
.B(n_16),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_188),
.B(n_17),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_189),
.B(n_17),
.Y(n_190)
);


endmodule