module real_jpeg_17926_n_8 (n_5, n_4, n_0, n_1, n_2, n_6, n_7, n_3, n_8);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_8;

wire n_17;
wire n_43;
wire n_37;
wire n_21;
wire n_33;
wire n_35;
wire n_50;
wire n_38;
wire n_29;
wire n_49;
wire n_10;
wire n_31;
wire n_9;
wire n_52;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_44;
wire n_46;
wire n_23;
wire n_51;
wire n_11;
wire n_14;
wire n_47;
wire n_45;
wire n_25;
wire n_42;
wire n_22;
wire n_18;
wire n_40;
wire n_36;
wire n_39;
wire n_41;
wire n_27;
wire n_32;
wire n_20;
wire n_19;
wire n_26;
wire n_48;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

OAI221xp5_ASAP7_75t_L g8 ( 
.A1(n_0),
.A2(n_9),
.B1(n_32),
.B2(n_33),
.C(n_34),
.Y(n_8)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

AOI222xp33_ASAP7_75t_SL g34 ( 
.A1(n_0),
.A2(n_35),
.B1(n_40),
.B2(n_46),
.C1(n_50),
.C2(n_51),
.Y(n_34)
);

INVx2_ASAP7_75t_SL g39 ( 
.A(n_0),
.Y(n_39)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_1),
.B(n_30),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_2),
.B(n_5),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_2),
.B(n_19),
.Y(n_20)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

AND2x2_ASAP7_75t_SL g31 ( 
.A(n_2),
.B(n_4),
.Y(n_31)
);

INVx2_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_3),
.B(n_22),
.Y(n_37)
);

OR2x4_ASAP7_75t_L g49 ( 
.A(n_3),
.B(n_22),
.Y(n_49)
);

INVx2_ASAP7_75t_R g14 ( 
.A(n_4),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_4),
.B(n_16),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_4),
.B(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_5),
.B(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_5),
.B(n_20),
.Y(n_45)
);

CKINVDCx14_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_10),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_SL g10 ( 
.A(n_11),
.B(n_27),
.Y(n_10)
);

AOI21xp5_ASAP7_75t_L g11 ( 
.A1(n_12),
.A2(n_21),
.B(n_24),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_13),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_15),
.Y(n_13)
);

AND2x2_ASAP7_75t_SL g29 ( 
.A(n_14),
.B(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_14),
.B(n_43),
.Y(n_52)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

NAND3xp33_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_18),
.C(n_20),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_21),
.A2(n_28),
.B1(n_29),
.B2(n_31),
.Y(n_27)
);

AND2x4_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_23),
.Y(n_21)
);

OR2x4_ASAP7_75t_L g25 ( 
.A(n_22),
.B(n_23),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_26),
.Y(n_24)
);

INVx2_ASAP7_75t_SL g28 ( 
.A(n_25),
.Y(n_28)
);

AOI22x1_ASAP7_75t_R g47 ( 
.A1(n_29),
.A2(n_31),
.B1(n_37),
.B2(n_48),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_36),
.B(n_38),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_38),
.B(n_49),
.Y(n_50)
);

BUFx12f_ASAP7_75t_SL g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_45),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);


endmodule