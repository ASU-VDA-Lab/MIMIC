module fake_ariane_3232_n_2935 (n_295, n_356, n_556, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_516, n_332, n_581, n_294, n_197, n_463, n_176, n_34, n_404, n_172, n_347, n_423, n_183, n_469, n_479, n_373, n_299, n_541, n_499, n_12, n_564, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_421, n_96, n_549, n_522, n_319, n_49, n_20, n_416, n_283, n_50, n_187, n_525, n_367, n_345, n_374, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_443, n_586, n_57, n_424, n_528, n_584, n_387, n_406, n_117, n_139, n_524, n_85, n_130, n_349, n_391, n_466, n_346, n_214, n_348, n_552, n_2, n_462, n_32, n_410, n_379, n_445, n_515, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_441, n_568, n_385, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_23, n_399, n_554, n_520, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_473, n_186, n_202, n_145, n_193, n_500, n_59, n_336, n_315, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_339, n_487, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_446, n_553, n_143, n_566, n_578, n_152, n_405, n_557, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_559, n_401, n_485, n_267, n_495, n_504, n_483, n_335, n_435, n_350, n_291, n_344, n_381, n_426, n_433, n_481, n_398, n_62, n_210, n_200, n_529, n_502, n_166, n_253, n_561, n_218, n_79, n_3, n_271, n_465, n_486, n_507, n_247, n_569, n_567, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_547, n_420, n_562, n_518, n_439, n_222, n_478, n_510, n_256, n_326, n_227, n_48, n_188, n_323, n_550, n_330, n_400, n_11, n_129, n_126, n_282, n_328, n_368, n_277, n_248, n_301, n_467, n_432, n_545, n_536, n_293, n_228, n_325, n_276, n_93, n_427, n_108, n_587, n_497, n_303, n_442, n_168, n_81, n_1, n_206, n_352, n_538, n_576, n_511, n_238, n_365, n_429, n_455, n_588, n_136, n_334, n_192, n_488, n_300, n_533, n_505, n_14, n_163, n_88, n_141, n_390, n_498, n_104, n_501, n_438, n_314, n_16, n_440, n_273, n_305, n_539, n_312, n_233, n_56, n_60, n_388, n_333, n_449, n_413, n_392, n_376, n_512, n_579, n_459, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_237, n_175, n_453, n_74, n_491, n_19, n_40, n_181, n_570, n_53, n_260, n_362, n_543, n_310, n_236, n_565, n_281, n_24, n_7, n_461, n_209, n_262, n_490, n_17, n_225, n_235, n_464, n_575, n_546, n_297, n_503, n_290, n_527, n_46, n_84, n_371, n_199, n_107, n_217, n_452, n_178, n_42, n_551, n_308, n_417, n_201, n_70, n_572, n_343, n_10, n_414, n_571, n_287, n_302, n_380, n_6, n_582, n_94, n_284, n_4, n_448, n_249, n_534, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_278, n_255, n_560, n_450, n_257, n_148, n_451, n_475, n_135, n_409, n_171, n_519, n_384, n_468, n_61, n_526, n_102, n_182, n_482, n_316, n_196, n_125, n_43, n_577, n_407, n_13, n_27, n_254, n_476, n_460, n_219, n_55, n_535, n_231, n_366, n_555, n_234, n_492, n_574, n_280, n_215, n_252, n_161, n_454, n_298, n_532, n_68, n_415, n_78, n_63, n_99, n_540, n_216, n_544, n_5, n_514, n_418, n_537, n_223, n_403, n_25, n_83, n_389, n_513, n_288, n_179, n_395, n_195, n_213, n_110, n_304, n_67, n_509, n_583, n_306, n_313, n_92, n_430, n_493, n_203, n_378, n_436, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_585, n_337, n_437, n_111, n_21, n_274, n_472, n_296, n_265, n_208, n_456, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_521, n_51, n_496, n_76, n_342, n_26, n_246, n_517, n_530, n_0, n_428, n_159, n_358, n_105, n_580, n_30, n_494, n_131, n_263, n_434, n_360, n_563, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_542, n_548, n_523, n_268, n_266, n_470, n_457, n_164, n_157, n_184, n_177, n_477, n_364, n_258, n_425, n_431, n_508, n_118, n_121, n_411, n_484, n_353, n_22, n_241, n_29, n_357, n_412, n_447, n_191, n_382, n_489, n_80, n_480, n_211, n_97, n_408, n_322, n_251, n_506, n_558, n_116, n_397, n_471, n_351, n_39, n_393, n_474, n_359, n_155, n_573, n_127, n_531, n_2935);

input n_295;
input n_356;
input n_556;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_516;
input n_332;
input n_581;
input n_294;
input n_197;
input n_463;
input n_176;
input n_34;
input n_404;
input n_172;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_373;
input n_299;
input n_541;
input n_499;
input n_12;
input n_564;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_549;
input n_522;
input n_319;
input n_49;
input n_20;
input n_416;
input n_283;
input n_50;
input n_187;
input n_525;
input n_367;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_443;
input n_586;
input n_57;
input n_424;
input n_528;
input n_584;
input n_387;
input n_406;
input n_117;
input n_139;
input n_524;
input n_85;
input n_130;
input n_349;
input n_391;
input n_466;
input n_346;
input n_214;
input n_348;
input n_552;
input n_2;
input n_462;
input n_32;
input n_410;
input n_379;
input n_445;
input n_515;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_568;
input n_385;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_23;
input n_399;
input n_554;
input n_520;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_202;
input n_145;
input n_193;
input n_500;
input n_59;
input n_336;
input n_315;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_487;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_446;
input n_553;
input n_143;
input n_566;
input n_578;
input n_152;
input n_405;
input n_557;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_559;
input n_401;
input n_485;
input n_267;
input n_495;
input n_504;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_344;
input n_381;
input n_426;
input n_433;
input n_481;
input n_398;
input n_62;
input n_210;
input n_200;
input n_529;
input n_502;
input n_166;
input n_253;
input n_561;
input n_218;
input n_79;
input n_3;
input n_271;
input n_465;
input n_486;
input n_507;
input n_247;
input n_569;
input n_567;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_547;
input n_420;
input n_562;
input n_518;
input n_439;
input n_222;
input n_478;
input n_510;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_550;
input n_330;
input n_400;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_545;
input n_536;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_427;
input n_108;
input n_587;
input n_497;
input n_303;
input n_442;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_538;
input n_576;
input n_511;
input n_238;
input n_365;
input n_429;
input n_455;
input n_588;
input n_136;
input n_334;
input n_192;
input n_488;
input n_300;
input n_533;
input n_505;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_498;
input n_104;
input n_501;
input n_438;
input n_314;
input n_16;
input n_440;
input n_273;
input n_305;
input n_539;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_449;
input n_413;
input n_392;
input n_376;
input n_512;
input n_579;
input n_459;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_237;
input n_175;
input n_453;
input n_74;
input n_491;
input n_19;
input n_40;
input n_181;
input n_570;
input n_53;
input n_260;
input n_362;
input n_543;
input n_310;
input n_236;
input n_565;
input n_281;
input n_24;
input n_7;
input n_461;
input n_209;
input n_262;
input n_490;
input n_17;
input n_225;
input n_235;
input n_464;
input n_575;
input n_546;
input n_297;
input n_503;
input n_290;
input n_527;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_217;
input n_452;
input n_178;
input n_42;
input n_551;
input n_308;
input n_417;
input n_201;
input n_70;
input n_572;
input n_343;
input n_10;
input n_414;
input n_571;
input n_287;
input n_302;
input n_380;
input n_6;
input n_582;
input n_94;
input n_284;
input n_4;
input n_448;
input n_249;
input n_534;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_278;
input n_255;
input n_560;
input n_450;
input n_257;
input n_148;
input n_451;
input n_475;
input n_135;
input n_409;
input n_171;
input n_519;
input n_384;
input n_468;
input n_61;
input n_526;
input n_102;
input n_182;
input n_482;
input n_316;
input n_196;
input n_125;
input n_43;
input n_577;
input n_407;
input n_13;
input n_27;
input n_254;
input n_476;
input n_460;
input n_219;
input n_55;
input n_535;
input n_231;
input n_366;
input n_555;
input n_234;
input n_492;
input n_574;
input n_280;
input n_215;
input n_252;
input n_161;
input n_454;
input n_298;
input n_532;
input n_68;
input n_415;
input n_78;
input n_63;
input n_99;
input n_540;
input n_216;
input n_544;
input n_5;
input n_514;
input n_418;
input n_537;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_513;
input n_288;
input n_179;
input n_395;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_509;
input n_583;
input n_306;
input n_313;
input n_92;
input n_430;
input n_493;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_585;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_472;
input n_296;
input n_265;
input n_208;
input n_456;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_521;
input n_51;
input n_496;
input n_76;
input n_342;
input n_26;
input n_246;
input n_517;
input n_530;
input n_0;
input n_428;
input n_159;
input n_358;
input n_105;
input n_580;
input n_30;
input n_494;
input n_131;
input n_263;
input n_434;
input n_360;
input n_563;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_542;
input n_548;
input n_523;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_425;
input n_431;
input n_508;
input n_118;
input n_121;
input n_411;
input n_484;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_412;
input n_447;
input n_191;
input n_382;
input n_489;
input n_80;
input n_480;
input n_211;
input n_97;
input n_408;
input n_322;
input n_251;
input n_506;
input n_558;
input n_116;
input n_397;
input n_471;
input n_351;
input n_39;
input n_393;
input n_474;
input n_359;
input n_155;
input n_573;
input n_127;
input n_531;

output n_2935;

wire n_2752;
wire n_913;
wire n_1681;
wire n_2163;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_2484;
wire n_2866;
wire n_1174;
wire n_2346;
wire n_1469;
wire n_691;
wire n_1353;
wire n_2679;
wire n_1355;
wire n_2131;
wire n_2559;
wire n_2500;
wire n_2509;
wire n_1383;
wire n_2182;
wire n_603;
wire n_2135;
wire n_2334;
wire n_2680;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_2879;
wire n_610;
wire n_1713;
wire n_1436;
wire n_2407;
wire n_690;
wire n_2818;
wire n_1109;
wire n_1430;
wire n_2537;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_1238;
wire n_2694;
wire n_2011;
wire n_2729;
wire n_1515;
wire n_1837;
wire n_817;
wire n_924;
wire n_781;
wire n_2013;
wire n_2786;
wire n_1566;
wire n_2837;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_2446;
wire n_1096;
wire n_1379;
wire n_2436;
wire n_2376;
wire n_2367;
wire n_2671;
wire n_2790;
wire n_1706;
wire n_2207;
wire n_2461;
wire n_2702;
wire n_2731;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_2238;
wire n_2529;
wire n_2374;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_2380;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_2646;
wire n_1298;
wire n_737;
wire n_2653;
wire n_1745;
wire n_2873;
wire n_1366;
wire n_2084;
wire n_2278;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_2482;
wire n_1682;
wire n_2750;
wire n_1836;
wire n_870;
wire n_2547;
wire n_1453;
wire n_945;
wire n_958;
wire n_2554;
wire n_2248;
wire n_813;
wire n_1985;
wire n_2288;
wire n_2621;
wire n_2908;
wire n_995;
wire n_2579;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_2323;
wire n_1073;
wire n_2844;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_738;
wire n_1690;
wire n_2221;
wire n_2807;
wire n_672;
wire n_740;
wire n_1283;
wire n_2317;
wire n_2838;
wire n_1974;
wire n_2906;
wire n_1736;
wire n_1018;
wire n_2342;
wire n_2200;
wire n_2781;
wire n_2442;
wire n_2735;
wire n_953;
wire n_1364;
wire n_2390;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_2634;
wire n_2709;
wire n_625;
wire n_2322;
wire n_2746;
wire n_1107;
wire n_2832;
wire n_1688;
wire n_989;
wire n_645;
wire n_1944;
wire n_2233;
wire n_2370;
wire n_2663;
wire n_2914;
wire n_1988;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_1428;
wire n_1284;
wire n_2878;
wire n_1241;
wire n_821;
wire n_770;
wire n_1514;
wire n_2539;
wire n_1528;
wire n_901;
wire n_2782;
wire n_2078;
wire n_1145;
wire n_971;
wire n_2359;
wire n_2201;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_2232;
wire n_1847;
wire n_2458;
wire n_2779;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_2227;
wire n_2301;
wire n_1539;
wire n_2859;
wire n_2847;
wire n_884;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_1636;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_1977;
wire n_693;
wire n_863;
wire n_2650;
wire n_1254;
wire n_929;
wire n_2433;
wire n_1703;
wire n_899;
wire n_2332;
wire n_2391;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_2571;
wire n_2427;
wire n_2885;
wire n_661;
wire n_2098;
wire n_2616;
wire n_1751;
wire n_2874;
wire n_2867;
wire n_1917;
wire n_2456;
wire n_2769;
wire n_1924;
wire n_1560;
wire n_1654;
wire n_2341;
wire n_2899;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_2575;
wire n_2722;
wire n_1396;
wire n_1230;
wire n_612;
wire n_1840;
wire n_2739;
wire n_1597;
wire n_1771;
wire n_2902;
wire n_1544;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2685;
wire n_2094;
wire n_2512;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_2382;
wire n_2043;
wire n_780;
wire n_2349;
wire n_1918;
wire n_2788;
wire n_1443;
wire n_1021;
wire n_2595;
wire n_1465;
wire n_2686;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_2727;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_1121;
wire n_1416;
wire n_2909;
wire n_1461;
wire n_2717;
wire n_1391;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_2527;
wire n_1112;
wire n_1159;
wire n_700;
wire n_772;
wire n_1216;
wire n_2759;
wire n_1245;
wire n_2743;
wire n_1669;
wire n_1675;
wire n_2466;
wire n_676;
wire n_2038;
wire n_2263;
wire n_2800;
wire n_2568;
wire n_2116;
wire n_2271;
wire n_2145;
wire n_2326;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_2806;
wire n_1716;
wire n_1872;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_1108;
wire n_851;
wire n_1590;
wire n_1351;
wire n_2216;
wire n_1274;
wire n_2426;
wire n_652;
wire n_1819;
wire n_947;
wire n_2134;
wire n_1260;
wire n_930;
wire n_1179;
wire n_2703;
wire n_1442;
wire n_696;
wire n_2926;
wire n_2620;
wire n_798;
wire n_1833;
wire n_1691;
wire n_916;
wire n_1386;
wire n_2810;
wire n_912;
wire n_1884;
wire n_1555;
wire n_1842;
wire n_2549;
wire n_2499;
wire n_1253;
wire n_1468;
wire n_762;
wire n_1661;
wire n_2791;
wire n_2683;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_2855;
wire n_2166;
wire n_2848;
wire n_1692;
wire n_2611;
wire n_1562;
wire n_2748;
wire n_2185;
wire n_2398;
wire n_1376;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_2925;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_2415;
wire n_2693;
wire n_2877;
wire n_2922;
wire n_2871;
wire n_2930;
wire n_2745;
wire n_2087;
wire n_931;
wire n_1491;
wire n_669;
wire n_2628;
wire n_619;
wire n_1083;
wire n_967;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1787;
wire n_2462;
wire n_1389;
wire n_2155;
wire n_2659;
wire n_615;
wire n_1139;
wire n_2836;
wire n_2439;
wire n_2864;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_2172;
wire n_2601;
wire n_892;
wire n_1880;
wire n_959;
wire n_2365;
wire n_2257;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_2219;
wire n_1855;
wire n_2100;
wire n_2333;
wire n_1623;
wire n_990;
wire n_1903;
wire n_867;
wire n_2147;
wire n_2435;
wire n_1226;
wire n_2224;
wire n_944;
wire n_1932;
wire n_749;
wire n_1780;
wire n_2825;
wire n_2888;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_2167;
wire n_2293;
wire n_2753;
wire n_1340;
wire n_2668;
wire n_1240;
wire n_2921;
wire n_1087;
wire n_2701;
wire n_2400;
wire n_632;
wire n_650;
wire n_2388;
wire n_2273;
wire n_2712;
wire n_1433;
wire n_1911;
wire n_2567;
wire n_2557;
wire n_2695;
wire n_2898;
wire n_1908;
wire n_1825;
wire n_1155;
wire n_2598;
wire n_1071;
wire n_2755;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_2795;
wire n_2682;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_2762;
wire n_964;
wire n_1627;
wire n_2220;
wire n_2294;
wire n_2274;
wire n_2895;
wire n_2903;
wire n_974;
wire n_1731;
wire n_799;
wire n_1147;
wire n_2829;
wire n_2378;
wire n_2467;
wire n_2768;
wire n_1914;
wire n_965;
wire n_2253;
wire n_934;
wire n_2213;
wire n_1447;
wire n_2363;
wire n_1220;
wire n_2019;
wire n_698;
wire n_2728;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_2924;
wire n_1209;
wire n_1563;
wire n_1020;
wire n_646;
wire n_2507;
wire n_2142;
wire n_1633;
wire n_2625;
wire n_2896;
wire n_1913;
wire n_2069;
wire n_2495;
wire n_1058;
wire n_2328;
wire n_2434;
wire n_1042;
wire n_1234;
wire n_2311;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_2287;
wire n_836;
wire n_2223;
wire n_1279;
wire n_2473;
wire n_2144;
wire n_2511;
wire n_1029;
wire n_2649;
wire n_1247;
wire n_760;
wire n_2438;
wire n_1568;
wire n_2919;
wire n_1483;
wire n_1363;
wire n_2681;
wire n_1111;
wire n_970;
wire n_1689;
wire n_2535;
wire n_713;
wire n_1255;
wire n_2632;
wire n_1646;
wire n_598;
wire n_2262;
wire n_2565;
wire n_1237;
wire n_927;
wire n_1095;
wire n_1728;
wire n_2335;
wire n_706;
wire n_2120;
wire n_2631;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_2860;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_2697;
wire n_1387;
wire n_1263;
wire n_1817;
wire n_2404;
wire n_2168;
wire n_2757;
wire n_2312;
wire n_670;
wire n_2677;
wire n_1826;
wire n_2834;
wire n_2483;
wire n_1951;
wire n_2490;
wire n_1032;
wire n_1217;
wire n_2558;
wire n_1496;
wire n_637;
wire n_1592;
wire n_2812;
wire n_2662;
wire n_1259;
wire n_2801;
wire n_1177;
wire n_2655;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_2718;
wire n_720;
wire n_926;
wire n_1943;
wire n_2687;
wire n_2296;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_2765;
wire n_1163;
wire n_2640;
wire n_2811;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_2241;
wire n_2373;
wire n_1173;
wire n_2350;
wire n_1068;
wire n_1198;
wire n_2531;
wire n_1570;
wire n_2099;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2617;
wire n_2481;
wire n_2129;
wire n_855;
wire n_2327;
wire n_808;
wire n_1365;
wire n_2476;
wire n_2814;
wire n_2059;
wire n_2437;
wire n_2636;
wire n_1439;
wire n_814;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_2841;
wire n_1611;
wire n_2122;
wire n_2399;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_2932;
wire n_1423;
wire n_2117;
wire n_600;
wire n_1609;
wire n_1053;
wire n_2822;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_1906;
wire n_1899;
wire n_2195;
wire n_2194;
wire n_1467;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_2267;
wire n_1105;
wire n_604;
wire n_677;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_681;
wire n_874;
wire n_2286;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_2783;
wire n_2599;
wire n_590;
wire n_699;
wire n_2075;
wire n_727;
wire n_1726;
wire n_2523;
wire n_1945;
wire n_1015;
wire n_2418;
wire n_1377;
wire n_1162;
wire n_1614;
wire n_2031;
wire n_2496;
wire n_2118;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_2853;
wire n_1098;
wire n_1490;
wire n_2338;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_2802;
wire n_729;
wire n_887;
wire n_2057;
wire n_2218;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_2593;
wire n_1693;
wire n_2125;
wire n_2716;
wire n_1132;
wire n_1156;
wire n_2741;
wire n_2184;
wire n_2714;
wire n_1823;
wire n_2861;
wire n_2780;
wire n_1120;
wire n_1202;
wire n_627;
wire n_2254;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_2618;
wire n_1402;
wire n_957;
wire n_1242;
wire n_2774;
wire n_2707;
wire n_2754;
wire n_2849;
wire n_1607;
wire n_1489;
wire n_2799;
wire n_1218;
wire n_2756;
wire n_2217;
wire n_2226;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_2763;
wire n_2256;
wire n_1189;
wire n_1089;
wire n_1859;
wire n_2660;
wire n_1502;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_2732;
wire n_1883;
wire n_2516;
wire n_2776;
wire n_2555;
wire n_1969;
wire n_2708;
wire n_735;
wire n_1005;
wire n_2379;
wire n_1294;
wire n_2661;
wire n_1667;
wire n_888;
wire n_845;
wire n_2894;
wire n_2300;
wire n_1649;
wire n_2452;
wire n_1677;
wire n_2470;
wire n_1927;
wire n_1297;
wire n_2827;
wire n_1708;
wire n_1222;
wire n_2284;
wire n_1844;
wire n_2283;
wire n_2526;
wire n_1957;
wire n_1953;
wire n_2643;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_1919;
wire n_710;
wire n_1791;
wire n_2508;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_2594;
wire n_2266;
wire n_2449;
wire n_890;
wire n_842;
wire n_1898;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_1373;
wire n_1081;
wire n_1975;
wire n_742;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_2119;
wire n_1719;
wire n_2742;
wire n_769;
wire n_1797;
wire n_2366;
wire n_2493;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_832;
wire n_744;
wire n_1895;
wire n_2821;
wire n_2690;
wire n_2474;
wire n_2623;
wire n_1800;
wire n_982;
wire n_915;
wire n_1075;
wire n_2008;
wire n_1331;
wire n_1890;
wire n_2904;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_1860;
wire n_1734;
wire n_2460;
wire n_2840;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_2448;
wire n_2211;
wire n_2292;
wire n_2480;
wire n_606;
wire n_951;
wire n_2772;
wire n_1700;
wire n_862;
wire n_2637;
wire n_659;
wire n_1332;
wire n_2306;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_2424;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2414;
wire n_2082;
wire n_2893;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_2389;
wire n_1309;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_2737;
wire n_1867;
wire n_852;
wire n_1394;
wire n_2916;
wire n_2576;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_2696;
wire n_2140;
wire n_1748;
wire n_1301;
wire n_873;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_2468;
wire n_1400;
wire n_2035;
wire n_2614;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_2581;
wire n_1783;
wire n_608;
wire n_2494;
wire n_1538;
wire n_2831;
wire n_2457;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_1993;
wire n_1545;
wire n_2629;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_2540;
wire n_1605;
wire n_1078;
wire n_2486;
wire n_1897;
wire n_2520;
wire n_2137;
wire n_1161;
wire n_2489;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_1191;
wire n_618;
wire n_2492;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_2337;
wire n_2265;
wire n_687;
wire n_2900;
wire n_797;
wire n_2026;
wire n_2912;
wire n_1786;
wire n_2627;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_2106;
wire n_1406;
wire n_595;
wire n_1405;
wire n_2684;
wire n_2726;
wire n_602;
wire n_2622;
wire n_2272;
wire n_1757;
wire n_592;
wire n_1499;
wire n_1318;
wire n_854;
wire n_2091;
wire n_1632;
wire n_1769;
wire n_1929;
wire n_1950;
wire n_2264;
wire n_2691;
wire n_805;
wire n_2032;
wire n_2090;
wire n_2929;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_2785;
wire n_1596;
wire n_2348;
wire n_2656;
wire n_1281;
wire n_2364;
wire n_1997;
wire n_2574;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_1856;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_2016;
wire n_2667;
wire n_2725;
wire n_2928;
wire n_943;
wire n_1118;
wire n_678;
wire n_2905;
wire n_2884;
wire n_651;
wire n_2850;
wire n_1874;
wire n_1293;
wire n_961;
wire n_1046;
wire n_1807;
wire n_1123;
wire n_726;
wire n_1657;
wire n_878;
wire n_2857;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_2307;
wire n_1488;
wire n_985;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_2730;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_2412;
wire n_2720;
wire n_1352;
wire n_2405;
wire n_2815;
wire n_1824;
wire n_643;
wire n_2606;
wire n_2700;
wire n_1492;
wire n_2383;
wire n_2764;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_2633;
wire n_2416;
wire n_819;
wire n_2386;
wire n_2907;
wire n_1971;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_2353;
wire n_2528;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_2325;
wire n_1130;
wire n_1450;
wire n_2022;
wire n_756;
wire n_2298;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_2408;
wire n_2698;
wire n_2320;
wire n_979;
wire n_2329;
wire n_2570;
wire n_1642;
wire n_2417;
wire n_2789;
wire n_2525;
wire n_1815;
wire n_2813;
wire n_897;
wire n_2546;
wire n_949;
wire n_2454;
wire n_1493;
wire n_2890;
wire n_2911;
wire n_807;
wire n_891;
wire n_1659;
wire n_885;
wire n_2354;
wire n_1864;
wire n_2760;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_2368;
wire n_802;
wire n_1151;
wire n_960;
wire n_2352;
wire n_2502;
wire n_1256;
wire n_714;
wire n_2170;
wire n_790;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_725;
wire n_2377;
wire n_1577;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_2652;
wire n_1133;
wire n_883;
wire n_1852;
wire n_801;
wire n_1286;
wire n_2612;
wire n_818;
wire n_1685;
wire n_779;
wire n_2410;
wire n_2314;
wire n_2477;
wire n_2279;
wire n_594;
wire n_2222;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2133;
wire n_2203;
wire n_833;
wire n_1426;
wire n_2250;
wire n_2497;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_2506;
wire n_1472;
wire n_2413;
wire n_1593;
wire n_2610;
wire n_1050;
wire n_2626;
wire n_2158;
wire n_2578;
wire n_2607;
wire n_2285;
wire n_2892;
wire n_1288;
wire n_1201;
wire n_2605;
wire n_858;
wire n_2796;
wire n_1185;
wire n_2475;
wire n_2804;
wire n_2173;
wire n_2715;
wire n_1035;
wire n_1143;
wire n_2665;
wire n_2070;
wire n_2136;
wire n_2771;
wire n_1090;
wire n_2403;
wire n_1367;
wire n_2044;
wire n_928;
wire n_1153;
wire n_1103;
wire n_825;
wire n_732;
wire n_2619;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_2854;
wire n_1291;
wire n_2020;
wire n_748;
wire n_2310;
wire n_1045;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_2711;
wire n_1881;
wire n_2635;
wire n_988;
wire n_914;
wire n_689;
wire n_1116;
wire n_1958;
wire n_2747;
wire n_1511;
wire n_2177;
wire n_2713;
wire n_1422;
wire n_2766;
wire n_1965;
wire n_644;
wire n_1197;
wire n_2820;
wire n_2613;
wire n_1165;
wire n_2934;
wire n_1641;
wire n_2845;
wire n_1517;
wire n_2036;
wire n_843;
wire n_2647;
wire n_638;
wire n_2003;
wire n_2533;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_2343;
wire n_775;
wire n_667;
wire n_2419;
wire n_1049;
wire n_2330;
wire n_2826;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_2777;
wire n_2450;
wire n_2411;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_2309;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_2431;
wire n_1773;
wire n_1440;
wire n_2666;
wire n_1370;
wire n_1603;
wire n_728;
wire n_2401;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_2588;
wire n_2863;
wire n_2331;
wire n_935;
wire n_2886;
wire n_2478;
wire n_685;
wire n_911;
wire n_2658;
wire n_623;
wire n_2608;
wire n_2920;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_1534;
wire n_1948;
wire n_2767;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_2396;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_2692;
wire n_601;
wire n_683;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_2862;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_2553;
wire n_2645;
wire n_907;
wire n_2749;
wire n_1454;
wire n_2592;
wire n_660;
wire n_2459;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_2566;
wire n_2751;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_673;
wire n_2842;
wire n_2833;
wire n_2196;
wire n_1038;
wire n_2371;
wire n_1978;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_593;
wire n_1695;
wire n_2560;
wire n_1164;
wire n_2313;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_2609;
wire n_2561;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_1653;
wire n_872;
wire n_2882;
wire n_2303;
wire n_2669;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_629;
wire n_1739;
wire n_2642;
wire n_1814;
wire n_2154;
wire n_2441;
wire n_2236;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_2688;
wire n_692;
wire n_2624;
wire n_2054;
wire n_1857;
wire n_2315;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_2498;
wire n_800;
wire n_2638;
wire n_2046;
wire n_1910;
wire n_1816;
wire n_2803;
wire n_1756;
wire n_2887;
wire n_1606;
wire n_2189;
wire n_621;
wire n_2648;
wire n_1587;
wire n_2093;
wire n_2340;
wire n_2018;
wire n_2672;
wire n_1772;
wire n_2444;
wire n_2602;
wire n_1014;
wire n_724;
wire n_2204;
wire n_2931;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_1311;
wire n_2199;
wire n_2881;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_875;
wire n_1617;
wire n_2455;
wire n_827;
wire n_2600;
wire n_2231;
wire n_697;
wire n_2828;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_2305;
wire n_880;
wire n_793;
wire n_2114;
wire n_2927;
wire n_1175;
wire n_2289;
wire n_2530;
wire n_2299;
wire n_751;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_2883;
wire n_1221;
wire n_1785;
wire n_1262;
wire n_792;
wire n_1942;
wire n_2180;
wire n_1579;
wire n_2809;
wire n_2181;
wire n_2014;
wire n_975;
wire n_1645;
wire n_923;
wire n_1124;
wire n_1381;
wire n_2870;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_2889;
wire n_2276;
wire n_1805;
wire n_2282;
wire n_981;
wire n_2910;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_2503;
wire n_2270;
wire n_2443;
wire n_1407;
wire n_2465;
wire n_1204;
wire n_2865;
wire n_1554;
wire n_994;
wire n_2428;
wire n_2586;
wire n_1360;
wire n_973;
wire n_2858;
wire n_972;
wire n_2251;
wire n_2923;
wire n_2843;
wire n_856;
wire n_2572;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_1679;
wire n_2872;
wire n_2126;
wire n_1952;
wire n_2425;
wire n_2394;
wire n_1858;
wire n_1678;
wire n_2589;
wire n_1482;
wire n_1361;
wire n_2356;
wire n_1601;
wire n_1057;
wire n_2487;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_2534;
wire n_2488;
wire n_1509;
wire n_828;
wire n_1411;
wire n_1359;
wire n_1721;
wire n_2564;
wire n_2591;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_2197;
wire n_783;
wire n_2550;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_2385;
wire n_2387;
wire n_1008;
wire n_1024;
wire n_830;
wire n_2291;
wire n_2816;
wire n_1980;
wire n_2518;
wire n_987;
wire n_936;
wire n_2510;
wire n_1620;
wire n_2501;
wire n_2542;
wire n_1385;
wire n_1525;
wire n_2793;
wire n_1998;
wire n_2165;
wire n_2675;
wire n_2604;
wire n_1775;
wire n_908;
wire n_788;
wire n_2639;
wire n_1036;
wire n_2169;
wire n_2603;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_2630;
wire n_591;
wire n_2794;
wire n_969;
wire n_2028;
wire n_1663;
wire n_919;
wire n_2901;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_2773;
wire n_2817;
wire n_1926;
wire n_2402;
wire n_1458;
wire n_679;
wire n_1630;
wire n_663;
wire n_1720;
wire n_2409;
wire n_2176;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_1358;
wire n_1200;
wire n_826;
wire n_2808;
wire n_2453;
wire n_2344;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_940;
wire n_2392;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_2543;
wire n_2321;
wire n_1077;
wire n_2597;
wire n_607;
wire n_956;
wire n_1930;
wire n_765;
wire n_1809;
wire n_2787;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_2805;
wire n_1268;
wire n_2676;
wire n_2758;
wire n_2395;
wire n_917;
wire n_2868;
wire n_2723;
wire n_1271;
wire n_2096;
wire n_2440;
wire n_2556;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_2770;
wire n_631;
wire n_1170;
wire n_2724;
wire n_2258;
wire n_1261;
wire n_2471;
wire n_702;
wire n_857;
wire n_898;
wire n_1067;
wire n_968;
wire n_1235;
wire n_1323;
wire n_2584;
wire n_2375;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_2212;
wire n_731;
wire n_1813;
wire n_2268;
wire n_1452;
wire n_2835;
wire n_1573;
wire n_2734;
wire n_668;
wire n_2569;
wire n_758;
wire n_2252;
wire n_2111;
wire n_2420;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_816;
wire n_2897;
wire n_1322;
wire n_2583;
wire n_2918;
wire n_1473;
wire n_835;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_2651;
wire n_753;
wire n_2445;
wire n_2733;
wire n_1770;
wire n_701;
wire n_1003;
wire n_2469;
wire n_1125;
wire n_2103;
wire n_2358;
wire n_1865;
wire n_1710;
wire n_2522;
wire n_2641;
wire n_2463;
wire n_1344;
wire n_2355;
wire n_1390;
wire n_2580;
wire n_2699;
wire n_1792;
wire n_2062;
wire n_1141;
wire n_1629;
wire n_1640;
wire n_822;
wire n_1094;
wire n_1459;
wire n_840;
wire n_2153;
wire n_2324;
wire n_1510;
wire n_2710;
wire n_2505;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_2397;
wire n_2521;
wire n_1727;
wire n_2740;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_2721;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_2615;
wire n_614;
wire n_2775;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_2351;
wire n_2260;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_2206;
wire n_2784;
wire n_2541;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_2347;
wire n_1152;
wire n_2657;
wire n_2538;
wire n_2034;
wire n_1845;
wire n_2447;
wire n_1934;
wire n_2101;
wire n_2577;
wire n_921;
wire n_2362;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_2372;
wire n_2552;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_2422;
wire n_2704;
wire n_1334;
wire n_654;
wire n_2290;
wire n_2933;
wire n_2856;
wire n_2088;
wire n_1275;
wire n_904;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2429;
wire n_2108;
wire n_2736;
wire n_1039;
wire n_2246;
wire n_1150;
wire n_977;
wire n_2339;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2532;
wire n_2191;
wire n_1497;
wire n_1866;
wire n_2472;
wire n_2664;
wire n_2705;
wire n_2056;
wire n_2852;
wire n_1136;
wire n_2515;
wire n_1782;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_2519;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_2360;
wire n_723;
wire n_1393;
wire n_2240;
wire n_658;
wire n_630;
wire n_1369;
wire n_2846;
wire n_1781;
wire n_709;
wire n_2917;
wire n_2544;
wire n_809;
wire n_2085;
wire n_2432;
wire n_1686;
wire n_1964;
wire n_881;
wire n_1477;
wire n_1777;
wire n_2188;
wire n_1019;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_2430;
wire n_2504;
wire n_910;
wire n_741;
wire n_1410;
wire n_2297;
wire n_939;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_1223;
wire n_2545;
wire n_1768;
wire n_2513;
wire n_2193;
wire n_2369;
wire n_1199;
wire n_865;
wire n_1983;
wire n_1273;
wire n_1041;
wire n_2451;
wire n_2115;
wire n_2913;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_2587;
wire n_1347;
wire n_2839;
wire n_860;
wire n_1043;
wire n_2869;
wire n_1923;
wire n_2670;
wire n_1764;
wire n_2674;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_2644;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_2148;
wire n_933;
wire n_1779;
wire n_2562;
wire n_596;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_656;
wire n_2673;
wire n_664;
wire n_1591;
wire n_2585;
wire n_1229;
wire n_1683;
wire n_2582;
wire n_2548;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_2381;
wire n_2744;
wire n_1967;
wire n_2384;
wire n_2678;
wire n_2179;
wire n_1280;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_2485;
wire n_1063;
wire n_2205;
wire n_2183;
wire n_2275;
wire n_991;
wire n_2563;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2761;
wire n_2357;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_2875;
wire n_1639;
wire n_2209;
wire n_2421;
wire n_1302;
wire n_1000;
wire n_626;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_2792;
wire n_1634;
wire n_2596;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_2269;
wire n_937;
wire n_1474;
wire n_2081;
wire n_2536;
wire n_2524;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_1211;
wire n_1368;
wire n_996;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_2891;
wire n_2318;
wire n_1827;
wire n_866;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1722;
wire n_1001;
wire n_2361;
wire n_1115;
wire n_2229;
wire n_2819;
wire n_2880;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_2551;
wire n_719;
wire n_1102;
wire n_2255;
wire n_1129;
wire n_1252;
wire n_2239;
wire n_1464;
wire n_1296;
wire n_773;
wire n_2798;
wire n_2316;
wire n_2464;
wire n_1010;
wire n_2830;
wire n_882;
wire n_2706;
wire n_2304;
wire n_1249;
wire n_803;
wire n_1871;
wire n_2514;
wire n_718;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_2573;
wire n_2336;
wire n_1662;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_2915;
wire n_2654;
wire n_2491;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_2517;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_2259;
wire n_849;
wire n_2095;
wire n_2719;
wire n_2738;
wire n_1820;
wire n_2590;
wire n_2876;
wire n_2797;
wire n_1251;
wire n_1989;
wire n_1421;
wire n_2208;
wire n_2423;
wire n_2689;
wire n_2778;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_2479;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2824;
wire n_2037;
wire n_1308;
wire n_796;
wire n_2851;
wire n_2823;
wire n_2345;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_145),
.Y(n_589)
);

CKINVDCx20_ASAP7_75t_R g590 ( 
.A(n_582),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_275),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_405),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_356),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_560),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_111),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_415),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_341),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_400),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_304),
.Y(n_599)
);

CKINVDCx20_ASAP7_75t_R g600 ( 
.A(n_67),
.Y(n_600)
);

INVx1_ASAP7_75t_SL g601 ( 
.A(n_231),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_291),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_519),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_129),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_190),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_78),
.Y(n_606)
);

HB1xp67_ASAP7_75t_L g607 ( 
.A(n_414),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_147),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_360),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_534),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_237),
.Y(n_611)
);

BUFx2_ASAP7_75t_SL g612 ( 
.A(n_516),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_541),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_540),
.Y(n_614)
);

CKINVDCx20_ASAP7_75t_R g615 ( 
.A(n_349),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_296),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_103),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_324),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_349),
.Y(n_619)
);

BUFx2_ASAP7_75t_SL g620 ( 
.A(n_52),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_478),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_145),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_478),
.Y(n_623)
);

INVx2_ASAP7_75t_SL g624 ( 
.A(n_553),
.Y(n_624)
);

CKINVDCx20_ASAP7_75t_R g625 ( 
.A(n_66),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_285),
.Y(n_626)
);

CKINVDCx20_ASAP7_75t_R g627 ( 
.A(n_58),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_585),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_441),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_38),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_479),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_194),
.Y(n_632)
);

CKINVDCx20_ASAP7_75t_R g633 ( 
.A(n_190),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_406),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_84),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_460),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_90),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_269),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_530),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_207),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_558),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_102),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_384),
.Y(n_643)
);

INVxp67_ASAP7_75t_L g644 ( 
.A(n_86),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_304),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_517),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_58),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_557),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_178),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_421),
.Y(n_650)
);

CKINVDCx20_ASAP7_75t_R g651 ( 
.A(n_362),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_142),
.Y(n_652)
);

INVx2_ASAP7_75t_SL g653 ( 
.A(n_369),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_71),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_527),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_22),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_39),
.Y(n_657)
);

CKINVDCx14_ASAP7_75t_R g658 ( 
.A(n_283),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_536),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_581),
.Y(n_660)
);

BUFx3_ASAP7_75t_L g661 ( 
.A(n_51),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_465),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_1),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_553),
.Y(n_664)
);

INVx1_ASAP7_75t_SL g665 ( 
.A(n_169),
.Y(n_665)
);

CKINVDCx20_ASAP7_75t_R g666 ( 
.A(n_501),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_362),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_108),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_170),
.Y(n_669)
);

INVx1_ASAP7_75t_SL g670 ( 
.A(n_374),
.Y(n_670)
);

BUFx10_ASAP7_75t_L g671 ( 
.A(n_504),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_547),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_360),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_61),
.Y(n_674)
);

BUFx10_ASAP7_75t_L g675 ( 
.A(n_520),
.Y(n_675)
);

BUFx10_ASAP7_75t_L g676 ( 
.A(n_515),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_523),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_452),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_79),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_484),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_385),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_214),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_53),
.Y(n_683)
);

CKINVDCx20_ASAP7_75t_R g684 ( 
.A(n_447),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_22),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_535),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_493),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_178),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_586),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_529),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_188),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_275),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_321),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_558),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_138),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_555),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_223),
.Y(n_697)
);

CKINVDCx14_ASAP7_75t_R g698 ( 
.A(n_523),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_172),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_182),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_522),
.Y(n_701)
);

BUFx5_ASAP7_75t_L g702 ( 
.A(n_216),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_416),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_295),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_3),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_569),
.Y(n_706)
);

BUFx10_ASAP7_75t_L g707 ( 
.A(n_45),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_329),
.Y(n_708)
);

BUFx10_ASAP7_75t_L g709 ( 
.A(n_410),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_366),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_217),
.Y(n_711)
);

BUFx10_ASAP7_75t_L g712 ( 
.A(n_361),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_332),
.Y(n_713)
);

INVx1_ASAP7_75t_SL g714 ( 
.A(n_327),
.Y(n_714)
);

CKINVDCx16_ASAP7_75t_R g715 ( 
.A(n_303),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_229),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_239),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_524),
.Y(n_718)
);

BUFx3_ASAP7_75t_L g719 ( 
.A(n_449),
.Y(n_719)
);

CKINVDCx14_ASAP7_75t_R g720 ( 
.A(n_274),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_257),
.Y(n_721)
);

HB1xp67_ASAP7_75t_L g722 ( 
.A(n_109),
.Y(n_722)
);

INVx1_ASAP7_75t_SL g723 ( 
.A(n_269),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_365),
.Y(n_724)
);

HB1xp67_ASAP7_75t_L g725 ( 
.A(n_576),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_56),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_184),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_559),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_225),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_268),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_439),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_358),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_62),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_124),
.Y(n_734)
);

BUFx3_ASAP7_75t_L g735 ( 
.A(n_140),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_384),
.Y(n_736)
);

INVx1_ASAP7_75t_SL g737 ( 
.A(n_231),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_490),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_465),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_42),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_567),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_547),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_194),
.Y(n_743)
);

INVxp67_ASAP7_75t_SL g744 ( 
.A(n_470),
.Y(n_744)
);

BUFx3_ASAP7_75t_L g745 ( 
.A(n_259),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_548),
.Y(n_746)
);

INVx1_ASAP7_75t_SL g747 ( 
.A(n_317),
.Y(n_747)
);

INVx2_ASAP7_75t_SL g748 ( 
.A(n_426),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_260),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_575),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_351),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_550),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_33),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_401),
.Y(n_754)
);

CKINVDCx20_ASAP7_75t_R g755 ( 
.A(n_338),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_181),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_185),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_507),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_389),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_460),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_507),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_6),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_3),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_411),
.Y(n_764)
);

BUFx5_ASAP7_75t_L g765 ( 
.A(n_207),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_563),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_20),
.Y(n_767)
);

CKINVDCx11_ASAP7_75t_R g768 ( 
.A(n_40),
.Y(n_768)
);

BUFx10_ASAP7_75t_L g769 ( 
.A(n_532),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_463),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_420),
.Y(n_771)
);

BUFx6f_ASAP7_75t_L g772 ( 
.A(n_264),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_476),
.Y(n_773)
);

CKINVDCx20_ASAP7_75t_R g774 ( 
.A(n_459),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_385),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_383),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_292),
.Y(n_777)
);

BUFx3_ASAP7_75t_L g778 ( 
.A(n_107),
.Y(n_778)
);

CKINVDCx14_ASAP7_75t_R g779 ( 
.A(n_355),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_364),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_116),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_329),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_122),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_277),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_376),
.Y(n_785)
);

CKINVDCx20_ASAP7_75t_R g786 ( 
.A(n_71),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_533),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_401),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_24),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_96),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_88),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_111),
.Y(n_792)
);

CKINVDCx11_ASAP7_75t_R g793 ( 
.A(n_236),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_126),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_412),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_157),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_241),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_363),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_224),
.Y(n_799)
);

BUFx10_ASAP7_75t_L g800 ( 
.A(n_200),
.Y(n_800)
);

CKINVDCx20_ASAP7_75t_R g801 ( 
.A(n_240),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_552),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_110),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_310),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_57),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_531),
.Y(n_806)
);

BUFx2_ASAP7_75t_L g807 ( 
.A(n_311),
.Y(n_807)
);

CKINVDCx20_ASAP7_75t_R g808 ( 
.A(n_271),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_388),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_296),
.Y(n_810)
);

CKINVDCx16_ASAP7_75t_R g811 ( 
.A(n_323),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_47),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_12),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_336),
.Y(n_814)
);

BUFx3_ASAP7_75t_L g815 ( 
.A(n_518),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_246),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_515),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_5),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_374),
.Y(n_819)
);

CKINVDCx14_ASAP7_75t_R g820 ( 
.A(n_88),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_492),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_574),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_237),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_113),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_540),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_286),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_588),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_494),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_448),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_505),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_389),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_221),
.Y(n_832)
);

BUFx2_ASAP7_75t_SL g833 ( 
.A(n_491),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_427),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_510),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_98),
.Y(n_836)
);

CKINVDCx14_ASAP7_75t_R g837 ( 
.A(n_177),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_270),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_474),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_199),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_578),
.Y(n_841)
);

BUFx5_ASAP7_75t_L g842 ( 
.A(n_9),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_542),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_420),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_470),
.Y(n_845)
);

INVx1_ASAP7_75t_SL g846 ( 
.A(n_46),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_33),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_413),
.Y(n_848)
);

BUFx6f_ASAP7_75t_L g849 ( 
.A(n_441),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_357),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_96),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_555),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_47),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_249),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_322),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_564),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_89),
.Y(n_857)
);

INVx2_ASAP7_75t_SL g858 ( 
.A(n_27),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_451),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_169),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_54),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_283),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_68),
.Y(n_863)
);

CKINVDCx20_ASAP7_75t_R g864 ( 
.A(n_561),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_433),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_266),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_550),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_97),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_387),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_126),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_379),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_268),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_173),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_580),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_529),
.Y(n_875)
);

CKINVDCx20_ASAP7_75t_R g876 ( 
.A(n_562),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_491),
.Y(n_877)
);

BUFx10_ASAP7_75t_L g878 ( 
.A(n_526),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_78),
.Y(n_879)
);

INVx1_ASAP7_75t_SL g880 ( 
.A(n_393),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_483),
.Y(n_881)
);

INVx1_ASAP7_75t_SL g882 ( 
.A(n_68),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_41),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_239),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_454),
.Y(n_885)
);

CKINVDCx20_ASAP7_75t_R g886 ( 
.A(n_527),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_222),
.Y(n_887)
);

BUFx3_ASAP7_75t_L g888 ( 
.A(n_24),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_456),
.Y(n_889)
);

BUFx5_ASAP7_75t_L g890 ( 
.A(n_521),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_539),
.Y(n_891)
);

CKINVDCx20_ASAP7_75t_R g892 ( 
.A(n_458),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_437),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_545),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_363),
.Y(n_895)
);

INVxp67_ASAP7_75t_L g896 ( 
.A(n_551),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_366),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_215),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_423),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_528),
.Y(n_900)
);

CKINVDCx20_ASAP7_75t_R g901 ( 
.A(n_250),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_123),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_213),
.Y(n_903)
);

BUFx6f_ASAP7_75t_L g904 ( 
.A(n_504),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_424),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_66),
.Y(n_906)
);

INVx1_ASAP7_75t_SL g907 ( 
.A(n_42),
.Y(n_907)
);

BUFx10_ASAP7_75t_L g908 ( 
.A(n_189),
.Y(n_908)
);

CKINVDCx20_ASAP7_75t_R g909 ( 
.A(n_306),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_306),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_9),
.Y(n_911)
);

CKINVDCx20_ASAP7_75t_R g912 ( 
.A(n_473),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_563),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_583),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_577),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_483),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_171),
.Y(n_917)
);

CKINVDCx20_ASAP7_75t_R g918 ( 
.A(n_399),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_44),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_286),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_192),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_114),
.Y(n_922)
);

INVx1_ASAP7_75t_SL g923 ( 
.A(n_556),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_102),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_387),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_142),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_579),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_95),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_442),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_180),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_500),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_315),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_165),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_160),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_566),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_246),
.Y(n_936)
);

INVx3_ASAP7_75t_L g937 ( 
.A(n_32),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_147),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_267),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_254),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_150),
.Y(n_941)
);

INVx2_ASAP7_75t_SL g942 ( 
.A(n_62),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_411),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_484),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_546),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_549),
.Y(n_946)
);

BUFx6f_ASAP7_75t_L g947 ( 
.A(n_85),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_584),
.Y(n_948)
);

BUFx8_ASAP7_75t_SL g949 ( 
.A(n_400),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_543),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_517),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_382),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_554),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_587),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_538),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_195),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_136),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_532),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_5),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_473),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_218),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_544),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_463),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_165),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_226),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_28),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_461),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_55),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_184),
.Y(n_969)
);

INVx2_ASAP7_75t_SL g970 ( 
.A(n_255),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_421),
.Y(n_971)
);

BUFx6f_ASAP7_75t_L g972 ( 
.A(n_486),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_407),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_85),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_494),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_242),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_274),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_535),
.Y(n_978)
);

BUFx6f_ASAP7_75t_L g979 ( 
.A(n_570),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_198),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_331),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_543),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_77),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_254),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_568),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_99),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_417),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_292),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_573),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_443),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_571),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_72),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_144),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_471),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_157),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_148),
.Y(n_996)
);

INVx2_ASAP7_75t_SL g997 ( 
.A(n_337),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_464),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_514),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_100),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_46),
.Y(n_1001)
);

INVx1_ASAP7_75t_SL g1002 ( 
.A(n_312),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_261),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_238),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_127),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_36),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_114),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_224),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_222),
.Y(n_1009)
);

CKINVDCx20_ASAP7_75t_R g1010 ( 
.A(n_14),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_525),
.Y(n_1011)
);

INVxp67_ASAP7_75t_L g1012 ( 
.A(n_35),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_154),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_297),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_398),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_121),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_65),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_409),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_35),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_537),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_472),
.Y(n_1021)
);

BUFx3_ASAP7_75t_L g1022 ( 
.A(n_299),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_19),
.Y(n_1023)
);

BUFx3_ASAP7_75t_L g1024 ( 
.A(n_572),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_373),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_290),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_383),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_179),
.Y(n_1028)
);

BUFx10_ASAP7_75t_L g1029 ( 
.A(n_423),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_702),
.Y(n_1030)
);

INVxp67_ASAP7_75t_SL g1031 ( 
.A(n_937),
.Y(n_1031)
);

CKINVDCx20_ASAP7_75t_R g1032 ( 
.A(n_658),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_702),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_702),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_702),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_702),
.Y(n_1036)
);

CKINVDCx20_ASAP7_75t_R g1037 ( 
.A(n_698),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_702),
.Y(n_1038)
);

INVxp67_ASAP7_75t_SL g1039 ( 
.A(n_937),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_702),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_702),
.Y(n_1041)
);

HB1xp67_ASAP7_75t_L g1042 ( 
.A(n_807),
.Y(n_1042)
);

BUFx3_ASAP7_75t_L g1043 ( 
.A(n_1024),
.Y(n_1043)
);

HB1xp67_ASAP7_75t_L g1044 ( 
.A(n_807),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_702),
.Y(n_1045)
);

BUFx6f_ASAP7_75t_L g1046 ( 
.A(n_979),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_765),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_765),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_765),
.Y(n_1049)
);

INVxp67_ASAP7_75t_SL g1050 ( 
.A(n_937),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_765),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_765),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_765),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_765),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_765),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_765),
.Y(n_1056)
);

INVxp67_ASAP7_75t_SL g1057 ( 
.A(n_937),
.Y(n_1057)
);

INVxp67_ASAP7_75t_SL g1058 ( 
.A(n_719),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_842),
.Y(n_1059)
);

INVxp33_ASAP7_75t_SL g1060 ( 
.A(n_607),
.Y(n_1060)
);

CKINVDCx14_ASAP7_75t_R g1061 ( 
.A(n_720),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_842),
.Y(n_1062)
);

CKINVDCx20_ASAP7_75t_R g1063 ( 
.A(n_779),
.Y(n_1063)
);

INVxp33_ASAP7_75t_SL g1064 ( 
.A(n_722),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_719),
.Y(n_1065)
);

CKINVDCx16_ASAP7_75t_R g1066 ( 
.A(n_820),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_842),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_842),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_719),
.Y(n_1069)
);

CKINVDCx20_ASAP7_75t_R g1070 ( 
.A(n_837),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_778),
.Y(n_1071)
);

CKINVDCx14_ASAP7_75t_R g1072 ( 
.A(n_768),
.Y(n_1072)
);

INVxp67_ASAP7_75t_L g1073 ( 
.A(n_612),
.Y(n_1073)
);

CKINVDCx20_ASAP7_75t_R g1074 ( 
.A(n_949),
.Y(n_1074)
);

INVxp67_ASAP7_75t_L g1075 ( 
.A(n_612),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_842),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_778),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_778),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_842),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_888),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_888),
.Y(n_1081)
);

INVxp67_ASAP7_75t_SL g1082 ( 
.A(n_888),
.Y(n_1082)
);

INVxp67_ASAP7_75t_L g1083 ( 
.A(n_620),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_1022),
.Y(n_1084)
);

INVxp67_ASAP7_75t_SL g1085 ( 
.A(n_1022),
.Y(n_1085)
);

CKINVDCx14_ASAP7_75t_R g1086 ( 
.A(n_793),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_842),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_842),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_842),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_890),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_890),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_890),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_890),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_890),
.Y(n_1094)
);

INVxp67_ASAP7_75t_L g1095 ( 
.A(n_620),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_890),
.Y(n_1096)
);

INVxp67_ASAP7_75t_SL g1097 ( 
.A(n_1022),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_890),
.Y(n_1098)
);

CKINVDCx20_ASAP7_75t_R g1099 ( 
.A(n_590),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_715),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_890),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_890),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_741),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_741),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_1099),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_1074),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_1033),
.Y(n_1107)
);

AND2x4_ASAP7_75t_L g1108 ( 
.A(n_1043),
.B(n_1031),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_1046),
.Y(n_1109)
);

NOR2xp33_ASAP7_75t_L g1110 ( 
.A(n_1039),
.B(n_725),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_1033),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_1072),
.Y(n_1112)
);

INVx2_ASAP7_75t_SL g1113 ( 
.A(n_1043),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_1046),
.Y(n_1114)
);

BUFx6f_ASAP7_75t_L g1115 ( 
.A(n_1046),
.Y(n_1115)
);

INVx3_ASAP7_75t_L g1116 ( 
.A(n_1030),
.Y(n_1116)
);

BUFx6f_ASAP7_75t_L g1117 ( 
.A(n_1046),
.Y(n_1117)
);

BUFx6f_ASAP7_75t_L g1118 ( 
.A(n_1046),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1034),
.Y(n_1119)
);

AND2x4_ASAP7_75t_L g1120 ( 
.A(n_1050),
.B(n_1057),
.Y(n_1120)
);

INVx6_ASAP7_75t_L g1121 ( 
.A(n_1066),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_1034),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_1035),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_1030),
.Y(n_1124)
);

BUFx6f_ASAP7_75t_L g1125 ( 
.A(n_1054),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_1054),
.Y(n_1126)
);

BUFx8_ASAP7_75t_L g1127 ( 
.A(n_1086),
.Y(n_1127)
);

AND2x4_ASAP7_75t_L g1128 ( 
.A(n_1103),
.B(n_661),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_1103),
.B(n_915),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_1104),
.B(n_915),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1035),
.Y(n_1131)
);

OA21x2_ASAP7_75t_L g1132 ( 
.A1(n_1104),
.A2(n_1038),
.B(n_1036),
.Y(n_1132)
);

INVx6_ASAP7_75t_L g1133 ( 
.A(n_1058),
.Y(n_1133)
);

NOR2x1_ASAP7_75t_L g1134 ( 
.A(n_1065),
.B(n_1024),
.Y(n_1134)
);

INVx2_ASAP7_75t_SL g1135 ( 
.A(n_1069),
.Y(n_1135)
);

BUFx2_ASAP7_75t_L g1136 ( 
.A(n_1100),
.Y(n_1136)
);

AND2x2_ASAP7_75t_L g1137 ( 
.A(n_1082),
.B(n_661),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_1079),
.Y(n_1138)
);

AOI22xp5_ASAP7_75t_L g1139 ( 
.A1(n_1060),
.A2(n_615),
.B1(n_625),
.B2(n_600),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_1079),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1036),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_1032),
.Y(n_1142)
);

CKINVDCx11_ASAP7_75t_R g1143 ( 
.A(n_1037),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_1063),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_1085),
.B(n_935),
.Y(n_1145)
);

AND2x4_ASAP7_75t_L g1146 ( 
.A(n_1097),
.B(n_1071),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_1077),
.B(n_935),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_1089),
.Y(n_1148)
);

CKINVDCx6p67_ASAP7_75t_R g1149 ( 
.A(n_1070),
.Y(n_1149)
);

HB1xp67_ASAP7_75t_L g1150 ( 
.A(n_1100),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_1089),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1038),
.Y(n_1152)
);

HB1xp67_ASAP7_75t_L g1153 ( 
.A(n_1042),
.Y(n_1153)
);

BUFx6f_ASAP7_75t_L g1154 ( 
.A(n_1092),
.Y(n_1154)
);

OAI21x1_ASAP7_75t_L g1155 ( 
.A1(n_1092),
.A2(n_948),
.B(n_750),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_1098),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_1098),
.Y(n_1157)
);

AND2x4_ASAP7_75t_L g1158 ( 
.A(n_1078),
.B(n_735),
.Y(n_1158)
);

AND2x4_ASAP7_75t_L g1159 ( 
.A(n_1080),
.B(n_735),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_1040),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1040),
.Y(n_1161)
);

AND2x2_ASAP7_75t_L g1162 ( 
.A(n_1081),
.B(n_1084),
.Y(n_1162)
);

INVx2_ASAP7_75t_SL g1163 ( 
.A(n_1041),
.Y(n_1163)
);

BUFx6f_ASAP7_75t_L g1164 ( 
.A(n_1041),
.Y(n_1164)
);

CKINVDCx20_ASAP7_75t_R g1165 ( 
.A(n_1061),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_1045),
.Y(n_1166)
);

NOR2xp33_ASAP7_75t_R g1167 ( 
.A(n_1112),
.B(n_628),
.Y(n_1167)
);

NOR2x1p5_ASAP7_75t_L g1168 ( 
.A(n_1149),
.B(n_745),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1162),
.Y(n_1169)
);

INVxp67_ASAP7_75t_SL g1170 ( 
.A(n_1113),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_1106),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1162),
.Y(n_1172)
);

AND2x2_ASAP7_75t_L g1173 ( 
.A(n_1120),
.B(n_1073),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_1105),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_1143),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_1127),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_1127),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1162),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_1127),
.Y(n_1179)
);

CKINVDCx8_ASAP7_75t_R g1180 ( 
.A(n_1142),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1135),
.Y(n_1181)
);

NOR2xp33_ASAP7_75t_R g1182 ( 
.A(n_1165),
.B(n_660),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_1127),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_1144),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_1149),
.Y(n_1185)
);

NOR2xp33_ASAP7_75t_SL g1186 ( 
.A(n_1121),
.B(n_1064),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_1149),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_1136),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_1136),
.Y(n_1189)
);

XOR2xp5_ASAP7_75t_L g1190 ( 
.A(n_1139),
.B(n_1044),
.Y(n_1190)
);

INVxp33_ASAP7_75t_L g1191 ( 
.A(n_1153),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1135),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1135),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_1121),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_1121),
.Y(n_1195)
);

CKINVDCx16_ASAP7_75t_R g1196 ( 
.A(n_1150),
.Y(n_1196)
);

NOR2xp33_ASAP7_75t_R g1197 ( 
.A(n_1121),
.B(n_689),
.Y(n_1197)
);

INVx2_ASAP7_75t_SL g1198 ( 
.A(n_1133),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_1121),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_1150),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_1139),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1133),
.B(n_1075),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_1153),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_1133),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1133),
.Y(n_1205)
);

INVx6_ASAP7_75t_L g1206 ( 
.A(n_1133),
.Y(n_1206)
);

INVx2_ASAP7_75t_SL g1207 ( 
.A(n_1108),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_1120),
.Y(n_1208)
);

BUFx10_ASAP7_75t_L g1209 ( 
.A(n_1108),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1116),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_1110),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_1113),
.Y(n_1212)
);

INVx3_ASAP7_75t_L g1213 ( 
.A(n_1132),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_1113),
.Y(n_1214)
);

AND2x2_ASAP7_75t_L g1215 ( 
.A(n_1120),
.B(n_1083),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_1124),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_1137),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_1137),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_1137),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_1120),
.Y(n_1220)
);

OAI21x1_ASAP7_75t_L g1221 ( 
.A1(n_1155),
.A2(n_1047),
.B(n_1045),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1116),
.Y(n_1222)
);

NOR2xp33_ASAP7_75t_R g1223 ( 
.A(n_1116),
.B(n_706),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_1108),
.Y(n_1224)
);

BUFx6f_ASAP7_75t_L g1225 ( 
.A(n_1213),
.Y(n_1225)
);

AND3x1_ASAP7_75t_L g1226 ( 
.A(n_1186),
.B(n_593),
.C(n_591),
.Y(n_1226)
);

BUFx4f_ASAP7_75t_L g1227 ( 
.A(n_1206),
.Y(n_1227)
);

NOR2xp33_ASAP7_75t_L g1228 ( 
.A(n_1211),
.B(n_1108),
.Y(n_1228)
);

AND2x2_ASAP7_75t_L g1229 ( 
.A(n_1173),
.B(n_1146),
.Y(n_1229)
);

AND2x4_ASAP7_75t_L g1230 ( 
.A(n_1194),
.B(n_1195),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1216),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1216),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1210),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1222),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_1184),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1213),
.Y(n_1236)
);

AND2x2_ASAP7_75t_L g1237 ( 
.A(n_1173),
.B(n_1146),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_1213),
.Y(n_1238)
);

NAND3xp33_ASAP7_75t_L g1239 ( 
.A(n_1208),
.B(n_1095),
.C(n_1145),
.Y(n_1239)
);

INVxp67_ASAP7_75t_L g1240 ( 
.A(n_1188),
.Y(n_1240)
);

INVx3_ASAP7_75t_L g1241 ( 
.A(n_1206),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_1221),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1221),
.Y(n_1243)
);

BUFx4f_ASAP7_75t_L g1244 ( 
.A(n_1206),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_1205),
.Y(n_1245)
);

INVx2_ASAP7_75t_L g1246 ( 
.A(n_1181),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1192),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1193),
.Y(n_1248)
);

INVxp67_ASAP7_75t_SL g1249 ( 
.A(n_1198),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1207),
.Y(n_1250)
);

INVx2_ASAP7_75t_SL g1251 ( 
.A(n_1209),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1207),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_1198),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1169),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1172),
.Y(n_1255)
);

OR2x2_ASAP7_75t_L g1256 ( 
.A(n_1196),
.B(n_1203),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1178),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_SL g1258 ( 
.A(n_1208),
.B(n_1146),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1206),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_1171),
.Y(n_1260)
);

INVx3_ASAP7_75t_L g1261 ( 
.A(n_1209),
.Y(n_1261)
);

BUFx2_ASAP7_75t_L g1262 ( 
.A(n_1203),
.Y(n_1262)
);

CKINVDCx5p33_ASAP7_75t_R g1263 ( 
.A(n_1171),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1209),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_1220),
.Y(n_1265)
);

BUFx6f_ASAP7_75t_L g1266 ( 
.A(n_1204),
.Y(n_1266)
);

AND2x2_ASAP7_75t_L g1267 ( 
.A(n_1215),
.B(n_1146),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1220),
.Y(n_1268)
);

INVx2_ASAP7_75t_L g1269 ( 
.A(n_1204),
.Y(n_1269)
);

OR2x2_ASAP7_75t_L g1270 ( 
.A(n_1217),
.B(n_1145),
.Y(n_1270)
);

INVx2_ASAP7_75t_L g1271 ( 
.A(n_1202),
.Y(n_1271)
);

INVx2_ASAP7_75t_SL g1272 ( 
.A(n_1199),
.Y(n_1272)
);

INVx4_ASAP7_75t_L g1273 ( 
.A(n_1224),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1215),
.Y(n_1274)
);

AOI22xp5_ASAP7_75t_L g1275 ( 
.A1(n_1224),
.A2(n_1128),
.B1(n_811),
.B2(n_715),
.Y(n_1275)
);

AND2x4_ASAP7_75t_L g1276 ( 
.A(n_1168),
.B(n_1128),
.Y(n_1276)
);

AO21x2_ASAP7_75t_L g1277 ( 
.A1(n_1223),
.A2(n_1155),
.B(n_1130),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1170),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1212),
.B(n_1163),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1218),
.Y(n_1280)
);

AOI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1219),
.A2(n_1128),
.B1(n_1132),
.B2(n_1134),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1214),
.Y(n_1282)
);

NOR2xp33_ASAP7_75t_L g1283 ( 
.A(n_1191),
.B(n_811),
.Y(n_1283)
);

BUFx6f_ASAP7_75t_L g1284 ( 
.A(n_1176),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_SL g1285 ( 
.A(n_1197),
.B(n_1128),
.Y(n_1285)
);

NAND3xp33_ASAP7_75t_L g1286 ( 
.A(n_1200),
.B(n_1189),
.C(n_1174),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_1174),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1201),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1201),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1180),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1167),
.B(n_1163),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_1176),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1180),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1177),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1190),
.Y(n_1295)
);

INVx2_ASAP7_75t_L g1296 ( 
.A(n_1179),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1182),
.B(n_1163),
.Y(n_1297)
);

NOR2xp33_ASAP7_75t_L g1298 ( 
.A(n_1183),
.B(n_1158),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1185),
.B(n_1152),
.Y(n_1299)
);

INVx4_ASAP7_75t_L g1300 ( 
.A(n_1187),
.Y(n_1300)
);

BUFx10_ASAP7_75t_L g1301 ( 
.A(n_1175),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_SL g1302 ( 
.A(n_1175),
.B(n_1129),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1229),
.B(n_1129),
.Y(n_1303)
);

AND2x2_ASAP7_75t_SL g1304 ( 
.A(n_1226),
.B(n_1130),
.Y(n_1304)
);

AND2x4_ASAP7_75t_L g1305 ( 
.A(n_1230),
.B(n_1158),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1229),
.B(n_1237),
.Y(n_1306)
);

NOR2xp33_ASAP7_75t_L g1307 ( 
.A(n_1228),
.B(n_1107),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1237),
.B(n_1158),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_1238),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1267),
.B(n_1158),
.Y(n_1310)
);

INVx2_ASAP7_75t_SL g1311 ( 
.A(n_1256),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1267),
.B(n_1159),
.Y(n_1312)
);

NOR2xp33_ASAP7_75t_L g1313 ( 
.A(n_1265),
.B(n_1107),
.Y(n_1313)
);

BUFx12f_ASAP7_75t_L g1314 ( 
.A(n_1301),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_SL g1315 ( 
.A(n_1266),
.B(n_1111),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1269),
.B(n_1159),
.Y(n_1316)
);

OR2x2_ASAP7_75t_L g1317 ( 
.A(n_1256),
.B(n_1159),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1269),
.B(n_1159),
.Y(n_1318)
);

NOR2xp33_ASAP7_75t_SL g1319 ( 
.A(n_1235),
.B(n_627),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1271),
.B(n_1132),
.Y(n_1320)
);

AOI22xp5_ASAP7_75t_L g1321 ( 
.A1(n_1268),
.A2(n_633),
.B1(n_666),
.B2(n_651),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1254),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_SL g1323 ( 
.A(n_1266),
.B(n_1111),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_L g1324 ( 
.A1(n_1274),
.A2(n_755),
.B1(n_774),
.B2(n_684),
.Y(n_1324)
);

AOI22xp5_ASAP7_75t_L g1325 ( 
.A1(n_1268),
.A2(n_786),
.B1(n_808),
.B2(n_801),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1271),
.B(n_1132),
.Y(n_1326)
);

BUFx3_ASAP7_75t_L g1327 ( 
.A(n_1235),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1274),
.B(n_1132),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1270),
.B(n_1147),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1270),
.B(n_1147),
.Y(n_1330)
);

AND2x2_ASAP7_75t_L g1331 ( 
.A(n_1262),
.B(n_864),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1279),
.B(n_1119),
.Y(n_1332)
);

OAI21xp33_ASAP7_75t_L g1333 ( 
.A1(n_1282),
.A2(n_744),
.B(n_614),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_SL g1334 ( 
.A(n_1266),
.B(n_876),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_SL g1335 ( 
.A(n_1266),
.B(n_886),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1266),
.B(n_1119),
.Y(n_1336)
);

NOR2xp33_ASAP7_75t_L g1337 ( 
.A(n_1265),
.B(n_1122),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1272),
.B(n_1122),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1272),
.B(n_1123),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_SL g1340 ( 
.A(n_1230),
.B(n_892),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_SL g1341 ( 
.A(n_1230),
.B(n_901),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1254),
.B(n_1123),
.Y(n_1342)
);

INVx3_ASAP7_75t_L g1343 ( 
.A(n_1227),
.Y(n_1343)
);

CKINVDCx5p33_ASAP7_75t_R g1344 ( 
.A(n_1260),
.Y(n_1344)
);

AOI22xp5_ASAP7_75t_L g1345 ( 
.A1(n_1280),
.A2(n_1273),
.B1(n_1258),
.B2(n_1282),
.Y(n_1345)
);

NAND3xp33_ASAP7_75t_L g1346 ( 
.A(n_1283),
.B(n_1263),
.C(n_1260),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1255),
.B(n_1257),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_SL g1348 ( 
.A(n_1225),
.B(n_1131),
.Y(n_1348)
);

NOR2xp33_ASAP7_75t_L g1349 ( 
.A(n_1280),
.B(n_1131),
.Y(n_1349)
);

INVx3_ASAP7_75t_L g1350 ( 
.A(n_1227),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_SL g1351 ( 
.A(n_1225),
.B(n_1227),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1255),
.B(n_1141),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1238),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1231),
.Y(n_1354)
);

A2O1A1Ixp33_ASAP7_75t_L g1355 ( 
.A1(n_1250),
.A2(n_1155),
.B(n_1141),
.C(n_1152),
.Y(n_1355)
);

AOI221xp5_ASAP7_75t_L g1356 ( 
.A1(n_1262),
.A2(n_918),
.B1(n_909),
.B2(n_1010),
.C(n_912),
.Y(n_1356)
);

AOI22xp5_ASAP7_75t_L g1357 ( 
.A1(n_1273),
.A2(n_665),
.B1(n_670),
.B2(n_601),
.Y(n_1357)
);

NAND3xp33_ASAP7_75t_L g1358 ( 
.A(n_1263),
.B(n_896),
.C(n_644),
.Y(n_1358)
);

INVx2_ASAP7_75t_SL g1359 ( 
.A(n_1287),
.Y(n_1359)
);

AOI22xp33_ASAP7_75t_L g1360 ( 
.A1(n_1257),
.A2(n_653),
.B1(n_748),
.B2(n_624),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1250),
.B(n_1161),
.Y(n_1361)
);

NOR2xp33_ASAP7_75t_L g1362 ( 
.A(n_1273),
.B(n_1161),
.Y(n_1362)
);

INVx1_ASAP7_75t_SL g1363 ( 
.A(n_1287),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1233),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_SL g1365 ( 
.A(n_1225),
.B(n_1160),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1231),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1252),
.B(n_1160),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1233),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1252),
.B(n_1160),
.Y(n_1369)
);

NOR3xp33_ASAP7_75t_L g1370 ( 
.A(n_1286),
.B(n_1012),
.C(n_723),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1264),
.B(n_1166),
.Y(n_1371)
);

NOR2xp33_ASAP7_75t_L g1372 ( 
.A(n_1239),
.B(n_1164),
.Y(n_1372)
);

AND2x4_ASAP7_75t_L g1373 ( 
.A(n_1276),
.B(n_1134),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1234),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1234),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_SL g1376 ( 
.A(n_1251),
.B(n_1291),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1264),
.B(n_1166),
.Y(n_1377)
);

BUFx2_ASAP7_75t_L g1378 ( 
.A(n_1240),
.Y(n_1378)
);

NOR2xp33_ASAP7_75t_L g1379 ( 
.A(n_1299),
.B(n_1164),
.Y(n_1379)
);

INVx3_ASAP7_75t_L g1380 ( 
.A(n_1244),
.Y(n_1380)
);

AOI22xp33_ASAP7_75t_L g1381 ( 
.A1(n_1281),
.A2(n_653),
.B1(n_748),
.B2(n_624),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1246),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1251),
.B(n_1261),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_1232),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1246),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_SL g1386 ( 
.A(n_1261),
.B(n_1164),
.Y(n_1386)
);

BUFx6f_ASAP7_75t_L g1387 ( 
.A(n_1225),
.Y(n_1387)
);

NOR2xp33_ASAP7_75t_L g1388 ( 
.A(n_1288),
.B(n_1164),
.Y(n_1388)
);

NOR2xp33_ASAP7_75t_L g1389 ( 
.A(n_1288),
.B(n_1164),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1289),
.B(n_671),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1261),
.B(n_1166),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1278),
.B(n_1116),
.Y(n_1392)
);

INVx2_ASAP7_75t_SL g1393 ( 
.A(n_1284),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_SL g1394 ( 
.A(n_1297),
.B(n_1164),
.Y(n_1394)
);

AOI22xp5_ASAP7_75t_L g1395 ( 
.A1(n_1298),
.A2(n_737),
.B1(n_747),
.B2(n_714),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1247),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_SL g1397 ( 
.A(n_1284),
.B(n_589),
.Y(n_1397)
);

INVx2_ASAP7_75t_L g1398 ( 
.A(n_1232),
.Y(n_1398)
);

NOR2xp67_ASAP7_75t_L g1399 ( 
.A(n_1300),
.B(n_948),
.Y(n_1399)
);

HB1xp67_ASAP7_75t_L g1400 ( 
.A(n_1276),
.Y(n_1400)
);

CKINVDCx5p33_ASAP7_75t_R g1401 ( 
.A(n_1301),
.Y(n_1401)
);

INVx4_ASAP7_75t_L g1402 ( 
.A(n_1244),
.Y(n_1402)
);

OR2x2_ASAP7_75t_SL g1403 ( 
.A(n_1284),
.B(n_595),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1278),
.B(n_1148),
.Y(n_1404)
);

AOI22xp5_ASAP7_75t_L g1405 ( 
.A1(n_1285),
.A2(n_1293),
.B1(n_1290),
.B2(n_1276),
.Y(n_1405)
);

AOI21xp5_ASAP7_75t_L g1406 ( 
.A1(n_1307),
.A2(n_1362),
.B(n_1365),
.Y(n_1406)
);

NOR2xp33_ASAP7_75t_SL g1407 ( 
.A(n_1344),
.B(n_1300),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1331),
.B(n_1289),
.Y(n_1408)
);

AOI21xp5_ASAP7_75t_L g1409 ( 
.A1(n_1307),
.A2(n_1243),
.B(n_1242),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1329),
.B(n_1275),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1330),
.B(n_1284),
.Y(n_1411)
);

BUFx2_ASAP7_75t_L g1412 ( 
.A(n_1378),
.Y(n_1412)
);

INVx3_ASAP7_75t_L g1413 ( 
.A(n_1402),
.Y(n_1413)
);

AOI21xp5_ASAP7_75t_L g1414 ( 
.A1(n_1362),
.A2(n_1243),
.B(n_1242),
.Y(n_1414)
);

AOI21xp5_ASAP7_75t_L g1415 ( 
.A1(n_1336),
.A2(n_1249),
.B(n_1236),
.Y(n_1415)
);

AOI21xp5_ASAP7_75t_L g1416 ( 
.A1(n_1365),
.A2(n_1236),
.B(n_1225),
.Y(n_1416)
);

INVx2_ASAP7_75t_SL g1417 ( 
.A(n_1327),
.Y(n_1417)
);

AOI21xp5_ASAP7_75t_L g1418 ( 
.A1(n_1379),
.A2(n_1244),
.B(n_1247),
.Y(n_1418)
);

BUFx3_ASAP7_75t_L g1419 ( 
.A(n_1314),
.Y(n_1419)
);

OR2x6_ASAP7_75t_L g1420 ( 
.A(n_1311),
.B(n_1284),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1322),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1303),
.B(n_1292),
.Y(n_1422)
);

OAI22xp5_ASAP7_75t_L g1423 ( 
.A1(n_1306),
.A2(n_1248),
.B1(n_1253),
.B2(n_1292),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_SL g1424 ( 
.A(n_1327),
.B(n_1359),
.Y(n_1424)
);

AOI21xp5_ASAP7_75t_L g1425 ( 
.A1(n_1379),
.A2(n_1361),
.B(n_1332),
.Y(n_1425)
);

AND2x4_ASAP7_75t_L g1426 ( 
.A(n_1305),
.B(n_1290),
.Y(n_1426)
);

NOR2xp33_ASAP7_75t_L g1427 ( 
.A(n_1363),
.B(n_1293),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_SL g1428 ( 
.A(n_1346),
.B(n_1300),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1390),
.B(n_1294),
.Y(n_1429)
);

BUFx4f_ASAP7_75t_L g1430 ( 
.A(n_1314),
.Y(n_1430)
);

NOR2xp33_ASAP7_75t_L g1431 ( 
.A(n_1334),
.B(n_1302),
.Y(n_1431)
);

O2A1O1Ixp33_ASAP7_75t_SL g1432 ( 
.A1(n_1315),
.A2(n_1248),
.B(n_1259),
.C(n_1253),
.Y(n_1432)
);

AOI21xp5_ASAP7_75t_L g1433 ( 
.A1(n_1391),
.A2(n_1277),
.B(n_1259),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1304),
.B(n_1296),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1304),
.B(n_1349),
.Y(n_1435)
);

NOR2xp33_ASAP7_75t_SL g1436 ( 
.A(n_1319),
.B(n_1301),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1349),
.B(n_1296),
.Y(n_1437)
);

AOI21xp5_ASAP7_75t_L g1438 ( 
.A1(n_1342),
.A2(n_1277),
.B(n_1245),
.Y(n_1438)
);

NOR2xp33_ASAP7_75t_L g1439 ( 
.A(n_1335),
.B(n_1294),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1308),
.B(n_1295),
.Y(n_1440)
);

NOR2xp33_ASAP7_75t_L g1441 ( 
.A(n_1321),
.B(n_1295),
.Y(n_1441)
);

AOI21xp33_ASAP7_75t_L g1442 ( 
.A1(n_1395),
.A2(n_1245),
.B(n_1241),
.Y(n_1442)
);

AOI21xp5_ASAP7_75t_L g1443 ( 
.A1(n_1352),
.A2(n_1277),
.B(n_1241),
.Y(n_1443)
);

AOI21xp5_ASAP7_75t_L g1444 ( 
.A1(n_1367),
.A2(n_1369),
.B(n_1348),
.Y(n_1444)
);

AOI21xp5_ASAP7_75t_L g1445 ( 
.A1(n_1348),
.A2(n_1241),
.B(n_1126),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1310),
.B(n_846),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_SL g1447 ( 
.A(n_1402),
.B(n_592),
.Y(n_1447)
);

OAI21xp5_ASAP7_75t_L g1448 ( 
.A1(n_1328),
.A2(n_1157),
.B(n_1156),
.Y(n_1448)
);

AOI21xp5_ASAP7_75t_L g1449 ( 
.A1(n_1351),
.A2(n_1126),
.B(n_1124),
.Y(n_1449)
);

AOI22xp5_ASAP7_75t_L g1450 ( 
.A1(n_1356),
.A2(n_882),
.B1(n_907),
.B2(n_880),
.Y(n_1450)
);

AOI21xp5_ASAP7_75t_L g1451 ( 
.A1(n_1351),
.A2(n_1126),
.B(n_1124),
.Y(n_1451)
);

AND2x4_ASAP7_75t_L g1452 ( 
.A(n_1305),
.B(n_591),
.Y(n_1452)
);

AOI21xp5_ASAP7_75t_L g1453 ( 
.A1(n_1315),
.A2(n_1140),
.B(n_1138),
.Y(n_1453)
);

AOI33xp33_ASAP7_75t_L g1454 ( 
.A1(n_1360),
.A2(n_596),
.A3(n_594),
.B1(n_605),
.B2(n_598),
.B3(n_593),
.Y(n_1454)
);

AOI21xp5_ASAP7_75t_L g1455 ( 
.A1(n_1355),
.A2(n_1140),
.B(n_1138),
.Y(n_1455)
);

AND2x4_ASAP7_75t_L g1456 ( 
.A(n_1400),
.B(n_594),
.Y(n_1456)
);

NOR2xp33_ASAP7_75t_L g1457 ( 
.A(n_1325),
.B(n_923),
.Y(n_1457)
);

AOI22xp5_ASAP7_75t_L g1458 ( 
.A1(n_1324),
.A2(n_1002),
.B1(n_597),
.B2(n_603),
.Y(n_1458)
);

AOI21xp5_ASAP7_75t_L g1459 ( 
.A1(n_1323),
.A2(n_1140),
.B(n_1138),
.Y(n_1459)
);

OR2x2_ASAP7_75t_L g1460 ( 
.A(n_1317),
.B(n_833),
.Y(n_1460)
);

AOI22xp5_ASAP7_75t_L g1461 ( 
.A1(n_1324),
.A2(n_604),
.B1(n_606),
.B2(n_602),
.Y(n_1461)
);

HB1xp67_ASAP7_75t_L g1462 ( 
.A(n_1373),
.Y(n_1462)
);

AOI21xp5_ASAP7_75t_L g1463 ( 
.A1(n_1323),
.A2(n_1151),
.B(n_1148),
.Y(n_1463)
);

AOI21xp5_ASAP7_75t_L g1464 ( 
.A1(n_1371),
.A2(n_1151),
.B(n_1148),
.Y(n_1464)
);

INVxp67_ASAP7_75t_L g1465 ( 
.A(n_1340),
.Y(n_1465)
);

NOR3xp33_ASAP7_75t_L g1466 ( 
.A(n_1358),
.B(n_598),
.C(n_596),
.Y(n_1466)
);

BUFx12f_ASAP7_75t_L g1467 ( 
.A(n_1401),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1312),
.B(n_1151),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_SL g1469 ( 
.A(n_1345),
.B(n_611),
.Y(n_1469)
);

OAI21xp5_ASAP7_75t_L g1470 ( 
.A1(n_1388),
.A2(n_1157),
.B(n_1156),
.Y(n_1470)
);

AOI21xp5_ASAP7_75t_L g1471 ( 
.A1(n_1377),
.A2(n_1157),
.B(n_1156),
.Y(n_1471)
);

AOI22xp33_ASAP7_75t_L g1472 ( 
.A1(n_1381),
.A2(n_675),
.B1(n_676),
.B2(n_671),
.Y(n_1472)
);

HB1xp67_ASAP7_75t_L g1473 ( 
.A(n_1373),
.Y(n_1473)
);

HB1xp67_ASAP7_75t_L g1474 ( 
.A(n_1403),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1396),
.Y(n_1475)
);

AND2x2_ASAP7_75t_SL g1476 ( 
.A(n_1381),
.B(n_610),
.Y(n_1476)
);

AOI21xp5_ASAP7_75t_L g1477 ( 
.A1(n_1347),
.A2(n_1154),
.B(n_1125),
.Y(n_1477)
);

INVxp67_ASAP7_75t_L g1478 ( 
.A(n_1341),
.Y(n_1478)
);

AOI21xp5_ASAP7_75t_L g1479 ( 
.A1(n_1313),
.A2(n_1154),
.B(n_1125),
.Y(n_1479)
);

O2A1O1Ixp5_ASAP7_75t_L g1480 ( 
.A1(n_1397),
.A2(n_609),
.B(n_610),
.C(n_605),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1313),
.B(n_858),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_SL g1482 ( 
.A(n_1357),
.B(n_616),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_SL g1483 ( 
.A(n_1343),
.B(n_617),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1364),
.Y(n_1484)
);

AOI21xp5_ASAP7_75t_L g1485 ( 
.A1(n_1383),
.A2(n_1154),
.B(n_1125),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1337),
.B(n_858),
.Y(n_1486)
);

NOR2xp33_ASAP7_75t_L g1487 ( 
.A(n_1405),
.B(n_619),
.Y(n_1487)
);

BUFx6f_ASAP7_75t_L g1488 ( 
.A(n_1387),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_SL g1489 ( 
.A(n_1343),
.B(n_622),
.Y(n_1489)
);

AOI21xp5_ASAP7_75t_L g1490 ( 
.A1(n_1337),
.A2(n_1154),
.B(n_1125),
.Y(n_1490)
);

CKINVDCx5p33_ASAP7_75t_R g1491 ( 
.A(n_1393),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1368),
.Y(n_1492)
);

INVx3_ASAP7_75t_L g1493 ( 
.A(n_1350),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1360),
.B(n_671),
.Y(n_1494)
);

AOI21xp5_ASAP7_75t_L g1495 ( 
.A1(n_1386),
.A2(n_1339),
.B(n_1338),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1374),
.Y(n_1496)
);

INVx3_ASAP7_75t_L g1497 ( 
.A(n_1350),
.Y(n_1497)
);

AOI21xp5_ASAP7_75t_L g1498 ( 
.A1(n_1320),
.A2(n_1154),
.B(n_1125),
.Y(n_1498)
);

AOI21xp5_ASAP7_75t_L g1499 ( 
.A1(n_1326),
.A2(n_1154),
.B(n_1125),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1375),
.Y(n_1500)
);

AOI21xp5_ASAP7_75t_L g1501 ( 
.A1(n_1387),
.A2(n_1048),
.B(n_1047),
.Y(n_1501)
);

AOI21xp5_ASAP7_75t_L g1502 ( 
.A1(n_1387),
.A2(n_1049),
.B(n_1048),
.Y(n_1502)
);

NOR2xp33_ASAP7_75t_L g1503 ( 
.A(n_1333),
.B(n_623),
.Y(n_1503)
);

BUFx12f_ASAP7_75t_L g1504 ( 
.A(n_1467),
.Y(n_1504)
);

HB1xp67_ASAP7_75t_L g1505 ( 
.A(n_1412),
.Y(n_1505)
);

AOI21xp5_ASAP7_75t_L g1506 ( 
.A1(n_1414),
.A2(n_1387),
.B(n_1376),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1410),
.B(n_1388),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_SL g1508 ( 
.A(n_1437),
.B(n_1399),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1421),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1475),
.Y(n_1510)
);

INVx3_ASAP7_75t_L g1511 ( 
.A(n_1413),
.Y(n_1511)
);

BUFx3_ASAP7_75t_L g1512 ( 
.A(n_1430),
.Y(n_1512)
);

O2A1O1Ixp33_ASAP7_75t_L g1513 ( 
.A1(n_1435),
.A2(n_1370),
.B(n_1318),
.C(n_1316),
.Y(n_1513)
);

A2O1A1Ixp33_ASAP7_75t_SL g1514 ( 
.A1(n_1495),
.A2(n_1389),
.B(n_1372),
.C(n_613),
.Y(n_1514)
);

OAI22xp5_ASAP7_75t_L g1515 ( 
.A1(n_1406),
.A2(n_1389),
.B1(n_1382),
.B2(n_1385),
.Y(n_1515)
);

OAI22xp5_ASAP7_75t_L g1516 ( 
.A1(n_1476),
.A2(n_1406),
.B1(n_1422),
.B2(n_1481),
.Y(n_1516)
);

INVx11_ASAP7_75t_L g1517 ( 
.A(n_1430),
.Y(n_1517)
);

NOR2xp33_ASAP7_75t_L g1518 ( 
.A(n_1427),
.B(n_1372),
.Y(n_1518)
);

O2A1O1Ixp5_ASAP7_75t_L g1519 ( 
.A1(n_1469),
.A2(n_1394),
.B(n_1353),
.C(n_1309),
.Y(n_1519)
);

NOR2xp33_ASAP7_75t_L g1520 ( 
.A(n_1426),
.B(n_1354),
.Y(n_1520)
);

AND2x6_ASAP7_75t_L g1521 ( 
.A(n_1413),
.B(n_1354),
.Y(n_1521)
);

AOI21xp5_ASAP7_75t_L g1522 ( 
.A1(n_1414),
.A2(n_1353),
.B(n_1309),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_SL g1523 ( 
.A(n_1436),
.B(n_1380),
.Y(n_1523)
);

OAI221xp5_ASAP7_75t_L g1524 ( 
.A1(n_1457),
.A2(n_997),
.B1(n_970),
.B2(n_942),
.C(n_618),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1484),
.Y(n_1525)
);

OR2x6_ASAP7_75t_L g1526 ( 
.A(n_1426),
.B(n_1462),
.Y(n_1526)
);

O2A1O1Ixp33_ASAP7_75t_L g1527 ( 
.A1(n_1434),
.A2(n_970),
.B(n_997),
.C(n_942),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1492),
.Y(n_1528)
);

AOI21x1_ASAP7_75t_L g1529 ( 
.A1(n_1498),
.A2(n_1499),
.B(n_1438),
.Y(n_1529)
);

AOI21xp5_ASAP7_75t_L g1530 ( 
.A1(n_1409),
.A2(n_1404),
.B(n_1392),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1496),
.Y(n_1531)
);

OAI22xp5_ASAP7_75t_L g1532 ( 
.A1(n_1411),
.A2(n_1380),
.B1(n_1384),
.B2(n_1366),
.Y(n_1532)
);

OAI22xp5_ASAP7_75t_L g1533 ( 
.A1(n_1487),
.A2(n_1366),
.B1(n_1398),
.B2(n_1384),
.Y(n_1533)
);

CKINVDCx5p33_ASAP7_75t_R g1534 ( 
.A(n_1419),
.Y(n_1534)
);

AND2x4_ASAP7_75t_L g1535 ( 
.A(n_1473),
.B(n_1398),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1500),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1440),
.B(n_632),
.Y(n_1537)
);

AND2x4_ASAP7_75t_L g1538 ( 
.A(n_1417),
.B(n_609),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_SL g1539 ( 
.A(n_1407),
.B(n_671),
.Y(n_1539)
);

XOR2xp5_ASAP7_75t_L g1540 ( 
.A(n_1474),
.B(n_634),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1408),
.B(n_635),
.Y(n_1541)
);

AND2x4_ASAP7_75t_L g1542 ( 
.A(n_1420),
.B(n_1491),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_SL g1543 ( 
.A(n_1439),
.B(n_1429),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1441),
.B(n_636),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1456),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1456),
.Y(n_1546)
);

NOR2xp33_ASAP7_75t_L g1547 ( 
.A(n_1431),
.B(n_637),
.Y(n_1547)
);

NOR2xp33_ASAP7_75t_L g1548 ( 
.A(n_1465),
.B(n_638),
.Y(n_1548)
);

OAI21xp5_ASAP7_75t_L g1549 ( 
.A1(n_1409),
.A2(n_1051),
.B(n_1049),
.Y(n_1549)
);

NOR2xp33_ASAP7_75t_L g1550 ( 
.A(n_1478),
.B(n_1482),
.Y(n_1550)
);

NAND3xp33_ASAP7_75t_L g1551 ( 
.A(n_1503),
.B(n_849),
.C(n_772),
.Y(n_1551)
);

BUFx6f_ASAP7_75t_L g1552 ( 
.A(n_1488),
.Y(n_1552)
);

CKINVDCx5p33_ASAP7_75t_R g1553 ( 
.A(n_1424),
.Y(n_1553)
);

AOI21xp5_ASAP7_75t_L g1554 ( 
.A1(n_1425),
.A2(n_750),
.B(n_1109),
.Y(n_1554)
);

INVx5_ASAP7_75t_L g1555 ( 
.A(n_1420),
.Y(n_1555)
);

AOI21xp5_ASAP7_75t_L g1556 ( 
.A1(n_1418),
.A2(n_1114),
.B(n_1109),
.Y(n_1556)
);

OAI22xp5_ASAP7_75t_L g1557 ( 
.A1(n_1486),
.A2(n_1460),
.B1(n_1423),
.B2(n_1472),
.Y(n_1557)
);

BUFx3_ASAP7_75t_L g1558 ( 
.A(n_1420),
.Y(n_1558)
);

AOI21xp5_ASAP7_75t_L g1559 ( 
.A1(n_1443),
.A2(n_1114),
.B(n_1109),
.Y(n_1559)
);

OR2x2_ASAP7_75t_L g1560 ( 
.A(n_1452),
.B(n_833),
.Y(n_1560)
);

OR2x2_ASAP7_75t_L g1561 ( 
.A(n_1452),
.B(n_745),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1454),
.Y(n_1562)
);

BUFx6f_ASAP7_75t_L g1563 ( 
.A(n_1488),
.Y(n_1563)
);

AOI21xp5_ASAP7_75t_L g1564 ( 
.A1(n_1498),
.A2(n_1114),
.B(n_599),
.Y(n_1564)
);

NOR2xp33_ASAP7_75t_L g1565 ( 
.A(n_1446),
.B(n_639),
.Y(n_1565)
);

O2A1O1Ixp33_ASAP7_75t_L g1566 ( 
.A1(n_1428),
.A2(n_618),
.B(n_626),
.C(n_613),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1494),
.B(n_641),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_SL g1568 ( 
.A(n_1493),
.B(n_675),
.Y(n_1568)
);

INVx3_ASAP7_75t_L g1569 ( 
.A(n_1488),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1450),
.B(n_645),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1468),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_SL g1572 ( 
.A(n_1493),
.B(n_675),
.Y(n_1572)
);

INVx4_ASAP7_75t_L g1573 ( 
.A(n_1497),
.Y(n_1573)
);

NOR2xp33_ASAP7_75t_L g1574 ( 
.A(n_1458),
.B(n_646),
.Y(n_1574)
);

AOI21xp5_ASAP7_75t_L g1575 ( 
.A1(n_1499),
.A2(n_599),
.B(n_595),
.Y(n_1575)
);

AOI21xp5_ASAP7_75t_L g1576 ( 
.A1(n_1479),
.A2(n_621),
.B(n_608),
.Y(n_1576)
);

NOR2xp33_ASAP7_75t_L g1577 ( 
.A(n_1461),
.B(n_648),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1480),
.Y(n_1578)
);

AOI21x1_ASAP7_75t_L g1579 ( 
.A1(n_1455),
.A2(n_1052),
.B(n_1051),
.Y(n_1579)
);

AND2x4_ASAP7_75t_L g1580 ( 
.A(n_1497),
.B(n_626),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1466),
.B(n_675),
.Y(n_1581)
);

OAI21xp33_ASAP7_75t_SL g1582 ( 
.A1(n_1483),
.A2(n_630),
.B(n_629),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1432),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_SL g1584 ( 
.A(n_1442),
.B(n_676),
.Y(n_1584)
);

OAI21xp33_ASAP7_75t_L g1585 ( 
.A1(n_1447),
.A2(n_815),
.B(n_679),
.Y(n_1585)
);

INVx1_ASAP7_75t_SL g1586 ( 
.A(n_1489),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_SL g1587 ( 
.A(n_1415),
.B(n_676),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1448),
.Y(n_1588)
);

NOR2xp33_ASAP7_75t_L g1589 ( 
.A(n_1501),
.B(n_649),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1470),
.Y(n_1590)
);

HB1xp67_ASAP7_75t_L g1591 ( 
.A(n_1501),
.Y(n_1591)
);

CKINVDCx5p33_ASAP7_75t_R g1592 ( 
.A(n_1502),
.Y(n_1592)
);

NOR2xp33_ASAP7_75t_R g1593 ( 
.A(n_1502),
.B(n_676),
.Y(n_1593)
);

NOR2xp33_ASAP7_75t_L g1594 ( 
.A(n_1445),
.B(n_652),
.Y(n_1594)
);

NOR2xp33_ASAP7_75t_L g1595 ( 
.A(n_1449),
.B(n_663),
.Y(n_1595)
);

BUFx2_ASAP7_75t_L g1596 ( 
.A(n_1490),
.Y(n_1596)
);

HB1xp67_ASAP7_75t_L g1597 ( 
.A(n_1479),
.Y(n_1597)
);

A2O1A1Ixp33_ASAP7_75t_L g1598 ( 
.A1(n_1444),
.A2(n_815),
.B(n_630),
.C(n_631),
.Y(n_1598)
);

CKINVDCx20_ASAP7_75t_R g1599 ( 
.A(n_1451),
.Y(n_1599)
);

OA21x2_ASAP7_75t_L g1600 ( 
.A1(n_1433),
.A2(n_1053),
.B(n_1052),
.Y(n_1600)
);

INVx3_ASAP7_75t_L g1601 ( 
.A(n_1416),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_SL g1602 ( 
.A(n_1453),
.B(n_707),
.Y(n_1602)
);

INVx2_ASAP7_75t_L g1603 ( 
.A(n_1459),
.Y(n_1603)
);

AOI21xp5_ASAP7_75t_L g1604 ( 
.A1(n_1477),
.A2(n_621),
.B(n_608),
.Y(n_1604)
);

NAND3xp33_ASAP7_75t_L g1605 ( 
.A(n_1455),
.B(n_849),
.C(n_772),
.Y(n_1605)
);

NAND2x1p5_ASAP7_75t_L g1606 ( 
.A(n_1555),
.B(n_1485),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1509),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1518),
.B(n_629),
.Y(n_1608)
);

OA21x2_ASAP7_75t_L g1609 ( 
.A1(n_1529),
.A2(n_1471),
.B(n_1464),
.Y(n_1609)
);

NOR2xp33_ASAP7_75t_L g1610 ( 
.A(n_1547),
.B(n_664),
.Y(n_1610)
);

OAI21x1_ASAP7_75t_L g1611 ( 
.A1(n_1559),
.A2(n_1463),
.B(n_1055),
.Y(n_1611)
);

CKINVDCx11_ASAP7_75t_R g1612 ( 
.A(n_1504),
.Y(n_1612)
);

NAND2xp33_ASAP7_75t_R g1613 ( 
.A(n_1534),
.B(n_827),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1507),
.B(n_631),
.Y(n_1614)
);

AO31x2_ASAP7_75t_L g1615 ( 
.A1(n_1515),
.A2(n_1530),
.A3(n_1588),
.B(n_1522),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1510),
.Y(n_1616)
);

A2O1A1Ixp33_ASAP7_75t_L g1617 ( 
.A1(n_1574),
.A2(n_643),
.B(n_647),
.C(n_640),
.Y(n_1617)
);

OAI21xp5_ASAP7_75t_L g1618 ( 
.A1(n_1516),
.A2(n_643),
.B(n_640),
.Y(n_1618)
);

A2O1A1Ixp33_ASAP7_75t_L g1619 ( 
.A1(n_1577),
.A2(n_647),
.B(n_654),
.C(n_650),
.Y(n_1619)
);

OAI21xp5_ASAP7_75t_L g1620 ( 
.A1(n_1516),
.A2(n_654),
.B(n_650),
.Y(n_1620)
);

NOR2xp33_ASAP7_75t_L g1621 ( 
.A(n_1505),
.B(n_667),
.Y(n_1621)
);

OAI22xp5_ASAP7_75t_L g1622 ( 
.A1(n_1544),
.A2(n_655),
.B1(n_662),
.B2(n_657),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1525),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1571),
.B(n_655),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1528),
.B(n_657),
.Y(n_1625)
);

OAI21x1_ASAP7_75t_L g1626 ( 
.A1(n_1579),
.A2(n_1506),
.B(n_1601),
.Y(n_1626)
);

OAI21x1_ASAP7_75t_L g1627 ( 
.A1(n_1601),
.A2(n_1055),
.B(n_1053),
.Y(n_1627)
);

NAND3x1_ASAP7_75t_L g1628 ( 
.A(n_1550),
.B(n_673),
.C(n_662),
.Y(n_1628)
);

AOI21xp5_ASAP7_75t_L g1629 ( 
.A1(n_1597),
.A2(n_656),
.B(n_642),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1531),
.Y(n_1630)
);

A2O1A1Ixp33_ASAP7_75t_L g1631 ( 
.A1(n_1589),
.A2(n_677),
.B(n_682),
.C(n_673),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1536),
.Y(n_1632)
);

OA21x2_ASAP7_75t_L g1633 ( 
.A1(n_1605),
.A2(n_1059),
.B(n_1056),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1535),
.Y(n_1634)
);

OA21x2_ASAP7_75t_L g1635 ( 
.A1(n_1605),
.A2(n_1059),
.B(n_1056),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_SL g1636 ( 
.A(n_1592),
.B(n_707),
.Y(n_1636)
);

BUFx6f_ASAP7_75t_L g1637 ( 
.A(n_1512),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1535),
.Y(n_1638)
);

AOI21x1_ASAP7_75t_L g1639 ( 
.A1(n_1596),
.A2(n_682),
.B(n_677),
.Y(n_1639)
);

AOI21xp5_ASAP7_75t_L g1640 ( 
.A1(n_1514),
.A2(n_1583),
.B(n_1549),
.Y(n_1640)
);

BUFx12f_ASAP7_75t_L g1641 ( 
.A(n_1553),
.Y(n_1641)
);

NOR2xp33_ASAP7_75t_L g1642 ( 
.A(n_1586),
.B(n_668),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1543),
.Y(n_1643)
);

BUFx2_ASAP7_75t_L g1644 ( 
.A(n_1542),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1546),
.Y(n_1645)
);

AOI21xp5_ASAP7_75t_L g1646 ( 
.A1(n_1549),
.A2(n_656),
.B(n_642),
.Y(n_1646)
);

INVx3_ASAP7_75t_SL g1647 ( 
.A(n_1542),
.Y(n_1647)
);

OAI21x1_ASAP7_75t_L g1648 ( 
.A1(n_1564),
.A2(n_1067),
.B(n_1062),
.Y(n_1648)
);

BUFx10_ASAP7_75t_L g1649 ( 
.A(n_1580),
.Y(n_1649)
);

AO31x2_ASAP7_75t_L g1650 ( 
.A1(n_1533),
.A2(n_785),
.A3(n_791),
.B(n_659),
.Y(n_1650)
);

AND2x4_ASAP7_75t_L g1651 ( 
.A(n_1526),
.B(n_687),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1520),
.B(n_687),
.Y(n_1652)
);

OAI21xp5_ASAP7_75t_L g1653 ( 
.A1(n_1513),
.A2(n_690),
.B(n_688),
.Y(n_1653)
);

AOI21xp5_ASAP7_75t_L g1654 ( 
.A1(n_1590),
.A2(n_785),
.B(n_659),
.Y(n_1654)
);

OAI21xp5_ASAP7_75t_L g1655 ( 
.A1(n_1557),
.A2(n_690),
.B(n_688),
.Y(n_1655)
);

INVx4_ASAP7_75t_L g1656 ( 
.A(n_1517),
.Y(n_1656)
);

INVx2_ASAP7_75t_SL g1657 ( 
.A(n_1538),
.Y(n_1657)
);

BUFx4_ASAP7_75t_SL g1658 ( 
.A(n_1560),
.Y(n_1658)
);

AOI21xp5_ASAP7_75t_L g1659 ( 
.A1(n_1532),
.A2(n_803),
.B(n_791),
.Y(n_1659)
);

A2O1A1Ixp33_ASAP7_75t_L g1660 ( 
.A1(n_1565),
.A2(n_697),
.B(n_699),
.C(n_695),
.Y(n_1660)
);

OAI21x1_ASAP7_75t_L g1661 ( 
.A1(n_1554),
.A2(n_1603),
.B(n_1556),
.Y(n_1661)
);

NOR4xp25_ASAP7_75t_L g1662 ( 
.A(n_1524),
.B(n_1557),
.C(n_1527),
.D(n_1566),
.Y(n_1662)
);

NAND2x1p5_ASAP7_75t_L g1663 ( 
.A(n_1555),
.B(n_695),
.Y(n_1663)
);

OAI21x1_ASAP7_75t_L g1664 ( 
.A1(n_1575),
.A2(n_1067),
.B(n_1062),
.Y(n_1664)
);

NAND3xp33_ASAP7_75t_L g1665 ( 
.A(n_1598),
.B(n_699),
.C(n_697),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1580),
.Y(n_1666)
);

AOI21xp5_ASAP7_75t_L g1667 ( 
.A1(n_1508),
.A2(n_829),
.B(n_803),
.Y(n_1667)
);

OAI21x1_ASAP7_75t_L g1668 ( 
.A1(n_1600),
.A2(n_1076),
.B(n_1068),
.Y(n_1668)
);

INVx3_ASAP7_75t_L g1669 ( 
.A(n_1552),
.Y(n_1669)
);

OAI21x1_ASAP7_75t_L g1670 ( 
.A1(n_1600),
.A2(n_1519),
.B(n_1604),
.Y(n_1670)
);

OAI21x1_ASAP7_75t_L g1671 ( 
.A1(n_1576),
.A2(n_1076),
.B(n_1068),
.Y(n_1671)
);

INVxp67_ASAP7_75t_SL g1672 ( 
.A(n_1591),
.Y(n_1672)
);

NOR4xp25_ASAP7_75t_L g1673 ( 
.A(n_1562),
.B(n_708),
.C(n_717),
.D(n_713),
.Y(n_1673)
);

OAI21x1_ASAP7_75t_SL g1674 ( 
.A1(n_1573),
.A2(n_899),
.B(n_829),
.Y(n_1674)
);

AOI21xp5_ASAP7_75t_L g1675 ( 
.A1(n_1587),
.A2(n_931),
.B(n_899),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1538),
.B(n_707),
.Y(n_1676)
);

AO21x2_ASAP7_75t_L g1677 ( 
.A1(n_1551),
.A2(n_713),
.B(n_708),
.Y(n_1677)
);

AOI211x1_ASAP7_75t_L g1678 ( 
.A1(n_1541),
.A2(n_721),
.B(n_726),
.C(n_717),
.Y(n_1678)
);

OAI21x1_ASAP7_75t_L g1679 ( 
.A1(n_1602),
.A2(n_1088),
.B(n_1087),
.Y(n_1679)
);

AOI21xp5_ASAP7_75t_L g1680 ( 
.A1(n_1551),
.A2(n_932),
.B(n_931),
.Y(n_1680)
);

AOI21x1_ASAP7_75t_L g1681 ( 
.A1(n_1584),
.A2(n_726),
.B(n_721),
.Y(n_1681)
);

OR2x2_ASAP7_75t_L g1682 ( 
.A(n_1545),
.B(n_736),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1555),
.B(n_736),
.Y(n_1683)
);

NOR2xp67_ASAP7_75t_L g1684 ( 
.A(n_1569),
.B(n_565),
.Y(n_1684)
);

OAI21x1_ASAP7_75t_SL g1685 ( 
.A1(n_1573),
.A2(n_940),
.B(n_932),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1558),
.Y(n_1686)
);

AO22x2_ASAP7_75t_L g1687 ( 
.A1(n_1540),
.A2(n_762),
.B1(n_764),
.B2(n_758),
.Y(n_1687)
);

NOR2xp33_ASAP7_75t_L g1688 ( 
.A(n_1586),
.B(n_669),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1607),
.B(n_1569),
.Y(n_1689)
);

INVx3_ASAP7_75t_L g1690 ( 
.A(n_1626),
.Y(n_1690)
);

OAI21x1_ASAP7_75t_L g1691 ( 
.A1(n_1670),
.A2(n_1578),
.B(n_1511),
.Y(n_1691)
);

O2A1O1Ixp33_ASAP7_75t_L g1692 ( 
.A1(n_1610),
.A2(n_1567),
.B(n_1539),
.C(n_1570),
.Y(n_1692)
);

INVx2_ASAP7_75t_L g1693 ( 
.A(n_1615),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1616),
.Y(n_1694)
);

OAI21x1_ASAP7_75t_L g1695 ( 
.A1(n_1661),
.A2(n_1511),
.B(n_1523),
.Y(n_1695)
);

A2O1A1Ixp33_ASAP7_75t_L g1696 ( 
.A1(n_1655),
.A2(n_1585),
.B(n_1594),
.C(n_1595),
.Y(n_1696)
);

AOI22xp33_ASAP7_75t_L g1697 ( 
.A1(n_1687),
.A2(n_1581),
.B1(n_1593),
.B2(n_1561),
.Y(n_1697)
);

OAI21x1_ASAP7_75t_L g1698 ( 
.A1(n_1668),
.A2(n_1572),
.B(n_1568),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1630),
.B(n_1552),
.Y(n_1699)
);

INVx3_ASAP7_75t_L g1700 ( 
.A(n_1609),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1615),
.Y(n_1701)
);

OAI22xp5_ASAP7_75t_L g1702 ( 
.A1(n_1655),
.A2(n_1537),
.B1(n_1599),
.B2(n_762),
.Y(n_1702)
);

AOI22xp33_ASAP7_75t_L g1703 ( 
.A1(n_1687),
.A2(n_1526),
.B1(n_1582),
.B2(n_1548),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1643),
.B(n_1521),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1632),
.Y(n_1705)
);

INVx1_ASAP7_75t_SL g1706 ( 
.A(n_1644),
.Y(n_1706)
);

BUFx2_ASAP7_75t_L g1707 ( 
.A(n_1672),
.Y(n_1707)
);

AO21x2_ASAP7_75t_L g1708 ( 
.A1(n_1618),
.A2(n_764),
.B(n_758),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1623),
.Y(n_1709)
);

OAI21x1_ASAP7_75t_L g1710 ( 
.A1(n_1606),
.A2(n_1088),
.B(n_1087),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1615),
.Y(n_1711)
);

AO21x2_ASAP7_75t_L g1712 ( 
.A1(n_1618),
.A2(n_770),
.B(n_767),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1620),
.B(n_1552),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1650),
.Y(n_1714)
);

OAI21x1_ASAP7_75t_SL g1715 ( 
.A1(n_1620),
.A2(n_971),
.B(n_940),
.Y(n_1715)
);

INVx2_ASAP7_75t_L g1716 ( 
.A(n_1609),
.Y(n_1716)
);

OAI21x1_ASAP7_75t_L g1717 ( 
.A1(n_1606),
.A2(n_1091),
.B(n_1090),
.Y(n_1717)
);

INVx4_ASAP7_75t_L g1718 ( 
.A(n_1647),
.Y(n_1718)
);

AOI21x1_ASAP7_75t_L g1719 ( 
.A1(n_1639),
.A2(n_770),
.B(n_767),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1650),
.Y(n_1720)
);

AND2x4_ASAP7_75t_L g1721 ( 
.A(n_1669),
.B(n_1563),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1650),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1651),
.B(n_1563),
.Y(n_1723)
);

OR2x2_ASAP7_75t_L g1724 ( 
.A(n_1608),
.B(n_1683),
.Y(n_1724)
);

AND2x6_ASAP7_75t_L g1725 ( 
.A(n_1634),
.B(n_1563),
.Y(n_1725)
);

OA21x2_ASAP7_75t_L g1726 ( 
.A1(n_1640),
.A2(n_773),
.B(n_771),
.Y(n_1726)
);

AOI21xp33_ASAP7_75t_SL g1727 ( 
.A1(n_1673),
.A2(n_773),
.B(n_771),
.Y(n_1727)
);

OAI21x1_ASAP7_75t_L g1728 ( 
.A1(n_1627),
.A2(n_1091),
.B(n_1090),
.Y(n_1728)
);

BUFx6f_ASAP7_75t_L g1729 ( 
.A(n_1633),
.Y(n_1729)
);

NAND3xp33_ASAP7_75t_L g1730 ( 
.A(n_1653),
.B(n_782),
.C(n_777),
.Y(n_1730)
);

AO31x2_ASAP7_75t_L g1731 ( 
.A1(n_1629),
.A2(n_980),
.A3(n_981),
.B(n_971),
.Y(n_1731)
);

A2O1A1Ixp33_ASAP7_75t_L g1732 ( 
.A1(n_1653),
.A2(n_782),
.B(n_783),
.C(n_777),
.Y(n_1732)
);

OAI21x1_ASAP7_75t_L g1733 ( 
.A1(n_1611),
.A2(n_1094),
.B(n_1093),
.Y(n_1733)
);

OA21x2_ASAP7_75t_L g1734 ( 
.A1(n_1659),
.A2(n_787),
.B(n_783),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1651),
.B(n_787),
.Y(n_1735)
);

AO32x2_ASAP7_75t_L g1736 ( 
.A1(n_1622),
.A2(n_1521),
.A3(n_1526),
.B1(n_712),
.B2(n_769),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1638),
.Y(n_1737)
);

AND2x4_ASAP7_75t_L g1738 ( 
.A(n_1669),
.B(n_1521),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1625),
.Y(n_1739)
);

INVx3_ASAP7_75t_L g1740 ( 
.A(n_1633),
.Y(n_1740)
);

AOI22xp33_ASAP7_75t_L g1741 ( 
.A1(n_1622),
.A2(n_709),
.B1(n_712),
.B2(n_707),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1645),
.Y(n_1742)
);

BUFx3_ASAP7_75t_L g1743 ( 
.A(n_1686),
.Y(n_1743)
);

OA21x2_ASAP7_75t_L g1744 ( 
.A1(n_1654),
.A2(n_796),
.B(n_794),
.Y(n_1744)
);

OAI21x1_ASAP7_75t_L g1745 ( 
.A1(n_1648),
.A2(n_1094),
.B(n_1093),
.Y(n_1745)
);

OAI22xp5_ASAP7_75t_L g1746 ( 
.A1(n_1665),
.A2(n_1678),
.B1(n_1631),
.B2(n_1628),
.Y(n_1746)
);

OAI21x1_ASAP7_75t_L g1747 ( 
.A1(n_1664),
.A2(n_1101),
.B(n_1096),
.Y(n_1747)
);

A2O1A1Ixp33_ASAP7_75t_L g1748 ( 
.A1(n_1642),
.A2(n_796),
.B(n_798),
.C(n_794),
.Y(n_1748)
);

AND2x4_ASAP7_75t_L g1749 ( 
.A(n_1743),
.B(n_1666),
.Y(n_1749)
);

BUFx6f_ASAP7_75t_L g1750 ( 
.A(n_1738),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1742),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1694),
.B(n_1625),
.Y(n_1752)
);

INVx2_ASAP7_75t_L g1753 ( 
.A(n_1742),
.Y(n_1753)
);

A2O1A1Ixp33_ASAP7_75t_L g1754 ( 
.A1(n_1696),
.A2(n_1688),
.B(n_1636),
.C(n_1619),
.Y(n_1754)
);

NAND2xp33_ASAP7_75t_SL g1755 ( 
.A(n_1718),
.B(n_1656),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1694),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1705),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1705),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1707),
.B(n_1614),
.Y(n_1759)
);

AO21x2_ASAP7_75t_L g1760 ( 
.A1(n_1714),
.A2(n_1673),
.B(n_1646),
.Y(n_1760)
);

INVx2_ASAP7_75t_L g1761 ( 
.A(n_1716),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1709),
.Y(n_1762)
);

A2O1A1Ixp33_ASAP7_75t_L g1763 ( 
.A1(n_1692),
.A2(n_1617),
.B(n_1660),
.C(n_1614),
.Y(n_1763)
);

INVx2_ASAP7_75t_L g1764 ( 
.A(n_1716),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1709),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1706),
.B(n_1624),
.Y(n_1766)
);

OAI22x1_ASAP7_75t_L g1767 ( 
.A1(n_1724),
.A2(n_1663),
.B1(n_1657),
.B2(n_1683),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1706),
.B(n_1624),
.Y(n_1768)
);

OAI21x1_ASAP7_75t_L g1769 ( 
.A1(n_1700),
.A2(n_1635),
.B(n_1671),
.Y(n_1769)
);

NAND2x1p5_ASAP7_75t_L g1770 ( 
.A(n_1707),
.B(n_1635),
.Y(n_1770)
);

AOI21xp5_ASAP7_75t_L g1771 ( 
.A1(n_1730),
.A2(n_1662),
.B(n_1665),
.Y(n_1771)
);

OAI21x1_ASAP7_75t_L g1772 ( 
.A1(n_1700),
.A2(n_1679),
.B(n_1680),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1737),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1724),
.B(n_1652),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1737),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1714),
.Y(n_1776)
);

INVx4_ASAP7_75t_SL g1777 ( 
.A(n_1725),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1699),
.B(n_1689),
.Y(n_1778)
);

NOR2xp33_ASAP7_75t_L g1779 ( 
.A(n_1718),
.B(n_1641),
.Y(n_1779)
);

AO31x2_ASAP7_75t_L g1780 ( 
.A1(n_1722),
.A2(n_1667),
.A3(n_1675),
.B(n_1652),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1720),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1716),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1720),
.Y(n_1783)
);

AOI21xp5_ASAP7_75t_L g1784 ( 
.A1(n_1730),
.A2(n_1662),
.B(n_1677),
.Y(n_1784)
);

BUFx6f_ASAP7_75t_L g1785 ( 
.A(n_1738),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1742),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1739),
.B(n_1621),
.Y(n_1787)
);

AO21x2_ASAP7_75t_L g1788 ( 
.A1(n_1722),
.A2(n_1685),
.B(n_1674),
.Y(n_1788)
);

INVx2_ASAP7_75t_L g1789 ( 
.A(n_1693),
.Y(n_1789)
);

OAI21x1_ASAP7_75t_L g1790 ( 
.A1(n_1700),
.A2(n_1681),
.B(n_1663),
.Y(n_1790)
);

OAI21xp5_ASAP7_75t_L g1791 ( 
.A1(n_1702),
.A2(n_867),
.B(n_857),
.Y(n_1791)
);

OAI22xp5_ASAP7_75t_L g1792 ( 
.A1(n_1702),
.A2(n_1637),
.B1(n_1682),
.B2(n_798),
.Y(n_1792)
);

INVx2_ASAP7_75t_L g1793 ( 
.A(n_1693),
.Y(n_1793)
);

OAI21xp5_ASAP7_75t_L g1794 ( 
.A1(n_1732),
.A2(n_1748),
.B(n_1727),
.Y(n_1794)
);

AO21x2_ASAP7_75t_L g1795 ( 
.A1(n_1722),
.A2(n_1677),
.B(n_1684),
.Y(n_1795)
);

BUFx2_ASAP7_75t_L g1796 ( 
.A(n_1743),
.Y(n_1796)
);

BUFx8_ASAP7_75t_L g1797 ( 
.A(n_1736),
.Y(n_1797)
);

HB1xp67_ASAP7_75t_L g1798 ( 
.A(n_1756),
.Y(n_1798)
);

BUFx3_ASAP7_75t_L g1799 ( 
.A(n_1796),
.Y(n_1799)
);

NAND2x1p5_ASAP7_75t_L g1800 ( 
.A(n_1796),
.B(n_1740),
.Y(n_1800)
);

INVx2_ASAP7_75t_L g1801 ( 
.A(n_1761),
.Y(n_1801)
);

INVx2_ASAP7_75t_L g1802 ( 
.A(n_1761),
.Y(n_1802)
);

BUFx6f_ASAP7_75t_L g1803 ( 
.A(n_1761),
.Y(n_1803)
);

INVx2_ASAP7_75t_SL g1804 ( 
.A(n_1750),
.Y(n_1804)
);

OR2x2_ASAP7_75t_L g1805 ( 
.A(n_1759),
.B(n_1711),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1756),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1764),
.Y(n_1807)
);

INVx2_ASAP7_75t_L g1808 ( 
.A(n_1764),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1757),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1757),
.Y(n_1810)
);

INVx2_ASAP7_75t_L g1811 ( 
.A(n_1764),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1758),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1758),
.Y(n_1813)
);

OAI21xp5_ASAP7_75t_L g1814 ( 
.A1(n_1771),
.A2(n_1746),
.B(n_1727),
.Y(n_1814)
);

OAI21xp5_ASAP7_75t_SL g1815 ( 
.A1(n_1754),
.A2(n_1697),
.B(n_1703),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1773),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1759),
.B(n_1752),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1752),
.B(n_1711),
.Y(n_1818)
);

AO21x2_ASAP7_75t_L g1819 ( 
.A1(n_1782),
.A2(n_1701),
.B(n_1693),
.Y(n_1819)
);

AND2x4_ASAP7_75t_L g1820 ( 
.A(n_1777),
.B(n_1690),
.Y(n_1820)
);

INVx2_ASAP7_75t_L g1821 ( 
.A(n_1782),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1773),
.Y(n_1822)
);

OAI21xp5_ASAP7_75t_L g1823 ( 
.A1(n_1784),
.A2(n_1746),
.B(n_1726),
.Y(n_1823)
);

OAI21x1_ASAP7_75t_L g1824 ( 
.A1(n_1769),
.A2(n_1700),
.B(n_1690),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1775),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1782),
.Y(n_1826)
);

INVx2_ASAP7_75t_L g1827 ( 
.A(n_1789),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_L g1828 ( 
.A(n_1775),
.B(n_1739),
.Y(n_1828)
);

OAI21x1_ASAP7_75t_L g1829 ( 
.A1(n_1769),
.A2(n_1690),
.B(n_1691),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1762),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1766),
.B(n_1701),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1762),
.Y(n_1832)
);

HB1xp67_ASAP7_75t_L g1833 ( 
.A(n_1778),
.Y(n_1833)
);

INVx3_ASAP7_75t_L g1834 ( 
.A(n_1750),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1778),
.B(n_1701),
.Y(n_1835)
);

HB1xp67_ASAP7_75t_L g1836 ( 
.A(n_1765),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1765),
.Y(n_1837)
);

INVx2_ASAP7_75t_L g1838 ( 
.A(n_1789),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1776),
.Y(n_1839)
);

BUFx2_ASAP7_75t_L g1840 ( 
.A(n_1750),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1776),
.Y(n_1841)
);

OR2x2_ASAP7_75t_L g1842 ( 
.A(n_1768),
.B(n_1743),
.Y(n_1842)
);

HB1xp67_ASAP7_75t_L g1843 ( 
.A(n_1781),
.Y(n_1843)
);

BUFx2_ASAP7_75t_L g1844 ( 
.A(n_1750),
.Y(n_1844)
);

AO21x2_ASAP7_75t_L g1845 ( 
.A1(n_1789),
.A2(n_1704),
.B(n_1691),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1781),
.Y(n_1846)
);

INVx2_ASAP7_75t_L g1847 ( 
.A(n_1793),
.Y(n_1847)
);

AND2x4_ASAP7_75t_L g1848 ( 
.A(n_1777),
.B(n_1750),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1783),
.Y(n_1849)
);

INVx2_ASAP7_75t_L g1850 ( 
.A(n_1793),
.Y(n_1850)
);

HB1xp67_ASAP7_75t_L g1851 ( 
.A(n_1783),
.Y(n_1851)
);

INVx2_ASAP7_75t_L g1852 ( 
.A(n_1803),
.Y(n_1852)
);

OAI211xp5_ASAP7_75t_SL g1853 ( 
.A1(n_1814),
.A2(n_1787),
.B(n_812),
.C(n_813),
.Y(n_1853)
);

AOI22xp33_ASAP7_75t_L g1854 ( 
.A1(n_1823),
.A2(n_1797),
.B1(n_1814),
.B2(n_1708),
.Y(n_1854)
);

BUFx3_ASAP7_75t_L g1855 ( 
.A(n_1842),
.Y(n_1855)
);

AOI22xp33_ASAP7_75t_L g1856 ( 
.A1(n_1823),
.A2(n_1797),
.B1(n_1708),
.B2(n_1712),
.Y(n_1856)
);

NAND3xp33_ASAP7_75t_L g1857 ( 
.A(n_1815),
.B(n_1797),
.C(n_1791),
.Y(n_1857)
);

BUFx3_ASAP7_75t_L g1858 ( 
.A(n_1842),
.Y(n_1858)
);

OAI22xp33_ASAP7_75t_L g1859 ( 
.A1(n_1815),
.A2(n_1767),
.B1(n_1817),
.B2(n_1726),
.Y(n_1859)
);

OR2x6_ASAP7_75t_L g1860 ( 
.A(n_1848),
.B(n_1785),
.Y(n_1860)
);

AOI221xp5_ASAP7_75t_SL g1861 ( 
.A1(n_1817),
.A2(n_812),
.B1(n_814),
.B2(n_813),
.C(n_805),
.Y(n_1861)
);

AOI22xp5_ASAP7_75t_L g1862 ( 
.A1(n_1831),
.A2(n_1797),
.B1(n_1767),
.B2(n_1792),
.Y(n_1862)
);

AOI22xp33_ASAP7_75t_L g1863 ( 
.A1(n_1831),
.A2(n_1708),
.B1(n_1712),
.B2(n_1726),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1843),
.Y(n_1864)
);

OAI21x1_ASAP7_75t_L g1865 ( 
.A1(n_1824),
.A2(n_1793),
.B(n_1690),
.Y(n_1865)
);

OAI21x1_ASAP7_75t_L g1866 ( 
.A1(n_1824),
.A2(n_1770),
.B(n_1772),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1798),
.Y(n_1867)
);

INVx3_ASAP7_75t_L g1868 ( 
.A(n_1799),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1843),
.Y(n_1869)
);

AOI22xp33_ASAP7_75t_L g1870 ( 
.A1(n_1805),
.A2(n_1708),
.B1(n_1712),
.B2(n_1726),
.Y(n_1870)
);

OAI22xp33_ASAP7_75t_L g1871 ( 
.A1(n_1842),
.A2(n_1785),
.B1(n_1794),
.B2(n_1774),
.Y(n_1871)
);

OAI21x1_ASAP7_75t_L g1872 ( 
.A1(n_1824),
.A2(n_1770),
.B(n_1772),
.Y(n_1872)
);

OAI221xp5_ASAP7_75t_L g1873 ( 
.A1(n_1818),
.A2(n_1763),
.B1(n_1741),
.B2(n_821),
.C(n_825),
.Y(n_1873)
);

AOI222xp33_ASAP7_75t_L g1874 ( 
.A1(n_1818),
.A2(n_1735),
.B1(n_1676),
.B2(n_825),
.C1(n_814),
.C2(n_830),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1833),
.B(n_1689),
.Y(n_1875)
);

CKINVDCx8_ASAP7_75t_R g1876 ( 
.A(n_1848),
.Y(n_1876)
);

AND2x4_ASAP7_75t_L g1877 ( 
.A(n_1848),
.B(n_1777),
.Y(n_1877)
);

AOI222xp33_ASAP7_75t_L g1878 ( 
.A1(n_1828),
.A2(n_1735),
.B1(n_831),
.B2(n_821),
.C1(n_835),
.C2(n_830),
.Y(n_1878)
);

AND2x2_ASAP7_75t_L g1879 ( 
.A(n_1833),
.B(n_1749),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1798),
.Y(n_1880)
);

AND2x4_ASAP7_75t_L g1881 ( 
.A(n_1848),
.B(n_1777),
.Y(n_1881)
);

OAI21x1_ASAP7_75t_L g1882 ( 
.A1(n_1829),
.A2(n_1770),
.B(n_1790),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1851),
.Y(n_1883)
);

INVx2_ASAP7_75t_L g1884 ( 
.A(n_1865),
.Y(n_1884)
);

OR2x2_ASAP7_75t_L g1885 ( 
.A(n_1864),
.B(n_1805),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_L g1886 ( 
.A(n_1867),
.B(n_1836),
.Y(n_1886)
);

OR2x2_ASAP7_75t_L g1887 ( 
.A(n_1864),
.B(n_1869),
.Y(n_1887)
);

INVx2_ASAP7_75t_L g1888 ( 
.A(n_1865),
.Y(n_1888)
);

OR2x2_ASAP7_75t_L g1889 ( 
.A(n_1869),
.B(n_1805),
.Y(n_1889)
);

INVx2_ASAP7_75t_L g1890 ( 
.A(n_1855),
.Y(n_1890)
);

INVx2_ASAP7_75t_L g1891 ( 
.A(n_1855),
.Y(n_1891)
);

AND2x2_ASAP7_75t_L g1892 ( 
.A(n_1879),
.B(n_1799),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1883),
.Y(n_1893)
);

INVxp67_ASAP7_75t_SL g1894 ( 
.A(n_1859),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_L g1895 ( 
.A(n_1880),
.B(n_1836),
.Y(n_1895)
);

BUFx3_ASAP7_75t_L g1896 ( 
.A(n_1876),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1883),
.B(n_1851),
.Y(n_1897)
);

AOI22xp33_ASAP7_75t_L g1898 ( 
.A1(n_1853),
.A2(n_1712),
.B1(n_1760),
.B2(n_1713),
.Y(n_1898)
);

OAI21xp5_ASAP7_75t_L g1899 ( 
.A1(n_1857),
.A2(n_831),
.B(n_805),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1875),
.Y(n_1900)
);

INVx2_ASAP7_75t_L g1901 ( 
.A(n_1858),
.Y(n_1901)
);

INVx2_ASAP7_75t_L g1902 ( 
.A(n_1858),
.Y(n_1902)
);

AND2x2_ASAP7_75t_L g1903 ( 
.A(n_1879),
.B(n_1799),
.Y(n_1903)
);

INVx2_ASAP7_75t_L g1904 ( 
.A(n_1852),
.Y(n_1904)
);

INVx2_ASAP7_75t_L g1905 ( 
.A(n_1852),
.Y(n_1905)
);

INVx2_ASAP7_75t_SL g1906 ( 
.A(n_1868),
.Y(n_1906)
);

HB1xp67_ASAP7_75t_L g1907 ( 
.A(n_1868),
.Y(n_1907)
);

INVxp67_ASAP7_75t_SL g1908 ( 
.A(n_1868),
.Y(n_1908)
);

CKINVDCx20_ASAP7_75t_R g1909 ( 
.A(n_1876),
.Y(n_1909)
);

INVx2_ASAP7_75t_L g1910 ( 
.A(n_1866),
.Y(n_1910)
);

INVx2_ASAP7_75t_L g1911 ( 
.A(n_1866),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1871),
.Y(n_1912)
);

AND2x2_ASAP7_75t_L g1913 ( 
.A(n_1860),
.B(n_1799),
.Y(n_1913)
);

AND2x2_ASAP7_75t_L g1914 ( 
.A(n_1860),
.B(n_1800),
.Y(n_1914)
);

INVxp67_ASAP7_75t_L g1915 ( 
.A(n_1896),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1887),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1887),
.Y(n_1917)
);

AND2x2_ASAP7_75t_L g1918 ( 
.A(n_1896),
.B(n_1860),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1887),
.Y(n_1919)
);

AND2x4_ASAP7_75t_L g1920 ( 
.A(n_1896),
.B(n_1877),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1893),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1893),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1885),
.Y(n_1923)
);

HB1xp67_ASAP7_75t_L g1924 ( 
.A(n_1890),
.Y(n_1924)
);

AND2x2_ASAP7_75t_L g1925 ( 
.A(n_1896),
.B(n_1860),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1894),
.B(n_1861),
.Y(n_1926)
);

AND2x4_ASAP7_75t_L g1927 ( 
.A(n_1909),
.B(n_1877),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1885),
.Y(n_1928)
);

NAND3xp33_ASAP7_75t_L g1929 ( 
.A(n_1894),
.B(n_1854),
.C(n_1878),
.Y(n_1929)
);

AND2x2_ASAP7_75t_L g1930 ( 
.A(n_1913),
.B(n_1877),
.Y(n_1930)
);

AND2x2_ASAP7_75t_L g1931 ( 
.A(n_1913),
.B(n_1881),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_L g1932 ( 
.A(n_1900),
.B(n_1828),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1885),
.Y(n_1933)
);

OR2x2_ASAP7_75t_L g1934 ( 
.A(n_1900),
.B(n_1806),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1889),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1889),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_SL g1937 ( 
.A(n_1909),
.B(n_1881),
.Y(n_1937)
);

BUFx2_ASAP7_75t_L g1938 ( 
.A(n_1890),
.Y(n_1938)
);

INVx2_ASAP7_75t_L g1939 ( 
.A(n_1884),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1889),
.Y(n_1940)
);

AND2x2_ASAP7_75t_L g1941 ( 
.A(n_1913),
.B(n_1881),
.Y(n_1941)
);

NOR3xp33_ASAP7_75t_L g1942 ( 
.A(n_1899),
.B(n_1873),
.C(n_1882),
.Y(n_1942)
);

NOR2xp33_ASAP7_75t_L g1943 ( 
.A(n_1890),
.B(n_1612),
.Y(n_1943)
);

OAI22xp5_ASAP7_75t_L g1944 ( 
.A1(n_1898),
.A2(n_1856),
.B1(n_1862),
.B2(n_1800),
.Y(n_1944)
);

INVx2_ASAP7_75t_L g1945 ( 
.A(n_1884),
.Y(n_1945)
);

AND2x2_ASAP7_75t_L g1946 ( 
.A(n_1892),
.B(n_1840),
.Y(n_1946)
);

AND2x2_ASAP7_75t_L g1947 ( 
.A(n_1892),
.B(n_1840),
.Y(n_1947)
);

INVx2_ASAP7_75t_L g1948 ( 
.A(n_1938),
.Y(n_1948)
);

AND4x1_ASAP7_75t_L g1949 ( 
.A(n_1942),
.B(n_1899),
.C(n_1874),
.D(n_1779),
.Y(n_1949)
);

NAND2xp5_ASAP7_75t_L g1950 ( 
.A(n_1926),
.B(n_1915),
.Y(n_1950)
);

HB1xp67_ASAP7_75t_L g1951 ( 
.A(n_1924),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_L g1952 ( 
.A(n_1938),
.B(n_1891),
.Y(n_1952)
);

AND2x2_ASAP7_75t_L g1953 ( 
.A(n_1930),
.B(n_1901),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1921),
.Y(n_1954)
);

NAND3xp33_ASAP7_75t_L g1955 ( 
.A(n_1929),
.B(n_844),
.C(n_835),
.Y(n_1955)
);

AOI22xp33_ASAP7_75t_L g1956 ( 
.A1(n_1944),
.A2(n_1912),
.B1(n_1898),
.B2(n_1870),
.Y(n_1956)
);

OR2x6_ASAP7_75t_L g1957 ( 
.A(n_1943),
.B(n_1891),
.Y(n_1957)
);

AND2x2_ASAP7_75t_L g1958 ( 
.A(n_1930),
.B(n_1902),
.Y(n_1958)
);

HB1xp67_ASAP7_75t_L g1959 ( 
.A(n_1916),
.Y(n_1959)
);

AOI22xp5_ASAP7_75t_L g1960 ( 
.A1(n_1927),
.A2(n_1912),
.B1(n_1863),
.B2(n_1760),
.Y(n_1960)
);

INVx2_ASAP7_75t_L g1961 ( 
.A(n_1939),
.Y(n_1961)
);

AND2x2_ASAP7_75t_L g1962 ( 
.A(n_1931),
.B(n_1891),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1921),
.Y(n_1963)
);

OAI21xp5_ASAP7_75t_L g1964 ( 
.A1(n_1918),
.A2(n_1902),
.B(n_1901),
.Y(n_1964)
);

AOI22xp33_ASAP7_75t_L g1965 ( 
.A1(n_1939),
.A2(n_1901),
.B1(n_1902),
.B2(n_1910),
.Y(n_1965)
);

AND2x2_ASAP7_75t_L g1966 ( 
.A(n_1931),
.B(n_1892),
.Y(n_1966)
);

INVx2_ASAP7_75t_L g1967 ( 
.A(n_1945),
.Y(n_1967)
);

INVx3_ASAP7_75t_L g1968 ( 
.A(n_1920),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1922),
.Y(n_1969)
);

BUFx2_ASAP7_75t_L g1970 ( 
.A(n_1920),
.Y(n_1970)
);

OAI31xp33_ASAP7_75t_L g1971 ( 
.A1(n_1918),
.A2(n_1911),
.A3(n_1910),
.B(n_1888),
.Y(n_1971)
);

AOI22xp33_ASAP7_75t_L g1972 ( 
.A1(n_1945),
.A2(n_1910),
.B1(n_1911),
.B2(n_1760),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1922),
.Y(n_1973)
);

OR2x2_ASAP7_75t_L g1974 ( 
.A(n_1923),
.B(n_1897),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1916),
.Y(n_1975)
);

OR2x2_ASAP7_75t_L g1976 ( 
.A(n_1923),
.B(n_1897),
.Y(n_1976)
);

INVx2_ASAP7_75t_SL g1977 ( 
.A(n_1927),
.Y(n_1977)
);

AOI221xp5_ASAP7_75t_L g1978 ( 
.A1(n_1928),
.A2(n_1911),
.B1(n_1888),
.B2(n_1884),
.C(n_845),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1954),
.Y(n_1979)
);

AND2x2_ASAP7_75t_L g1980 ( 
.A(n_1966),
.B(n_1941),
.Y(n_1980)
);

INVx2_ASAP7_75t_SL g1981 ( 
.A(n_1968),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1954),
.Y(n_1982)
);

INVx2_ASAP7_75t_L g1983 ( 
.A(n_1970),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_L g1984 ( 
.A(n_1977),
.B(n_1928),
.Y(n_1984)
);

AND2x2_ASAP7_75t_L g1985 ( 
.A(n_1966),
.B(n_1927),
.Y(n_1985)
);

AND2x2_ASAP7_75t_L g1986 ( 
.A(n_1970),
.B(n_1941),
.Y(n_1986)
);

AND2x2_ASAP7_75t_L g1987 ( 
.A(n_1968),
.B(n_1920),
.Y(n_1987)
);

NAND2xp33_ASAP7_75t_SL g1988 ( 
.A(n_1977),
.B(n_1937),
.Y(n_1988)
);

AND2x2_ASAP7_75t_L g1989 ( 
.A(n_1968),
.B(n_1953),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_L g1990 ( 
.A(n_1950),
.B(n_1933),
.Y(n_1990)
);

AND2x2_ASAP7_75t_L g1991 ( 
.A(n_1968),
.B(n_1933),
.Y(n_1991)
);

OR2x2_ASAP7_75t_L g1992 ( 
.A(n_1974),
.B(n_1935),
.Y(n_1992)
);

NOR3xp33_ASAP7_75t_L g1993 ( 
.A(n_1955),
.B(n_1925),
.C(n_1919),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_L g1994 ( 
.A(n_1951),
.B(n_1935),
.Y(n_1994)
);

INVxp67_ASAP7_75t_SL g1995 ( 
.A(n_1949),
.Y(n_1995)
);

NOR3xp33_ASAP7_75t_SL g1996 ( 
.A(n_1952),
.B(n_1919),
.C(n_1917),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1963),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_L g1998 ( 
.A(n_1949),
.B(n_1936),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1963),
.Y(n_1999)
);

NAND4xp25_ASAP7_75t_L g2000 ( 
.A(n_1948),
.B(n_1917),
.C(n_1940),
.D(n_1936),
.Y(n_2000)
);

OAI211xp5_ASAP7_75t_SL g2001 ( 
.A1(n_1948),
.A2(n_1940),
.B(n_1908),
.C(n_1906),
.Y(n_2001)
);

NOR3xp33_ASAP7_75t_L g2002 ( 
.A(n_1955),
.B(n_1925),
.C(n_1888),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1969),
.Y(n_2003)
);

OAI21xp5_ASAP7_75t_L g2004 ( 
.A1(n_1960),
.A2(n_1978),
.B(n_1964),
.Y(n_2004)
);

AND2x4_ASAP7_75t_L g2005 ( 
.A(n_1957),
.B(n_1946),
.Y(n_2005)
);

OAI21xp5_ASAP7_75t_L g2006 ( 
.A1(n_1960),
.A2(n_1908),
.B(n_1932),
.Y(n_2006)
);

INVx2_ASAP7_75t_L g2007 ( 
.A(n_1948),
.Y(n_2007)
);

NOR3xp33_ASAP7_75t_SL g2008 ( 
.A(n_1975),
.B(n_1755),
.C(n_1886),
.Y(n_2008)
);

INVx2_ASAP7_75t_L g2009 ( 
.A(n_1961),
.Y(n_2009)
);

INVxp67_ASAP7_75t_L g2010 ( 
.A(n_1957),
.Y(n_2010)
);

AND2x2_ASAP7_75t_L g2011 ( 
.A(n_1953),
.B(n_1946),
.Y(n_2011)
);

INVxp67_ASAP7_75t_L g2012 ( 
.A(n_1957),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_L g2013 ( 
.A(n_1958),
.B(n_1934),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1969),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1973),
.Y(n_2015)
);

INVx2_ASAP7_75t_SL g2016 ( 
.A(n_1957),
.Y(n_2016)
);

OR2x2_ASAP7_75t_L g2017 ( 
.A(n_1974),
.B(n_1934),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_L g2018 ( 
.A(n_1958),
.B(n_1962),
.Y(n_2018)
);

NAND4xp25_ASAP7_75t_L g2019 ( 
.A(n_1975),
.B(n_1947),
.C(n_1718),
.D(n_1903),
.Y(n_2019)
);

INVx2_ASAP7_75t_SL g2020 ( 
.A(n_1957),
.Y(n_2020)
);

INVx1_ASAP7_75t_SL g2021 ( 
.A(n_1962),
.Y(n_2021)
);

AND2x2_ASAP7_75t_L g2022 ( 
.A(n_1959),
.B(n_1947),
.Y(n_2022)
);

AND2x2_ASAP7_75t_L g2023 ( 
.A(n_1986),
.B(n_1976),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_2007),
.Y(n_2024)
);

AND2x2_ASAP7_75t_L g2025 ( 
.A(n_1986),
.B(n_1976),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_2007),
.Y(n_2026)
);

INVx2_ASAP7_75t_L g2027 ( 
.A(n_1987),
.Y(n_2027)
);

OR2x2_ASAP7_75t_L g2028 ( 
.A(n_2021),
.B(n_1973),
.Y(n_2028)
);

AND2x2_ASAP7_75t_L g2029 ( 
.A(n_1985),
.B(n_1903),
.Y(n_2029)
);

AND2x2_ASAP7_75t_SL g2030 ( 
.A(n_1998),
.B(n_1656),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_L g2031 ( 
.A(n_1996),
.B(n_1956),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_SL g2032 ( 
.A(n_1988),
.B(n_2016),
.Y(n_2032)
);

NAND2xp5_ASAP7_75t_L g2033 ( 
.A(n_1995),
.B(n_1961),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1983),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1983),
.Y(n_2035)
);

AND2x2_ASAP7_75t_L g2036 ( 
.A(n_1980),
.B(n_1903),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_1979),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_L g2038 ( 
.A(n_1993),
.B(n_1961),
.Y(n_2038)
);

AND2x2_ASAP7_75t_L g2039 ( 
.A(n_1980),
.B(n_1906),
.Y(n_2039)
);

AND2x2_ASAP7_75t_L g2040 ( 
.A(n_1989),
.B(n_1906),
.Y(n_2040)
);

NAND2xp5_ASAP7_75t_L g2041 ( 
.A(n_2000),
.B(n_1991),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_L g2042 ( 
.A(n_1991),
.B(n_1967),
.Y(n_2042)
);

OR2x2_ASAP7_75t_L g2043 ( 
.A(n_2018),
.B(n_1886),
.Y(n_2043)
);

OR2x2_ASAP7_75t_L g2044 ( 
.A(n_2013),
.B(n_1895),
.Y(n_2044)
);

AND2x4_ASAP7_75t_L g2045 ( 
.A(n_1987),
.B(n_1907),
.Y(n_2045)
);

AND2x2_ASAP7_75t_L g2046 ( 
.A(n_1989),
.B(n_1907),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_SL g2047 ( 
.A(n_1988),
.B(n_1965),
.Y(n_2047)
);

INVx1_ASAP7_75t_SL g2048 ( 
.A(n_2016),
.Y(n_2048)
);

OR2x2_ASAP7_75t_L g2049 ( 
.A(n_1984),
.B(n_1895),
.Y(n_2049)
);

INVx2_ASAP7_75t_L g2050 ( 
.A(n_2005),
.Y(n_2050)
);

OR2x2_ASAP7_75t_L g2051 ( 
.A(n_1990),
.B(n_1967),
.Y(n_2051)
);

OR2x2_ASAP7_75t_L g2052 ( 
.A(n_2017),
.B(n_1967),
.Y(n_2052)
);

AND2x2_ASAP7_75t_L g2053 ( 
.A(n_2005),
.B(n_1914),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_1982),
.Y(n_2054)
);

AND2x2_ASAP7_75t_L g2055 ( 
.A(n_2005),
.B(n_1914),
.Y(n_2055)
);

OR2x2_ASAP7_75t_L g2056 ( 
.A(n_1992),
.B(n_1972),
.Y(n_2056)
);

OR2x2_ASAP7_75t_L g2057 ( 
.A(n_1994),
.B(n_1904),
.Y(n_2057)
);

AND2x2_ASAP7_75t_L g2058 ( 
.A(n_2011),
.B(n_1914),
.Y(n_2058)
);

INVx1_ASAP7_75t_SL g2059 ( 
.A(n_2020),
.Y(n_2059)
);

INVx1_ASAP7_75t_SL g2060 ( 
.A(n_2020),
.Y(n_2060)
);

AND2x2_ASAP7_75t_L g2061 ( 
.A(n_2011),
.B(n_1904),
.Y(n_2061)
);

OR2x2_ASAP7_75t_L g2062 ( 
.A(n_2022),
.B(n_1904),
.Y(n_2062)
);

OR2x6_ASAP7_75t_L g2063 ( 
.A(n_2010),
.B(n_1637),
.Y(n_2063)
);

NOR3x1_ASAP7_75t_L g2064 ( 
.A(n_2019),
.B(n_844),
.C(n_840),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_1997),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_L g2066 ( 
.A(n_2022),
.B(n_1971),
.Y(n_2066)
);

NAND2xp5_ASAP7_75t_L g2067 ( 
.A(n_1999),
.B(n_2003),
.Y(n_2067)
);

AND2x2_ASAP7_75t_L g2068 ( 
.A(n_2008),
.B(n_1905),
.Y(n_2068)
);

NAND2xp5_ASAP7_75t_L g2069 ( 
.A(n_2014),
.B(n_840),
.Y(n_2069)
);

AND2x2_ASAP7_75t_L g2070 ( 
.A(n_1981),
.B(n_1905),
.Y(n_2070)
);

AND2x2_ASAP7_75t_L g2071 ( 
.A(n_1981),
.B(n_1905),
.Y(n_2071)
);

AND2x2_ASAP7_75t_L g2072 ( 
.A(n_2012),
.B(n_1718),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_2015),
.Y(n_2073)
);

OR2x2_ASAP7_75t_L g2074 ( 
.A(n_2006),
.B(n_1806),
.Y(n_2074)
);

AND2x4_ASAP7_75t_L g2075 ( 
.A(n_2002),
.B(n_1809),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_2009),
.Y(n_2076)
);

HB1xp67_ASAP7_75t_L g2077 ( 
.A(n_2004),
.Y(n_2077)
);

INVx2_ASAP7_75t_L g2078 ( 
.A(n_2009),
.Y(n_2078)
);

BUFx2_ASAP7_75t_L g2079 ( 
.A(n_2001),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_2007),
.Y(n_2080)
);

NAND2x1p5_ASAP7_75t_L g2081 ( 
.A(n_2016),
.B(n_1637),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_2007),
.Y(n_2082)
);

NAND2xp5_ASAP7_75t_L g2083 ( 
.A(n_1996),
.B(n_845),
.Y(n_2083)
);

OR2x2_ASAP7_75t_L g2084 ( 
.A(n_2021),
.B(n_1809),
.Y(n_2084)
);

NAND2xp5_ASAP7_75t_L g2085 ( 
.A(n_1996),
.B(n_847),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_2007),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_2042),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_2042),
.Y(n_2088)
);

INVx2_ASAP7_75t_SL g2089 ( 
.A(n_2050),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_2052),
.Y(n_2090)
);

O2A1O1Ixp33_ASAP7_75t_L g2091 ( 
.A1(n_2047),
.A2(n_2032),
.B(n_2077),
.C(n_2083),
.Y(n_2091)
);

OAI22xp5_ASAP7_75t_L g2092 ( 
.A1(n_2047),
.A2(n_1800),
.B1(n_1834),
.B2(n_1812),
.Y(n_2092)
);

OAI22xp33_ASAP7_75t_L g2093 ( 
.A1(n_2031),
.A2(n_1803),
.B1(n_1804),
.B2(n_1613),
.Y(n_2093)
);

OAI21xp33_ASAP7_75t_L g2094 ( 
.A1(n_2032),
.A2(n_2041),
.B(n_2031),
.Y(n_2094)
);

AOI21xp33_ASAP7_75t_L g2095 ( 
.A1(n_2077),
.A2(n_981),
.B(n_980),
.Y(n_2095)
);

AOI211x1_ASAP7_75t_L g2096 ( 
.A1(n_2041),
.A2(n_848),
.B(n_854),
.C(n_847),
.Y(n_2096)
);

NAND2xp5_ASAP7_75t_L g2097 ( 
.A(n_2023),
.B(n_848),
.Y(n_2097)
);

NOR2xp33_ASAP7_75t_L g2098 ( 
.A(n_2083),
.B(n_854),
.Y(n_2098)
);

INVx2_ASAP7_75t_L g2099 ( 
.A(n_2036),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_2034),
.Y(n_2100)
);

AOI22xp5_ASAP7_75t_L g2101 ( 
.A1(n_2033),
.A2(n_862),
.B1(n_866),
.B2(n_863),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_2035),
.Y(n_2102)
);

AND2x2_ASAP7_75t_L g2103 ( 
.A(n_2025),
.B(n_1810),
.Y(n_2103)
);

OAI211xp5_ASAP7_75t_SL g2104 ( 
.A1(n_2033),
.A2(n_862),
.B(n_863),
.C(n_857),
.Y(n_2104)
);

INVx2_ASAP7_75t_L g2105 ( 
.A(n_2029),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_2051),
.Y(n_2106)
);

AOI22xp5_ASAP7_75t_L g2107 ( 
.A1(n_2038),
.A2(n_867),
.B1(n_871),
.B2(n_866),
.Y(n_2107)
);

INVx2_ASAP7_75t_L g2108 ( 
.A(n_2027),
.Y(n_2108)
);

INVx2_ASAP7_75t_SL g2109 ( 
.A(n_2046),
.Y(n_2109)
);

INVx2_ASAP7_75t_L g2110 ( 
.A(n_2039),
.Y(n_2110)
);

OAI22xp5_ASAP7_75t_L g2111 ( 
.A1(n_2079),
.A2(n_1800),
.B1(n_1834),
.B2(n_1812),
.Y(n_2111)
);

NAND2xp5_ASAP7_75t_L g2112 ( 
.A(n_2048),
.B(n_871),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_2078),
.Y(n_2113)
);

AOI21xp5_ASAP7_75t_L g2114 ( 
.A1(n_2085),
.A2(n_2066),
.B(n_2038),
.Y(n_2114)
);

INVx2_ASAP7_75t_L g2115 ( 
.A(n_2081),
.Y(n_2115)
);

OAI21xp33_ASAP7_75t_L g2116 ( 
.A1(n_2066),
.A2(n_873),
.B(n_872),
.Y(n_2116)
);

AOI31xp33_ASAP7_75t_L g2117 ( 
.A1(n_2085),
.A2(n_2048),
.A3(n_2060),
.B(n_2059),
.Y(n_2117)
);

AOI22xp5_ASAP7_75t_L g2118 ( 
.A1(n_2024),
.A2(n_885),
.B1(n_891),
.B2(n_872),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_2069),
.Y(n_2119)
);

NAND2xp5_ASAP7_75t_L g2120 ( 
.A(n_2059),
.B(n_873),
.Y(n_2120)
);

NOR2xp33_ASAP7_75t_L g2121 ( 
.A(n_2030),
.B(n_885),
.Y(n_2121)
);

INVxp67_ASAP7_75t_SL g2122 ( 
.A(n_2064),
.Y(n_2122)
);

HB1xp67_ASAP7_75t_L g2123 ( 
.A(n_2060),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_2069),
.Y(n_2124)
);

OR2x2_ASAP7_75t_L g2125 ( 
.A(n_2043),
.B(n_1810),
.Y(n_2125)
);

OAI21xp5_ASAP7_75t_L g2126 ( 
.A1(n_2056),
.A2(n_893),
.B(n_891),
.Y(n_2126)
);

AOI21xp33_ASAP7_75t_SL g2127 ( 
.A1(n_2030),
.A2(n_900),
.B(n_893),
.Y(n_2127)
);

AND2x2_ASAP7_75t_L g2128 ( 
.A(n_2053),
.B(n_1813),
.Y(n_2128)
);

AND2x2_ASAP7_75t_L g2129 ( 
.A(n_2055),
.B(n_1813),
.Y(n_2129)
);

OR2x2_ASAP7_75t_L g2130 ( 
.A(n_2044),
.B(n_1816),
.Y(n_2130)
);

OAI22xp5_ASAP7_75t_L g2131 ( 
.A1(n_2058),
.A2(n_1834),
.B1(n_1816),
.B2(n_1825),
.Y(n_2131)
);

NOR2xp33_ASAP7_75t_L g2132 ( 
.A(n_2028),
.B(n_900),
.Y(n_2132)
);

AOI211xp5_ASAP7_75t_L g2133 ( 
.A1(n_2068),
.A2(n_903),
.B(n_906),
.C(n_902),
.Y(n_2133)
);

OAI21xp33_ASAP7_75t_SL g2134 ( 
.A1(n_2040),
.A2(n_1872),
.B(n_1882),
.Y(n_2134)
);

OAI22xp5_ASAP7_75t_L g2135 ( 
.A1(n_2062),
.A2(n_1834),
.B1(n_1822),
.B2(n_1825),
.Y(n_2135)
);

INVx2_ASAP7_75t_L g2136 ( 
.A(n_2081),
.Y(n_2136)
);

NAND2xp5_ASAP7_75t_SL g2137 ( 
.A(n_2045),
.B(n_1820),
.Y(n_2137)
);

OAI21xp5_ASAP7_75t_L g2138 ( 
.A1(n_2086),
.A2(n_903),
.B(n_902),
.Y(n_2138)
);

INVxp67_ASAP7_75t_L g2139 ( 
.A(n_2072),
.Y(n_2139)
);

NAND2xp5_ASAP7_75t_L g2140 ( 
.A(n_2026),
.B(n_906),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_2080),
.Y(n_2141)
);

INVx2_ASAP7_75t_SL g2142 ( 
.A(n_2045),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_2082),
.Y(n_2143)
);

OAI31xp33_ASAP7_75t_L g2144 ( 
.A1(n_2076),
.A2(n_921),
.A3(n_990),
.B(n_962),
.Y(n_2144)
);

INVx1_ASAP7_75t_L g2145 ( 
.A(n_2067),
.Y(n_2145)
);

INVx1_ASAP7_75t_SL g2146 ( 
.A(n_2049),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_2067),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_2037),
.Y(n_2148)
);

OAI21xp33_ASAP7_75t_SL g2149 ( 
.A1(n_2054),
.A2(n_1872),
.B(n_1822),
.Y(n_2149)
);

OA21x2_ASAP7_75t_L g2150 ( 
.A1(n_2065),
.A2(n_2073),
.B(n_2071),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_2084),
.Y(n_2151)
);

INVx1_ASAP7_75t_SL g2152 ( 
.A(n_2057),
.Y(n_2152)
);

AOI22xp5_ASAP7_75t_L g2153 ( 
.A1(n_2075),
.A2(n_926),
.B1(n_941),
.B2(n_917),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_2075),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_2061),
.Y(n_2155)
);

OAI22xp33_ASAP7_75t_L g2156 ( 
.A1(n_2074),
.A2(n_1803),
.B1(n_1804),
.B2(n_1840),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_2070),
.Y(n_2157)
);

OAI22xp5_ASAP7_75t_L g2158 ( 
.A1(n_2063),
.A2(n_1834),
.B1(n_1830),
.B2(n_1832),
.Y(n_2158)
);

INVx2_ASAP7_75t_L g2159 ( 
.A(n_2063),
.Y(n_2159)
);

AOI21xp5_ASAP7_75t_L g2160 ( 
.A1(n_2063),
.A2(n_921),
.B(n_917),
.Y(n_2160)
);

AOI32xp33_ASAP7_75t_L g2161 ( 
.A1(n_2031),
.A2(n_945),
.A3(n_951),
.B1(n_941),
.B2(n_926),
.Y(n_2161)
);

INVx2_ASAP7_75t_L g2162 ( 
.A(n_2036),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_2042),
.Y(n_2163)
);

AOI32xp33_ASAP7_75t_L g2164 ( 
.A1(n_2031),
.A2(n_952),
.A3(n_953),
.B1(n_951),
.B2(n_945),
.Y(n_2164)
);

OAI322xp33_ASAP7_75t_L g2165 ( 
.A1(n_2047),
.A2(n_960),
.A3(n_968),
.B1(n_978),
.B2(n_952),
.C1(n_956),
.C2(n_961),
.Y(n_2165)
);

OAI21xp33_ASAP7_75t_SL g2166 ( 
.A1(n_2047),
.A2(n_955),
.B(n_953),
.Y(n_2166)
);

INVxp67_ASAP7_75t_L g2167 ( 
.A(n_2032),
.Y(n_2167)
);

AOI22xp33_ASAP7_75t_L g2168 ( 
.A1(n_2077),
.A2(n_1725),
.B1(n_1845),
.B2(n_1744),
.Y(n_2168)
);

HB1xp67_ASAP7_75t_L g2169 ( 
.A(n_2050),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_2042),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_2042),
.Y(n_2171)
);

INVxp67_ASAP7_75t_L g2172 ( 
.A(n_2032),
.Y(n_2172)
);

NAND2xp5_ASAP7_75t_L g2173 ( 
.A(n_2023),
.B(n_955),
.Y(n_2173)
);

OAI22xp33_ASAP7_75t_L g2174 ( 
.A1(n_2117),
.A2(n_1803),
.B1(n_1804),
.B2(n_1844),
.Y(n_2174)
);

INVx2_ASAP7_75t_L g2175 ( 
.A(n_2150),
.Y(n_2175)
);

NAND2xp5_ASAP7_75t_L g2176 ( 
.A(n_2167),
.B(n_956),
.Y(n_2176)
);

OAI21xp5_ASAP7_75t_L g2177 ( 
.A1(n_2172),
.A2(n_974),
.B(n_964),
.Y(n_2177)
);

OAI32xp33_ASAP7_75t_L g2178 ( 
.A1(n_2094),
.A2(n_962),
.A3(n_963),
.B1(n_961),
.B2(n_960),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_2123),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_2150),
.Y(n_2180)
);

NAND2xp5_ASAP7_75t_L g2181 ( 
.A(n_2096),
.B(n_963),
.Y(n_2181)
);

NAND2xp5_ASAP7_75t_L g2182 ( 
.A(n_2146),
.B(n_964),
.Y(n_2182)
);

NAND2xp5_ASAP7_75t_L g2183 ( 
.A(n_2127),
.B(n_966),
.Y(n_2183)
);

OAI21xp33_ASAP7_75t_SL g2184 ( 
.A1(n_2145),
.A2(n_968),
.B(n_966),
.Y(n_2184)
);

OAI21xp5_ASAP7_75t_L g2185 ( 
.A1(n_2091),
.A2(n_983),
.B(n_974),
.Y(n_2185)
);

OAI21xp33_ASAP7_75t_L g2186 ( 
.A1(n_2094),
.A2(n_976),
.B(n_969),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_2169),
.Y(n_2187)
);

INVx1_ASAP7_75t_SL g2188 ( 
.A(n_2152),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_2097),
.Y(n_2189)
);

AOI22xp5_ASAP7_75t_L g2190 ( 
.A1(n_2114),
.A2(n_1699),
.B1(n_976),
.B2(n_978),
.Y(n_2190)
);

OR2x2_ASAP7_75t_L g2191 ( 
.A(n_2090),
.B(n_969),
.Y(n_2191)
);

AOI21xp33_ASAP7_75t_L g2192 ( 
.A1(n_2166),
.A2(n_1017),
.B(n_986),
.Y(n_2192)
);

AOI22xp33_ASAP7_75t_L g2193 ( 
.A1(n_2126),
.A2(n_1725),
.B1(n_1845),
.B2(n_712),
.Y(n_2193)
);

INVx2_ASAP7_75t_L g2194 ( 
.A(n_2089),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_2173),
.Y(n_2195)
);

AND2x2_ASAP7_75t_L g2196 ( 
.A(n_2109),
.B(n_1844),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_2112),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_2120),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_2098),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_2106),
.Y(n_2200)
);

NAND2xp33_ASAP7_75t_SL g2201 ( 
.A(n_2142),
.B(n_672),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_2108),
.Y(n_2202)
);

INVx1_ASAP7_75t_L g2203 ( 
.A(n_2155),
.Y(n_2203)
);

OAI322xp33_ASAP7_75t_L g2204 ( 
.A1(n_2154),
.A2(n_993),
.A3(n_986),
.B1(n_995),
.B2(n_999),
.C1(n_990),
.C2(n_983),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_2118),
.Y(n_2205)
);

OAI21xp5_ASAP7_75t_L g2206 ( 
.A1(n_2101),
.A2(n_995),
.B(n_993),
.Y(n_2206)
);

AND2x2_ASAP7_75t_L g2207 ( 
.A(n_2105),
.B(n_1844),
.Y(n_2207)
);

OAI221xp5_ASAP7_75t_SL g2208 ( 
.A1(n_2134),
.A2(n_1018),
.B1(n_1021),
.B2(n_1015),
.C(n_999),
.Y(n_2208)
);

INVxp67_ASAP7_75t_SL g2209 ( 
.A(n_2121),
.Y(n_2209)
);

NAND2xp5_ASAP7_75t_L g2210 ( 
.A(n_2161),
.B(n_1015),
.Y(n_2210)
);

NAND2xp5_ASAP7_75t_L g2211 ( 
.A(n_2164),
.B(n_1018),
.Y(n_2211)
);

NOR2xp33_ASAP7_75t_L g2212 ( 
.A(n_2165),
.B(n_1021),
.Y(n_2212)
);

AOI22xp5_ASAP7_75t_L g2213 ( 
.A1(n_2104),
.A2(n_712),
.B1(n_769),
.B2(n_709),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_2118),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_2140),
.Y(n_2215)
);

NAND2xp33_ASAP7_75t_L g2216 ( 
.A(n_2110),
.B(n_1023),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_2132),
.Y(n_2217)
);

AOI21xp5_ASAP7_75t_L g2218 ( 
.A1(n_2116),
.A2(n_1025),
.B(n_1023),
.Y(n_2218)
);

INVxp33_ASAP7_75t_L g2219 ( 
.A(n_2099),
.Y(n_2219)
);

INVx2_ASAP7_75t_L g2220 ( 
.A(n_2162),
.Y(n_2220)
);

INVxp67_ASAP7_75t_L g2221 ( 
.A(n_2122),
.Y(n_2221)
);

AOI222xp33_ASAP7_75t_L g2222 ( 
.A1(n_2113),
.A2(n_1027),
.B1(n_1025),
.B2(n_878),
.C1(n_769),
.C2(n_908),
.Y(n_2222)
);

AND2x2_ASAP7_75t_L g2223 ( 
.A(n_2157),
.B(n_2139),
.Y(n_2223)
);

NAND2xp5_ASAP7_75t_L g2224 ( 
.A(n_2087),
.B(n_1027),
.Y(n_2224)
);

NAND2xp5_ASAP7_75t_L g2225 ( 
.A(n_2088),
.B(n_1017),
.Y(n_2225)
);

OAI211xp5_ASAP7_75t_SL g2226 ( 
.A1(n_2163),
.A2(n_769),
.B(n_800),
.C(n_709),
.Y(n_2226)
);

INVx1_ASAP7_75t_SL g2227 ( 
.A(n_2119),
.Y(n_2227)
);

OAI21xp33_ASAP7_75t_L g2228 ( 
.A1(n_2151),
.A2(n_1832),
.B(n_1830),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_2101),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_2153),
.Y(n_2230)
);

OR2x2_ASAP7_75t_L g2231 ( 
.A(n_2170),
.B(n_1837),
.Y(n_2231)
);

OAI22xp33_ASAP7_75t_L g2232 ( 
.A1(n_2107),
.A2(n_1803),
.B1(n_1785),
.B2(n_1837),
.Y(n_2232)
);

OR2x2_ASAP7_75t_L g2233 ( 
.A(n_2171),
.B(n_1839),
.Y(n_2233)
);

INVxp67_ASAP7_75t_L g2234 ( 
.A(n_2159),
.Y(n_2234)
);

NAND2xp5_ASAP7_75t_L g2235 ( 
.A(n_2124),
.B(n_674),
.Y(n_2235)
);

INVx1_ASAP7_75t_L g2236 ( 
.A(n_2153),
.Y(n_2236)
);

AND2x4_ASAP7_75t_L g2237 ( 
.A(n_2100),
.B(n_1839),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_2102),
.Y(n_2238)
);

INVxp67_ASAP7_75t_L g2239 ( 
.A(n_2147),
.Y(n_2239)
);

AOI21xp5_ASAP7_75t_L g2240 ( 
.A1(n_2116),
.A2(n_680),
.B(n_678),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_2141),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_2143),
.Y(n_2242)
);

AND2x2_ASAP7_75t_SL g2243 ( 
.A(n_2148),
.B(n_1658),
.Y(n_2243)
);

OR2x2_ASAP7_75t_L g2244 ( 
.A(n_2130),
.B(n_1841),
.Y(n_2244)
);

AOI22xp5_ASAP7_75t_L g2245 ( 
.A1(n_2107),
.A2(n_1723),
.B1(n_800),
.B2(n_908),
.Y(n_2245)
);

OAI22xp5_ASAP7_75t_L g2246 ( 
.A1(n_2137),
.A2(n_1820),
.B1(n_1846),
.B2(n_1841),
.Y(n_2246)
);

NAND2xp5_ASAP7_75t_L g2247 ( 
.A(n_2133),
.B(n_681),
.Y(n_2247)
);

INVx1_ASAP7_75t_L g2248 ( 
.A(n_2138),
.Y(n_2248)
);

BUFx3_ASAP7_75t_L g2249 ( 
.A(n_2115),
.Y(n_2249)
);

OAI21xp33_ASAP7_75t_L g2250 ( 
.A1(n_2103),
.A2(n_1849),
.B(n_1846),
.Y(n_2250)
);

AOI32xp33_ASAP7_75t_L g2251 ( 
.A1(n_2149),
.A2(n_686),
.A3(n_691),
.B1(n_685),
.B2(n_683),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_2125),
.Y(n_2252)
);

NOR2xp33_ASAP7_75t_L g2253 ( 
.A(n_2136),
.B(n_692),
.Y(n_2253)
);

AOI32xp33_ASAP7_75t_L g2254 ( 
.A1(n_2092),
.A2(n_2111),
.A3(n_2093),
.B1(n_2156),
.B2(n_2158),
.Y(n_2254)
);

OR2x2_ASAP7_75t_L g2255 ( 
.A(n_2128),
.B(n_1849),
.Y(n_2255)
);

AOI22xp33_ASAP7_75t_L g2256 ( 
.A1(n_2168),
.A2(n_1725),
.B1(n_1845),
.B2(n_800),
.Y(n_2256)
);

NAND2xp5_ASAP7_75t_L g2257 ( 
.A(n_2144),
.B(n_693),
.Y(n_2257)
);

OAI32xp33_ASAP7_75t_L g2258 ( 
.A1(n_2129),
.A2(n_700),
.A3(n_701),
.B1(n_696),
.B2(n_694),
.Y(n_2258)
);

O2A1O1Ixp33_ASAP7_75t_L g2259 ( 
.A1(n_2095),
.A2(n_1715),
.B(n_800),
.C(n_878),
.Y(n_2259)
);

AND2x4_ASAP7_75t_L g2260 ( 
.A(n_2160),
.B(n_1820),
.Y(n_2260)
);

AOI22xp5_ASAP7_75t_L g2261 ( 
.A1(n_2135),
.A2(n_878),
.B1(n_908),
.B2(n_709),
.Y(n_2261)
);

AOI221xp5_ASAP7_75t_L g2262 ( 
.A1(n_2131),
.A2(n_705),
.B1(n_710),
.B2(n_704),
.C(n_703),
.Y(n_2262)
);

AOI21xp5_ASAP7_75t_L g2263 ( 
.A1(n_2091),
.A2(n_716),
.B(n_711),
.Y(n_2263)
);

NAND2x1p5_ASAP7_75t_L g2264 ( 
.A(n_2142),
.B(n_1723),
.Y(n_2264)
);

AND2x2_ASAP7_75t_L g2265 ( 
.A(n_2167),
.B(n_1835),
.Y(n_2265)
);

OAI22xp33_ASAP7_75t_L g2266 ( 
.A1(n_2117),
.A2(n_1803),
.B1(n_1785),
.B2(n_1821),
.Y(n_2266)
);

OAI22xp5_ASAP7_75t_L g2267 ( 
.A1(n_2167),
.A2(n_1820),
.B1(n_1848),
.B2(n_1785),
.Y(n_2267)
);

NAND2xp5_ASAP7_75t_L g2268 ( 
.A(n_2167),
.B(n_718),
.Y(n_2268)
);

NAND3xp33_ASAP7_75t_L g2269 ( 
.A(n_2167),
.B(n_727),
.C(n_724),
.Y(n_2269)
);

OAI22xp5_ASAP7_75t_L g2270 ( 
.A1(n_2167),
.A2(n_1820),
.B1(n_1749),
.B2(n_1803),
.Y(n_2270)
);

OAI21xp33_ASAP7_75t_L g2271 ( 
.A1(n_2094),
.A2(n_729),
.B(n_728),
.Y(n_2271)
);

AOI22xp5_ASAP7_75t_L g2272 ( 
.A1(n_2094),
.A2(n_908),
.B1(n_1029),
.B2(n_878),
.Y(n_2272)
);

INVxp67_ASAP7_75t_SL g2273 ( 
.A(n_2167),
.Y(n_2273)
);

OAI22xp5_ASAP7_75t_L g2274 ( 
.A1(n_2167),
.A2(n_1749),
.B1(n_1803),
.B2(n_1835),
.Y(n_2274)
);

AOI322xp5_ASAP7_75t_L g2275 ( 
.A1(n_2094),
.A2(n_1835),
.A3(n_1713),
.B1(n_1821),
.B2(n_1736),
.C1(n_1807),
.C2(n_1802),
.Y(n_2275)
);

O2A1O1Ixp33_ASAP7_75t_L g2276 ( 
.A1(n_2091),
.A2(n_1715),
.B(n_1029),
.C(n_1734),
.Y(n_2276)
);

OR2x2_ASAP7_75t_L g2277 ( 
.A(n_2123),
.B(n_0),
.Y(n_2277)
);

OR2x2_ASAP7_75t_L g2278 ( 
.A(n_2123),
.B(n_0),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_2123),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_2123),
.Y(n_2280)
);

INVxp67_ASAP7_75t_L g2281 ( 
.A(n_2123),
.Y(n_2281)
);

AND2x2_ASAP7_75t_L g2282 ( 
.A(n_2167),
.B(n_730),
.Y(n_2282)
);

OAI31xp33_ASAP7_75t_L g2283 ( 
.A1(n_2094),
.A2(n_1736),
.A3(n_1738),
.B(n_1749),
.Y(n_2283)
);

AOI22xp5_ASAP7_75t_L g2284 ( 
.A1(n_2094),
.A2(n_1029),
.B1(n_1845),
.B2(n_1738),
.Y(n_2284)
);

NAND2xp5_ASAP7_75t_SL g2285 ( 
.A(n_2167),
.B(n_1029),
.Y(n_2285)
);

A2O1A1Ixp33_ASAP7_75t_L g2286 ( 
.A1(n_2091),
.A2(n_732),
.B(n_733),
.C(n_731),
.Y(n_2286)
);

AOI22xp5_ASAP7_75t_L g2287 ( 
.A1(n_2094),
.A2(n_1845),
.B1(n_738),
.B2(n_739),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_2123),
.Y(n_2288)
);

INVxp67_ASAP7_75t_L g2289 ( 
.A(n_2123),
.Y(n_2289)
);

OAI22xp33_ASAP7_75t_L g2290 ( 
.A1(n_2117),
.A2(n_1821),
.B1(n_1734),
.B2(n_1802),
.Y(n_2290)
);

NAND2xp5_ASAP7_75t_L g2291 ( 
.A(n_2167),
.B(n_734),
.Y(n_2291)
);

AOI222xp33_ASAP7_75t_L g2292 ( 
.A1(n_2094),
.A2(n_746),
.B1(n_742),
.B2(n_749),
.C1(n_743),
.C2(n_740),
.Y(n_2292)
);

NAND2xp5_ASAP7_75t_L g2293 ( 
.A(n_2167),
.B(n_751),
.Y(n_2293)
);

OAI21xp5_ASAP7_75t_L g2294 ( 
.A1(n_2167),
.A2(n_753),
.B(n_752),
.Y(n_2294)
);

NAND2xp5_ASAP7_75t_L g2295 ( 
.A(n_2167),
.B(n_754),
.Y(n_2295)
);

INVx1_ASAP7_75t_L g2296 ( 
.A(n_2123),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_2123),
.Y(n_2297)
);

INVx1_ASAP7_75t_L g2298 ( 
.A(n_2123),
.Y(n_2298)
);

AOI321xp33_ASAP7_75t_L g2299 ( 
.A1(n_2091),
.A2(n_1736),
.A3(n_1721),
.B1(n_1821),
.B2(n_1807),
.C(n_1802),
.Y(n_2299)
);

OR2x2_ASAP7_75t_L g2300 ( 
.A(n_2123),
.B(n_1),
.Y(n_2300)
);

OAI32xp33_ASAP7_75t_L g2301 ( 
.A1(n_2167),
.A2(n_759),
.A3(n_760),
.B1(n_757),
.B2(n_756),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_2123),
.Y(n_2302)
);

AOI22xp5_ASAP7_75t_L g2303 ( 
.A1(n_2094),
.A2(n_763),
.B1(n_766),
.B2(n_761),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_2123),
.Y(n_2304)
);

NAND2xp5_ASAP7_75t_L g2305 ( 
.A(n_2167),
.B(n_775),
.Y(n_2305)
);

NAND2xp5_ASAP7_75t_L g2306 ( 
.A(n_2167),
.B(n_776),
.Y(n_2306)
);

O2A1O1Ixp33_ASAP7_75t_L g2307 ( 
.A1(n_2091),
.A2(n_1734),
.B(n_1744),
.C(n_781),
.Y(n_2307)
);

INVx1_ASAP7_75t_L g2308 ( 
.A(n_2123),
.Y(n_2308)
);

AOI22xp5_ASAP7_75t_L g2309 ( 
.A1(n_2094),
.A2(n_780),
.B1(n_788),
.B2(n_784),
.Y(n_2309)
);

AND2x2_ASAP7_75t_L g2310 ( 
.A(n_2167),
.B(n_789),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_2123),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_2123),
.Y(n_2312)
);

OAI32xp33_ASAP7_75t_L g2313 ( 
.A1(n_2167),
.A2(n_795),
.A3(n_797),
.B1(n_792),
.B2(n_790),
.Y(n_2313)
);

BUFx2_ASAP7_75t_L g2314 ( 
.A(n_2123),
.Y(n_2314)
);

INVx2_ASAP7_75t_SL g2315 ( 
.A(n_2169),
.Y(n_2315)
);

NAND2xp5_ASAP7_75t_L g2316 ( 
.A(n_2167),
.B(n_799),
.Y(n_2316)
);

INVx2_ASAP7_75t_L g2317 ( 
.A(n_2150),
.Y(n_2317)
);

INVx2_ASAP7_75t_L g2318 ( 
.A(n_2150),
.Y(n_2318)
);

OAI22xp5_ASAP7_75t_L g2319 ( 
.A1(n_2167),
.A2(n_802),
.B1(n_806),
.B2(n_804),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_2123),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_2123),
.Y(n_2321)
);

INVx2_ASAP7_75t_L g2322 ( 
.A(n_2150),
.Y(n_2322)
);

OAI322xp33_ASAP7_75t_L g2323 ( 
.A1(n_2167),
.A2(n_816),
.A3(n_809),
.B1(n_817),
.B2(n_819),
.C1(n_818),
.C2(n_810),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_2314),
.Y(n_2324)
);

INVxp67_ASAP7_75t_L g2325 ( 
.A(n_2273),
.Y(n_2325)
);

OAI22xp5_ASAP7_75t_L g2326 ( 
.A1(n_2188),
.A2(n_823),
.B1(n_826),
.B2(n_824),
.Y(n_2326)
);

NAND2xp5_ASAP7_75t_L g2327 ( 
.A(n_2315),
.B(n_828),
.Y(n_2327)
);

OR2x2_ASAP7_75t_L g2328 ( 
.A(n_2187),
.B(n_2),
.Y(n_2328)
);

AOI21xp5_ASAP7_75t_L g2329 ( 
.A1(n_2180),
.A2(n_2317),
.B(n_2175),
.Y(n_2329)
);

INVx2_ASAP7_75t_L g2330 ( 
.A(n_2277),
.Y(n_2330)
);

INVx1_ASAP7_75t_L g2331 ( 
.A(n_2318),
.Y(n_2331)
);

AOI22xp5_ASAP7_75t_L g2332 ( 
.A1(n_2322),
.A2(n_832),
.B1(n_836),
.B2(n_834),
.Y(n_2332)
);

INVx1_ASAP7_75t_SL g2333 ( 
.A(n_2201),
.Y(n_2333)
);

NOR2xp33_ASAP7_75t_L g2334 ( 
.A(n_2323),
.B(n_838),
.Y(n_2334)
);

AND2x2_ASAP7_75t_L g2335 ( 
.A(n_2194),
.B(n_839),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_2278),
.Y(n_2336)
);

INVx1_ASAP7_75t_L g2337 ( 
.A(n_2300),
.Y(n_2337)
);

AOI32xp33_ASAP7_75t_L g2338 ( 
.A1(n_2227),
.A2(n_851),
.A3(n_852),
.B1(n_850),
.B2(n_843),
.Y(n_2338)
);

INVx2_ASAP7_75t_L g2339 ( 
.A(n_2264),
.Y(n_2339)
);

AOI222xp33_ASAP7_75t_L g2340 ( 
.A1(n_2221),
.A2(n_2184),
.B1(n_2229),
.B2(n_2236),
.C1(n_2230),
.C2(n_2214),
.Y(n_2340)
);

INVx1_ASAP7_75t_L g2341 ( 
.A(n_2181),
.Y(n_2341)
);

INVx1_ASAP7_75t_L g2342 ( 
.A(n_2216),
.Y(n_2342)
);

INVx2_ASAP7_75t_L g2343 ( 
.A(n_2260),
.Y(n_2343)
);

INVxp67_ASAP7_75t_L g2344 ( 
.A(n_2212),
.Y(n_2344)
);

OR2x2_ASAP7_75t_L g2345 ( 
.A(n_2179),
.B(n_2),
.Y(n_2345)
);

OAI21xp33_ASAP7_75t_SL g2346 ( 
.A1(n_2303),
.A2(n_1829),
.B(n_1790),
.Y(n_2346)
);

INVx1_ASAP7_75t_L g2347 ( 
.A(n_2183),
.Y(n_2347)
);

A2O1A1Ixp33_ASAP7_75t_L g2348 ( 
.A1(n_2251),
.A2(n_879),
.B(n_897),
.C(n_861),
.Y(n_2348)
);

AOI211xp5_ASAP7_75t_L g2349 ( 
.A1(n_2219),
.A2(n_855),
.B(n_856),
.C(n_853),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_2279),
.Y(n_2350)
);

AOI221xp5_ASAP7_75t_L g2351 ( 
.A1(n_2290),
.A2(n_859),
.B1(n_868),
.B2(n_865),
.C(n_860),
.Y(n_2351)
);

NAND2xp5_ASAP7_75t_L g2352 ( 
.A(n_2282),
.B(n_869),
.Y(n_2352)
);

INVx1_ASAP7_75t_L g2353 ( 
.A(n_2280),
.Y(n_2353)
);

INVx1_ASAP7_75t_L g2354 ( 
.A(n_2288),
.Y(n_2354)
);

AOI222xp33_ASAP7_75t_L g2355 ( 
.A1(n_2184),
.A2(n_881),
.B1(n_870),
.B2(n_883),
.C1(n_877),
.C2(n_875),
.Y(n_2355)
);

NAND2x1p5_ASAP7_75t_L g2356 ( 
.A(n_2249),
.B(n_772),
.Y(n_2356)
);

AND2x2_ASAP7_75t_L g2357 ( 
.A(n_2243),
.B(n_2220),
.Y(n_2357)
);

INVx2_ASAP7_75t_L g2358 ( 
.A(n_2260),
.Y(n_2358)
);

NAND2xp33_ASAP7_75t_L g2359 ( 
.A(n_2296),
.B(n_884),
.Y(n_2359)
);

AO22x1_ASAP7_75t_L g2360 ( 
.A1(n_2297),
.A2(n_889),
.B1(n_894),
.B2(n_887),
.Y(n_2360)
);

AOI322xp5_ASAP7_75t_L g2361 ( 
.A1(n_2303),
.A2(n_898),
.A3(n_905),
.B1(n_911),
.B2(n_913),
.C1(n_910),
.C2(n_895),
.Y(n_2361)
);

AOI33xp33_ASAP7_75t_L g2362 ( 
.A1(n_2298),
.A2(n_7),
.A3(n_10),
.B1(n_4),
.B2(n_6),
.B3(n_8),
.Y(n_2362)
);

OR2x2_ASAP7_75t_L g2363 ( 
.A(n_2302),
.B(n_4),
.Y(n_2363)
);

AOI22xp5_ASAP7_75t_L g2364 ( 
.A1(n_2253),
.A2(n_919),
.B1(n_920),
.B2(n_916),
.Y(n_2364)
);

AOI21xp33_ASAP7_75t_L g2365 ( 
.A1(n_2222),
.A2(n_2178),
.B(n_2307),
.Y(n_2365)
);

AOI21xp33_ASAP7_75t_L g2366 ( 
.A1(n_2234),
.A2(n_924),
.B(n_922),
.Y(n_2366)
);

INVx2_ASAP7_75t_SL g2367 ( 
.A(n_2304),
.Y(n_2367)
);

AOI221x1_ASAP7_75t_L g2368 ( 
.A1(n_2271),
.A2(n_904),
.B1(n_947),
.B2(n_849),
.C(n_772),
.Y(n_2368)
);

NAND2xp5_ASAP7_75t_L g2369 ( 
.A(n_2310),
.B(n_925),
.Y(n_2369)
);

INVx1_ASAP7_75t_L g2370 ( 
.A(n_2308),
.Y(n_2370)
);

INVx1_ASAP7_75t_L g2371 ( 
.A(n_2311),
.Y(n_2371)
);

INVx1_ASAP7_75t_L g2372 ( 
.A(n_2312),
.Y(n_2372)
);

OAI22xp5_ASAP7_75t_L g2373 ( 
.A1(n_2281),
.A2(n_929),
.B1(n_930),
.B2(n_928),
.Y(n_2373)
);

AOI221xp5_ASAP7_75t_L g2374 ( 
.A1(n_2208),
.A2(n_936),
.B1(n_938),
.B2(n_934),
.C(n_933),
.Y(n_2374)
);

INVx3_ASAP7_75t_L g2375 ( 
.A(n_2320),
.Y(n_2375)
);

NAND2xp5_ASAP7_75t_L g2376 ( 
.A(n_2292),
.B(n_939),
.Y(n_2376)
);

OR2x2_ASAP7_75t_L g2377 ( 
.A(n_2321),
.B(n_7),
.Y(n_2377)
);

OAI221xp5_ASAP7_75t_L g2378 ( 
.A1(n_2299),
.A2(n_946),
.B1(n_950),
.B2(n_944),
.C(n_943),
.Y(n_2378)
);

INVx2_ASAP7_75t_L g2379 ( 
.A(n_2191),
.Y(n_2379)
);

XOR2xp5_ASAP7_75t_L g2380 ( 
.A(n_2213),
.B(n_2190),
.Y(n_2380)
);

NAND2xp5_ASAP7_75t_L g2381 ( 
.A(n_2289),
.B(n_957),
.Y(n_2381)
);

A2O1A1Ixp33_ASAP7_75t_L g2382 ( 
.A1(n_2263),
.A2(n_984),
.B(n_996),
.C(n_965),
.Y(n_2382)
);

AOI22xp5_ASAP7_75t_L g2383 ( 
.A1(n_2213),
.A2(n_959),
.B1(n_967),
.B2(n_958),
.Y(n_2383)
);

OR2x2_ASAP7_75t_L g2384 ( 
.A(n_2200),
.B(n_8),
.Y(n_2384)
);

INVxp67_ASAP7_75t_L g2385 ( 
.A(n_2209),
.Y(n_2385)
);

OR2x2_ASAP7_75t_L g2386 ( 
.A(n_2268),
.B(n_10),
.Y(n_2386)
);

OAI22xp5_ASAP7_75t_L g2387 ( 
.A1(n_2309),
.A2(n_975),
.B1(n_977),
.B2(n_973),
.Y(n_2387)
);

AOI21xp5_ASAP7_75t_L g2388 ( 
.A1(n_2286),
.A2(n_2185),
.B(n_2186),
.Y(n_2388)
);

NAND2xp5_ASAP7_75t_L g2389 ( 
.A(n_2248),
.B(n_982),
.Y(n_2389)
);

INVx1_ASAP7_75t_L g2390 ( 
.A(n_2182),
.Y(n_2390)
);

INVx2_ASAP7_75t_L g2391 ( 
.A(n_2265),
.Y(n_2391)
);

NAND2xp5_ASAP7_75t_L g2392 ( 
.A(n_2202),
.B(n_987),
.Y(n_2392)
);

NAND2xp5_ASAP7_75t_L g2393 ( 
.A(n_2252),
.B(n_988),
.Y(n_2393)
);

NAND3xp33_ASAP7_75t_L g2394 ( 
.A(n_2287),
.B(n_994),
.C(n_992),
.Y(n_2394)
);

INVx1_ASAP7_75t_L g2395 ( 
.A(n_2210),
.Y(n_2395)
);

AOI21xp33_ASAP7_75t_L g2396 ( 
.A1(n_2276),
.A2(n_1000),
.B(n_998),
.Y(n_2396)
);

INVx1_ASAP7_75t_L g2397 ( 
.A(n_2211),
.Y(n_2397)
);

AND2x2_ASAP7_75t_L g2398 ( 
.A(n_2223),
.B(n_2196),
.Y(n_2398)
);

INVx1_ASAP7_75t_L g2399 ( 
.A(n_2204),
.Y(n_2399)
);

OAI221xp5_ASAP7_75t_L g2400 ( 
.A1(n_2283),
.A2(n_1004),
.B1(n_1005),
.B2(n_1003),
.C(n_1001),
.Y(n_2400)
);

AOI21xp33_ASAP7_75t_SL g2401 ( 
.A1(n_2319),
.A2(n_1016),
.B(n_1007),
.Y(n_2401)
);

AOI222xp33_ASAP7_75t_L g2402 ( 
.A1(n_2205),
.A2(n_1011),
.B1(n_1008),
.B2(n_1013),
.C1(n_1009),
.C2(n_1006),
.Y(n_2402)
);

INVx2_ASAP7_75t_L g2403 ( 
.A(n_2217),
.Y(n_2403)
);

OAI21xp5_ASAP7_75t_L g2404 ( 
.A1(n_2239),
.A2(n_1019),
.B(n_1014),
.Y(n_2404)
);

INVx1_ASAP7_75t_SL g2405 ( 
.A(n_2247),
.Y(n_2405)
);

INVx1_ASAP7_75t_L g2406 ( 
.A(n_2235),
.Y(n_2406)
);

NAND2xp5_ASAP7_75t_L g2407 ( 
.A(n_2272),
.B(n_1020),
.Y(n_2407)
);

AOI22xp5_ASAP7_75t_L g2408 ( 
.A1(n_2197),
.A2(n_1028),
.B1(n_1026),
.B2(n_1744),
.Y(n_2408)
);

AOI221xp5_ASAP7_75t_L g2409 ( 
.A1(n_2238),
.A2(n_904),
.B1(n_947),
.B2(n_849),
.C(n_772),
.Y(n_2409)
);

INVx1_ASAP7_75t_L g2410 ( 
.A(n_2199),
.Y(n_2410)
);

OAI22xp33_ASAP7_75t_L g2411 ( 
.A1(n_2291),
.A2(n_1734),
.B1(n_1807),
.B2(n_1801),
.Y(n_2411)
);

AOI22xp33_ASAP7_75t_L g2412 ( 
.A1(n_2198),
.A2(n_1725),
.B1(n_1744),
.B2(n_1788),
.Y(n_2412)
);

A2O1A1Ixp33_ASAP7_75t_SL g2413 ( 
.A1(n_2241),
.A2(n_13),
.B(n_11),
.C(n_12),
.Y(n_2413)
);

INVxp33_ASAP7_75t_L g2414 ( 
.A(n_2293),
.Y(n_2414)
);

NAND3xp33_ASAP7_75t_L g2415 ( 
.A(n_2262),
.B(n_849),
.C(n_772),
.Y(n_2415)
);

AOI22xp5_ASAP7_75t_L g2416 ( 
.A1(n_2245),
.A2(n_1649),
.B1(n_1721),
.B2(n_1725),
.Y(n_2416)
);

AND2x2_ASAP7_75t_L g2417 ( 
.A(n_2207),
.B(n_1829),
.Y(n_2417)
);

AOI22xp33_ASAP7_75t_L g2418 ( 
.A1(n_2189),
.A2(n_1725),
.B1(n_1788),
.B2(n_904),
.Y(n_2418)
);

AOI221xp5_ASAP7_75t_L g2419 ( 
.A1(n_2242),
.A2(n_849),
.B1(n_972),
.B2(n_947),
.C(n_904),
.Y(n_2419)
);

INVx1_ASAP7_75t_L g2420 ( 
.A(n_2176),
.Y(n_2420)
);

INVx1_ASAP7_75t_L g2421 ( 
.A(n_2257),
.Y(n_2421)
);

AOI32xp33_ASAP7_75t_L g2422 ( 
.A1(n_2266),
.A2(n_1736),
.A3(n_1698),
.B1(n_1721),
.B2(n_1740),
.Y(n_2422)
);

NOR2xp33_ASAP7_75t_SL g2423 ( 
.A(n_2269),
.B(n_1649),
.Y(n_2423)
);

HB1xp67_ASAP7_75t_L g2424 ( 
.A(n_2203),
.Y(n_2424)
);

INVx1_ASAP7_75t_L g2425 ( 
.A(n_2195),
.Y(n_2425)
);

INVx1_ASAP7_75t_L g2426 ( 
.A(n_2224),
.Y(n_2426)
);

INVx2_ASAP7_75t_L g2427 ( 
.A(n_2255),
.Y(n_2427)
);

NAND2xp5_ASAP7_75t_L g2428 ( 
.A(n_2294),
.B(n_11),
.Y(n_2428)
);

NAND2xp5_ASAP7_75t_SL g2429 ( 
.A(n_2174),
.B(n_904),
.Y(n_2429)
);

OAI221xp5_ASAP7_75t_SL g2430 ( 
.A1(n_2254),
.A2(n_2275),
.B1(n_2284),
.B2(n_2261),
.C(n_2233),
.Y(n_2430)
);

INVx1_ASAP7_75t_L g2431 ( 
.A(n_2225),
.Y(n_2431)
);

AND2x2_ASAP7_75t_L g2432 ( 
.A(n_2295),
.B(n_13),
.Y(n_2432)
);

NAND2xp5_ASAP7_75t_L g2433 ( 
.A(n_2305),
.B(n_14),
.Y(n_2433)
);

INVx2_ASAP7_75t_L g2434 ( 
.A(n_2244),
.Y(n_2434)
);

INVx1_ASAP7_75t_L g2435 ( 
.A(n_2206),
.Y(n_2435)
);

AOI32xp33_ASAP7_75t_L g2436 ( 
.A1(n_2226),
.A2(n_1736),
.A3(n_1698),
.B1(n_1721),
.B2(n_1740),
.Y(n_2436)
);

INVx1_ASAP7_75t_L g2437 ( 
.A(n_2306),
.Y(n_2437)
);

INVx1_ASAP7_75t_L g2438 ( 
.A(n_2316),
.Y(n_2438)
);

OAI21xp5_ASAP7_75t_L g2439 ( 
.A1(n_2261),
.A2(n_1717),
.B(n_1710),
.Y(n_2439)
);

INVx1_ASAP7_75t_SL g2440 ( 
.A(n_2215),
.Y(n_2440)
);

NAND2xp5_ASAP7_75t_L g2441 ( 
.A(n_2177),
.B(n_15),
.Y(n_2441)
);

NAND2xp5_ASAP7_75t_SL g2442 ( 
.A(n_2232),
.B(n_904),
.Y(n_2442)
);

NAND3x1_ASAP7_75t_L g2443 ( 
.A(n_2375),
.B(n_2240),
.C(n_2301),
.Y(n_2443)
);

O2A1O1Ixp33_ASAP7_75t_L g2444 ( 
.A1(n_2413),
.A2(n_2285),
.B(n_2313),
.C(n_2258),
.Y(n_2444)
);

NOR2xp33_ASAP7_75t_L g2445 ( 
.A(n_2325),
.B(n_2231),
.Y(n_2445)
);

NAND2xp5_ASAP7_75t_L g2446 ( 
.A(n_2360),
.B(n_2237),
.Y(n_2446)
);

AOI221xp5_ASAP7_75t_L g2447 ( 
.A1(n_2329),
.A2(n_2256),
.B1(n_2237),
.B2(n_2192),
.C(n_2228),
.Y(n_2447)
);

NAND3xp33_ASAP7_75t_L g2448 ( 
.A(n_2338),
.B(n_2259),
.C(n_2193),
.Y(n_2448)
);

OR2x2_ASAP7_75t_L g2449 ( 
.A(n_2324),
.B(n_2250),
.Y(n_2449)
);

AOI322xp5_ASAP7_75t_L g2450 ( 
.A1(n_2331),
.A2(n_2218),
.A3(n_2246),
.B1(n_2274),
.B2(n_2267),
.C1(n_2270),
.C2(n_1826),
.Y(n_2450)
);

OAI221xp5_ASAP7_75t_SL g2451 ( 
.A1(n_2385),
.A2(n_1808),
.B1(n_1826),
.B2(n_1811),
.C(n_1801),
.Y(n_2451)
);

OAI322xp33_ASAP7_75t_L g2452 ( 
.A1(n_2350),
.A2(n_972),
.A3(n_947),
.B1(n_20),
.B2(n_17),
.C1(n_19),
.C2(n_15),
.Y(n_2452)
);

INVx1_ASAP7_75t_L g2453 ( 
.A(n_2424),
.Y(n_2453)
);

NOR2xp33_ASAP7_75t_L g2454 ( 
.A(n_2414),
.B(n_2333),
.Y(n_2454)
);

INVx1_ASAP7_75t_L g2455 ( 
.A(n_2362),
.Y(n_2455)
);

AOI211xp5_ASAP7_75t_L g2456 ( 
.A1(n_2357),
.A2(n_972),
.B(n_947),
.C(n_18),
.Y(n_2456)
);

AOI22xp5_ASAP7_75t_L g2457 ( 
.A1(n_2330),
.A2(n_1725),
.B1(n_1788),
.B2(n_972),
.Y(n_2457)
);

OAI21xp5_ASAP7_75t_SL g2458 ( 
.A1(n_2398),
.A2(n_972),
.B(n_947),
.Y(n_2458)
);

AOI22xp5_ASAP7_75t_L g2459 ( 
.A1(n_2406),
.A2(n_972),
.B1(n_1808),
.B2(n_1801),
.Y(n_2459)
);

NAND2xp5_ASAP7_75t_L g2460 ( 
.A(n_2336),
.B(n_16),
.Y(n_2460)
);

AND2x2_ASAP7_75t_L g2461 ( 
.A(n_2367),
.B(n_16),
.Y(n_2461)
);

AOI22xp33_ASAP7_75t_L g2462 ( 
.A1(n_2341),
.A2(n_1808),
.B1(n_1826),
.B2(n_1811),
.Y(n_2462)
);

OAI222xp33_ASAP7_75t_L g2463 ( 
.A1(n_2430),
.A2(n_1719),
.B1(n_1811),
.B2(n_1847),
.C1(n_1838),
.C2(n_1827),
.Y(n_2463)
);

AOI221xp5_ASAP7_75t_L g2464 ( 
.A1(n_2400),
.A2(n_979),
.B1(n_874),
.B2(n_914),
.C(n_841),
.Y(n_2464)
);

OAI22xp5_ASAP7_75t_L g2465 ( 
.A1(n_2391),
.A2(n_1827),
.B1(n_1847),
.B2(n_1838),
.Y(n_2465)
);

OAI21xp5_ASAP7_75t_L g2466 ( 
.A1(n_2388),
.A2(n_1717),
.B(n_1710),
.Y(n_2466)
);

INVxp67_ASAP7_75t_L g2467 ( 
.A(n_2423),
.Y(n_2467)
);

INVx1_ASAP7_75t_L g2468 ( 
.A(n_2384),
.Y(n_2468)
);

OAI211xp5_ASAP7_75t_L g2469 ( 
.A1(n_2375),
.A2(n_21),
.B(n_17),
.C(n_18),
.Y(n_2469)
);

A2O1A1Ixp33_ASAP7_75t_L g2470 ( 
.A1(n_2378),
.A2(n_2436),
.B(n_2337),
.C(n_2382),
.Y(n_2470)
);

O2A1O1Ixp33_ASAP7_75t_L g2471 ( 
.A1(n_2359),
.A2(n_25),
.B(n_21),
.C(n_23),
.Y(n_2471)
);

AOI22xp5_ASAP7_75t_L g2472 ( 
.A1(n_2437),
.A2(n_1521),
.B1(n_1795),
.B2(n_1827),
.Y(n_2472)
);

NAND4xp25_ASAP7_75t_L g2473 ( 
.A(n_2440),
.B(n_26),
.C(n_23),
.D(n_25),
.Y(n_2473)
);

AOI221xp5_ASAP7_75t_L g2474 ( 
.A1(n_2365),
.A2(n_979),
.B1(n_954),
.B2(n_927),
.C(n_822),
.Y(n_2474)
);

NAND4xp25_ASAP7_75t_SL g2475 ( 
.A(n_2353),
.B(n_28),
.C(n_26),
.D(n_27),
.Y(n_2475)
);

AOI32xp33_ASAP7_75t_L g2476 ( 
.A1(n_2339),
.A2(n_1740),
.A3(n_31),
.B1(n_29),
.B2(n_30),
.Y(n_2476)
);

OAI211xp5_ASAP7_75t_SL g2477 ( 
.A1(n_2354),
.A2(n_31),
.B(n_29),
.C(n_30),
.Y(n_2477)
);

AOI22xp33_ASAP7_75t_L g2478 ( 
.A1(n_2405),
.A2(n_1729),
.B1(n_1795),
.B2(n_1819),
.Y(n_2478)
);

OAI21xp5_ASAP7_75t_L g2479 ( 
.A1(n_2370),
.A2(n_1719),
.B(n_1695),
.Y(n_2479)
);

OAI221xp5_ASAP7_75t_SL g2480 ( 
.A1(n_2343),
.A2(n_1850),
.B1(n_1847),
.B2(n_1838),
.C(n_36),
.Y(n_2480)
);

AOI221xp5_ASAP7_75t_L g2481 ( 
.A1(n_2438),
.A2(n_979),
.B1(n_991),
.B2(n_985),
.C(n_989),
.Y(n_2481)
);

INVx1_ASAP7_75t_L g2482 ( 
.A(n_2345),
.Y(n_2482)
);

AOI211xp5_ASAP7_75t_L g2483 ( 
.A1(n_2371),
.A2(n_37),
.B(n_32),
.C(n_34),
.Y(n_2483)
);

NAND2xp5_ASAP7_75t_SL g2484 ( 
.A(n_2402),
.B(n_2358),
.Y(n_2484)
);

AOI211xp5_ASAP7_75t_L g2485 ( 
.A1(n_2372),
.A2(n_38),
.B(n_34),
.C(n_37),
.Y(n_2485)
);

OAI22xp33_ASAP7_75t_L g2486 ( 
.A1(n_2383),
.A2(n_1729),
.B1(n_1850),
.B2(n_1786),
.Y(n_2486)
);

OAI221xp5_ASAP7_75t_L g2487 ( 
.A1(n_2383),
.A2(n_1850),
.B1(n_1729),
.B2(n_1786),
.C(n_979),
.Y(n_2487)
);

NOR3xp33_ASAP7_75t_L g2488 ( 
.A(n_2415),
.B(n_39),
.C(n_40),
.Y(n_2488)
);

AOI21xp5_ASAP7_75t_L g2489 ( 
.A1(n_2376),
.A2(n_44),
.B(n_43),
.Y(n_2489)
);

AOI21xp5_ASAP7_75t_L g2490 ( 
.A1(n_2326),
.A2(n_45),
.B(n_43),
.Y(n_2490)
);

OAI21xp5_ASAP7_75t_SL g2491 ( 
.A1(n_2410),
.A2(n_41),
.B(n_48),
.Y(n_2491)
);

NAND4xp25_ASAP7_75t_L g2492 ( 
.A(n_2425),
.B(n_2332),
.C(n_2340),
.D(n_2403),
.Y(n_2492)
);

AOI221xp5_ASAP7_75t_L g2493 ( 
.A1(n_2351),
.A2(n_979),
.B1(n_1729),
.B2(n_1795),
.C(n_50),
.Y(n_2493)
);

AOI22xp5_ASAP7_75t_L g2494 ( 
.A1(n_2421),
.A2(n_1729),
.B1(n_1819),
.B2(n_1753),
.Y(n_2494)
);

OAI221xp5_ASAP7_75t_L g2495 ( 
.A1(n_2346),
.A2(n_1729),
.B1(n_1753),
.B2(n_1751),
.C(n_50),
.Y(n_2495)
);

O2A1O1Ixp33_ASAP7_75t_L g2496 ( 
.A1(n_2401),
.A2(n_51),
.B(n_48),
.C(n_49),
.Y(n_2496)
);

NAND4xp75_ASAP7_75t_L g2497 ( 
.A(n_2368),
.B(n_53),
.C(n_49),
.D(n_52),
.Y(n_2497)
);

AOI221xp5_ASAP7_75t_L g2498 ( 
.A1(n_2399),
.A2(n_2346),
.B1(n_2394),
.B2(n_2380),
.C(n_2401),
.Y(n_2498)
);

NAND3xp33_ASAP7_75t_L g2499 ( 
.A(n_2349),
.B(n_54),
.C(n_55),
.Y(n_2499)
);

NAND3xp33_ASAP7_75t_SL g2500 ( 
.A(n_2328),
.B(n_56),
.C(n_57),
.Y(n_2500)
);

INVxp67_ASAP7_75t_L g2501 ( 
.A(n_2334),
.Y(n_2501)
);

AOI221xp5_ASAP7_75t_L g2502 ( 
.A1(n_2392),
.A2(n_61),
.B1(n_59),
.B2(n_60),
.C(n_63),
.Y(n_2502)
);

NAND2xp5_ASAP7_75t_L g2503 ( 
.A(n_2335),
.B(n_59),
.Y(n_2503)
);

OAI221xp5_ASAP7_75t_L g2504 ( 
.A1(n_2422),
.A2(n_1751),
.B1(n_64),
.B2(n_60),
.C(n_63),
.Y(n_2504)
);

OA22x2_ASAP7_75t_L g2505 ( 
.A1(n_2434),
.A2(n_67),
.B1(n_64),
.B2(n_65),
.Y(n_2505)
);

NAND4xp25_ASAP7_75t_L g2506 ( 
.A(n_2427),
.B(n_72),
.C(n_69),
.D(n_70),
.Y(n_2506)
);

OAI21xp33_ASAP7_75t_L g2507 ( 
.A1(n_2389),
.A2(n_1695),
.B(n_1728),
.Y(n_2507)
);

NAND3xp33_ASAP7_75t_L g2508 ( 
.A(n_2409),
.B(n_69),
.C(n_70),
.Y(n_2508)
);

AOI221xp5_ASAP7_75t_L g2509 ( 
.A1(n_2393),
.A2(n_75),
.B1(n_73),
.B2(n_74),
.C(n_76),
.Y(n_2509)
);

A2O1A1Ixp33_ASAP7_75t_L g2510 ( 
.A1(n_2364),
.A2(n_75),
.B(n_73),
.C(n_74),
.Y(n_2510)
);

INVx1_ASAP7_75t_L g2511 ( 
.A(n_2363),
.Y(n_2511)
);

O2A1O1Ixp33_ASAP7_75t_SL g2512 ( 
.A1(n_2327),
.A2(n_79),
.B(n_76),
.C(n_77),
.Y(n_2512)
);

NAND3xp33_ASAP7_75t_L g2513 ( 
.A(n_2419),
.B(n_80),
.C(n_81),
.Y(n_2513)
);

OAI211xp5_ASAP7_75t_SL g2514 ( 
.A1(n_2429),
.A2(n_82),
.B(n_80),
.C(n_81),
.Y(n_2514)
);

NAND3xp33_ASAP7_75t_SL g2515 ( 
.A(n_2377),
.B(n_2356),
.C(n_2342),
.Y(n_2515)
);

AOI21xp5_ASAP7_75t_L g2516 ( 
.A1(n_2348),
.A2(n_82),
.B(n_83),
.Y(n_2516)
);

OAI21xp33_ASAP7_75t_L g2517 ( 
.A1(n_2381),
.A2(n_2435),
.B(n_2426),
.Y(n_2517)
);

OAI21xp5_ASAP7_75t_SL g2518 ( 
.A1(n_2344),
.A2(n_83),
.B(n_84),
.Y(n_2518)
);

AOI22xp5_ASAP7_75t_L g2519 ( 
.A1(n_2352),
.A2(n_1819),
.B1(n_1728),
.B2(n_1747),
.Y(n_2519)
);

INVx1_ASAP7_75t_L g2520 ( 
.A(n_2441),
.Y(n_2520)
);

AOI322xp5_ASAP7_75t_L g2521 ( 
.A1(n_2390),
.A2(n_1731),
.A3(n_1780),
.B1(n_92),
.B2(n_89),
.C1(n_91),
.C2(n_86),
.Y(n_2521)
);

XOR2x2_ASAP7_75t_L g2522 ( 
.A(n_2369),
.B(n_87),
.Y(n_2522)
);

OAI221xp5_ASAP7_75t_L g2523 ( 
.A1(n_2439),
.A2(n_91),
.B1(n_87),
.B2(n_90),
.C(n_92),
.Y(n_2523)
);

AOI222xp33_ASAP7_75t_L g2524 ( 
.A1(n_2347),
.A2(n_1731),
.B1(n_95),
.B2(n_98),
.C1(n_93),
.C2(n_94),
.Y(n_2524)
);

AOI21xp5_ASAP7_75t_L g2525 ( 
.A1(n_2404),
.A2(n_93),
.B(n_94),
.Y(n_2525)
);

O2A1O1Ixp33_ASAP7_75t_L g2526 ( 
.A1(n_2428),
.A2(n_100),
.B(n_97),
.C(n_99),
.Y(n_2526)
);

OAI321xp33_ASAP7_75t_L g2527 ( 
.A1(n_2431),
.A2(n_1731),
.A3(n_104),
.B1(n_106),
.B2(n_101),
.C(n_103),
.Y(n_2527)
);

AOI221xp5_ASAP7_75t_L g2528 ( 
.A1(n_2420),
.A2(n_105),
.B1(n_101),
.B2(n_104),
.C(n_106),
.Y(n_2528)
);

NOR4xp25_ASAP7_75t_L g2529 ( 
.A(n_2395),
.B(n_108),
.C(n_105),
.D(n_107),
.Y(n_2529)
);

AO21x1_ASAP7_75t_L g2530 ( 
.A1(n_2373),
.A2(n_109),
.B(n_110),
.Y(n_2530)
);

NAND2xp5_ASAP7_75t_SL g2531 ( 
.A(n_2355),
.B(n_112),
.Y(n_2531)
);

OR2x2_ASAP7_75t_L g2532 ( 
.A(n_2386),
.B(n_112),
.Y(n_2532)
);

OAI31xp33_ASAP7_75t_L g2533 ( 
.A1(n_2397),
.A2(n_116),
.A3(n_113),
.B(n_115),
.Y(n_2533)
);

HB1xp67_ASAP7_75t_L g2534 ( 
.A(n_2432),
.Y(n_2534)
);

OA21x2_ASAP7_75t_L g2535 ( 
.A1(n_2366),
.A2(n_115),
.B(n_117),
.Y(n_2535)
);

A2O1A1Ixp33_ASAP7_75t_SL g2536 ( 
.A1(n_2387),
.A2(n_119),
.B(n_117),
.C(n_118),
.Y(n_2536)
);

NAND2xp5_ASAP7_75t_L g2537 ( 
.A(n_2361),
.B(n_118),
.Y(n_2537)
);

OR2x2_ASAP7_75t_L g2538 ( 
.A(n_2433),
.B(n_119),
.Y(n_2538)
);

AND2x2_ASAP7_75t_L g2539 ( 
.A(n_2417),
.B(n_120),
.Y(n_2539)
);

OR2x2_ASAP7_75t_L g2540 ( 
.A(n_2407),
.B(n_120),
.Y(n_2540)
);

OAI21xp5_ASAP7_75t_SL g2541 ( 
.A1(n_2416),
.A2(n_121),
.B(n_122),
.Y(n_2541)
);

INVx1_ASAP7_75t_L g2542 ( 
.A(n_2379),
.Y(n_2542)
);

AOI211xp5_ASAP7_75t_SL g2543 ( 
.A1(n_2396),
.A2(n_125),
.B(n_123),
.C(n_124),
.Y(n_2543)
);

INVx1_ASAP7_75t_L g2544 ( 
.A(n_2408),
.Y(n_2544)
);

NAND2xp5_ASAP7_75t_L g2545 ( 
.A(n_2374),
.B(n_2418),
.Y(n_2545)
);

NAND3xp33_ASAP7_75t_L g2546 ( 
.A(n_2442),
.B(n_125),
.C(n_127),
.Y(n_2546)
);

NOR2xp33_ASAP7_75t_SL g2547 ( 
.A(n_2411),
.B(n_128),
.Y(n_2547)
);

AOI211xp5_ASAP7_75t_SL g2548 ( 
.A1(n_2408),
.A2(n_130),
.B(n_128),
.C(n_129),
.Y(n_2548)
);

AOI211xp5_ASAP7_75t_SL g2549 ( 
.A1(n_2412),
.A2(n_132),
.B(n_130),
.C(n_131),
.Y(n_2549)
);

NOR3xp33_ASAP7_75t_L g2550 ( 
.A(n_2360),
.B(n_131),
.C(n_132),
.Y(n_2550)
);

AOI221xp5_ASAP7_75t_L g2551 ( 
.A1(n_2329),
.A2(n_135),
.B1(n_133),
.B2(n_134),
.C(n_136),
.Y(n_2551)
);

A2O1A1Ixp33_ASAP7_75t_L g2552 ( 
.A1(n_2329),
.A2(n_135),
.B(n_133),
.C(n_134),
.Y(n_2552)
);

NAND2xp5_ASAP7_75t_L g2553 ( 
.A(n_2360),
.B(n_137),
.Y(n_2553)
);

INVx1_ASAP7_75t_L g2554 ( 
.A(n_2424),
.Y(n_2554)
);

OAI21xp5_ASAP7_75t_L g2555 ( 
.A1(n_2325),
.A2(n_1733),
.B(n_1745),
.Y(n_2555)
);

AND2x2_ASAP7_75t_L g2556 ( 
.A(n_2398),
.B(n_137),
.Y(n_2556)
);

NOR2xp33_ASAP7_75t_L g2557 ( 
.A(n_2325),
.B(n_138),
.Y(n_2557)
);

AOI322xp5_ASAP7_75t_L g2558 ( 
.A1(n_2331),
.A2(n_1731),
.A3(n_1780),
.B1(n_146),
.B2(n_141),
.C1(n_144),
.C2(n_139),
.Y(n_2558)
);

AOI21xp5_ASAP7_75t_L g2559 ( 
.A1(n_2413),
.A2(n_139),
.B(n_140),
.Y(n_2559)
);

NOR4xp75_ASAP7_75t_SL g2560 ( 
.A(n_2327),
.B(n_146),
.C(n_141),
.D(n_143),
.Y(n_2560)
);

NAND2xp5_ASAP7_75t_SL g2561 ( 
.A(n_2324),
.B(n_143),
.Y(n_2561)
);

AOI22xp5_ASAP7_75t_L g2562 ( 
.A1(n_2333),
.A2(n_1819),
.B1(n_1747),
.B2(n_1745),
.Y(n_2562)
);

NAND4xp25_ASAP7_75t_L g2563 ( 
.A(n_2357),
.B(n_150),
.C(n_148),
.D(n_149),
.Y(n_2563)
);

AO21x1_ASAP7_75t_L g2564 ( 
.A1(n_2329),
.A2(n_149),
.B(n_151),
.Y(n_2564)
);

O2A1O1Ixp33_ASAP7_75t_L g2565 ( 
.A1(n_2413),
.A2(n_153),
.B(n_151),
.C(n_152),
.Y(n_2565)
);

OAI21xp33_ASAP7_75t_L g2566 ( 
.A1(n_2357),
.A2(n_152),
.B(n_153),
.Y(n_2566)
);

NAND3xp33_ASAP7_75t_L g2567 ( 
.A(n_2325),
.B(n_154),
.C(n_155),
.Y(n_2567)
);

NAND3xp33_ASAP7_75t_SL g2568 ( 
.A(n_2333),
.B(n_155),
.C(n_156),
.Y(n_2568)
);

NOR3xp33_ASAP7_75t_L g2569 ( 
.A(n_2360),
.B(n_156),
.C(n_158),
.Y(n_2569)
);

OAI211xp5_ASAP7_75t_L g2570 ( 
.A1(n_2325),
.A2(n_160),
.B(n_158),
.C(n_159),
.Y(n_2570)
);

NAND3xp33_ASAP7_75t_SL g2571 ( 
.A(n_2333),
.B(n_159),
.C(n_161),
.Y(n_2571)
);

OAI21xp5_ASAP7_75t_L g2572 ( 
.A1(n_2325),
.A2(n_1733),
.B(n_161),
.Y(n_2572)
);

AOI22xp5_ASAP7_75t_L g2573 ( 
.A1(n_2333),
.A2(n_1819),
.B1(n_1731),
.B2(n_1780),
.Y(n_2573)
);

AOI211xp5_ASAP7_75t_SL g2574 ( 
.A1(n_2325),
.A2(n_164),
.B(n_162),
.C(n_163),
.Y(n_2574)
);

NOR3xp33_ASAP7_75t_L g2575 ( 
.A(n_2360),
.B(n_162),
.C(n_163),
.Y(n_2575)
);

NAND2xp5_ASAP7_75t_SL g2576 ( 
.A(n_2324),
.B(n_164),
.Y(n_2576)
);

AOI21xp33_ASAP7_75t_L g2577 ( 
.A1(n_2414),
.A2(n_166),
.B(n_167),
.Y(n_2577)
);

AOI22xp33_ASAP7_75t_L g2578 ( 
.A1(n_2341),
.A2(n_1731),
.B1(n_1101),
.B2(n_1102),
.Y(n_2578)
);

NOR3xp33_ASAP7_75t_L g2579 ( 
.A(n_2360),
.B(n_166),
.C(n_167),
.Y(n_2579)
);

AOI22xp33_ASAP7_75t_L g2580 ( 
.A1(n_2341),
.A2(n_1102),
.B1(n_1096),
.B2(n_1780),
.Y(n_2580)
);

AOI221xp5_ASAP7_75t_L g2581 ( 
.A1(n_2329),
.A2(n_171),
.B1(n_168),
.B2(n_170),
.C(n_172),
.Y(n_2581)
);

AOI21xp5_ASAP7_75t_L g2582 ( 
.A1(n_2413),
.A2(n_168),
.B(n_173),
.Y(n_2582)
);

NAND4xp25_ASAP7_75t_SL g2583 ( 
.A(n_2324),
.B(n_176),
.C(n_174),
.D(n_175),
.Y(n_2583)
);

AOI22xp33_ASAP7_75t_L g2584 ( 
.A1(n_2341),
.A2(n_1780),
.B1(n_1117),
.B2(n_1118),
.Y(n_2584)
);

OAI21xp33_ASAP7_75t_L g2585 ( 
.A1(n_2357),
.A2(n_174),
.B(n_175),
.Y(n_2585)
);

OAI21xp5_ASAP7_75t_SL g2586 ( 
.A1(n_2325),
.A2(n_176),
.B(n_177),
.Y(n_2586)
);

AOI22xp5_ASAP7_75t_L g2587 ( 
.A1(n_2333),
.A2(n_181),
.B1(n_179),
.B2(n_180),
.Y(n_2587)
);

NOR2xp67_ASAP7_75t_L g2588 ( 
.A(n_2325),
.B(n_182),
.Y(n_2588)
);

AOI321xp33_ASAP7_75t_L g2589 ( 
.A1(n_2329),
.A2(n_186),
.A3(n_188),
.B1(n_183),
.B2(n_185),
.C(n_187),
.Y(n_2589)
);

NOR2xp33_ASAP7_75t_L g2590 ( 
.A(n_2325),
.B(n_183),
.Y(n_2590)
);

AOI21xp5_ASAP7_75t_L g2591 ( 
.A1(n_2413),
.A2(n_186),
.B(n_187),
.Y(n_2591)
);

OAI21xp5_ASAP7_75t_SL g2592 ( 
.A1(n_2454),
.A2(n_189),
.B(n_191),
.Y(n_2592)
);

AOI22xp5_ASAP7_75t_L g2593 ( 
.A1(n_2539),
.A2(n_193),
.B1(n_191),
.B2(n_192),
.Y(n_2593)
);

AND2x2_ASAP7_75t_L g2594 ( 
.A(n_2556),
.B(n_193),
.Y(n_2594)
);

INVx1_ASAP7_75t_L g2595 ( 
.A(n_2534),
.Y(n_2595)
);

AOI221x1_ASAP7_75t_L g2596 ( 
.A1(n_2492),
.A2(n_197),
.B1(n_195),
.B2(n_196),
.C(n_198),
.Y(n_2596)
);

NOR2xp33_ASAP7_75t_L g2597 ( 
.A(n_2568),
.B(n_196),
.Y(n_2597)
);

AOI22xp5_ASAP7_75t_L g2598 ( 
.A1(n_2520),
.A2(n_200),
.B1(n_197),
.B2(n_199),
.Y(n_2598)
);

AOI22xp5_ASAP7_75t_L g2599 ( 
.A1(n_2484),
.A2(n_2571),
.B1(n_2482),
.B2(n_2511),
.Y(n_2599)
);

INVx1_ASAP7_75t_L g2600 ( 
.A(n_2505),
.Y(n_2600)
);

OAI322xp33_ASAP7_75t_L g2601 ( 
.A1(n_2467),
.A2(n_2554),
.A3(n_2453),
.B1(n_2547),
.B2(n_2449),
.C1(n_2446),
.C2(n_2445),
.Y(n_2601)
);

AOI22xp5_ASAP7_75t_L g2602 ( 
.A1(n_2564),
.A2(n_203),
.B1(n_201),
.B2(n_202),
.Y(n_2602)
);

INVx1_ASAP7_75t_L g2603 ( 
.A(n_2505),
.Y(n_2603)
);

OAI22xp33_ASAP7_75t_L g2604 ( 
.A1(n_2492),
.A2(n_203),
.B1(n_201),
.B2(n_202),
.Y(n_2604)
);

NAND2xp5_ASAP7_75t_L g2605 ( 
.A(n_2574),
.B(n_204),
.Y(n_2605)
);

OAI221xp5_ASAP7_75t_L g2606 ( 
.A1(n_2565),
.A2(n_206),
.B1(n_204),
.B2(n_205),
.C(n_208),
.Y(n_2606)
);

OAI22xp33_ASAP7_75t_SL g2607 ( 
.A1(n_2468),
.A2(n_208),
.B1(n_205),
.B2(n_206),
.Y(n_2607)
);

OAI22xp5_ASAP7_75t_L g2608 ( 
.A1(n_2587),
.A2(n_211),
.B1(n_209),
.B2(n_210),
.Y(n_2608)
);

INVx1_ASAP7_75t_L g2609 ( 
.A(n_2588),
.Y(n_2609)
);

AOI21xp33_ASAP7_75t_SL g2610 ( 
.A1(n_2444),
.A2(n_209),
.B(n_210),
.Y(n_2610)
);

AOI321xp33_ASAP7_75t_L g2611 ( 
.A1(n_2498),
.A2(n_213),
.A3(n_215),
.B1(n_211),
.B2(n_212),
.C(n_214),
.Y(n_2611)
);

INVx1_ASAP7_75t_L g2612 ( 
.A(n_2532),
.Y(n_2612)
);

INVxp67_ASAP7_75t_L g2613 ( 
.A(n_2497),
.Y(n_2613)
);

AOI211xp5_ASAP7_75t_L g2614 ( 
.A1(n_2455),
.A2(n_217),
.B(n_212),
.C(n_216),
.Y(n_2614)
);

INVxp67_ASAP7_75t_L g2615 ( 
.A(n_2461),
.Y(n_2615)
);

OAI21xp33_ASAP7_75t_L g2616 ( 
.A1(n_2517),
.A2(n_218),
.B(n_219),
.Y(n_2616)
);

AOI22xp33_ASAP7_75t_L g2617 ( 
.A1(n_2544),
.A2(n_1117),
.B1(n_1118),
.B2(n_1115),
.Y(n_2617)
);

INVx2_ASAP7_75t_L g2618 ( 
.A(n_2522),
.Y(n_2618)
);

BUFx2_ASAP7_75t_L g2619 ( 
.A(n_2443),
.Y(n_2619)
);

INVx1_ASAP7_75t_L g2620 ( 
.A(n_2589),
.Y(n_2620)
);

AOI31xp33_ASAP7_75t_L g2621 ( 
.A1(n_2557),
.A2(n_221),
.A3(n_219),
.B(n_220),
.Y(n_2621)
);

OAI21xp5_ASAP7_75t_L g2622 ( 
.A1(n_2552),
.A2(n_220),
.B(n_223),
.Y(n_2622)
);

NOR3xp33_ASAP7_75t_SL g2623 ( 
.A(n_2515),
.B(n_225),
.C(n_226),
.Y(n_2623)
);

AOI21xp5_ASAP7_75t_L g2624 ( 
.A1(n_2559),
.A2(n_2591),
.B(n_2582),
.Y(n_2624)
);

INVx1_ASAP7_75t_L g2625 ( 
.A(n_2538),
.Y(n_2625)
);

INVx1_ASAP7_75t_L g2626 ( 
.A(n_2530),
.Y(n_2626)
);

AOI21xp5_ASAP7_75t_L g2627 ( 
.A1(n_2561),
.A2(n_227),
.B(n_228),
.Y(n_2627)
);

AOI22xp33_ASAP7_75t_L g2628 ( 
.A1(n_2531),
.A2(n_1117),
.B1(n_1118),
.B2(n_1115),
.Y(n_2628)
);

OAI21xp5_ASAP7_75t_L g2629 ( 
.A1(n_2491),
.A2(n_227),
.B(n_228),
.Y(n_2629)
);

AOI22xp33_ASAP7_75t_L g2630 ( 
.A1(n_2495),
.A2(n_1117),
.B1(n_1118),
.B2(n_1115),
.Y(n_2630)
);

AOI221xp5_ASAP7_75t_L g2631 ( 
.A1(n_2463),
.A2(n_232),
.B1(n_229),
.B2(n_230),
.C(n_233),
.Y(n_2631)
);

OAI32xp33_ASAP7_75t_L g2632 ( 
.A1(n_2542),
.A2(n_233),
.A3(n_230),
.B1(n_232),
.B2(n_234),
.Y(n_2632)
);

INVx1_ASAP7_75t_L g2633 ( 
.A(n_2553),
.Y(n_2633)
);

AOI22xp33_ASAP7_75t_L g2634 ( 
.A1(n_2504),
.A2(n_1117),
.B1(n_1118),
.B2(n_1115),
.Y(n_2634)
);

NOR2xp33_ASAP7_75t_L g2635 ( 
.A(n_2473),
.B(n_234),
.Y(n_2635)
);

OAI322xp33_ASAP7_75t_L g2636 ( 
.A1(n_2545),
.A2(n_235),
.A3(n_236),
.B1(n_238),
.B2(n_240),
.C1(n_241),
.C2(n_242),
.Y(n_2636)
);

NAND5xp2_ASAP7_75t_L g2637 ( 
.A(n_2447),
.B(n_244),
.C(n_235),
.D(n_243),
.E(n_245),
.Y(n_2637)
);

NAND2xp5_ASAP7_75t_L g2638 ( 
.A(n_2529),
.B(n_243),
.Y(n_2638)
);

OAI22xp33_ASAP7_75t_L g2639 ( 
.A1(n_2549),
.A2(n_2548),
.B1(n_2543),
.B2(n_2460),
.Y(n_2639)
);

OAI21xp5_ASAP7_75t_L g2640 ( 
.A1(n_2518),
.A2(n_244),
.B(n_245),
.Y(n_2640)
);

INVx1_ASAP7_75t_L g2641 ( 
.A(n_2535),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_2535),
.Y(n_2642)
);

OAI22xp33_ASAP7_75t_L g2643 ( 
.A1(n_2537),
.A2(n_249),
.B1(n_247),
.B2(n_248),
.Y(n_2643)
);

NAND2xp5_ASAP7_75t_L g2644 ( 
.A(n_2550),
.B(n_247),
.Y(n_2644)
);

A2O1A1Ixp33_ASAP7_75t_L g2645 ( 
.A1(n_2526),
.A2(n_251),
.B(n_248),
.C(n_250),
.Y(n_2645)
);

OAI221xp5_ASAP7_75t_SL g2646 ( 
.A1(n_2450),
.A2(n_253),
.B1(n_251),
.B2(n_252),
.C(n_255),
.Y(n_2646)
);

A2O1A1Ixp33_ASAP7_75t_L g2647 ( 
.A1(n_2496),
.A2(n_256),
.B(n_252),
.C(n_253),
.Y(n_2647)
);

OAI211xp5_ASAP7_75t_SL g2648 ( 
.A1(n_2470),
.A2(n_258),
.B(n_256),
.C(n_257),
.Y(n_2648)
);

AOI32xp33_ASAP7_75t_L g2649 ( 
.A1(n_2477),
.A2(n_260),
.A3(n_258),
.B1(n_259),
.B2(n_261),
.Y(n_2649)
);

OR2x2_ASAP7_75t_L g2650 ( 
.A(n_2576),
.B(n_262),
.Y(n_2650)
);

NOR2x1_ASAP7_75t_L g2651 ( 
.A(n_2583),
.B(n_262),
.Y(n_2651)
);

INVx1_ASAP7_75t_L g2652 ( 
.A(n_2503),
.Y(n_2652)
);

AOI221xp5_ASAP7_75t_SL g2653 ( 
.A1(n_2474),
.A2(n_265),
.B1(n_263),
.B2(n_264),
.C(n_266),
.Y(n_2653)
);

AOI221xp5_ASAP7_75t_L g2654 ( 
.A1(n_2507),
.A2(n_267),
.B1(n_263),
.B2(n_265),
.C(n_270),
.Y(n_2654)
);

AOI22xp33_ASAP7_75t_SL g2655 ( 
.A1(n_2448),
.A2(n_273),
.B1(n_271),
.B2(n_272),
.Y(n_2655)
);

OAI222xp33_ASAP7_75t_L g2656 ( 
.A1(n_2480),
.A2(n_272),
.B1(n_273),
.B2(n_276),
.C1(n_277),
.C2(n_278),
.Y(n_2656)
);

O2A1O1Ixp33_ASAP7_75t_L g2657 ( 
.A1(n_2536),
.A2(n_279),
.B(n_276),
.C(n_278),
.Y(n_2657)
);

AOI221xp5_ASAP7_75t_L g2658 ( 
.A1(n_2493),
.A2(n_281),
.B1(n_279),
.B2(n_280),
.C(n_282),
.Y(n_2658)
);

OAI21xp5_ASAP7_75t_SL g2659 ( 
.A1(n_2586),
.A2(n_280),
.B(n_281),
.Y(n_2659)
);

OAI22xp5_ASAP7_75t_L g2660 ( 
.A1(n_2590),
.A2(n_285),
.B1(n_282),
.B2(n_284),
.Y(n_2660)
);

OAI21xp33_ASAP7_75t_SL g2661 ( 
.A1(n_2476),
.A2(n_284),
.B(n_287),
.Y(n_2661)
);

NOR2x1_ASAP7_75t_L g2662 ( 
.A(n_2567),
.B(n_287),
.Y(n_2662)
);

AOI211x1_ASAP7_75t_L g2663 ( 
.A1(n_2523),
.A2(n_290),
.B(n_288),
.C(n_289),
.Y(n_2663)
);

AOI22xp33_ASAP7_75t_L g2664 ( 
.A1(n_2501),
.A2(n_1118),
.B1(n_1117),
.B2(n_1115),
.Y(n_2664)
);

AOI211xp5_ASAP7_75t_L g2665 ( 
.A1(n_2572),
.A2(n_291),
.B(n_288),
.C(n_289),
.Y(n_2665)
);

AOI322xp5_ASAP7_75t_L g2666 ( 
.A1(n_2500),
.A2(n_2569),
.A3(n_2579),
.B1(n_2575),
.B2(n_2585),
.C1(n_2566),
.C2(n_2488),
.Y(n_2666)
);

OAI211xp5_ASAP7_75t_SL g2667 ( 
.A1(n_2458),
.A2(n_295),
.B(n_293),
.C(n_294),
.Y(n_2667)
);

AOI221xp5_ASAP7_75t_L g2668 ( 
.A1(n_2541),
.A2(n_297),
.B1(n_293),
.B2(n_294),
.C(n_298),
.Y(n_2668)
);

AOI31xp33_ASAP7_75t_L g2669 ( 
.A1(n_2551),
.A2(n_2581),
.A3(n_2456),
.B(n_2540),
.Y(n_2669)
);

NAND2xp5_ASAP7_75t_L g2670 ( 
.A(n_2483),
.B(n_298),
.Y(n_2670)
);

INVx1_ASAP7_75t_L g2671 ( 
.A(n_2512),
.Y(n_2671)
);

O2A1O1Ixp33_ASAP7_75t_L g2672 ( 
.A1(n_2469),
.A2(n_301),
.B(n_299),
.C(n_300),
.Y(n_2672)
);

AOI32xp33_ASAP7_75t_L g2673 ( 
.A1(n_2514),
.A2(n_302),
.A3(n_300),
.B1(n_301),
.B2(n_303),
.Y(n_2673)
);

AOI22xp33_ASAP7_75t_L g2674 ( 
.A1(n_2478),
.A2(n_1115),
.B1(n_307),
.B2(n_302),
.Y(n_2674)
);

AOI321xp33_ASAP7_75t_L g2675 ( 
.A1(n_2487),
.A2(n_305),
.A3(n_307),
.B1(n_308),
.B2(n_309),
.C(n_310),
.Y(n_2675)
);

NAND2xp5_ASAP7_75t_L g2676 ( 
.A(n_2485),
.B(n_305),
.Y(n_2676)
);

AOI21xp33_ASAP7_75t_L g2677 ( 
.A1(n_2546),
.A2(n_308),
.B(n_309),
.Y(n_2677)
);

NAND2xp33_ASAP7_75t_L g2678 ( 
.A(n_2499),
.B(n_311),
.Y(n_2678)
);

OAI31xp33_ASAP7_75t_SL g2679 ( 
.A1(n_2570),
.A2(n_314),
.A3(n_312),
.B(n_313),
.Y(n_2679)
);

AOI22xp5_ASAP7_75t_L g2680 ( 
.A1(n_2615),
.A2(n_2475),
.B1(n_2563),
.B2(n_2506),
.Y(n_2680)
);

NAND2x1p5_ASAP7_75t_L g2681 ( 
.A(n_2595),
.B(n_2490),
.Y(n_2681)
);

INVx1_ASAP7_75t_L g2682 ( 
.A(n_2594),
.Y(n_2682)
);

INVxp67_ASAP7_75t_L g2683 ( 
.A(n_2651),
.Y(n_2683)
);

AND2x2_ASAP7_75t_L g2684 ( 
.A(n_2619),
.B(n_2525),
.Y(n_2684)
);

O2A1O1Ixp33_ASAP7_75t_L g2685 ( 
.A1(n_2638),
.A2(n_2471),
.B(n_2510),
.C(n_2577),
.Y(n_2685)
);

OAI22xp5_ASAP7_75t_L g2686 ( 
.A1(n_2606),
.A2(n_2562),
.B1(n_2489),
.B2(n_2516),
.Y(n_2686)
);

AOI22xp5_ASAP7_75t_SL g2687 ( 
.A1(n_2624),
.A2(n_2560),
.B1(n_2466),
.B2(n_2533),
.Y(n_2687)
);

AOI221x1_ASAP7_75t_L g2688 ( 
.A1(n_2610),
.A2(n_2508),
.B1(n_2513),
.B2(n_2479),
.C(n_2555),
.Y(n_2688)
);

AOI211xp5_ASAP7_75t_L g2689 ( 
.A1(n_2601),
.A2(n_2452),
.B(n_2464),
.C(n_2481),
.Y(n_2689)
);

AND2x2_ASAP7_75t_L g2690 ( 
.A(n_2623),
.B(n_2502),
.Y(n_2690)
);

AOI22xp33_ASAP7_75t_L g2691 ( 
.A1(n_2609),
.A2(n_2494),
.B1(n_2486),
.B2(n_2519),
.Y(n_2691)
);

INVx1_ASAP7_75t_L g2692 ( 
.A(n_2641),
.Y(n_2692)
);

O2A1O1Ixp33_ASAP7_75t_L g2693 ( 
.A1(n_2604),
.A2(n_2626),
.B(n_2657),
.C(n_2642),
.Y(n_2693)
);

INVx1_ASAP7_75t_L g2694 ( 
.A(n_2621),
.Y(n_2694)
);

INVx2_ASAP7_75t_SL g2695 ( 
.A(n_2650),
.Y(n_2695)
);

AOI32xp33_ASAP7_75t_L g2696 ( 
.A1(n_2671),
.A2(n_2528),
.A3(n_2509),
.B1(n_2527),
.B2(n_2465),
.Y(n_2696)
);

OAI22xp5_ASAP7_75t_L g2697 ( 
.A1(n_2655),
.A2(n_2451),
.B1(n_2459),
.B2(n_2457),
.Y(n_2697)
);

INVx1_ASAP7_75t_L g2698 ( 
.A(n_2621),
.Y(n_2698)
);

AOI21xp5_ASAP7_75t_L g2699 ( 
.A1(n_2592),
.A2(n_2524),
.B(n_2578),
.Y(n_2699)
);

AOI22xp5_ASAP7_75t_L g2700 ( 
.A1(n_2600),
.A2(n_2580),
.B1(n_2472),
.B2(n_2573),
.Y(n_2700)
);

INVx2_ASAP7_75t_L g2701 ( 
.A(n_2618),
.Y(n_2701)
);

INVx1_ASAP7_75t_L g2702 ( 
.A(n_2603),
.Y(n_2702)
);

INVx1_ASAP7_75t_L g2703 ( 
.A(n_2605),
.Y(n_2703)
);

OR2x2_ASAP7_75t_L g2704 ( 
.A(n_2620),
.B(n_2462),
.Y(n_2704)
);

AND2x2_ASAP7_75t_L g2705 ( 
.A(n_2629),
.B(n_2558),
.Y(n_2705)
);

OAI211xp5_ASAP7_75t_SL g2706 ( 
.A1(n_2599),
.A2(n_2633),
.B(n_2661),
.C(n_2613),
.Y(n_2706)
);

AOI221x1_ASAP7_75t_SL g2707 ( 
.A1(n_2639),
.A2(n_2521),
.B1(n_2584),
.B2(n_315),
.C(n_313),
.Y(n_2707)
);

INVx1_ASAP7_75t_SL g2708 ( 
.A(n_2670),
.Y(n_2708)
);

O2A1O1Ixp33_ASAP7_75t_L g2709 ( 
.A1(n_2659),
.A2(n_317),
.B(n_314),
.C(n_316),
.Y(n_2709)
);

AND2x2_ASAP7_75t_L g2710 ( 
.A(n_2640),
.B(n_316),
.Y(n_2710)
);

INVx1_ASAP7_75t_L g2711 ( 
.A(n_2596),
.Y(n_2711)
);

OAI21xp33_ASAP7_75t_L g2712 ( 
.A1(n_2679),
.A2(n_318),
.B(n_319),
.Y(n_2712)
);

AOI21xp5_ASAP7_75t_L g2713 ( 
.A1(n_2627),
.A2(n_318),
.B(n_319),
.Y(n_2713)
);

AOI21xp5_ASAP7_75t_L g2714 ( 
.A1(n_2672),
.A2(n_320),
.B(n_321),
.Y(n_2714)
);

O2A1O1Ixp33_ASAP7_75t_L g2715 ( 
.A1(n_2648),
.A2(n_323),
.B(n_320),
.C(n_322),
.Y(n_2715)
);

OAI22xp5_ASAP7_75t_L g2716 ( 
.A1(n_2646),
.A2(n_326),
.B1(n_324),
.B2(n_325),
.Y(n_2716)
);

INVx1_ASAP7_75t_L g2717 ( 
.A(n_2612),
.Y(n_2717)
);

AOI22xp5_ASAP7_75t_L g2718 ( 
.A1(n_2597),
.A2(n_327),
.B1(n_325),
.B2(n_326),
.Y(n_2718)
);

AND2x2_ASAP7_75t_L g2719 ( 
.A(n_2635),
.B(n_328),
.Y(n_2719)
);

OAI21xp5_ASAP7_75t_L g2720 ( 
.A1(n_2602),
.A2(n_328),
.B(n_330),
.Y(n_2720)
);

AOI211xp5_ASAP7_75t_L g2721 ( 
.A1(n_2656),
.A2(n_332),
.B(n_330),
.C(n_331),
.Y(n_2721)
);

AOI21xp33_ASAP7_75t_L g2722 ( 
.A1(n_2625),
.A2(n_333),
.B(n_334),
.Y(n_2722)
);

OAI22xp5_ASAP7_75t_L g2723 ( 
.A1(n_2614),
.A2(n_335),
.B1(n_333),
.B2(n_334),
.Y(n_2723)
);

INVx2_ASAP7_75t_L g2724 ( 
.A(n_2663),
.Y(n_2724)
);

OAI21xp5_ASAP7_75t_L g2725 ( 
.A1(n_2662),
.A2(n_335),
.B(n_336),
.Y(n_2725)
);

AOI22xp33_ASAP7_75t_L g2726 ( 
.A1(n_2652),
.A2(n_339),
.B1(n_337),
.B2(n_338),
.Y(n_2726)
);

INVx1_ASAP7_75t_L g2727 ( 
.A(n_2611),
.Y(n_2727)
);

BUFx2_ASAP7_75t_L g2728 ( 
.A(n_2622),
.Y(n_2728)
);

OAI221xp5_ASAP7_75t_L g2729 ( 
.A1(n_2665),
.A2(n_339),
.B1(n_340),
.B2(n_341),
.C(n_342),
.Y(n_2729)
);

AOI21xp33_ASAP7_75t_L g2730 ( 
.A1(n_2678),
.A2(n_340),
.B(n_342),
.Y(n_2730)
);

AOI221x1_ASAP7_75t_L g2731 ( 
.A1(n_2607),
.A2(n_2616),
.B1(n_2660),
.B2(n_2677),
.C(n_2645),
.Y(n_2731)
);

OAI211xp5_ASAP7_75t_L g2732 ( 
.A1(n_2654),
.A2(n_345),
.B(n_343),
.C(n_344),
.Y(n_2732)
);

INVxp67_ASAP7_75t_L g2733 ( 
.A(n_2637),
.Y(n_2733)
);

AOI321xp33_ASAP7_75t_L g2734 ( 
.A1(n_2628),
.A2(n_343),
.A3(n_344),
.B1(n_345),
.B2(n_346),
.C(n_347),
.Y(n_2734)
);

INVx2_ASAP7_75t_SL g2735 ( 
.A(n_2676),
.Y(n_2735)
);

O2A1O1Ixp33_ASAP7_75t_L g2736 ( 
.A1(n_2647),
.A2(n_348),
.B(n_346),
.C(n_347),
.Y(n_2736)
);

NOR3xp33_ASAP7_75t_L g2737 ( 
.A(n_2643),
.B(n_348),
.C(n_350),
.Y(n_2737)
);

NAND2x1p5_ASAP7_75t_L g2738 ( 
.A(n_2717),
.B(n_2598),
.Y(n_2738)
);

AOI22xp33_ASAP7_75t_L g2739 ( 
.A1(n_2703),
.A2(n_2631),
.B1(n_2630),
.B2(n_2674),
.Y(n_2739)
);

AOI22xp5_ASAP7_75t_L g2740 ( 
.A1(n_2702),
.A2(n_2608),
.B1(n_2668),
.B2(n_2658),
.Y(n_2740)
);

XNOR2xp5_ASAP7_75t_L g2741 ( 
.A(n_2680),
.B(n_2593),
.Y(n_2741)
);

INVx1_ASAP7_75t_L g2742 ( 
.A(n_2711),
.Y(n_2742)
);

XOR2xp5_ASAP7_75t_L g2743 ( 
.A(n_2680),
.B(n_2644),
.Y(n_2743)
);

AOI32xp33_ASAP7_75t_L g2744 ( 
.A1(n_2684),
.A2(n_2692),
.A3(n_2706),
.B1(n_2690),
.B2(n_2727),
.Y(n_2744)
);

XNOR2x1_ASAP7_75t_L g2745 ( 
.A(n_2682),
.B(n_2701),
.Y(n_2745)
);

OAI22x1_ASAP7_75t_SL g2746 ( 
.A1(n_2695),
.A2(n_2653),
.B1(n_2666),
.B2(n_2669),
.Y(n_2746)
);

NOR2xp33_ASAP7_75t_R g2747 ( 
.A(n_2694),
.B(n_2634),
.Y(n_2747)
);

OAI221xp5_ASAP7_75t_SL g2748 ( 
.A1(n_2693),
.A2(n_2683),
.B1(n_2696),
.B2(n_2689),
.C(n_2733),
.Y(n_2748)
);

AOI22xp5_ASAP7_75t_L g2749 ( 
.A1(n_2686),
.A2(n_2667),
.B1(n_2664),
.B2(n_2617),
.Y(n_2749)
);

AOI22xp5_ASAP7_75t_L g2750 ( 
.A1(n_2712),
.A2(n_2669),
.B1(n_2649),
.B2(n_2673),
.Y(n_2750)
);

CKINVDCx6p67_ASAP7_75t_R g2751 ( 
.A(n_2719),
.Y(n_2751)
);

OAI21xp5_ASAP7_75t_L g2752 ( 
.A1(n_2709),
.A2(n_2632),
.B(n_2675),
.Y(n_2752)
);

OAI32xp33_ASAP7_75t_L g2753 ( 
.A1(n_2681),
.A2(n_2636),
.A3(n_351),
.B1(n_352),
.B2(n_353),
.Y(n_2753)
);

AOI22xp5_ASAP7_75t_L g2754 ( 
.A1(n_2735),
.A2(n_353),
.B1(n_350),
.B2(n_352),
.Y(n_2754)
);

INVx1_ASAP7_75t_L g2755 ( 
.A(n_2698),
.Y(n_2755)
);

INVx1_ASAP7_75t_L g2756 ( 
.A(n_2728),
.Y(n_2756)
);

AND2x2_ASAP7_75t_L g2757 ( 
.A(n_2687),
.B(n_354),
.Y(n_2757)
);

NAND2xp5_ASAP7_75t_L g2758 ( 
.A(n_2724),
.B(n_354),
.Y(n_2758)
);

OAI22xp5_ASAP7_75t_L g2759 ( 
.A1(n_2718),
.A2(n_2726),
.B1(n_2729),
.B2(n_2721),
.Y(n_2759)
);

AOI22xp5_ASAP7_75t_L g2760 ( 
.A1(n_2708),
.A2(n_2705),
.B1(n_2710),
.B2(n_2716),
.Y(n_2760)
);

INVx1_ASAP7_75t_L g2761 ( 
.A(n_2715),
.Y(n_2761)
);

NAND2xp5_ASAP7_75t_L g2762 ( 
.A(n_2707),
.B(n_355),
.Y(n_2762)
);

NAND2xp5_ASAP7_75t_L g2763 ( 
.A(n_2714),
.B(n_356),
.Y(n_2763)
);

AOI221xp5_ASAP7_75t_SL g2764 ( 
.A1(n_2685),
.A2(n_357),
.B1(n_358),
.B2(n_359),
.C(n_361),
.Y(n_2764)
);

AOI21xp33_ASAP7_75t_L g2765 ( 
.A1(n_2704),
.A2(n_359),
.B(n_364),
.Y(n_2765)
);

AOI211xp5_ASAP7_75t_SL g2766 ( 
.A1(n_2730),
.A2(n_368),
.B(n_365),
.C(n_367),
.Y(n_2766)
);

INVx1_ASAP7_75t_L g2767 ( 
.A(n_2734),
.Y(n_2767)
);

AOI21xp5_ASAP7_75t_L g2768 ( 
.A1(n_2713),
.A2(n_367),
.B(n_368),
.Y(n_2768)
);

OAI21xp33_ASAP7_75t_L g2769 ( 
.A1(n_2720),
.A2(n_369),
.B(n_370),
.Y(n_2769)
);

INVx3_ASAP7_75t_L g2770 ( 
.A(n_2722),
.Y(n_2770)
);

NAND3xp33_ASAP7_75t_L g2771 ( 
.A(n_2718),
.B(n_370),
.C(n_371),
.Y(n_2771)
);

AOI31xp33_ASAP7_75t_L g2772 ( 
.A1(n_2725),
.A2(n_2723),
.A3(n_2732),
.B(n_2699),
.Y(n_2772)
);

OAI22xp33_ASAP7_75t_SL g2773 ( 
.A1(n_2697),
.A2(n_373),
.B1(n_371),
.B2(n_372),
.Y(n_2773)
);

NOR2xp67_ASAP7_75t_L g2774 ( 
.A(n_2756),
.B(n_2700),
.Y(n_2774)
);

AO22x2_ASAP7_75t_L g2775 ( 
.A1(n_2745),
.A2(n_2757),
.B1(n_2767),
.B2(n_2761),
.Y(n_2775)
);

INVx1_ASAP7_75t_L g2776 ( 
.A(n_2751),
.Y(n_2776)
);

OAI22xp33_ASAP7_75t_L g2777 ( 
.A1(n_2742),
.A2(n_2688),
.B1(n_2731),
.B2(n_2700),
.Y(n_2777)
);

INVx2_ASAP7_75t_L g2778 ( 
.A(n_2738),
.Y(n_2778)
);

INVx1_ASAP7_75t_L g2779 ( 
.A(n_2746),
.Y(n_2779)
);

INVx1_ASAP7_75t_L g2780 ( 
.A(n_2762),
.Y(n_2780)
);

INVx1_ASAP7_75t_L g2781 ( 
.A(n_2763),
.Y(n_2781)
);

INVx1_ASAP7_75t_L g2782 ( 
.A(n_2773),
.Y(n_2782)
);

INVxp67_ASAP7_75t_L g2783 ( 
.A(n_2758),
.Y(n_2783)
);

NOR2x1_ASAP7_75t_L g2784 ( 
.A(n_2755),
.B(n_2736),
.Y(n_2784)
);

INVx1_ASAP7_75t_L g2785 ( 
.A(n_2743),
.Y(n_2785)
);

AND2x2_ASAP7_75t_L g2786 ( 
.A(n_2764),
.B(n_2737),
.Y(n_2786)
);

INVx2_ASAP7_75t_L g2787 ( 
.A(n_2770),
.Y(n_2787)
);

OAI22xp33_ASAP7_75t_L g2788 ( 
.A1(n_2740),
.A2(n_2691),
.B1(n_376),
.B2(n_372),
.Y(n_2788)
);

INVx2_ASAP7_75t_L g2789 ( 
.A(n_2770),
.Y(n_2789)
);

NOR3xp33_ASAP7_75t_L g2790 ( 
.A(n_2748),
.B(n_375),
.C(n_377),
.Y(n_2790)
);

NOR2x1_ASAP7_75t_L g2791 ( 
.A(n_2771),
.B(n_375),
.Y(n_2791)
);

INVx1_ASAP7_75t_L g2792 ( 
.A(n_2750),
.Y(n_2792)
);

NOR2x1_ASAP7_75t_L g2793 ( 
.A(n_2741),
.B(n_377),
.Y(n_2793)
);

AOI22xp5_ASAP7_75t_L g2794 ( 
.A1(n_2780),
.A2(n_2769),
.B1(n_2759),
.B2(n_2760),
.Y(n_2794)
);

NAND2xp5_ASAP7_75t_L g2795 ( 
.A(n_2774),
.B(n_2766),
.Y(n_2795)
);

XNOR2xp5_ASAP7_75t_L g2796 ( 
.A(n_2775),
.B(n_2752),
.Y(n_2796)
);

NAND4xp75_ASAP7_75t_L g2797 ( 
.A(n_2784),
.B(n_2765),
.C(n_2768),
.D(n_2749),
.Y(n_2797)
);

NOR2xp33_ASAP7_75t_L g2798 ( 
.A(n_2777),
.B(n_2753),
.Y(n_2798)
);

NAND4xp75_ASAP7_75t_L g2799 ( 
.A(n_2779),
.B(n_2754),
.C(n_2744),
.D(n_2747),
.Y(n_2799)
);

INVx1_ASAP7_75t_L g2800 ( 
.A(n_2775),
.Y(n_2800)
);

XOR2x1_ASAP7_75t_L g2801 ( 
.A(n_2776),
.B(n_2772),
.Y(n_2801)
);

NOR2x1_ASAP7_75t_L g2802 ( 
.A(n_2778),
.B(n_2739),
.Y(n_2802)
);

NOR2xp67_ASAP7_75t_L g2803 ( 
.A(n_2782),
.B(n_378),
.Y(n_2803)
);

INVxp67_ASAP7_75t_SL g2804 ( 
.A(n_2793),
.Y(n_2804)
);

AOI22xp5_ASAP7_75t_L g2805 ( 
.A1(n_2787),
.A2(n_380),
.B1(n_378),
.B2(n_379),
.Y(n_2805)
);

INVx1_ASAP7_75t_L g2806 ( 
.A(n_2786),
.Y(n_2806)
);

NOR2x1_ASAP7_75t_L g2807 ( 
.A(n_2792),
.B(n_2789),
.Y(n_2807)
);

INVx1_ASAP7_75t_L g2808 ( 
.A(n_2791),
.Y(n_2808)
);

HB1xp67_ASAP7_75t_L g2809 ( 
.A(n_2785),
.Y(n_2809)
);

INVx1_ASAP7_75t_SL g2810 ( 
.A(n_2781),
.Y(n_2810)
);

XOR2xp5_ASAP7_75t_L g2811 ( 
.A(n_2796),
.B(n_2788),
.Y(n_2811)
);

NOR3xp33_ASAP7_75t_L g2812 ( 
.A(n_2800),
.B(n_2783),
.C(n_2790),
.Y(n_2812)
);

OAI22xp33_ASAP7_75t_SL g2813 ( 
.A1(n_2795),
.A2(n_382),
.B1(n_380),
.B2(n_381),
.Y(n_2813)
);

NAND2xp5_ASAP7_75t_L g2814 ( 
.A(n_2807),
.B(n_381),
.Y(n_2814)
);

AOI22xp33_ASAP7_75t_L g2815 ( 
.A1(n_2804),
.A2(n_390),
.B1(n_386),
.B2(n_388),
.Y(n_2815)
);

AOI22xp5_ASAP7_75t_L g2816 ( 
.A1(n_2798),
.A2(n_391),
.B1(n_386),
.B2(n_390),
.Y(n_2816)
);

OAI321xp33_ASAP7_75t_L g2817 ( 
.A1(n_2806),
.A2(n_391),
.A3(n_392),
.B1(n_393),
.B2(n_394),
.C(n_395),
.Y(n_2817)
);

NOR3xp33_ASAP7_75t_L g2818 ( 
.A(n_2809),
.B(n_392),
.C(n_394),
.Y(n_2818)
);

INVx1_ASAP7_75t_SL g2819 ( 
.A(n_2810),
.Y(n_2819)
);

AOI222xp33_ASAP7_75t_L g2820 ( 
.A1(n_2803),
.A2(n_395),
.B1(n_396),
.B2(n_397),
.C1(n_398),
.C2(n_399),
.Y(n_2820)
);

INVx1_ASAP7_75t_L g2821 ( 
.A(n_2802),
.Y(n_2821)
);

AOI211xp5_ASAP7_75t_L g2822 ( 
.A1(n_2808),
.A2(n_402),
.B(n_396),
.C(n_397),
.Y(n_2822)
);

OAI22xp5_ASAP7_75t_L g2823 ( 
.A1(n_2794),
.A2(n_404),
.B1(n_402),
.B2(n_403),
.Y(n_2823)
);

AOI22xp5_ASAP7_75t_L g2824 ( 
.A1(n_2799),
.A2(n_405),
.B1(n_403),
.B2(n_404),
.Y(n_2824)
);

OAI221xp5_ASAP7_75t_L g2825 ( 
.A1(n_2805),
.A2(n_406),
.B1(n_407),
.B2(n_408),
.C(n_409),
.Y(n_2825)
);

NOR2xp67_ASAP7_75t_L g2826 ( 
.A(n_2801),
.B(n_408),
.Y(n_2826)
);

AOI22xp5_ASAP7_75t_L g2827 ( 
.A1(n_2797),
.A2(n_410),
.B1(n_412),
.B2(n_413),
.Y(n_2827)
);

OA22x2_ASAP7_75t_L g2828 ( 
.A1(n_2794),
.A2(n_414),
.B1(n_415),
.B2(n_416),
.Y(n_2828)
);

OR3x2_ASAP7_75t_L g2829 ( 
.A(n_2800),
.B(n_417),
.C(n_418),
.Y(n_2829)
);

XNOR2xp5_ASAP7_75t_L g2830 ( 
.A(n_2811),
.B(n_418),
.Y(n_2830)
);

OAI22xp5_ASAP7_75t_SL g2831 ( 
.A1(n_2819),
.A2(n_419),
.B1(n_422),
.B2(n_424),
.Y(n_2831)
);

INVx1_ASAP7_75t_L g2832 ( 
.A(n_2821),
.Y(n_2832)
);

XNOR2x1_ASAP7_75t_L g2833 ( 
.A(n_2826),
.B(n_419),
.Y(n_2833)
);

XNOR2xp5_ASAP7_75t_L g2834 ( 
.A(n_2824),
.B(n_422),
.Y(n_2834)
);

XNOR2x1_ASAP7_75t_L g2835 ( 
.A(n_2828),
.B(n_425),
.Y(n_2835)
);

OR2x2_ASAP7_75t_L g2836 ( 
.A(n_2814),
.B(n_425),
.Y(n_2836)
);

INVx2_ASAP7_75t_L g2837 ( 
.A(n_2829),
.Y(n_2837)
);

OAI22xp5_ASAP7_75t_L g2838 ( 
.A1(n_2816),
.A2(n_426),
.B1(n_427),
.B2(n_428),
.Y(n_2838)
);

AND2x4_ASAP7_75t_L g2839 ( 
.A(n_2812),
.B(n_428),
.Y(n_2839)
);

OAI21xp5_ASAP7_75t_L g2840 ( 
.A1(n_2820),
.A2(n_429),
.B(n_430),
.Y(n_2840)
);

NOR2xp67_ASAP7_75t_L g2841 ( 
.A(n_2817),
.B(n_429),
.Y(n_2841)
);

AOI21xp5_ASAP7_75t_L g2842 ( 
.A1(n_2813),
.A2(n_2823),
.B(n_2825),
.Y(n_2842)
);

AND3x4_ASAP7_75t_L g2843 ( 
.A(n_2818),
.B(n_430),
.C(n_431),
.Y(n_2843)
);

NOR2xp67_ASAP7_75t_L g2844 ( 
.A(n_2827),
.B(n_431),
.Y(n_2844)
);

NAND3x1_ASAP7_75t_L g2845 ( 
.A(n_2822),
.B(n_432),
.C(n_433),
.Y(n_2845)
);

INVx1_ASAP7_75t_L g2846 ( 
.A(n_2815),
.Y(n_2846)
);

INVx1_ASAP7_75t_L g2847 ( 
.A(n_2821),
.Y(n_2847)
);

INVx2_ASAP7_75t_L g2848 ( 
.A(n_2821),
.Y(n_2848)
);

OR2x6_ASAP7_75t_L g2849 ( 
.A(n_2821),
.B(n_432),
.Y(n_2849)
);

INVxp33_ASAP7_75t_SL g2850 ( 
.A(n_2811),
.Y(n_2850)
);

INVx3_ASAP7_75t_L g2851 ( 
.A(n_2848),
.Y(n_2851)
);

AOI22xp5_ASAP7_75t_L g2852 ( 
.A1(n_2832),
.A2(n_2847),
.B1(n_2850),
.B2(n_2837),
.Y(n_2852)
);

BUFx12f_ASAP7_75t_L g2853 ( 
.A(n_2839),
.Y(n_2853)
);

INVx2_ASAP7_75t_L g2854 ( 
.A(n_2833),
.Y(n_2854)
);

XOR2x1_ASAP7_75t_L g2855 ( 
.A(n_2835),
.B(n_434),
.Y(n_2855)
);

NAND2xp33_ASAP7_75t_SL g2856 ( 
.A(n_2831),
.B(n_434),
.Y(n_2856)
);

XOR2x2_ASAP7_75t_L g2857 ( 
.A(n_2830),
.B(n_435),
.Y(n_2857)
);

NOR2xp33_ASAP7_75t_L g2858 ( 
.A(n_2849),
.B(n_435),
.Y(n_2858)
);

INVx1_ASAP7_75t_SL g2859 ( 
.A(n_2836),
.Y(n_2859)
);

INVx3_ASAP7_75t_L g2860 ( 
.A(n_2849),
.Y(n_2860)
);

INVx1_ASAP7_75t_L g2861 ( 
.A(n_2841),
.Y(n_2861)
);

NAND2xp5_ASAP7_75t_L g2862 ( 
.A(n_2844),
.B(n_436),
.Y(n_2862)
);

INVx3_ASAP7_75t_L g2863 ( 
.A(n_2845),
.Y(n_2863)
);

OAI22x1_ASAP7_75t_L g2864 ( 
.A1(n_2843),
.A2(n_436),
.B1(n_437),
.B2(n_438),
.Y(n_2864)
);

NAND2xp5_ASAP7_75t_L g2865 ( 
.A(n_2840),
.B(n_438),
.Y(n_2865)
);

AO21x2_ASAP7_75t_L g2866 ( 
.A1(n_2852),
.A2(n_2842),
.B(n_2834),
.Y(n_2866)
);

INVx1_ASAP7_75t_L g2867 ( 
.A(n_2851),
.Y(n_2867)
);

INVx2_ASAP7_75t_L g2868 ( 
.A(n_2855),
.Y(n_2868)
);

OAI22x1_ASAP7_75t_L g2869 ( 
.A1(n_2858),
.A2(n_2846),
.B1(n_2838),
.B2(n_442),
.Y(n_2869)
);

CKINVDCx20_ASAP7_75t_R g2870 ( 
.A(n_2857),
.Y(n_2870)
);

HB1xp67_ASAP7_75t_L g2871 ( 
.A(n_2864),
.Y(n_2871)
);

XNOR2xp5_ASAP7_75t_L g2872 ( 
.A(n_2859),
.B(n_439),
.Y(n_2872)
);

AOI22xp5_ASAP7_75t_L g2873 ( 
.A1(n_2861),
.A2(n_440),
.B1(n_443),
.B2(n_444),
.Y(n_2873)
);

AOI221xp5_ASAP7_75t_L g2874 ( 
.A1(n_2856),
.A2(n_2863),
.B1(n_2854),
.B2(n_2860),
.C(n_2865),
.Y(n_2874)
);

NOR2xp33_ASAP7_75t_L g2875 ( 
.A(n_2853),
.B(n_440),
.Y(n_2875)
);

OA21x2_ASAP7_75t_L g2876 ( 
.A1(n_2862),
.A2(n_444),
.B(n_445),
.Y(n_2876)
);

INVx1_ASAP7_75t_L g2877 ( 
.A(n_2851),
.Y(n_2877)
);

INVx1_ASAP7_75t_SL g2878 ( 
.A(n_2851),
.Y(n_2878)
);

INVx1_ASAP7_75t_L g2879 ( 
.A(n_2851),
.Y(n_2879)
);

AOI22xp5_ASAP7_75t_L g2880 ( 
.A1(n_2878),
.A2(n_445),
.B1(n_446),
.B2(n_447),
.Y(n_2880)
);

OAI22xp5_ASAP7_75t_SL g2881 ( 
.A1(n_2870),
.A2(n_446),
.B1(n_448),
.B2(n_449),
.Y(n_2881)
);

AOI22xp5_ASAP7_75t_L g2882 ( 
.A1(n_2867),
.A2(n_450),
.B1(n_451),
.B2(n_452),
.Y(n_2882)
);

INVxp67_ASAP7_75t_L g2883 ( 
.A(n_2868),
.Y(n_2883)
);

OAI211xp5_ASAP7_75t_L g2884 ( 
.A1(n_2874),
.A2(n_450),
.B(n_453),
.C(n_454),
.Y(n_2884)
);

XOR2xp5_ASAP7_75t_L g2885 ( 
.A(n_2877),
.B(n_453),
.Y(n_2885)
);

XOR2xp5_ASAP7_75t_L g2886 ( 
.A(n_2879),
.B(n_455),
.Y(n_2886)
);

INVx1_ASAP7_75t_L g2887 ( 
.A(n_2872),
.Y(n_2887)
);

OAI22xp5_ASAP7_75t_L g2888 ( 
.A1(n_2871),
.A2(n_455),
.B1(n_456),
.B2(n_457),
.Y(n_2888)
);

OAI31xp33_ASAP7_75t_L g2889 ( 
.A1(n_2875),
.A2(n_457),
.A3(n_458),
.B(n_459),
.Y(n_2889)
);

AND3x1_ASAP7_75t_L g2890 ( 
.A(n_2873),
.B(n_461),
.C(n_462),
.Y(n_2890)
);

INVx1_ASAP7_75t_L g2891 ( 
.A(n_2876),
.Y(n_2891)
);

NAND2x1p5_ASAP7_75t_L g2892 ( 
.A(n_2866),
.B(n_462),
.Y(n_2892)
);

OAI22xp5_ASAP7_75t_SL g2893 ( 
.A1(n_2869),
.A2(n_464),
.B1(n_466),
.B2(n_467),
.Y(n_2893)
);

OAI21xp5_ASAP7_75t_L g2894 ( 
.A1(n_2878),
.A2(n_466),
.B(n_467),
.Y(n_2894)
);

NAND3xp33_ASAP7_75t_L g2895 ( 
.A(n_2883),
.B(n_468),
.C(n_469),
.Y(n_2895)
);

OAI22xp5_ASAP7_75t_SL g2896 ( 
.A1(n_2893),
.A2(n_468),
.B1(n_469),
.B2(n_471),
.Y(n_2896)
);

BUFx2_ASAP7_75t_L g2897 ( 
.A(n_2892),
.Y(n_2897)
);

INVx2_ASAP7_75t_L g2898 ( 
.A(n_2891),
.Y(n_2898)
);

INVxp33_ASAP7_75t_L g2899 ( 
.A(n_2885),
.Y(n_2899)
);

CKINVDCx20_ASAP7_75t_R g2900 ( 
.A(n_2887),
.Y(n_2900)
);

XNOR2x1_ASAP7_75t_L g2901 ( 
.A(n_2890),
.B(n_472),
.Y(n_2901)
);

INVx1_ASAP7_75t_L g2902 ( 
.A(n_2886),
.Y(n_2902)
);

OAI22xp5_ASAP7_75t_SL g2903 ( 
.A1(n_2881),
.A2(n_474),
.B1(n_475),
.B2(n_476),
.Y(n_2903)
);

CKINVDCx20_ASAP7_75t_R g2904 ( 
.A(n_2894),
.Y(n_2904)
);

AOI22x1_ASAP7_75t_L g2905 ( 
.A1(n_2884),
.A2(n_475),
.B1(n_477),
.B2(n_479),
.Y(n_2905)
);

BUFx2_ASAP7_75t_L g2906 ( 
.A(n_2880),
.Y(n_2906)
);

OAI22xp5_ASAP7_75t_SL g2907 ( 
.A1(n_2900),
.A2(n_2897),
.B1(n_2904),
.B2(n_2898),
.Y(n_2907)
);

INVx1_ASAP7_75t_L g2908 ( 
.A(n_2901),
.Y(n_2908)
);

OAI22xp5_ASAP7_75t_SL g2909 ( 
.A1(n_2896),
.A2(n_2888),
.B1(n_2882),
.B2(n_2889),
.Y(n_2909)
);

OA22x2_ASAP7_75t_L g2910 ( 
.A1(n_2903),
.A2(n_477),
.B1(n_480),
.B2(n_481),
.Y(n_2910)
);

OAI22xp5_ASAP7_75t_SL g2911 ( 
.A1(n_2899),
.A2(n_480),
.B1(n_481),
.B2(n_482),
.Y(n_2911)
);

NAND2xp5_ASAP7_75t_L g2912 ( 
.A(n_2902),
.B(n_482),
.Y(n_2912)
);

OAI21xp33_ASAP7_75t_L g2913 ( 
.A1(n_2895),
.A2(n_485),
.B(n_486),
.Y(n_2913)
);

OAI22xp33_ASAP7_75t_L g2914 ( 
.A1(n_2906),
.A2(n_485),
.B1(n_487),
.B2(n_488),
.Y(n_2914)
);

AOI21xp33_ASAP7_75t_SL g2915 ( 
.A1(n_2905),
.A2(n_487),
.B(n_488),
.Y(n_2915)
);

OAI22xp5_ASAP7_75t_L g2916 ( 
.A1(n_2900),
.A2(n_489),
.B1(n_490),
.B2(n_492),
.Y(n_2916)
);

HB1xp67_ASAP7_75t_L g2917 ( 
.A(n_2898),
.Y(n_2917)
);

AOI21xp5_ASAP7_75t_L g2918 ( 
.A1(n_2907),
.A2(n_489),
.B(n_493),
.Y(n_2918)
);

OAI21xp5_ASAP7_75t_L g2919 ( 
.A1(n_2917),
.A2(n_495),
.B(n_496),
.Y(n_2919)
);

OAI22xp5_ASAP7_75t_L g2920 ( 
.A1(n_2908),
.A2(n_495),
.B1(n_496),
.B2(n_497),
.Y(n_2920)
);

NAND2xp5_ASAP7_75t_L g2921 ( 
.A(n_2915),
.B(n_497),
.Y(n_2921)
);

INVx1_ASAP7_75t_L g2922 ( 
.A(n_2912),
.Y(n_2922)
);

OAI22xp5_ASAP7_75t_L g2923 ( 
.A1(n_2910),
.A2(n_498),
.B1(n_499),
.B2(n_500),
.Y(n_2923)
);

AOI21xp5_ASAP7_75t_L g2924 ( 
.A1(n_2909),
.A2(n_498),
.B(n_499),
.Y(n_2924)
);

OA22x2_ASAP7_75t_L g2925 ( 
.A1(n_2913),
.A2(n_501),
.B1(n_502),
.B2(n_503),
.Y(n_2925)
);

XNOR2xp5_ASAP7_75t_L g2926 ( 
.A(n_2911),
.B(n_502),
.Y(n_2926)
);

AOI21xp5_ASAP7_75t_SL g2927 ( 
.A1(n_2916),
.A2(n_503),
.B(n_505),
.Y(n_2927)
);

AOI222xp33_ASAP7_75t_L g2928 ( 
.A1(n_2923),
.A2(n_2914),
.B1(n_508),
.B2(n_509),
.C1(n_510),
.C2(n_511),
.Y(n_2928)
);

AOI21xp33_ASAP7_75t_L g2929 ( 
.A1(n_2922),
.A2(n_506),
.B(n_508),
.Y(n_2929)
);

AOI221xp5_ASAP7_75t_L g2930 ( 
.A1(n_2918),
.A2(n_506),
.B1(n_509),
.B2(n_511),
.C(n_512),
.Y(n_2930)
);

AOI21xp33_ASAP7_75t_SL g2931 ( 
.A1(n_2926),
.A2(n_512),
.B(n_513),
.Y(n_2931)
);

AOI22xp33_ASAP7_75t_L g2932 ( 
.A1(n_2930),
.A2(n_2925),
.B1(n_2921),
.B2(n_2924),
.Y(n_2932)
);

OAI21xp5_ASAP7_75t_L g2933 ( 
.A1(n_2932),
.A2(n_2931),
.B(n_2927),
.Y(n_2933)
);

AOI21xp33_ASAP7_75t_L g2934 ( 
.A1(n_2933),
.A2(n_2928),
.B(n_2919),
.Y(n_2934)
);

AOI211xp5_ASAP7_75t_L g2935 ( 
.A1(n_2934),
.A2(n_2929),
.B(n_2920),
.C(n_516),
.Y(n_2935)
);


endmodule