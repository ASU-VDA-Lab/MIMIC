module fake_jpeg_21593_n_242 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_242);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_242;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_207;
wire n_155;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_213;
wire n_153;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx16f_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

INVx13_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_3),
.B(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_16),
.B(n_6),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_32),
.B(n_16),
.Y(n_46)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_34),
.Y(n_77)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_37),
.Y(n_75)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx4_ASAP7_75t_SL g42 ( 
.A(n_26),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_15),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_46),
.B(n_48),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_45),
.A2(n_20),
.B1(n_19),
.B2(n_27),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_47),
.A2(n_50),
.B1(n_70),
.B2(n_72),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_32),
.B(n_19),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_45),
.A2(n_20),
.B1(n_27),
.B2(n_23),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_25),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_52),
.B(n_54),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_17),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_53),
.B(n_63),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_35),
.B(n_25),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_14),
.C(n_28),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_55),
.B(n_40),
.C(n_43),
.Y(n_78)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_57),
.Y(n_82)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_33),
.B(n_24),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_59),
.B(n_30),
.Y(n_90)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_61),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_17),
.Y(n_63)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_69),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_39),
.B(n_14),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_42),
.A2(n_20),
.B1(n_23),
.B2(n_24),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_40),
.B(n_14),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_15),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_42),
.A2(n_21),
.B1(n_29),
.B2(n_30),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_34),
.Y(n_73)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_42),
.A2(n_21),
.B1(n_29),
.B2(n_30),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_74),
.A2(n_22),
.B1(n_44),
.B2(n_28),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_78),
.B(n_105),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_57),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_80),
.B(n_90),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_85),
.Y(n_133)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_86),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_55),
.B(n_38),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_87),
.B(n_95),
.Y(n_112)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_64),
.Y(n_88)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_88),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_60),
.A2(n_29),
.B1(n_43),
.B2(n_34),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_89),
.A2(n_103),
.B1(n_76),
.B2(n_56),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_75),
.A2(n_31),
.B1(n_15),
.B2(n_22),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_91),
.A2(n_99),
.B1(n_104),
.B2(n_107),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_48),
.B(n_15),
.Y(n_92)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_92),
.Y(n_123)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_64),
.Y(n_94)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_94),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_62),
.B(n_43),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_53),
.B(n_44),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_101),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_63),
.B(n_28),
.Y(n_101)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_102),
.B(n_93),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_60),
.A2(n_22),
.B1(n_7),
.B2(n_8),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_62),
.B(n_0),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_59),
.B(n_5),
.C(n_12),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_56),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_106),
.B(n_66),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_75),
.A2(n_5),
.B1(n_12),
.B2(n_10),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_68),
.B(n_0),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_108),
.B(n_1),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_51),
.B(n_1),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_109),
.B(n_51),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_46),
.B(n_7),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_110),
.B(n_13),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_82),
.A2(n_76),
.B1(n_73),
.B2(n_58),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_111),
.A2(n_113),
.B1(n_125),
.B2(n_131),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_117),
.B(n_98),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_120),
.A2(n_91),
.B(n_107),
.Y(n_154)
);

INVxp33_ASAP7_75t_L g121 ( 
.A(n_84),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_121),
.B(n_124),
.Y(n_150)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_122),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_81),
.B(n_61),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_82),
.A2(n_65),
.B1(n_67),
.B2(n_77),
.Y(n_125)
);

INVxp33_ASAP7_75t_L g126 ( 
.A(n_108),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_126),
.B(n_102),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_97),
.B(n_68),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_128),
.B(n_129),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_97),
.B(n_77),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_79),
.Y(n_130)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_130),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_96),
.A2(n_67),
.B1(n_77),
.B2(n_66),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_87),
.A2(n_101),
.B1(n_100),
.B2(n_80),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_132),
.A2(n_104),
.B1(n_109),
.B2(n_95),
.Y(n_144)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_79),
.Y(n_134)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_134),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_135),
.B(n_136),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_87),
.B(n_1),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_83),
.Y(n_137)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_137),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_139),
.B(n_105),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_112),
.A2(n_106),
.B(n_104),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_141),
.A2(n_120),
.B(n_114),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_123),
.B(n_98),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_142),
.B(n_158),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_144),
.B(n_152),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_112),
.B(n_78),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_145),
.B(n_131),
.C(n_133),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_146),
.B(n_160),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_114),
.A2(n_95),
.B1(n_103),
.B2(n_109),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_149),
.A2(n_151),
.B1(n_113),
.B2(n_139),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_114),
.A2(n_83),
.B1(n_94),
.B2(n_88),
.Y(n_151)
);

OR2x2_ASAP7_75t_L g152 ( 
.A(n_132),
.B(n_136),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_154),
.A2(n_157),
.B(n_1),
.Y(n_181)
);

HB1xp67_ASAP7_75t_L g156 ( 
.A(n_127),
.Y(n_156)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_156),
.Y(n_180)
);

OR2x2_ASAP7_75t_L g157 ( 
.A(n_129),
.B(n_93),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_115),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_117),
.B(n_110),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_161),
.B(n_162),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_116),
.B(n_86),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_163),
.B(n_128),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_164),
.A2(n_168),
.B(n_144),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_167),
.B(n_173),
.Y(n_184)
);

AOI221xp5_ASAP7_75t_L g169 ( 
.A1(n_141),
.A2(n_118),
.B1(n_116),
.B2(n_138),
.C(n_133),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_169),
.B(n_174),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_158),
.B(n_137),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_171),
.B(n_172),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_150),
.B(n_140),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_150),
.B(n_127),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_157),
.A2(n_134),
.B1(n_130),
.B2(n_138),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_175),
.A2(n_179),
.B1(n_143),
.B2(n_152),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_146),
.B(n_120),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_176),
.B(n_177),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_140),
.B(n_119),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_178),
.B(n_145),
.C(n_149),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_157),
.A2(n_119),
.B1(n_115),
.B2(n_10),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_181),
.A2(n_182),
.B(n_160),
.Y(n_196)
);

AOI322xp5_ASAP7_75t_L g182 ( 
.A1(n_148),
.A2(n_8),
.A3(n_10),
.B1(n_12),
.B2(n_13),
.C1(n_3),
.C2(n_4),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_171),
.Y(n_183)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_183),
.Y(n_204)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_177),
.Y(n_185)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_185),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_165),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_186),
.B(n_189),
.Y(n_199)
);

CKINVDCx14_ASAP7_75t_R g200 ( 
.A(n_188),
.Y(n_200)
);

BUFx12f_ASAP7_75t_L g189 ( 
.A(n_180),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_180),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_190),
.B(n_196),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_192),
.B(n_174),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_178),
.B(n_164),
.C(n_168),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_194),
.B(n_170),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_181),
.A2(n_151),
.B(n_154),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_195),
.A2(n_197),
.B(n_198),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_175),
.A2(n_152),
.B(n_159),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_186),
.A2(n_165),
.B1(n_172),
.B2(n_143),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_201),
.A2(n_203),
.B1(n_197),
.B2(n_187),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_202),
.B(n_205),
.C(n_207),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_188),
.A2(n_167),
.B1(n_163),
.B2(n_147),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_192),
.B(n_194),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_198),
.B(n_195),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_193),
.B(n_170),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_210),
.B(n_166),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_211),
.B(n_166),
.C(n_148),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_200),
.A2(n_183),
.B1(n_185),
.B2(n_196),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_213),
.B(n_217),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_214),
.B(n_219),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_207),
.A2(n_184),
.B1(n_147),
.B2(n_191),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_215),
.A2(n_218),
.B1(n_220),
.B2(n_209),
.Y(n_221)
);

AOI31xp67_ASAP7_75t_L g216 ( 
.A1(n_208),
.A2(n_184),
.A3(n_193),
.B(n_176),
.Y(n_216)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_216),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_209),
.B(n_190),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_206),
.A2(n_179),
.B1(n_155),
.B2(n_159),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_221),
.B(n_222),
.Y(n_230)
);

BUFx24_ASAP7_75t_SL g222 ( 
.A(n_213),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_212),
.B(n_202),
.C(n_205),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_224),
.A2(n_225),
.B(n_211),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_220),
.A2(n_208),
.B1(n_203),
.B2(n_204),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_226),
.A2(n_212),
.B1(n_217),
.B2(n_216),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_228),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_229),
.B(n_224),
.C(n_223),
.Y(n_235)
);

O2A1O1Ixp5_ASAP7_75t_L g231 ( 
.A1(n_227),
.A2(n_215),
.B(n_204),
.C(n_199),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_231),
.A2(n_189),
.B(n_8),
.Y(n_236)
);

OAI221xp5_ASAP7_75t_L g232 ( 
.A1(n_227),
.A2(n_153),
.B1(n_155),
.B2(n_162),
.C(n_189),
.Y(n_232)
);

AOI21x1_ASAP7_75t_L g233 ( 
.A1(n_232),
.A2(n_189),
.B(n_153),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_233),
.B(n_2),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_235),
.B(n_236),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_234),
.A2(n_230),
.B(n_13),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_237),
.B(n_238),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_239),
.A2(n_2),
.B(n_4),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_241),
.B(n_240),
.Y(n_242)
);


endmodule