module fake_netlist_6_2968_n_890 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_890);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_890;

wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_881;
wire n_875;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_760;
wire n_741;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_828;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_384;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_342;
wire n_820;
wire n_783;
wire n_725;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_628;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_845;
wire n_255;
wire n_807;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_865;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_669;
wire n_200;
wire n_447;
wire n_872;
wire n_198;
wire n_222;
wire n_248;
wire n_300;
wire n_517;
wire n_718;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_544;
wire n_468;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_866;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_658;
wire n_616;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_822;
wire n_693;
wire n_631;
wire n_516;
wire n_720;
wire n_758;
wire n_525;
wire n_842;
wire n_611;
wire n_491;
wire n_878;
wire n_772;
wire n_656;
wire n_843;
wire n_797;
wire n_666;
wire n_371;
wire n_795;
wire n_770;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_197;
wire n_844;
wire n_343;
wire n_448;
wire n_886;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_888;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_887;
wire n_752;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_224;
wire n_839;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_779;
wire n_800;
wire n_460;
wire n_854;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_777;
wire n_407;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_552;
wire n_619;
wire n_885;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_792;
wire n_880;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_821;
wire n_325;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_806;
wire n_864;
wire n_879;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_707;
wire n_322;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_811;
wire n_882;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_775;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_835;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_816;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_205;
wire n_604;
wire n_848;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_862;
wire n_869;
wire n_351;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_637;
wire n_385;
wire n_295;
wire n_701;
wire n_817;
wire n_629;
wire n_388;
wire n_190;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_846;
wire n_501;
wire n_841;
wire n_531;
wire n_827;
wire n_508;
wire n_361;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_332;
wire n_336;
wire n_410;
wire n_398;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_678;
wire n_192;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_102),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_69),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_37),
.Y(n_191)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_65),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_149),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_178),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_166),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_17),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_108),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_181),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_7),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_16),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_184),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_27),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_97),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_107),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_179),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_82),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_28),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_73),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_110),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_154),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_98),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_169),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_95),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_123),
.Y(n_214)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_144),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_112),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_138),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_175),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_14),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_186),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_106),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_104),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_159),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_188),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_182),
.Y(n_225)
);

INVxp33_ASAP7_75t_L g226 ( 
.A(n_50),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_177),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_183),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_26),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_172),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_4),
.Y(n_231)
);

BUFx5_ASAP7_75t_L g232 ( 
.A(n_185),
.Y(n_232)
);

INVx2_ASAP7_75t_SL g233 ( 
.A(n_128),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_187),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_40),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_167),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_130),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_10),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_23),
.Y(n_239)
);

BUFx10_ASAP7_75t_L g240 ( 
.A(n_14),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_180),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_96),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_109),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_38),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_52),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_119),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_173),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_75),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_62),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_53),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_30),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_20),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_17),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_64),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_68),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_66),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_76),
.Y(n_257)
);

BUFx10_ASAP7_75t_L g258 ( 
.A(n_48),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_135),
.Y(n_259)
);

BUFx2_ASAP7_75t_L g260 ( 
.A(n_145),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_7),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_174),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_78),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_49),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_80),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_13),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_63),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_55),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_136),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_31),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_153),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_161),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_74),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_189),
.Y(n_274)
);

BUFx2_ASAP7_75t_L g275 ( 
.A(n_199),
.Y(n_275)
);

AND2x4_ASAP7_75t_L g276 ( 
.A(n_192),
.B(n_0),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_209),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_196),
.Y(n_278)
);

INVx2_ASAP7_75t_SL g279 ( 
.A(n_240),
.Y(n_279)
);

INVx4_ASAP7_75t_L g280 ( 
.A(n_209),
.Y(n_280)
);

INVxp33_ASAP7_75t_SL g281 ( 
.A(n_200),
.Y(n_281)
);

AND2x4_ASAP7_75t_L g282 ( 
.A(n_192),
.B(n_215),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_232),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_209),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_240),
.B(n_0),
.Y(n_285)
);

AND2x4_ASAP7_75t_L g286 ( 
.A(n_215),
.B(n_1),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_209),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_226),
.B(n_1),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_208),
.B(n_260),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_227),
.B(n_2),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_191),
.Y(n_291)
);

AND2x4_ASAP7_75t_L g292 ( 
.A(n_233),
.B(n_2),
.Y(n_292)
);

BUFx12f_ASAP7_75t_L g293 ( 
.A(n_258),
.Y(n_293)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_258),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_244),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_229),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_202),
.B(n_3),
.Y(n_297)
);

BUFx12f_ASAP7_75t_L g298 ( 
.A(n_207),
.Y(n_298)
);

INVx5_ASAP7_75t_L g299 ( 
.A(n_244),
.Y(n_299)
);

AND2x4_ASAP7_75t_L g300 ( 
.A(n_194),
.B(n_3),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_244),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_231),
.B(n_4),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_232),
.Y(n_303)
);

INVx4_ASAP7_75t_L g304 ( 
.A(n_244),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_271),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_252),
.B(n_5),
.Y(n_306)
);

INVx4_ASAP7_75t_L g307 ( 
.A(n_271),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_219),
.B(n_5),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_248),
.B(n_6),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_239),
.B(n_6),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_271),
.Y(n_311)
);

INVx5_ASAP7_75t_L g312 ( 
.A(n_271),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_197),
.Y(n_313)
);

AND2x4_ASAP7_75t_L g314 ( 
.A(n_198),
.B(n_8),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_201),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_204),
.B(n_8),
.Y(n_316)
);

BUFx2_ASAP7_75t_L g317 ( 
.A(n_238),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_253),
.B(n_9),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_214),
.Y(n_319)
);

BUFx8_ASAP7_75t_SL g320 ( 
.A(n_190),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_216),
.B(n_9),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_261),
.B(n_10),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_217),
.Y(n_323)
);

NOR2x1_ASAP7_75t_L g324 ( 
.A(n_218),
.B(n_29),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_222),
.B(n_11),
.Y(n_325)
);

BUFx12f_ASAP7_75t_L g326 ( 
.A(n_266),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_232),
.Y(n_327)
);

AND2x4_ASAP7_75t_L g328 ( 
.A(n_230),
.B(n_11),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_232),
.B(n_12),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_289),
.A2(n_211),
.B1(n_236),
.B2(n_251),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_317),
.B(n_193),
.Y(n_331)
);

OR2x6_ASAP7_75t_L g332 ( 
.A(n_298),
.B(n_245),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_287),
.Y(n_333)
);

OAI22xp33_ASAP7_75t_L g334 ( 
.A1(n_285),
.A2(n_318),
.B1(n_310),
.B2(n_329),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_289),
.A2(n_250),
.B1(n_272),
.B2(n_255),
.Y(n_335)
);

INVx3_ASAP7_75t_L g336 ( 
.A(n_277),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_294),
.B(n_195),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_294),
.B(n_203),
.Y(n_338)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_277),
.Y(n_339)
);

OR2x2_ASAP7_75t_L g340 ( 
.A(n_275),
.B(n_12),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_315),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_278),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_287),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_287),
.Y(n_344)
);

AND2x2_ASAP7_75t_L g345 ( 
.A(n_274),
.B(n_205),
.Y(n_345)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_282),
.B(n_206),
.Y(n_346)
);

OAI22xp33_ASAP7_75t_SL g347 ( 
.A1(n_329),
.A2(n_259),
.B1(n_264),
.B2(n_269),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_287),
.Y(n_348)
);

AO22x2_ASAP7_75t_L g349 ( 
.A1(n_276),
.A2(n_232),
.B1(n_15),
.B2(n_16),
.Y(n_349)
);

OAI22xp33_ASAP7_75t_L g350 ( 
.A1(n_285),
.A2(n_273),
.B1(n_270),
.B2(n_268),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_291),
.B(n_210),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_313),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_313),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_288),
.A2(n_267),
.B1(n_265),
.B2(n_263),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_279),
.B(n_212),
.Y(n_355)
);

OAI22xp33_ASAP7_75t_SL g356 ( 
.A1(n_310),
.A2(n_262),
.B1(n_257),
.B2(n_256),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_288),
.B(n_213),
.Y(n_357)
);

OAI22xp33_ASAP7_75t_SL g358 ( 
.A1(n_318),
.A2(n_254),
.B1(n_249),
.B2(n_247),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_297),
.B(n_220),
.Y(n_359)
);

INVx3_ASAP7_75t_L g360 ( 
.A(n_277),
.Y(n_360)
);

BUFx6f_ASAP7_75t_SL g361 ( 
.A(n_282),
.Y(n_361)
);

AO22x2_ASAP7_75t_L g362 ( 
.A1(n_276),
.A2(n_232),
.B1(n_15),
.B2(n_18),
.Y(n_362)
);

OAI22xp33_ASAP7_75t_SL g363 ( 
.A1(n_286),
.A2(n_321),
.B1(n_325),
.B2(n_281),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_290),
.A2(n_246),
.B1(n_243),
.B2(n_242),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_313),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_319),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_311),
.Y(n_367)
);

OAI22xp33_ASAP7_75t_SL g368 ( 
.A1(n_286),
.A2(n_241),
.B1(n_237),
.B2(n_235),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_308),
.B(n_221),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_284),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_311),
.Y(n_371)
);

AOI22x1_ASAP7_75t_SL g372 ( 
.A1(n_320),
.A2(n_234),
.B1(n_228),
.B2(n_225),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_290),
.A2(n_224),
.B1(n_223),
.B2(n_19),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g374 ( 
.A(n_322),
.B(n_32),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_309),
.A2(n_13),
.B1(n_18),
.B2(n_19),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_302),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_309),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_377)
);

AO22x2_ASAP7_75t_L g378 ( 
.A1(n_292),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_326),
.A2(n_24),
.B1(n_25),
.B2(n_27),
.Y(n_379)
);

OAI22xp33_ASAP7_75t_L g380 ( 
.A1(n_302),
.A2(n_306),
.B1(n_296),
.B2(n_325),
.Y(n_380)
);

OAI22xp33_ASAP7_75t_SL g381 ( 
.A1(n_321),
.A2(n_28),
.B1(n_33),
.B2(n_34),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_292),
.B(n_35),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_319),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_296),
.B(n_36),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_299),
.B(n_39),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_342),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_SL g387 ( 
.A(n_334),
.B(n_320),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_330),
.Y(n_388)
);

NOR2x1_ASAP7_75t_L g389 ( 
.A(n_350),
.B(n_280),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_341),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_336),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_336),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_339),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_339),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_360),
.Y(n_395)
);

AND2x4_ASAP7_75t_L g396 ( 
.A(n_384),
.B(n_300),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_360),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_352),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_353),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_365),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_366),
.Y(n_401)
);

INVxp67_ASAP7_75t_SL g402 ( 
.A(n_370),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_350),
.B(n_319),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_383),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_372),
.Y(n_405)
);

INVxp33_ASAP7_75t_L g406 ( 
.A(n_357),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_346),
.B(n_300),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_333),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_333),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_343),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_L g411 ( 
.A1(n_382),
.A2(n_328),
.B(n_314),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_346),
.B(n_314),
.Y(n_412)
);

AND2x4_ASAP7_75t_L g413 ( 
.A(n_382),
.B(n_328),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_343),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_344),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_344),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_348),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_348),
.Y(n_418)
);

NAND2x1p5_ASAP7_75t_L g419 ( 
.A(n_374),
.B(n_324),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_335),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_SL g421 ( 
.A(n_334),
.B(n_293),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_357),
.B(n_323),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_367),
.Y(n_423)
);

INVx1_ASAP7_75t_SL g424 ( 
.A(n_355),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_367),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_371),
.Y(n_426)
);

BUFx3_ASAP7_75t_L g427 ( 
.A(n_370),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_371),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_L g429 ( 
.A1(n_337),
.A2(n_327),
.B(n_283),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_370),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_370),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_338),
.B(n_299),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_361),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_361),
.Y(n_434)
);

INVxp67_ASAP7_75t_SL g435 ( 
.A(n_385),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_349),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_331),
.B(n_323),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_380),
.B(n_323),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_340),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_332),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_SL g441 ( 
.A(n_380),
.B(n_316),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_359),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_369),
.Y(n_443)
);

AND2x2_ASAP7_75t_L g444 ( 
.A(n_345),
.B(n_316),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_349),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_349),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_362),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_362),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_362),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_381),
.Y(n_450)
);

NOR2xp67_ASAP7_75t_L g451 ( 
.A(n_364),
.B(n_299),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_363),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_378),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_351),
.B(n_306),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_454),
.B(n_378),
.Y(n_455)
);

HB1xp67_ASAP7_75t_L g456 ( 
.A(n_452),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_435),
.B(n_354),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_454),
.B(n_407),
.Y(n_458)
);

BUFx3_ASAP7_75t_L g459 ( 
.A(n_386),
.Y(n_459)
);

INVxp33_ASAP7_75t_L g460 ( 
.A(n_439),
.Y(n_460)
);

OR2x2_ASAP7_75t_SL g461 ( 
.A(n_453),
.B(n_378),
.Y(n_461)
);

INVx1_ASAP7_75t_SL g462 ( 
.A(n_424),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_411),
.B(n_422),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_417),
.Y(n_464)
);

AND2x4_ASAP7_75t_L g465 ( 
.A(n_437),
.B(n_390),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g466 ( 
.A(n_407),
.B(n_412),
.Y(n_466)
);

OAI21xp5_ASAP7_75t_L g467 ( 
.A1(n_429),
.A2(n_347),
.B(n_368),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_417),
.Y(n_468)
);

HB1xp67_ASAP7_75t_L g469 ( 
.A(n_437),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_426),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_426),
.Y(n_471)
);

INVx3_ASAP7_75t_L g472 ( 
.A(n_408),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_422),
.B(n_356),
.Y(n_473)
);

OR2x2_ASAP7_75t_SL g474 ( 
.A(n_436),
.B(n_358),
.Y(n_474)
);

INVxp67_ASAP7_75t_L g475 ( 
.A(n_421),
.Y(n_475)
);

BUFx3_ASAP7_75t_L g476 ( 
.A(n_433),
.Y(n_476)
);

INVx3_ASAP7_75t_L g477 ( 
.A(n_409),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_406),
.B(n_373),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_410),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g480 ( 
.A(n_450),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_412),
.B(n_303),
.Y(n_481)
);

AND2x4_ASAP7_75t_L g482 ( 
.A(n_436),
.B(n_448),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_414),
.Y(n_483)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_415),
.Y(n_484)
);

INVx3_ASAP7_75t_SL g485 ( 
.A(n_405),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g486 ( 
.A(n_427),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_416),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_396),
.B(n_280),
.Y(n_488)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_444),
.B(n_375),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_418),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_444),
.B(n_332),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_413),
.B(n_332),
.Y(n_492)
);

HB1xp67_ASAP7_75t_L g493 ( 
.A(n_442),
.Y(n_493)
);

INVx3_ASAP7_75t_L g494 ( 
.A(n_423),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_396),
.B(n_304),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_425),
.Y(n_496)
);

AND2x4_ASAP7_75t_SL g497 ( 
.A(n_448),
.B(n_379),
.Y(n_497)
);

INVx2_ASAP7_75t_SL g498 ( 
.A(n_396),
.Y(n_498)
);

AND2x6_ASAP7_75t_L g499 ( 
.A(n_445),
.B(n_311),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_413),
.B(n_376),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_428),
.Y(n_501)
);

INVx4_ASAP7_75t_L g502 ( 
.A(n_427),
.Y(n_502)
);

HB1xp67_ASAP7_75t_L g503 ( 
.A(n_443),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_413),
.B(n_304),
.Y(n_504)
);

AND2x2_ASAP7_75t_SL g505 ( 
.A(n_441),
.B(n_307),
.Y(n_505)
);

BUFx3_ASAP7_75t_L g506 ( 
.A(n_434),
.Y(n_506)
);

INVxp67_ASAP7_75t_SL g507 ( 
.A(n_402),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_406),
.B(n_307),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_398),
.Y(n_509)
);

BUFx6f_ASAP7_75t_L g510 ( 
.A(n_430),
.Y(n_510)
);

AND2x6_ASAP7_75t_L g511 ( 
.A(n_446),
.B(n_311),
.Y(n_511)
);

BUFx3_ASAP7_75t_L g512 ( 
.A(n_399),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_403),
.B(n_299),
.Y(n_513)
);

AND2x4_ASAP7_75t_SL g514 ( 
.A(n_447),
.B(n_284),
.Y(n_514)
);

OAI21xp5_ASAP7_75t_L g515 ( 
.A1(n_403),
.A2(n_376),
.B(n_312),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_400),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_401),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_404),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_391),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_392),
.Y(n_520)
);

HB1xp67_ASAP7_75t_L g521 ( 
.A(n_438),
.Y(n_521)
);

INVxp67_ASAP7_75t_L g522 ( 
.A(n_387),
.Y(n_522)
);

HB1xp67_ASAP7_75t_L g523 ( 
.A(n_438),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_389),
.B(n_312),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_482),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_486),
.Y(n_526)
);

AND2x2_ASAP7_75t_SL g527 ( 
.A(n_463),
.B(n_449),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_482),
.Y(n_528)
);

BUFx10_ASAP7_75t_L g529 ( 
.A(n_497),
.Y(n_529)
);

NOR2x1_ASAP7_75t_SL g530 ( 
.A(n_502),
.B(n_432),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_482),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_483),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_458),
.B(n_419),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_458),
.B(n_419),
.Y(n_534)
);

AND2x4_ASAP7_75t_L g535 ( 
.A(n_498),
.B(n_451),
.Y(n_535)
);

OR2x2_ASAP7_75t_L g536 ( 
.A(n_462),
.B(n_393),
.Y(n_536)
);

BUFx3_ASAP7_75t_L g537 ( 
.A(n_476),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_521),
.B(n_431),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_483),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_469),
.B(n_388),
.Y(n_540)
);

AND2x4_ASAP7_75t_L g541 ( 
.A(n_498),
.B(n_394),
.Y(n_541)
);

NAND2xp33_ASAP7_75t_L g542 ( 
.A(n_457),
.B(n_523),
.Y(n_542)
);

AND2x4_ASAP7_75t_L g543 ( 
.A(n_465),
.B(n_395),
.Y(n_543)
);

OR2x6_ASAP7_75t_L g544 ( 
.A(n_522),
.B(n_377),
.Y(n_544)
);

INVx2_ASAP7_75t_SL g545 ( 
.A(n_493),
.Y(n_545)
);

INVxp33_ASAP7_75t_L g546 ( 
.A(n_503),
.Y(n_546)
);

AND2x4_ASAP7_75t_L g547 ( 
.A(n_465),
.B(n_397),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_481),
.B(n_388),
.Y(n_548)
);

BUFx2_ASAP7_75t_L g549 ( 
.A(n_475),
.Y(n_549)
);

OR2x6_ASAP7_75t_L g550 ( 
.A(n_492),
.B(n_440),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_485),
.Y(n_551)
);

AND2x2_ASAP7_75t_L g552 ( 
.A(n_460),
.B(n_466),
.Y(n_552)
);

AND2x6_ASAP7_75t_L g553 ( 
.A(n_455),
.B(n_284),
.Y(n_553)
);

INVx4_ASAP7_75t_L g554 ( 
.A(n_486),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_466),
.B(n_420),
.Y(n_555)
);

INVx1_ASAP7_75t_SL g556 ( 
.A(n_505),
.Y(n_556)
);

OR2x2_ASAP7_75t_L g557 ( 
.A(n_478),
.B(n_405),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_486),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_486),
.Y(n_559)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_489),
.B(n_420),
.Y(n_560)
);

AND2x2_ASAP7_75t_L g561 ( 
.A(n_489),
.B(n_440),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_481),
.B(n_295),
.Y(n_562)
);

BUFx3_ASAP7_75t_L g563 ( 
.A(n_476),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g564 ( 
.A(n_486),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_505),
.B(n_295),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_464),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_508),
.B(n_456),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_455),
.B(n_295),
.Y(n_568)
);

AND2x4_ASAP7_75t_L g569 ( 
.A(n_465),
.B(n_41),
.Y(n_569)
);

BUFx2_ASAP7_75t_L g570 ( 
.A(n_474),
.Y(n_570)
);

AND2x4_ASAP7_75t_L g571 ( 
.A(n_459),
.B(n_42),
.Y(n_571)
);

OR2x2_ASAP7_75t_L g572 ( 
.A(n_474),
.B(n_43),
.Y(n_572)
);

AND2x4_ASAP7_75t_L g573 ( 
.A(n_459),
.B(n_44),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_487),
.Y(n_574)
);

NAND2x1p5_ASAP7_75t_L g575 ( 
.A(n_502),
.B(n_301),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_487),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_496),
.Y(n_577)
);

INVx3_ASAP7_75t_L g578 ( 
.A(n_502),
.Y(n_578)
);

INVx3_ASAP7_75t_L g579 ( 
.A(n_510),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_496),
.Y(n_580)
);

INVxp67_ASAP7_75t_SL g581 ( 
.A(n_480),
.Y(n_581)
);

BUFx3_ASAP7_75t_L g582 ( 
.A(n_506),
.Y(n_582)
);

OR2x6_ASAP7_75t_L g583 ( 
.A(n_492),
.B(n_301),
.Y(n_583)
);

BUFx12f_ASAP7_75t_L g584 ( 
.A(n_551),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_566),
.Y(n_585)
);

CKINVDCx11_ASAP7_75t_R g586 ( 
.A(n_550),
.Y(n_586)
);

AND2x2_ASAP7_75t_L g587 ( 
.A(n_527),
.B(n_500),
.Y(n_587)
);

INVx1_ASAP7_75t_SL g588 ( 
.A(n_549),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_525),
.Y(n_589)
);

BUFx2_ASAP7_75t_L g590 ( 
.A(n_570),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_567),
.B(n_500),
.Y(n_591)
);

CKINVDCx16_ASAP7_75t_R g592 ( 
.A(n_560),
.Y(n_592)
);

INVx3_ASAP7_75t_L g593 ( 
.A(n_578),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_528),
.Y(n_594)
);

BUFx6f_ASAP7_75t_L g595 ( 
.A(n_526),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_531),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_532),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_539),
.Y(n_598)
);

INVx4_ASAP7_75t_L g599 ( 
.A(n_526),
.Y(n_599)
);

BUFx3_ASAP7_75t_L g600 ( 
.A(n_529),
.Y(n_600)
);

INVx8_ASAP7_75t_L g601 ( 
.A(n_569),
.Y(n_601)
);

AOI22xp33_ASAP7_75t_L g602 ( 
.A1(n_527),
.A2(n_556),
.B1(n_542),
.B2(n_572),
.Y(n_602)
);

BUFx6f_ASAP7_75t_L g603 ( 
.A(n_526),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_574),
.Y(n_604)
);

INVx2_ASAP7_75t_SL g605 ( 
.A(n_558),
.Y(n_605)
);

INVxp67_ASAP7_75t_SL g606 ( 
.A(n_578),
.Y(n_606)
);

BUFx3_ASAP7_75t_L g607 ( 
.A(n_529),
.Y(n_607)
);

INVx5_ASAP7_75t_L g608 ( 
.A(n_558),
.Y(n_608)
);

BUFx2_ASAP7_75t_SL g609 ( 
.A(n_558),
.Y(n_609)
);

INVx3_ASAP7_75t_L g610 ( 
.A(n_559),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_576),
.Y(n_611)
);

INVx3_ASAP7_75t_L g612 ( 
.A(n_559),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_577),
.Y(n_613)
);

INVx2_ASAP7_75t_SL g614 ( 
.A(n_559),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_556),
.B(n_491),
.Y(n_615)
);

INVx3_ASAP7_75t_L g616 ( 
.A(n_564),
.Y(n_616)
);

BUFx12f_ASAP7_75t_L g617 ( 
.A(n_550),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_567),
.B(n_473),
.Y(n_618)
);

INVx2_ASAP7_75t_SL g619 ( 
.A(n_564),
.Y(n_619)
);

CKINVDCx20_ASAP7_75t_R g620 ( 
.A(n_548),
.Y(n_620)
);

BUFx6f_ASAP7_75t_SL g621 ( 
.A(n_550),
.Y(n_621)
);

BUFx3_ASAP7_75t_L g622 ( 
.A(n_564),
.Y(n_622)
);

BUFx2_ASAP7_75t_SL g623 ( 
.A(n_554),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_580),
.Y(n_624)
);

BUFx4f_ASAP7_75t_L g625 ( 
.A(n_569),
.Y(n_625)
);

AOI22xp33_ASAP7_75t_L g626 ( 
.A1(n_542),
.A2(n_467),
.B1(n_515),
.B2(n_497),
.Y(n_626)
);

INVx4_ASAP7_75t_L g627 ( 
.A(n_554),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_579),
.Y(n_628)
);

INVx1_ASAP7_75t_SL g629 ( 
.A(n_540),
.Y(n_629)
);

BUFx12f_ASAP7_75t_L g630 ( 
.A(n_545),
.Y(n_630)
);

BUFx2_ASAP7_75t_R g631 ( 
.A(n_609),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_598),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_598),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_611),
.Y(n_634)
);

INVx3_ASAP7_75t_L g635 ( 
.A(n_627),
.Y(n_635)
);

OAI22xp5_ASAP7_75t_L g636 ( 
.A1(n_626),
.A2(n_548),
.B1(n_571),
.B2(n_573),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_611),
.Y(n_637)
);

AOI22xp33_ASAP7_75t_L g638 ( 
.A1(n_587),
.A2(n_555),
.B1(n_544),
.B2(n_561),
.Y(n_638)
);

AOI22xp33_ASAP7_75t_L g639 ( 
.A1(n_587),
.A2(n_544),
.B1(n_557),
.B2(n_552),
.Y(n_639)
);

AOI22xp33_ASAP7_75t_L g640 ( 
.A1(n_620),
.A2(n_544),
.B1(n_491),
.B2(n_534),
.Y(n_640)
);

INVx5_ASAP7_75t_L g641 ( 
.A(n_595),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_613),
.Y(n_642)
);

OAI22xp5_ASAP7_75t_L g643 ( 
.A1(n_591),
.A2(n_571),
.B1(n_573),
.B2(n_581),
.Y(n_643)
);

INVx6_ASAP7_75t_L g644 ( 
.A(n_630),
.Y(n_644)
);

BUFx2_ASAP7_75t_SL g645 ( 
.A(n_588),
.Y(n_645)
);

CKINVDCx11_ASAP7_75t_R g646 ( 
.A(n_584),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_597),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_613),
.Y(n_648)
);

CKINVDCx11_ASAP7_75t_R g649 ( 
.A(n_584),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_597),
.Y(n_650)
);

CKINVDCx20_ASAP7_75t_R g651 ( 
.A(n_592),
.Y(n_651)
);

AOI22xp33_ASAP7_75t_SL g652 ( 
.A1(n_592),
.A2(n_581),
.B1(n_534),
.B2(n_533),
.Y(n_652)
);

AOI22xp33_ASAP7_75t_SL g653 ( 
.A1(n_621),
.A2(n_533),
.B1(n_582),
.B2(n_563),
.Y(n_653)
);

NAND2x1p5_ASAP7_75t_L g654 ( 
.A(n_608),
.B(n_579),
.Y(n_654)
);

CKINVDCx11_ASAP7_75t_R g655 ( 
.A(n_630),
.Y(n_655)
);

AOI22xp5_ASAP7_75t_L g656 ( 
.A1(n_629),
.A2(n_535),
.B1(n_546),
.B2(n_543),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_597),
.Y(n_657)
);

INVx6_ASAP7_75t_L g658 ( 
.A(n_617),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_604),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_604),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_604),
.Y(n_661)
);

NOR2x1_ASAP7_75t_SL g662 ( 
.A(n_623),
.B(n_608),
.Y(n_662)
);

BUFx6f_ASAP7_75t_L g663 ( 
.A(n_595),
.Y(n_663)
);

BUFx2_ASAP7_75t_L g664 ( 
.A(n_590),
.Y(n_664)
);

AOI22xp33_ASAP7_75t_L g665 ( 
.A1(n_615),
.A2(n_553),
.B1(n_546),
.B2(n_543),
.Y(n_665)
);

BUFx6f_ASAP7_75t_L g666 ( 
.A(n_595),
.Y(n_666)
);

CKINVDCx20_ASAP7_75t_R g667 ( 
.A(n_586),
.Y(n_667)
);

OAI22xp33_ASAP7_75t_L g668 ( 
.A1(n_618),
.A2(n_536),
.B1(n_537),
.B2(n_485),
.Y(n_668)
);

AOI22xp33_ASAP7_75t_L g669 ( 
.A1(n_625),
.A2(n_553),
.B1(n_547),
.B2(n_541),
.Y(n_669)
);

INVx6_ASAP7_75t_L g670 ( 
.A(n_617),
.Y(n_670)
);

BUFx2_ASAP7_75t_L g671 ( 
.A(n_590),
.Y(n_671)
);

INVxp67_ASAP7_75t_SL g672 ( 
.A(n_606),
.Y(n_672)
);

AOI22xp33_ASAP7_75t_L g673 ( 
.A1(n_625),
.A2(n_553),
.B1(n_547),
.B2(n_541),
.Y(n_673)
);

OAI22xp5_ASAP7_75t_L g674 ( 
.A1(n_643),
.A2(n_625),
.B1(n_602),
.B2(n_601),
.Y(n_674)
);

OAI21xp33_ASAP7_75t_L g675 ( 
.A1(n_639),
.A2(n_638),
.B(n_640),
.Y(n_675)
);

OAI21xp5_ASAP7_75t_SL g676 ( 
.A1(n_636),
.A2(n_535),
.B(n_517),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_664),
.B(n_568),
.Y(n_677)
);

INVx4_ASAP7_75t_L g678 ( 
.A(n_641),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_647),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_632),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_633),
.Y(n_681)
);

INVx4_ASAP7_75t_L g682 ( 
.A(n_641),
.Y(n_682)
);

INVx4_ASAP7_75t_R g683 ( 
.A(n_631),
.Y(n_683)
);

HB1xp67_ASAP7_75t_L g684 ( 
.A(n_650),
.Y(n_684)
);

AOI22xp33_ASAP7_75t_L g685 ( 
.A1(n_636),
.A2(n_621),
.B1(n_601),
.B2(n_512),
.Y(n_685)
);

CKINVDCx8_ASAP7_75t_R g686 ( 
.A(n_645),
.Y(n_686)
);

OAI221xp5_ASAP7_75t_L g687 ( 
.A1(n_656),
.A2(n_506),
.B1(n_512),
.B2(n_517),
.C(n_518),
.Y(n_687)
);

AOI22xp33_ASAP7_75t_L g688 ( 
.A1(n_652),
.A2(n_621),
.B1(n_601),
.B2(n_553),
.Y(n_688)
);

OAI222xp33_ASAP7_75t_L g689 ( 
.A1(n_643),
.A2(n_565),
.B1(n_624),
.B2(n_538),
.C1(n_594),
.C2(n_596),
.Y(n_689)
);

AOI22xp33_ASAP7_75t_L g690 ( 
.A1(n_668),
.A2(n_601),
.B1(n_596),
.B2(n_509),
.Y(n_690)
);

AOI22xp33_ASAP7_75t_L g691 ( 
.A1(n_651),
.A2(n_601),
.B1(n_596),
.B2(n_509),
.Y(n_691)
);

AOI22xp33_ASAP7_75t_SL g692 ( 
.A1(n_658),
.A2(n_565),
.B1(n_624),
.B2(n_600),
.Y(n_692)
);

AOI22xp33_ASAP7_75t_L g693 ( 
.A1(n_653),
.A2(n_589),
.B1(n_583),
.B2(n_518),
.Y(n_693)
);

AOI22xp33_ASAP7_75t_SL g694 ( 
.A1(n_658),
.A2(n_607),
.B1(n_600),
.B2(n_594),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_634),
.Y(n_695)
);

OAI22xp5_ASAP7_75t_L g696 ( 
.A1(n_665),
.A2(n_607),
.B1(n_600),
.B2(n_538),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_637),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_642),
.Y(n_698)
);

INVx3_ASAP7_75t_L g699 ( 
.A(n_663),
.Y(n_699)
);

OAI22xp5_ASAP7_75t_L g700 ( 
.A1(n_669),
.A2(n_607),
.B1(n_583),
.B2(n_589),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_671),
.B(n_583),
.Y(n_701)
);

AOI22xp33_ASAP7_75t_SL g702 ( 
.A1(n_670),
.A2(n_623),
.B1(n_593),
.B2(n_585),
.Y(n_702)
);

AOI22xp33_ASAP7_75t_L g703 ( 
.A1(n_670),
.A2(n_516),
.B1(n_520),
.B2(n_519),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_648),
.Y(n_704)
);

AOI22xp33_ASAP7_75t_L g705 ( 
.A1(n_673),
.A2(n_516),
.B1(n_520),
.B2(n_519),
.Y(n_705)
);

AOI22xp33_ASAP7_75t_L g706 ( 
.A1(n_667),
.A2(n_504),
.B1(n_488),
.B2(n_495),
.Y(n_706)
);

OAI22xp33_ASAP7_75t_L g707 ( 
.A1(n_659),
.A2(n_585),
.B1(n_562),
.B2(n_627),
.Y(n_707)
);

OAI22xp5_ASAP7_75t_L g708 ( 
.A1(n_672),
.A2(n_461),
.B1(n_593),
.B2(n_627),
.Y(n_708)
);

OAI22xp5_ASAP7_75t_SL g709 ( 
.A1(n_644),
.A2(n_461),
.B1(n_599),
.B2(n_622),
.Y(n_709)
);

AOI22xp33_ASAP7_75t_L g710 ( 
.A1(n_644),
.A2(n_501),
.B1(n_562),
.B2(n_479),
.Y(n_710)
);

INVx2_ASAP7_75t_SL g711 ( 
.A(n_663),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_660),
.Y(n_712)
);

AOI22xp33_ASAP7_75t_L g713 ( 
.A1(n_661),
.A2(n_501),
.B1(n_479),
.B2(n_490),
.Y(n_713)
);

BUFx12f_ASAP7_75t_L g714 ( 
.A(n_646),
.Y(n_714)
);

INVx1_ASAP7_75t_SL g715 ( 
.A(n_631),
.Y(n_715)
);

AOI22xp33_ASAP7_75t_L g716 ( 
.A1(n_657),
.A2(n_490),
.B1(n_524),
.B2(n_511),
.Y(n_716)
);

BUFx2_ASAP7_75t_L g717 ( 
.A(n_663),
.Y(n_717)
);

INVx8_ASAP7_75t_L g718 ( 
.A(n_641),
.Y(n_718)
);

AOI22xp33_ASAP7_75t_SL g719 ( 
.A1(n_662),
.A2(n_641),
.B1(n_635),
.B2(n_593),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_655),
.B(n_628),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_649),
.Y(n_721)
);

AOI22xp33_ASAP7_75t_L g722 ( 
.A1(n_635),
.A2(n_511),
.B1(n_499),
.B2(n_513),
.Y(n_722)
);

AOI22xp33_ASAP7_75t_L g723 ( 
.A1(n_666),
.A2(n_511),
.B1(n_499),
.B2(n_628),
.Y(n_723)
);

OAI22xp5_ASAP7_75t_L g724 ( 
.A1(n_693),
.A2(n_593),
.B1(n_627),
.B2(n_654),
.Y(n_724)
);

AOI22xp5_ASAP7_75t_L g725 ( 
.A1(n_675),
.A2(n_514),
.B1(n_599),
.B2(n_614),
.Y(n_725)
);

NAND3xp33_ASAP7_75t_L g726 ( 
.A(n_706),
.B(n_628),
.C(n_666),
.Y(n_726)
);

AOI22xp33_ASAP7_75t_SL g727 ( 
.A1(n_674),
.A2(n_530),
.B1(n_609),
.B2(n_666),
.Y(n_727)
);

AOI22xp33_ASAP7_75t_L g728 ( 
.A1(n_685),
.A2(n_687),
.B1(n_690),
.B2(n_691),
.Y(n_728)
);

AOI22xp33_ASAP7_75t_SL g729 ( 
.A1(n_709),
.A2(n_628),
.B1(n_608),
.B2(n_622),
.Y(n_729)
);

OAI222xp33_ASAP7_75t_L g730 ( 
.A1(n_688),
.A2(n_692),
.B1(n_708),
.B2(n_694),
.C1(n_686),
.C2(n_700),
.Y(n_730)
);

AOI22xp33_ASAP7_75t_SL g731 ( 
.A1(n_696),
.A2(n_628),
.B1(n_608),
.B2(n_622),
.Y(n_731)
);

OAI22xp5_ASAP7_75t_L g732 ( 
.A1(n_703),
.A2(n_654),
.B1(n_575),
.B2(n_605),
.Y(n_732)
);

OAI22xp5_ASAP7_75t_L g733 ( 
.A1(n_694),
.A2(n_575),
.B1(n_614),
.B2(n_605),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_677),
.B(n_610),
.Y(n_734)
);

OAI22xp5_ASAP7_75t_L g735 ( 
.A1(n_692),
.A2(n_619),
.B1(n_616),
.B2(n_612),
.Y(n_735)
);

AOI22xp33_ASAP7_75t_L g736 ( 
.A1(n_705),
.A2(n_510),
.B1(n_477),
.B2(n_472),
.Y(n_736)
);

OAI22xp5_ASAP7_75t_L g737 ( 
.A1(n_715),
.A2(n_619),
.B1(n_616),
.B2(n_612),
.Y(n_737)
);

AOI22xp33_ASAP7_75t_SL g738 ( 
.A1(n_718),
.A2(n_608),
.B1(n_612),
.B2(n_610),
.Y(n_738)
);

AOI22xp33_ASAP7_75t_L g739 ( 
.A1(n_701),
.A2(n_510),
.B1(n_472),
.B2(n_477),
.Y(n_739)
);

AOI22xp33_ASAP7_75t_L g740 ( 
.A1(n_710),
.A2(n_510),
.B1(n_472),
.B2(n_477),
.Y(n_740)
);

AOI22xp33_ASAP7_75t_L g741 ( 
.A1(n_720),
.A2(n_510),
.B1(n_484),
.B2(n_494),
.Y(n_741)
);

INVx3_ASAP7_75t_L g742 ( 
.A(n_699),
.Y(n_742)
);

AOI22xp33_ASAP7_75t_L g743 ( 
.A1(n_714),
.A2(n_494),
.B1(n_484),
.B2(n_470),
.Y(n_743)
);

AOI22xp33_ASAP7_75t_L g744 ( 
.A1(n_680),
.A2(n_494),
.B1(n_484),
.B2(n_470),
.Y(n_744)
);

AOI22xp33_ASAP7_75t_L g745 ( 
.A1(n_681),
.A2(n_468),
.B1(n_471),
.B2(n_616),
.Y(n_745)
);

AOI22xp33_ASAP7_75t_L g746 ( 
.A1(n_695),
.A2(n_697),
.B1(n_698),
.B2(n_704),
.Y(n_746)
);

OAI22xp5_ASAP7_75t_L g747 ( 
.A1(n_676),
.A2(n_616),
.B1(n_612),
.B2(n_610),
.Y(n_747)
);

AOI22xp33_ASAP7_75t_L g748 ( 
.A1(n_702),
.A2(n_499),
.B1(n_511),
.B2(n_610),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_717),
.B(n_595),
.Y(n_749)
);

AOI22xp33_ASAP7_75t_L g750 ( 
.A1(n_702),
.A2(n_499),
.B1(n_511),
.B2(n_599),
.Y(n_750)
);

AOI22xp33_ASAP7_75t_SL g751 ( 
.A1(n_718),
.A2(n_608),
.B1(n_603),
.B2(n_595),
.Y(n_751)
);

AOI22xp33_ASAP7_75t_L g752 ( 
.A1(n_707),
.A2(n_511),
.B1(n_499),
.B2(n_599),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_679),
.B(n_603),
.Y(n_753)
);

AOI221xp5_ASAP7_75t_L g754 ( 
.A1(n_689),
.A2(n_514),
.B1(n_468),
.B2(n_471),
.C(n_464),
.Y(n_754)
);

AOI22xp5_ASAP7_75t_L g755 ( 
.A1(n_721),
.A2(n_507),
.B1(n_499),
.B2(n_603),
.Y(n_755)
);

AOI22xp33_ASAP7_75t_L g756 ( 
.A1(n_707),
.A2(n_603),
.B1(n_305),
.B2(n_301),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_712),
.B(n_603),
.Y(n_757)
);

AOI22xp33_ASAP7_75t_L g758 ( 
.A1(n_713),
.A2(n_305),
.B1(n_312),
.B2(n_47),
.Y(n_758)
);

AND2x2_ASAP7_75t_L g759 ( 
.A(n_699),
.B(n_45),
.Y(n_759)
);

AOI222xp33_ASAP7_75t_L g760 ( 
.A1(n_689),
.A2(n_305),
.B1(n_312),
.B2(n_54),
.C1(n_56),
.C2(n_57),
.Y(n_760)
);

OAI222xp33_ASAP7_75t_L g761 ( 
.A1(n_719),
.A2(n_46),
.B1(n_51),
.B2(n_58),
.C1(n_59),
.C2(n_60),
.Y(n_761)
);

AOI221xp5_ASAP7_75t_L g762 ( 
.A1(n_716),
.A2(n_61),
.B1(n_67),
.B2(n_70),
.C(n_71),
.Y(n_762)
);

NAND3xp33_ASAP7_75t_L g763 ( 
.A(n_760),
.B(n_684),
.C(n_719),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_746),
.B(n_684),
.Y(n_764)
);

NAND3xp33_ASAP7_75t_L g765 ( 
.A(n_726),
.B(n_722),
.C(n_723),
.Y(n_765)
);

AND2x2_ASAP7_75t_L g766 ( 
.A(n_746),
.B(n_711),
.Y(n_766)
);

AND2x2_ASAP7_75t_SL g767 ( 
.A(n_728),
.B(n_678),
.Y(n_767)
);

AOI22xp33_ASAP7_75t_L g768 ( 
.A1(n_762),
.A2(n_718),
.B1(n_682),
.B2(n_678),
.Y(n_768)
);

AND2x2_ASAP7_75t_L g769 ( 
.A(n_753),
.B(n_682),
.Y(n_769)
);

NAND3xp33_ASAP7_75t_L g770 ( 
.A(n_743),
.B(n_683),
.C(n_77),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_729),
.B(n_727),
.Y(n_771)
);

AND2x2_ASAP7_75t_L g772 ( 
.A(n_734),
.B(n_72),
.Y(n_772)
);

HB1xp67_ASAP7_75t_L g773 ( 
.A(n_757),
.Y(n_773)
);

AOI21xp5_ASAP7_75t_L g774 ( 
.A1(n_761),
.A2(n_79),
.B(n_81),
.Y(n_774)
);

OAI21xp5_ASAP7_75t_SL g775 ( 
.A1(n_730),
.A2(n_83),
.B(n_84),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_749),
.B(n_85),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_742),
.B(n_86),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_731),
.B(n_87),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_742),
.B(n_759),
.Y(n_779)
);

OAI21xp5_ASAP7_75t_SL g780 ( 
.A1(n_755),
.A2(n_88),
.B(n_89),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_725),
.B(n_90),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_735),
.B(n_91),
.Y(n_782)
);

OAI221xp5_ASAP7_75t_SL g783 ( 
.A1(n_756),
.A2(n_92),
.B1(n_93),
.B2(n_94),
.C(n_99),
.Y(n_783)
);

AND2x2_ASAP7_75t_SL g784 ( 
.A(n_752),
.B(n_100),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_754),
.B(n_101),
.Y(n_785)
);

NOR3xp33_ASAP7_75t_L g786 ( 
.A(n_737),
.B(n_103),
.C(n_105),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_745),
.B(n_111),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_745),
.B(n_113),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_747),
.B(n_114),
.Y(n_789)
);

OAI211xp5_ASAP7_75t_L g790 ( 
.A1(n_743),
.A2(n_115),
.B(n_116),
.C(n_117),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_773),
.Y(n_791)
);

NAND4xp75_ASAP7_75t_L g792 ( 
.A(n_774),
.B(n_751),
.C(n_738),
.D(n_750),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_779),
.B(n_724),
.Y(n_793)
);

NOR2x1_ASAP7_75t_L g794 ( 
.A(n_763),
.B(n_733),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_769),
.B(n_741),
.Y(n_795)
);

NAND3xp33_ASAP7_75t_L g796 ( 
.A(n_775),
.B(n_758),
.C(n_739),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_776),
.B(n_732),
.Y(n_797)
);

NAND3xp33_ASAP7_75t_L g798 ( 
.A(n_780),
.B(n_748),
.C(n_740),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_764),
.B(n_744),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_764),
.B(n_744),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_766),
.B(n_736),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_784),
.A2(n_118),
.B(n_120),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_766),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_769),
.B(n_121),
.Y(n_804)
);

NOR3xp33_ASAP7_75t_L g805 ( 
.A(n_770),
.B(n_122),
.C(n_124),
.Y(n_805)
);

INVx3_ASAP7_75t_L g806 ( 
.A(n_772),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_772),
.B(n_125),
.Y(n_807)
);

OA211x2_ASAP7_75t_L g808 ( 
.A1(n_771),
.A2(n_126),
.B(n_127),
.C(n_129),
.Y(n_808)
);

AOI221xp5_ASAP7_75t_L g809 ( 
.A1(n_763),
.A2(n_131),
.B1(n_132),
.B2(n_133),
.C(n_134),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_806),
.B(n_771),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_791),
.Y(n_811)
);

BUFx3_ASAP7_75t_L g812 ( 
.A(n_806),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_803),
.B(n_767),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_799),
.Y(n_814)
);

XNOR2x1_ASAP7_75t_L g815 ( 
.A(n_794),
.B(n_787),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_795),
.Y(n_816)
);

NAND4xp75_ASAP7_75t_L g817 ( 
.A(n_809),
.B(n_767),
.C(n_784),
.D(n_778),
.Y(n_817)
);

XNOR2xp5_ASAP7_75t_L g818 ( 
.A(n_792),
.B(n_807),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_800),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_793),
.Y(n_820)
);

NAND4xp75_ASAP7_75t_SL g821 ( 
.A(n_797),
.B(n_778),
.C(n_787),
.D(n_783),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_811),
.Y(n_822)
);

XNOR2x1_ASAP7_75t_L g823 ( 
.A(n_815),
.B(n_804),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_816),
.Y(n_824)
);

BUFx12f_ASAP7_75t_L g825 ( 
.A(n_812),
.Y(n_825)
);

AOI22xp5_ASAP7_75t_L g826 ( 
.A1(n_817),
.A2(n_796),
.B1(n_805),
.B2(n_798),
.Y(n_826)
);

OA22x2_ASAP7_75t_L g827 ( 
.A1(n_826),
.A2(n_818),
.B1(n_820),
.B2(n_815),
.Y(n_827)
);

HB1xp67_ASAP7_75t_L g828 ( 
.A(n_824),
.Y(n_828)
);

BUFx3_ASAP7_75t_L g829 ( 
.A(n_825),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_822),
.Y(n_830)
);

XNOR2x1_ASAP7_75t_L g831 ( 
.A(n_823),
.B(n_818),
.Y(n_831)
);

INVx3_ASAP7_75t_L g832 ( 
.A(n_829),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_828),
.Y(n_833)
);

INVxp67_ASAP7_75t_SL g834 ( 
.A(n_831),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_828),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_832),
.Y(n_836)
);

HB1xp67_ASAP7_75t_L g837 ( 
.A(n_835),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_832),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_837),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_836),
.Y(n_840)
);

AOI22xp5_ASAP7_75t_L g841 ( 
.A1(n_838),
.A2(n_827),
.B1(n_834),
.B2(n_826),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_837),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_841),
.B(n_832),
.Y(n_843)
);

AOI211xp5_ASAP7_75t_SL g844 ( 
.A1(n_839),
.A2(n_832),
.B(n_833),
.C(n_835),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_842),
.B(n_829),
.Y(n_845)
);

AOI221xp5_ASAP7_75t_L g846 ( 
.A1(n_840),
.A2(n_833),
.B1(n_835),
.B2(n_827),
.C(n_830),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_839),
.Y(n_847)
);

NAND4xp25_ASAP7_75t_L g848 ( 
.A(n_841),
.B(n_810),
.C(n_802),
.D(n_808),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_841),
.B(n_814),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_846),
.B(n_810),
.Y(n_850)
);

NOR2x1_ASAP7_75t_L g851 ( 
.A(n_843),
.B(n_821),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_845),
.B(n_816),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_847),
.Y(n_853)
);

OAI22xp5_ASAP7_75t_L g854 ( 
.A1(n_849),
.A2(n_819),
.B1(n_812),
.B2(n_813),
.Y(n_854)
);

OR2x2_ASAP7_75t_L g855 ( 
.A(n_848),
.B(n_844),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_847),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_847),
.Y(n_857)
);

NOR4xp25_ASAP7_75t_L g858 ( 
.A(n_855),
.B(n_790),
.C(n_782),
.D(n_785),
.Y(n_858)
);

AND4x1_ASAP7_75t_L g859 ( 
.A(n_851),
.B(n_786),
.C(n_781),
.D(n_798),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_853),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_856),
.Y(n_861)
);

A2O1A1Ixp33_ASAP7_75t_L g862 ( 
.A1(n_850),
.A2(n_857),
.B(n_852),
.C(n_854),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_853),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_853),
.Y(n_864)
);

NAND4xp75_ASAP7_75t_L g865 ( 
.A(n_851),
.B(n_777),
.C(n_789),
.D(n_788),
.Y(n_865)
);

OAI211xp5_ASAP7_75t_L g866 ( 
.A1(n_862),
.A2(n_768),
.B(n_819),
.C(n_765),
.Y(n_866)
);

A2O1A1Ixp33_ASAP7_75t_SL g867 ( 
.A1(n_860),
.A2(n_801),
.B(n_139),
.C(n_140),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_863),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_864),
.Y(n_869)
);

OR2x2_ASAP7_75t_L g870 ( 
.A(n_861),
.B(n_137),
.Y(n_870)
);

BUFx2_ASAP7_75t_L g871 ( 
.A(n_865),
.Y(n_871)
);

INVx1_ASAP7_75t_SL g872 ( 
.A(n_859),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_870),
.Y(n_873)
);

OAI22xp5_ASAP7_75t_L g874 ( 
.A1(n_872),
.A2(n_858),
.B1(n_142),
.B2(n_143),
.Y(n_874)
);

OAI22xp5_ASAP7_75t_L g875 ( 
.A1(n_871),
.A2(n_141),
.B1(n_146),
.B2(n_147),
.Y(n_875)
);

AOI22xp5_ASAP7_75t_L g876 ( 
.A1(n_866),
.A2(n_868),
.B1(n_869),
.B2(n_867),
.Y(n_876)
);

BUFx2_ASAP7_75t_L g877 ( 
.A(n_868),
.Y(n_877)
);

AOI22x1_ASAP7_75t_SL g878 ( 
.A1(n_872),
.A2(n_148),
.B1(n_150),
.B2(n_151),
.Y(n_878)
);

AOI22xp33_ASAP7_75t_L g879 ( 
.A1(n_871),
.A2(n_152),
.B1(n_155),
.B2(n_156),
.Y(n_879)
);

BUFx2_ASAP7_75t_L g880 ( 
.A(n_877),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_873),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_876),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_878),
.Y(n_883)
);

AOI22xp5_ASAP7_75t_L g884 ( 
.A1(n_882),
.A2(n_874),
.B1(n_875),
.B2(n_879),
.Y(n_884)
);

AOI22xp5_ASAP7_75t_L g885 ( 
.A1(n_883),
.A2(n_157),
.B1(n_158),
.B2(n_160),
.Y(n_885)
);

OR2x2_ASAP7_75t_L g886 ( 
.A(n_884),
.B(n_880),
.Y(n_886)
);

AO22x1_ASAP7_75t_L g887 ( 
.A1(n_886),
.A2(n_881),
.B1(n_885),
.B2(n_164),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_887),
.Y(n_888)
);

AOI221xp5_ASAP7_75t_L g889 ( 
.A1(n_888),
.A2(n_162),
.B1(n_163),
.B2(n_165),
.C(n_168),
.Y(n_889)
);

AOI211xp5_ASAP7_75t_L g890 ( 
.A1(n_889),
.A2(n_170),
.B(n_171),
.C(n_176),
.Y(n_890)
);


endmodule