module fake_jpeg_24027_n_334 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_334);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_334;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_3),
.B(n_16),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_33),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_33),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_22),
.B(n_0),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_42),
.B(n_48),
.Y(n_76)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_31),
.B(n_0),
.Y(n_46)
);

AND2x2_ASAP7_75t_SL g82 ( 
.A(n_46),
.B(n_50),
.Y(n_82)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_22),
.B(n_0),
.Y(n_48)
);

INVx6_ASAP7_75t_SL g49 ( 
.A(n_19),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_51),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_31),
.B(n_0),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_52),
.B(n_55),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_53),
.Y(n_87)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_43),
.A2(n_20),
.B1(n_18),
.B2(n_32),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_56),
.A2(n_57),
.B1(n_64),
.B2(n_66),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_43),
.A2(n_20),
.B1(n_18),
.B2(n_32),
.Y(n_57)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_60),
.B(n_65),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx11_ASAP7_75t_L g109 ( 
.A(n_61),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_25),
.Y(n_63)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_43),
.A2(n_20),
.B1(n_18),
.B2(n_32),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_43),
.A2(n_36),
.B1(n_24),
.B2(n_23),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_28),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_67),
.B(n_23),
.Y(n_122)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_68),
.B(n_75),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_40),
.A2(n_27),
.B1(n_35),
.B2(n_25),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_69),
.A2(n_85),
.B1(n_21),
.B2(n_28),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_48),
.B(n_29),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_70),
.B(n_72),
.Y(n_117)
);

BUFx4f_ASAP7_75t_SL g71 ( 
.A(n_44),
.Y(n_71)
);

INVx13_ASAP7_75t_L g111 ( 
.A(n_71),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_48),
.B(n_29),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_41),
.B(n_26),
.Y(n_73)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_78),
.B(n_27),
.Y(n_94)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_40),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_30),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_47),
.B(n_17),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_38),
.Y(n_88)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_81),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_47),
.A2(n_24),
.B1(n_23),
.B2(n_19),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_84),
.A2(n_23),
.B1(n_21),
.B2(n_34),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_47),
.A2(n_27),
.B1(n_26),
.B2(n_35),
.Y(n_85)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_39),
.Y(n_86)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_86),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_88),
.B(n_117),
.Y(n_158)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_91),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_82),
.B(n_37),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_92),
.B(n_93),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_37),
.Y(n_93)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_94),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_37),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_95),
.B(n_98),
.Y(n_134)
);

NAND3xp33_ASAP7_75t_L g96 ( 
.A(n_70),
.B(n_17),
.C(n_34),
.Y(n_96)
);

NAND3xp33_ASAP7_75t_L g151 ( 
.A(n_96),
.B(n_116),
.C(n_119),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_71),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_97),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_55),
.B(n_37),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_52),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_100),
.B(n_103),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_101),
.A2(n_77),
.B1(n_62),
.B2(n_38),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_60),
.B(n_39),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_102),
.B(n_105),
.Y(n_140)
);

A2O1A1Ixp33_ASAP7_75t_L g103 ( 
.A1(n_67),
.A2(n_41),
.B(n_49),
.C(n_23),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_65),
.B(n_39),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_68),
.B(n_51),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_106),
.B(n_108),
.Y(n_143)
);

INVx4_ASAP7_75t_SL g107 ( 
.A(n_53),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_107),
.B(n_110),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_76),
.B(n_51),
.Y(n_108)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_77),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_76),
.B(n_51),
.Y(n_114)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_114),
.Y(n_154)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_80),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_59),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_118),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_53),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_120),
.A2(n_49),
.B1(n_74),
.B2(n_54),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_75),
.B(n_49),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_121),
.B(n_122),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_115),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_124),
.B(n_125),
.Y(n_168)
);

INVxp33_ASAP7_75t_L g125 ( 
.A(n_94),
.Y(n_125)
);

BUFx2_ASAP7_75t_L g126 ( 
.A(n_107),
.Y(n_126)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_126),
.Y(n_160)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_109),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_128),
.B(n_133),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_92),
.A2(n_78),
.B1(n_79),
.B2(n_81),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_129),
.A2(n_135),
.B1(n_149),
.B2(n_152),
.Y(n_165)
);

AOI21xp33_ASAP7_75t_L g130 ( 
.A1(n_93),
.A2(n_72),
.B(n_30),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_130),
.A2(n_45),
.B(n_61),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_SL g132 ( 
.A(n_99),
.B(n_71),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_132),
.B(n_150),
.C(n_113),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_100),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_95),
.A2(n_74),
.B1(n_83),
.B2(n_58),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_123),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_136),
.B(n_137),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_97),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_122),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_138),
.B(n_144),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_142),
.A2(n_155),
.B1(n_111),
.B2(n_30),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_123),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_103),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_147),
.B(n_156),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_98),
.A2(n_58),
.B1(n_83),
.B2(n_54),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_106),
.B(n_71),
.C(n_39),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_102),
.A2(n_86),
.B1(n_62),
.B2(n_77),
.Y(n_152)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_99),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_105),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_157),
.A2(n_87),
.B1(n_111),
.B2(n_38),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_158),
.B(n_45),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_116),
.A2(n_38),
.B1(n_45),
.B2(n_30),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_159),
.A2(n_87),
.B1(n_119),
.B2(n_109),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_147),
.A2(n_114),
.B1(n_108),
.B2(n_88),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_161),
.A2(n_162),
.B1(n_178),
.B2(n_168),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_124),
.A2(n_104),
.B1(n_118),
.B2(n_110),
.Y(n_162)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_127),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_163),
.A2(n_189),
.B1(n_160),
.B2(n_186),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_141),
.A2(n_104),
.B(n_112),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_164),
.A2(n_173),
.B(n_193),
.Y(n_221)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_148),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_166),
.B(n_178),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_129),
.A2(n_117),
.B1(n_112),
.B2(n_113),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_167),
.A2(n_171),
.B1(n_183),
.B2(n_159),
.Y(n_194)
);

BUFx24_ASAP7_75t_SL g169 ( 
.A(n_156),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_169),
.B(n_174),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_170),
.B(n_134),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_135),
.A2(n_117),
.B1(n_87),
.B2(n_107),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_128),
.Y(n_174)
);

MAJx2_ASAP7_75t_L g175 ( 
.A(n_140),
.B(n_89),
.C(n_45),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_175),
.B(n_187),
.C(n_131),
.Y(n_213)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_149),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_179),
.A2(n_184),
.B1(n_185),
.B2(n_144),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_142),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_180),
.B(n_181),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_150),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_126),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_182),
.B(n_186),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_133),
.A2(n_89),
.B1(n_90),
.B2(n_111),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_126),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_146),
.B(n_157),
.C(n_132),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_152),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_188),
.B(n_191),
.Y(n_199)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_145),
.Y(n_189)
);

OAI21xp33_ASAP7_75t_L g190 ( 
.A1(n_143),
.A2(n_90),
.B(n_11),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_190),
.A2(n_138),
.B(n_136),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_140),
.B(n_61),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_194),
.A2(n_162),
.B1(n_165),
.B2(n_187),
.Y(n_225)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_172),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_196),
.B(n_202),
.Y(n_226)
);

OAI21xp33_ASAP7_75t_SL g230 ( 
.A1(n_197),
.A2(n_224),
.B(n_165),
.Y(n_230)
);

OAI32xp33_ASAP7_75t_L g198 ( 
.A1(n_161),
.A2(n_146),
.A3(n_154),
.B1(n_158),
.B2(n_134),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_198),
.B(n_9),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_177),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_200),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_201),
.B(n_8),
.Y(n_244)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_192),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_204),
.B(n_208),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_174),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_205),
.B(n_206),
.Y(n_235)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_179),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_207),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_191),
.B(n_158),
.Y(n_208)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_208),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_176),
.A2(n_154),
.B(n_153),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_209),
.A2(n_217),
.B(n_160),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_164),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_210),
.B(n_212),
.Y(n_237)
);

A2O1A1O1Ixp25_ASAP7_75t_L g211 ( 
.A1(n_193),
.A2(n_151),
.B(n_139),
.C(n_153),
.D(n_131),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_211),
.B(n_213),
.C(n_223),
.Y(n_234)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_171),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_188),
.A2(n_145),
.B1(n_97),
.B2(n_3),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_214),
.A2(n_220),
.B1(n_215),
.B2(n_197),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_173),
.B(n_1),
.Y(n_215)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_215),
.Y(n_246)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_167),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_216),
.B(n_219),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_181),
.A2(n_2),
.B(n_3),
.Y(n_217)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_163),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_180),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_170),
.B(n_2),
.C(n_5),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_225),
.A2(n_231),
.B1(n_244),
.B2(n_249),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_227),
.B(n_232),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_221),
.A2(n_166),
.B(n_182),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_228),
.A2(n_238),
.B(n_217),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_229),
.B(n_242),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_230),
.A2(n_206),
.B1(n_216),
.B2(n_243),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_212),
.A2(n_175),
.B1(n_189),
.B2(n_5),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_204),
.B(n_11),
.Y(n_232)
);

A2O1A1Ixp33_ASAP7_75t_L g256 ( 
.A1(n_233),
.A2(n_239),
.B(n_220),
.C(n_224),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_213),
.B(n_5),
.C(n_16),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_236),
.B(n_223),
.C(n_210),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_218),
.A2(n_6),
.B(n_7),
.Y(n_238)
);

A2O1A1Ixp33_ASAP7_75t_L g239 ( 
.A1(n_221),
.A2(n_6),
.B(n_8),
.C(n_9),
.Y(n_239)
);

CKINVDCx14_ASAP7_75t_R g242 ( 
.A(n_222),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_243),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_199),
.B(n_9),
.Y(n_247)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_247),
.Y(n_259)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_214),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_251),
.A2(n_253),
.B1(n_262),
.B2(n_265),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_240),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_252),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_240),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_255),
.B(n_266),
.Y(n_271)
);

CKINVDCx14_ASAP7_75t_R g277 ( 
.A(n_256),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_258),
.B(n_236),
.C(n_234),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_248),
.A2(n_199),
.B1(n_203),
.B2(n_202),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_260),
.A2(n_264),
.B1(n_231),
.B2(n_233),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_245),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_261),
.B(n_269),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_248),
.A2(n_209),
.B(n_196),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_237),
.A2(n_200),
.B1(n_198),
.B2(n_211),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_228),
.A2(n_205),
.B(n_201),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_226),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_226),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_267),
.B(n_269),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_227),
.B(n_195),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_268),
.B(n_232),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_235),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_260),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_270),
.B(n_276),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_272),
.A2(n_250),
.B1(n_259),
.B2(n_241),
.Y(n_294)
);

O2A1O1Ixp33_ASAP7_75t_L g273 ( 
.A1(n_254),
.A2(n_229),
.B(n_247),
.C(n_249),
.Y(n_273)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_273),
.Y(n_291)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_263),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_278),
.B(n_283),
.Y(n_301)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_262),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_279),
.B(n_280),
.Y(n_292)
);

BUFx24_ASAP7_75t_SL g280 ( 
.A(n_268),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_266),
.B(n_246),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_281),
.Y(n_297)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_265),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_282),
.B(n_286),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_257),
.B(n_234),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_285),
.B(n_287),
.C(n_258),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_259),
.B(n_246),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_284),
.B(n_257),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_288),
.B(n_296),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_290),
.B(n_295),
.C(n_274),
.Y(n_307)
);

BUFx12_ASAP7_75t_L g293 ( 
.A(n_275),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_293),
.B(n_298),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_294),
.A2(n_277),
.B1(n_281),
.B2(n_261),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_285),
.B(n_241),
.C(n_264),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_SL g296 ( 
.A(n_272),
.B(n_225),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_283),
.B(n_253),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_270),
.A2(n_251),
.B1(n_256),
.B2(n_239),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_299),
.A2(n_273),
.B1(n_291),
.B2(n_276),
.Y(n_304)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_302),
.Y(n_313)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_289),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_303),
.B(n_304),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_290),
.A2(n_297),
.B(n_271),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_306),
.B(n_301),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_307),
.B(n_309),
.C(n_311),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_297),
.A2(n_274),
.B(n_287),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_300),
.B(n_244),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_310),
.B(n_293),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_301),
.B(n_278),
.C(n_219),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_312),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_307),
.A2(n_296),
.B1(n_295),
.B2(n_288),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_316),
.A2(n_311),
.B1(n_308),
.B2(n_305),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_304),
.B(n_293),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_317),
.B(n_318),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_309),
.B(n_292),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_319),
.B(n_314),
.Y(n_323)
);

OAI21x1_ASAP7_75t_L g326 ( 
.A1(n_322),
.A2(n_323),
.B(n_324),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_315),
.B(n_313),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_321),
.Y(n_325)
);

OR2x2_ASAP7_75t_L g329 ( 
.A(n_325),
.B(n_327),
.Y(n_329)
);

A2O1A1Ixp33_ASAP7_75t_SL g327 ( 
.A1(n_320),
.A2(n_305),
.B(n_314),
.C(n_316),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g328 ( 
.A(n_326),
.B(n_322),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_328),
.A2(n_238),
.B(n_13),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_12),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_331),
.A2(n_329),
.B(n_13),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_332),
.A2(n_12),
.B1(n_14),
.B2(n_16),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_12),
.C(n_14),
.Y(n_334)
);


endmodule