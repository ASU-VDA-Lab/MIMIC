module fake_jpeg_3217_n_57 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_57);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_57;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

INVx6_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_7),
.B(n_3),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

CKINVDCx14_ASAP7_75t_R g11 ( 
.A(n_5),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_1),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_6),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

INVx6_ASAP7_75t_SL g18 ( 
.A(n_11),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_18),
.B(n_21),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_20),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_22),
.B(n_13),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_17),
.B(n_10),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_12),
.C(n_15),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_13),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_21),
.B(n_14),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_29),
.B(n_18),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_27),
.A2(n_20),
.B1(n_19),
.B2(n_16),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_33),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_32),
.Y(n_42)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_34),
.B(n_35),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_36),
.B(n_12),
.C(n_26),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_SL g37 ( 
.A1(n_31),
.A2(n_26),
.B(n_25),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_38),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g39 ( 
.A1(n_36),
.A2(n_25),
.B(n_8),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_30),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_43),
.B(n_45),
.Y(n_50)
);

FAx1_ASAP7_75t_SL g45 ( 
.A(n_42),
.B(n_8),
.CI(n_1),
.CON(n_45),
.SN(n_45)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_41),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_46),
.A2(n_40),
.B1(n_2),
.B2(n_0),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_0),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g49 ( 
.A(n_47),
.B(n_2),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_48),
.B(n_49),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_50),
.B(n_44),
.C(n_47),
.Y(n_51)
);

MAJx2_ASAP7_75t_L g53 ( 
.A(n_51),
.B(n_44),
.C(n_49),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_53),
.B(n_54),
.C(n_45),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_SL g54 ( 
.A1(n_52),
.A2(n_45),
.B(n_43),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_55),
.A2(n_43),
.B1(n_48),
.B2(n_4),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_56),
.B(n_7),
.Y(n_57)
);


endmodule