module real_aes_4582_n_249 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_942, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_246, n_248, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_249);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_942;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_249;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_905;
wire n_878;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_329;
wire n_852;
wire n_766;
wire n_919;
wire n_857;
wire n_461;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_923;
wire n_894;
wire n_429;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_767;
wire n_696;
wire n_889;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_932;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_918;
wire n_478;
wire n_356;
wire n_883;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_892;
wire n_495;
wire n_370;
wire n_938;
wire n_384;
wire n_744;
wire n_352;
wire n_935;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_906;
wire n_263;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_693;
wire n_281;
wire n_496;
wire n_468;
wire n_746;
wire n_284;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_523;
wire n_298;
wire n_909;
wire n_439;
wire n_576;
wire n_924;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_671;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_925;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_737;
wire n_581;
wire n_610;
wire n_936;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_940;
wire n_770;
wire n_808;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_417;
wire n_363;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_807;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_913;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_917;
wire n_361;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_296;
wire n_702;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_756;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_269;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_934;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_927;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_291;
wire n_907;
wire n_847;
wire n_779;
wire n_481;
wire n_691;
wire n_498;
wire n_765;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_487;
wire n_831;
wire n_653;
wire n_365;
wire n_899;
wire n_526;
wire n_290;
wire n_637;
wire n_928;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_922;
wire n_520;
wire n_633;
wire n_679;
wire n_926;
wire n_472;
wire n_866;
wire n_452;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_623;
wire n_721;
wire n_446;
wire n_681;
wire n_359;
wire n_456;
wire n_717;
wire n_712;
wire n_266;
wire n_312;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_639;
wire n_587;
wire n_811;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_888;
wire n_836;
wire n_793;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_921;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_842;
wire n_259;
wire n_849;
wire n_475;
wire n_554;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp5_ASAP7_75t_L g358 ( .A1(n_0), .A2(n_207), .B1(n_359), .B2(n_365), .Y(n_358) );
AOI22xp5_ASAP7_75t_L g755 ( .A1(n_1), .A2(n_53), .B1(n_718), .B2(n_721), .Y(n_755) );
HB1xp67_ASAP7_75t_L g261 ( .A(n_2), .Y(n_261) );
AND2x4_ASAP7_75t_L g687 ( .A(n_2), .B(n_239), .Y(n_687) );
AND2x4_ASAP7_75t_L g692 ( .A(n_2), .B(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g489 ( .A(n_3), .Y(n_489) );
INVx1_ASAP7_75t_L g443 ( .A(n_4), .Y(n_443) );
AOI22xp5_ASAP7_75t_L g390 ( .A1(n_5), .A2(n_40), .B1(n_326), .B2(n_391), .Y(n_390) );
AOI22xp5_ASAP7_75t_L g910 ( .A1(n_6), .A2(n_160), .B1(n_610), .B2(n_613), .Y(n_910) );
AOI22xp33_ASAP7_75t_L g469 ( .A1(n_7), .A2(n_216), .B1(n_299), .B2(n_470), .Y(n_469) );
AOI22xp33_ASAP7_75t_L g461 ( .A1(n_8), .A2(n_61), .B1(n_371), .B2(n_462), .Y(n_461) );
AOI22xp33_ASAP7_75t_L g642 ( .A1(n_9), .A2(n_21), .B1(n_430), .B2(n_431), .Y(n_642) );
AOI22xp33_ASAP7_75t_L g904 ( .A1(n_10), .A2(n_223), .B1(n_594), .B2(n_603), .Y(n_904) );
AOI21xp33_ASAP7_75t_L g596 ( .A1(n_11), .A2(n_597), .B(n_598), .Y(n_596) );
AOI22xp5_ASAP7_75t_L g652 ( .A1(n_12), .A2(n_105), .B1(n_466), .B2(n_468), .Y(n_652) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_13), .A2(n_172), .B1(n_612), .B2(n_613), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_14), .A2(n_20), .B1(n_526), .B2(n_527), .Y(n_525) );
AOI21xp5_ASAP7_75t_L g646 ( .A1(n_15), .A2(n_274), .B(n_647), .Y(n_646) );
AOI22xp33_ASAP7_75t_L g398 ( .A1(n_16), .A2(n_215), .B1(n_399), .B2(n_400), .Y(n_398) );
XNOR2x2_ASAP7_75t_L g481 ( .A(n_17), .B(n_482), .Y(n_481) );
AOI22xp5_ASAP7_75t_L g754 ( .A1(n_17), .A2(n_77), .B1(n_696), .B2(n_711), .Y(n_754) );
AOI22xp33_ASAP7_75t_L g662 ( .A1(n_18), .A2(n_245), .B1(n_604), .B2(n_610), .Y(n_662) );
AOI22xp33_ASAP7_75t_L g394 ( .A1(n_19), .A2(n_135), .B1(n_395), .B2(n_397), .Y(n_394) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_22), .A2(n_54), .B1(n_380), .B2(n_408), .Y(n_456) );
AOI22xp33_ASAP7_75t_L g902 ( .A1(n_23), .A2(n_205), .B1(n_593), .B2(n_903), .Y(n_902) );
AOI22xp33_ASAP7_75t_L g930 ( .A1(n_24), .A2(n_151), .B1(n_606), .B2(n_607), .Y(n_930) );
XNOR2x1_ASAP7_75t_L g268 ( .A(n_25), .B(n_269), .Y(n_268) );
AO22x1_ASAP7_75t_L g913 ( .A1(n_26), .A2(n_145), .B1(n_606), .B2(n_607), .Y(n_913) );
AOI22xp33_ASAP7_75t_SL g348 ( .A1(n_27), .A2(n_191), .B1(n_349), .B2(n_354), .Y(n_348) );
INVx1_ASAP7_75t_L g744 ( .A(n_28), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_29), .B(n_472), .Y(n_471) );
AOI22xp5_ASAP7_75t_L g574 ( .A1(n_30), .A2(n_130), .B1(n_407), .B2(n_575), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g465 ( .A1(n_31), .A2(n_244), .B1(n_466), .B2(n_468), .Y(n_465) );
AOI22xp33_ASAP7_75t_L g623 ( .A1(n_32), .A2(n_68), .B1(n_411), .B2(n_430), .Y(n_623) );
INVx1_ASAP7_75t_L g304 ( .A(n_33), .Y(n_304) );
AOI22xp33_ASAP7_75t_L g649 ( .A1(n_34), .A2(n_189), .B1(n_445), .B2(n_546), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g683 ( .A1(n_35), .A2(n_74), .B1(n_684), .B2(n_688), .Y(n_683) );
AOI22xp5_ASAP7_75t_L g559 ( .A1(n_36), .A2(n_71), .B1(n_560), .B2(n_561), .Y(n_559) );
INVx1_ASAP7_75t_SL g794 ( .A(n_37), .Y(n_794) );
AOI22xp33_ASAP7_75t_L g458 ( .A1(n_38), .A2(n_181), .B1(n_430), .B2(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g673 ( .A(n_39), .Y(n_673) );
AOI21xp5_ASAP7_75t_L g905 ( .A1(n_41), .A2(n_672), .B(n_906), .Y(n_905) );
NOR2xp33_ASAP7_75t_L g259 ( .A(n_42), .B(n_187), .Y(n_259) );
INVx1_ASAP7_75t_L g294 ( .A(n_42), .Y(n_294) );
INVxp67_ASAP7_75t_L g338 ( .A(n_42), .Y(n_338) );
AOI22xp33_ASAP7_75t_L g566 ( .A1(n_43), .A2(n_120), .B1(n_274), .B2(n_475), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g726 ( .A1(n_44), .A2(n_81), .B1(n_691), .B2(n_706), .Y(n_726) );
AOI22xp33_ASAP7_75t_L g605 ( .A1(n_45), .A2(n_58), .B1(n_606), .B2(n_607), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_46), .B(n_306), .Y(n_393) );
AOI22xp33_ASAP7_75t_L g671 ( .A1(n_47), .A2(n_134), .B1(n_594), .B2(n_672), .Y(n_671) );
AO22x1_ASAP7_75t_L g911 ( .A1(n_48), .A2(n_142), .B1(n_604), .B2(n_612), .Y(n_911) );
NAND2xp5_ASAP7_75t_SL g290 ( .A(n_49), .B(n_279), .Y(n_290) );
INVx1_ASAP7_75t_L g324 ( .A(n_50), .Y(n_324) );
AOI22xp33_ASAP7_75t_L g428 ( .A1(n_51), .A2(n_155), .B1(n_349), .B2(n_403), .Y(n_428) );
AOI22xp33_ASAP7_75t_L g426 ( .A1(n_52), .A2(n_76), .B1(n_377), .B2(n_380), .Y(n_426) );
AOI22xp33_ASAP7_75t_L g406 ( .A1(n_55), .A2(n_208), .B1(n_407), .B2(n_408), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g702 ( .A1(n_56), .A2(n_248), .B1(n_703), .B2(n_704), .Y(n_702) );
CKINVDCx20_ASAP7_75t_R g719 ( .A(n_57), .Y(n_719) );
AOI22xp33_ASAP7_75t_L g518 ( .A1(n_59), .A2(n_197), .B1(n_519), .B2(n_521), .Y(n_518) );
INVxp67_ASAP7_75t_R g746 ( .A(n_60), .Y(n_746) );
AOI22xp5_ASAP7_75t_L g499 ( .A1(n_62), .A2(n_232), .B1(n_411), .B2(n_500), .Y(n_499) );
AOI22xp33_ASAP7_75t_SL g370 ( .A1(n_63), .A2(n_230), .B1(n_371), .B2(n_373), .Y(n_370) );
INVx2_ASAP7_75t_L g256 ( .A(n_64), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g901 ( .A(n_65), .B(n_597), .Y(n_901) );
AOI22xp33_ASAP7_75t_L g486 ( .A1(n_66), .A2(n_126), .B1(n_377), .B2(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g686 ( .A(n_67), .Y(n_686) );
AND2x4_ASAP7_75t_L g689 ( .A(n_67), .B(n_256), .Y(n_689) );
INVx1_ASAP7_75t_SL g712 ( .A(n_67), .Y(n_712) );
AOI22xp33_ASAP7_75t_SL g542 ( .A1(n_69), .A2(n_247), .B1(n_543), .B2(n_544), .Y(n_542) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_70), .A2(n_97), .B1(n_591), .B2(n_593), .Y(n_667) );
INVx1_ASAP7_75t_L g387 ( .A(n_72), .Y(n_387) );
AOI22xp5_ASAP7_75t_L g729 ( .A1(n_72), .A2(n_180), .B1(n_696), .B2(n_711), .Y(n_729) );
BUFx6f_ASAP7_75t_L g279 ( .A(n_73), .Y(n_279) );
AOI22xp33_ASAP7_75t_L g621 ( .A1(n_75), .A2(n_80), .B1(n_407), .B2(n_408), .Y(n_621) );
AOI22xp33_ASAP7_75t_L g409 ( .A1(n_78), .A2(n_178), .B1(n_410), .B2(n_411), .Y(n_409) );
INVx1_ASAP7_75t_L g272 ( .A(n_79), .Y(n_272) );
AOI21x1_ASAP7_75t_SL g437 ( .A1(n_82), .A2(n_438), .B(n_442), .Y(n_437) );
AOI22xp33_ASAP7_75t_L g433 ( .A1(n_83), .A2(n_154), .B1(n_299), .B2(n_434), .Y(n_433) );
CKINVDCx16_ASAP7_75t_R g742 ( .A(n_84), .Y(n_742) );
AOI22xp33_ASAP7_75t_L g690 ( .A1(n_85), .A2(n_156), .B1(n_691), .B2(n_694), .Y(n_690) );
AOI22xp5_ASAP7_75t_L g402 ( .A1(n_86), .A2(n_157), .B1(n_403), .B2(n_404), .Y(n_402) );
AOI22xp33_ASAP7_75t_L g931 ( .A1(n_87), .A2(n_212), .B1(n_590), .B2(n_609), .Y(n_931) );
AOI22xp33_ASAP7_75t_L g435 ( .A1(n_88), .A2(n_113), .B1(n_397), .B2(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g283 ( .A(n_89), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_89), .B(n_186), .Y(n_335) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_90), .A2(n_110), .B1(n_609), .B2(n_612), .Y(n_663) );
INVx1_ASAP7_75t_L g495 ( .A(n_91), .Y(n_495) );
OAI22x1_ASAP7_75t_L g637 ( .A1(n_92), .A2(n_638), .B1(n_643), .B2(n_653), .Y(n_637) );
NAND5xp2_ASAP7_75t_SL g638 ( .A(n_92), .B(n_639), .C(n_640), .D(n_641), .E(n_642), .Y(n_638) );
AOI22xp33_ASAP7_75t_L g474 ( .A1(n_93), .A2(n_132), .B1(n_449), .B2(n_475), .Y(n_474) );
AOI22xp33_ASAP7_75t_L g429 ( .A1(n_94), .A2(n_164), .B1(n_430), .B2(n_431), .Y(n_429) );
AOI22xp33_ASAP7_75t_L g423 ( .A1(n_95), .A2(n_183), .B1(n_424), .B2(n_425), .Y(n_423) );
XNOR2x1_ASAP7_75t_L g586 ( .A(n_96), .B(n_587), .Y(n_586) );
AOI22xp5_ASAP7_75t_L g929 ( .A1(n_98), .A2(n_243), .B1(n_604), .B2(n_610), .Y(n_929) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_99), .B(n_533), .Y(n_666) );
INVx1_ASAP7_75t_L g713 ( .A(n_100), .Y(n_713) );
AOI22xp33_ASAP7_75t_L g725 ( .A1(n_101), .A2(n_159), .B1(n_684), .B2(n_704), .Y(n_725) );
INVx1_ASAP7_75t_L g907 ( .A(n_102), .Y(n_907) );
AOI221xp5_ASAP7_75t_SL g933 ( .A1(n_103), .A2(n_220), .B1(n_493), .B2(n_603), .C(n_934), .Y(n_933) );
AOI22xp5_ASAP7_75t_L g622 ( .A1(n_104), .A2(n_210), .B1(n_373), .B2(n_414), .Y(n_622) );
AOI22xp33_ASAP7_75t_L g640 ( .A1(n_106), .A2(n_173), .B1(n_371), .B2(n_373), .Y(n_640) );
CKINVDCx5p33_ASAP7_75t_R g935 ( .A(n_107), .Y(n_935) );
AOI221xp5_ASAP7_75t_L g936 ( .A1(n_108), .A2(n_168), .B1(n_591), .B2(n_593), .C(n_937), .Y(n_936) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_109), .A2(n_213), .B1(n_609), .B2(n_610), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g457 ( .A1(n_111), .A2(n_211), .B1(n_349), .B2(n_403), .Y(n_457) );
AOI22xp33_ASAP7_75t_L g522 ( .A1(n_112), .A2(n_165), .B1(n_523), .B2(n_524), .Y(n_522) );
INVx1_ASAP7_75t_L g535 ( .A(n_114), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_115), .B(n_493), .Y(n_595) );
AOI22xp5_ASAP7_75t_L g567 ( .A1(n_116), .A2(n_169), .B1(n_473), .B2(n_568), .Y(n_567) );
INVx1_ASAP7_75t_L g617 ( .A(n_117), .Y(n_617) );
AOI22xp5_ASAP7_75t_L g932 ( .A1(n_118), .A2(n_149), .B1(n_612), .B2(n_613), .Y(n_932) );
NAND2xp33_ASAP7_75t_L g554 ( .A(n_119), .B(n_487), .Y(n_554) );
AOI22xp33_ASAP7_75t_L g796 ( .A1(n_121), .A2(n_163), .B1(n_688), .B2(n_703), .Y(n_796) );
INVx1_ASAP7_75t_L g599 ( .A(n_122), .Y(n_599) );
AOI22xp33_ASAP7_75t_L g639 ( .A1(n_123), .A2(n_221), .B1(n_377), .B2(n_380), .Y(n_639) );
AOI22xp33_ASAP7_75t_L g329 ( .A1(n_124), .A2(n_182), .B1(n_330), .B2(n_339), .Y(n_329) );
AO22x1_ASAP7_75t_L g912 ( .A1(n_125), .A2(n_237), .B1(n_590), .B2(n_609), .Y(n_912) );
AOI22xp5_ASAP7_75t_L g641 ( .A1(n_127), .A2(n_200), .B1(n_349), .B2(n_403), .Y(n_641) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_128), .A2(n_141), .B1(n_462), .B2(n_502), .Y(n_501) );
AOI21xp33_ASAP7_75t_SL g530 ( .A1(n_129), .A2(n_531), .B(n_534), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g504 ( .A1(n_131), .A2(n_158), .B1(n_475), .B2(n_505), .Y(n_504) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_133), .A2(n_229), .B1(n_603), .B2(n_604), .Y(n_602) );
AOI22xp33_ASAP7_75t_SL g376 ( .A1(n_136), .A2(n_214), .B1(n_377), .B2(n_380), .Y(n_376) );
INVx1_ASAP7_75t_L g447 ( .A(n_137), .Y(n_447) );
AOI22xp33_ASAP7_75t_L g592 ( .A1(n_138), .A2(n_192), .B1(n_593), .B2(n_594), .Y(n_592) );
AOI22xp5_ASAP7_75t_L g513 ( .A1(n_139), .A2(n_162), .B1(n_514), .B2(n_517), .Y(n_513) );
INVx1_ASAP7_75t_L g648 ( .A(n_140), .Y(n_648) );
AOI22xp33_ASAP7_75t_L g620 ( .A1(n_143), .A2(n_144), .B1(n_380), .B2(n_403), .Y(n_620) );
INVx1_ASAP7_75t_L g716 ( .A(n_146), .Y(n_716) );
AOI22xp5_ASAP7_75t_L g730 ( .A1(n_147), .A2(n_219), .B1(n_718), .B2(n_721), .Y(n_730) );
AO22x1_ASAP7_75t_L g937 ( .A1(n_148), .A2(n_206), .B1(n_594), .B2(n_597), .Y(n_937) );
AOI22x1_ASAP7_75t_L g509 ( .A1(n_150), .A2(n_510), .B1(n_511), .B2(n_547), .Y(n_509) );
INVx1_ASAP7_75t_L g547 ( .A(n_150), .Y(n_547) );
OAI22x1_ASAP7_75t_L g579 ( .A1(n_150), .A2(n_510), .B1(n_511), .B2(n_547), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g661 ( .A1(n_152), .A2(n_218), .B1(n_590), .B2(n_613), .Y(n_661) );
INVx1_ASAP7_75t_L g297 ( .A(n_153), .Y(n_297) );
XNOR2x2_ASAP7_75t_L g898 ( .A(n_159), .B(n_899), .Y(n_898) );
AOI22xp33_ASAP7_75t_L g919 ( .A1(n_159), .A2(n_920), .B1(n_922), .B2(n_938), .Y(n_919) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_161), .B(n_339), .Y(n_537) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_166), .A2(n_194), .B1(n_590), .B2(n_591), .Y(n_589) );
INVx1_ASAP7_75t_L g628 ( .A(n_167), .Y(n_628) );
OA22x2_ASAP7_75t_L g277 ( .A1(n_170), .A2(n_187), .B1(n_278), .B2(n_279), .Y(n_277) );
INVx1_ASAP7_75t_L g320 ( .A(n_170), .Y(n_320) );
AOI22xp5_ASAP7_75t_L g571 ( .A1(n_171), .A2(n_184), .B1(n_572), .B2(n_573), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_174), .A2(n_195), .B1(n_399), .B2(n_507), .Y(n_506) );
AOI221xp5_ASAP7_75t_L g625 ( .A1(n_175), .A2(n_201), .B1(n_306), .B2(n_626), .C(n_627), .Y(n_625) );
INVx1_ASAP7_75t_L g670 ( .A(n_176), .Y(n_670) );
XNOR2x1_ASAP7_75t_L g420 ( .A(n_177), .B(n_421), .Y(n_420) );
AOI221x1_ASAP7_75t_L g555 ( .A1(n_179), .A2(n_222), .B1(n_500), .B2(n_556), .C(n_557), .Y(n_555) );
CKINVDCx6p67_ASAP7_75t_R g741 ( .A(n_185), .Y(n_741) );
INVx1_ASAP7_75t_L g296 ( .A(n_186), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_186), .B(n_318), .Y(n_345) );
OAI21xp33_ASAP7_75t_L g321 ( .A1(n_187), .A2(n_196), .B(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g557 ( .A(n_188), .B(n_520), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g705 ( .A1(n_190), .A2(n_246), .B1(n_691), .B2(n_706), .Y(n_705) );
AOI22xp33_ASAP7_75t_L g631 ( .A1(n_193), .A2(n_204), .B1(n_299), .B2(n_445), .Y(n_631) );
NOR2xp33_ASAP7_75t_L g260 ( .A(n_196), .B(n_233), .Y(n_260) );
INVx1_ASAP7_75t_L g285 ( .A(n_196), .Y(n_285) );
AOI22xp33_ASAP7_75t_L g664 ( .A1(n_198), .A2(n_228), .B1(n_606), .B2(n_607), .Y(n_664) );
AOI21xp33_ASAP7_75t_L g492 ( .A1(n_199), .A2(n_493), .B(n_494), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_202), .B(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g795 ( .A(n_203), .Y(n_795) );
AOI22xp33_ASAP7_75t_L g538 ( .A1(n_209), .A2(n_217), .B1(n_539), .B2(n_541), .Y(n_538) );
AOI22xp5_ASAP7_75t_L g412 ( .A1(n_224), .A2(n_236), .B1(n_413), .B2(n_414), .Y(n_412) );
NOR3xp33_ASAP7_75t_L g552 ( .A(n_225), .B(n_553), .C(n_558), .Y(n_552) );
AOI22xp5_ASAP7_75t_L g577 ( .A1(n_225), .A2(n_558), .B1(n_565), .B2(n_942), .Y(n_577) );
OAI21xp5_ASAP7_75t_L g578 ( .A1(n_225), .A2(n_553), .B(n_570), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g632 ( .A1(n_226), .A2(n_242), .B1(n_434), .B2(n_468), .Y(n_632) );
INVx1_ASAP7_75t_L g311 ( .A(n_227), .Y(n_311) );
INVx1_ASAP7_75t_L g452 ( .A(n_231), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_233), .B(n_289), .Y(n_288) );
AOI22xp33_ASAP7_75t_L g484 ( .A1(n_234), .A2(n_240), .B1(n_414), .B2(n_485), .Y(n_484) );
AOI21xp33_ASAP7_75t_L g668 ( .A1(n_235), .A2(n_603), .B(n_669), .Y(n_668) );
OAI22xp5_ASAP7_75t_L g922 ( .A1(n_238), .A2(n_923), .B1(n_924), .B2(n_925), .Y(n_922) );
CKINVDCx20_ASAP7_75t_R g923 ( .A(n_238), .Y(n_923) );
INVx1_ASAP7_75t_L g693 ( .A(n_239), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_241), .B(n_651), .Y(n_650) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_262), .B(n_674), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
BUFx3_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
HB1xp67_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
NAND3xp33_ASAP7_75t_L g253 ( .A(n_254), .B(n_257), .C(n_261), .Y(n_253) );
AND2x2_ASAP7_75t_L g916 ( .A(n_254), .B(n_917), .Y(n_916) );
AND2x2_ASAP7_75t_L g921 ( .A(n_254), .B(n_918), .Y(n_921) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
OA21x2_ASAP7_75t_L g939 ( .A1(n_255), .A2(n_712), .B(n_940), .Y(n_939) );
HB1xp67_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g685 ( .A(n_256), .B(n_686), .Y(n_685) );
AND3x4_ASAP7_75t_L g711 ( .A(n_256), .B(n_692), .C(n_712), .Y(n_711) );
NOR2xp33_ASAP7_75t_L g917 ( .A(n_257), .B(n_918), .Y(n_917) );
HB1xp67_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
AO21x2_ASAP7_75t_L g342 ( .A1(n_258), .A2(n_343), .B(n_344), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_259), .B(n_260), .Y(n_258) );
INVx1_ASAP7_75t_L g918 ( .A(n_261), .Y(n_918) );
XNOR2xp5_ASAP7_75t_L g262 ( .A(n_263), .B(n_582), .Y(n_262) );
AOI22xp5_ASAP7_75t_L g263 ( .A1(n_264), .A2(n_478), .B1(n_580), .B2(n_581), .Y(n_263) );
INVx1_ASAP7_75t_L g581 ( .A(n_264), .Y(n_581) );
AOI22xp5_ASAP7_75t_L g264 ( .A1(n_265), .A2(n_417), .B1(n_418), .B2(n_477), .Y(n_264) );
INVx1_ASAP7_75t_L g477 ( .A(n_265), .Y(n_477) );
OAI22xp5_ASAP7_75t_L g265 ( .A1(n_266), .A2(n_267), .B1(n_382), .B2(n_415), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
INVx2_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_346), .Y(n_269) );
NOR3xp33_ASAP7_75t_L g270 ( .A(n_271), .B(n_303), .C(n_323), .Y(n_270) );
OAI22xp5_ASAP7_75t_L g271 ( .A1(n_272), .A2(n_273), .B1(n_297), .B2(n_298), .Y(n_271) );
INVx2_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
BUFx3_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
INVx1_ASAP7_75t_L g396 ( .A(n_275), .Y(n_396) );
BUFx6f_ASAP7_75t_L g434 ( .A(n_275), .Y(n_434) );
BUFx3_ASAP7_75t_L g505 ( .A(n_275), .Y(n_505) );
AND2x4_ASAP7_75t_L g275 ( .A(n_276), .B(n_286), .Y(n_275) );
AND2x4_ASAP7_75t_L g308 ( .A(n_276), .B(n_309), .Y(n_308) );
AND2x4_ASAP7_75t_L g603 ( .A(n_276), .B(n_286), .Y(n_603) );
AND2x2_ASAP7_75t_L g672 ( .A(n_276), .B(n_309), .Y(n_672) );
AND2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_280), .Y(n_276) );
AND2x2_ASAP7_75t_L g302 ( .A(n_277), .B(n_281), .Y(n_302) );
AND2x2_ASAP7_75t_L g336 ( .A(n_277), .B(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g364 ( .A(n_277), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_278), .B(n_285), .Y(n_284) );
INVx2_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
NAND2xp33_ASAP7_75t_L g282 ( .A(n_279), .B(n_283), .Y(n_282) );
INVx3_ASAP7_75t_L g289 ( .A(n_279), .Y(n_289) );
NAND2xp33_ASAP7_75t_L g295 ( .A(n_279), .B(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g322 ( .A(n_279), .Y(n_322) );
HB1xp67_ASAP7_75t_L g334 ( .A(n_279), .Y(n_334) );
AND2x4_ASAP7_75t_L g363 ( .A(n_280), .B(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_282), .B(n_284), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_283), .B(n_320), .Y(n_319) );
OAI21xp5_ASAP7_75t_L g337 ( .A1(n_285), .A2(n_322), .B(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g301 ( .A(n_286), .B(n_302), .Y(n_301) );
AND2x4_ASAP7_75t_L g362 ( .A(n_286), .B(n_363), .Y(n_362) );
AND2x4_ASAP7_75t_L g593 ( .A(n_286), .B(n_302), .Y(n_593) );
AND2x4_ASAP7_75t_L g606 ( .A(n_286), .B(n_363), .Y(n_606) );
AND2x4_ASAP7_75t_L g286 ( .A(n_287), .B(n_291), .Y(n_286) );
INVx2_ASAP7_75t_L g310 ( .A(n_287), .Y(n_310) );
AND2x2_ASAP7_75t_L g332 ( .A(n_287), .B(n_333), .Y(n_332) );
AND2x4_ASAP7_75t_L g351 ( .A(n_287), .B(n_352), .Y(n_351) );
OR2x2_ASAP7_75t_L g357 ( .A(n_287), .B(n_353), .Y(n_357) );
AND2x4_ASAP7_75t_L g287 ( .A(n_288), .B(n_290), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_289), .B(n_294), .Y(n_293) );
INVxp67_ASAP7_75t_L g318 ( .A(n_289), .Y(n_318) );
NAND3xp33_ASAP7_75t_L g344 ( .A(n_290), .B(n_317), .C(n_345), .Y(n_344) );
AND2x4_ASAP7_75t_L g309 ( .A(n_291), .B(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
INVx1_ASAP7_75t_L g353 ( .A(n_292), .Y(n_353) );
AND2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_295), .Y(n_292) );
INVx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx2_ASAP7_75t_L g560 ( .A(n_300), .Y(n_560) );
INVx2_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
BUFx6f_ASAP7_75t_L g399 ( .A(n_301), .Y(n_399) );
BUFx3_ASAP7_75t_L g546 ( .A(n_301), .Y(n_546) );
AND2x2_ASAP7_75t_L g328 ( .A(n_302), .B(n_309), .Y(n_328) );
AND2x2_ASAP7_75t_L g350 ( .A(n_302), .B(n_351), .Y(n_350) );
AND2x4_ASAP7_75t_L g355 ( .A(n_302), .B(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g520 ( .A(n_302), .B(n_351), .Y(n_520) );
AND2x2_ASAP7_75t_L g597 ( .A(n_302), .B(n_309), .Y(n_597) );
AND2x4_ASAP7_75t_L g604 ( .A(n_302), .B(n_351), .Y(n_604) );
AND2x4_ASAP7_75t_L g610 ( .A(n_302), .B(n_379), .Y(n_610) );
OAI22xp5_ASAP7_75t_L g303 ( .A1(n_304), .A2(n_305), .B1(n_311), .B2(n_312), .Y(n_303) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx3_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx2_ASAP7_75t_L g436 ( .A(n_307), .Y(n_436) );
INVx2_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx2_ASAP7_75t_L g467 ( .A(n_308), .Y(n_467) );
BUFx6f_ASAP7_75t_L g493 ( .A(n_308), .Y(n_493) );
BUFx6f_ASAP7_75t_L g540 ( .A(n_308), .Y(n_540) );
BUFx3_ASAP7_75t_L g563 ( .A(n_308), .Y(n_563) );
AND2x4_ASAP7_75t_L g315 ( .A(n_309), .B(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g368 ( .A(n_309), .B(n_363), .Y(n_368) );
AND2x4_ASAP7_75t_L g594 ( .A(n_309), .B(n_316), .Y(n_594) );
AND2x4_ASAP7_75t_L g607 ( .A(n_309), .B(n_363), .Y(n_607) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx3_ASAP7_75t_L g397 ( .A(n_314), .Y(n_397) );
INVx2_ASAP7_75t_L g507 ( .A(n_314), .Y(n_507) );
INVx3_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
BUFx6f_ASAP7_75t_L g468 ( .A(n_315), .Y(n_468) );
BUFx6f_ASAP7_75t_L g561 ( .A(n_315), .Y(n_561) );
AND2x4_ASAP7_75t_L g375 ( .A(n_316), .B(n_351), .Y(n_375) );
AND2x4_ASAP7_75t_L g381 ( .A(n_316), .B(n_379), .Y(n_381) );
AND2x4_ASAP7_75t_L g612 ( .A(n_316), .B(n_351), .Y(n_612) );
AND2x4_ASAP7_75t_L g613 ( .A(n_316), .B(n_379), .Y(n_613) );
AND2x2_ASAP7_75t_L g316 ( .A(n_317), .B(n_321), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
OAI21xp33_ASAP7_75t_L g323 ( .A1(n_324), .A2(n_325), .B(n_329), .Y(n_323) );
INVx2_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx3_ASAP7_75t_SL g626 ( .A(n_327), .Y(n_626) );
INVx3_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx2_ASAP7_75t_L g441 ( .A(n_328), .Y(n_441) );
BUFx3_ASAP7_75t_L g533 ( .A(n_328), .Y(n_533) );
INVx2_ASAP7_75t_SL g536 ( .A(n_330), .Y(n_536) );
BUFx4f_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
BUFx2_ASAP7_75t_L g400 ( .A(n_331), .Y(n_400) );
INVx5_ASAP7_75t_L g446 ( .A(n_331), .Y(n_446) );
AND2x4_ASAP7_75t_L g331 ( .A(n_332), .B(n_336), .Y(n_331) );
AND2x2_ASAP7_75t_L g591 ( .A(n_332), .B(n_336), .Y(n_591) );
AND2x4_ASAP7_75t_L g903 ( .A(n_332), .B(n_336), .Y(n_903) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
INVx1_ASAP7_75t_L g343 ( .A(n_334), .Y(n_343) );
INVx4_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
NOR2xp33_ASAP7_75t_L g669 ( .A(n_340), .B(n_670), .Y(n_669) );
INVx3_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx4_ASAP7_75t_L g600 ( .A(n_341), .Y(n_600) );
INVx3_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
BUFx6f_ASAP7_75t_L g392 ( .A(n_342), .Y(n_392) );
NOR2xp33_ASAP7_75t_L g346 ( .A(n_347), .B(n_369), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_348), .B(n_358), .Y(n_347) );
BUFx8_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
BUFx6f_ASAP7_75t_L g414 ( .A(n_350), .Y(n_414) );
AND2x4_ASAP7_75t_L g372 ( .A(n_351), .B(n_363), .Y(n_372) );
AND2x4_ASAP7_75t_L g609 ( .A(n_351), .B(n_363), .Y(n_609) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
BUFx3_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
BUFx6f_ASAP7_75t_L g403 ( .A(n_355), .Y(n_403) );
BUFx12f_ASAP7_75t_L g485 ( .A(n_355), .Y(n_485) );
BUFx6f_ASAP7_75t_L g575 ( .A(n_355), .Y(n_575) );
AND2x4_ASAP7_75t_L g590 ( .A(n_356), .B(n_363), .Y(n_590) );
INVx2_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx2_ASAP7_75t_L g379 ( .A(n_357), .Y(n_379) );
BUFx4f_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g410 ( .A(n_361), .Y(n_410) );
INVx1_ASAP7_75t_L g523 ( .A(n_361), .Y(n_523) );
INVx3_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
BUFx6f_ASAP7_75t_L g430 ( .A(n_362), .Y(n_430) );
BUFx12f_ASAP7_75t_L g500 ( .A(n_362), .Y(n_500) );
AND2x4_ASAP7_75t_L g378 ( .A(n_363), .B(n_379), .Y(n_378) );
BUFx6f_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g460 ( .A(n_366), .Y(n_460) );
INVx2_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
BUFx6f_ASAP7_75t_L g411 ( .A(n_368), .Y(n_411) );
BUFx5_ASAP7_75t_L g431 ( .A(n_368), .Y(n_431) );
BUFx3_ASAP7_75t_L g572 ( .A(n_368), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_370), .B(n_376), .Y(n_369) );
BUFx6f_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
BUFx12f_ASAP7_75t_L g407 ( .A(n_372), .Y(n_407) );
BUFx6f_ASAP7_75t_L g502 ( .A(n_372), .Y(n_502) );
INVx4_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx2_ASAP7_75t_L g413 ( .A(n_374), .Y(n_413) );
INVx1_ASAP7_75t_L g425 ( .A(n_374), .Y(n_425) );
INVx4_ASAP7_75t_L g462 ( .A(n_374), .Y(n_462) );
INVx2_ASAP7_75t_L g528 ( .A(n_374), .Y(n_528) );
INVx4_ASAP7_75t_L g573 ( .A(n_374), .Y(n_573) );
INVx8_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
BUFx6f_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
BUFx6f_ASAP7_75t_L g408 ( .A(n_378), .Y(n_408) );
BUFx6f_ASAP7_75t_L g516 ( .A(n_378), .Y(n_516) );
BUFx6f_ASAP7_75t_L g556 ( .A(n_378), .Y(n_556) );
BUFx3_ASAP7_75t_L g517 ( .A(n_380), .Y(n_517) );
BUFx12f_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx6_ASAP7_75t_L g405 ( .A(n_381), .Y(n_405) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g416 ( .A(n_383), .Y(n_416) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
XNOR2xp5_ASAP7_75t_L g385 ( .A(n_386), .B(n_388), .Y(n_385) );
CKINVDCx5p33_ASAP7_75t_R g386 ( .A(n_387), .Y(n_386) );
NOR2x1_ASAP7_75t_L g388 ( .A(n_389), .B(n_401), .Y(n_388) );
NAND4xp25_ASAP7_75t_L g389 ( .A(n_390), .B(n_393), .C(n_394), .D(n_398), .Y(n_389) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx2_ASAP7_75t_SL g449 ( .A(n_392), .Y(n_449) );
INVx2_ASAP7_75t_L g497 ( .A(n_392), .Y(n_497) );
BUFx6f_ASAP7_75t_L g569 ( .A(n_392), .Y(n_569) );
NOR2xp33_ASAP7_75t_L g934 ( .A(n_392), .B(n_935), .Y(n_934) );
INVx2_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx2_ASAP7_75t_L g470 ( .A(n_396), .Y(n_470) );
NAND4xp25_ASAP7_75t_L g401 ( .A(n_402), .B(n_406), .C(n_409), .D(n_412), .Y(n_401) );
INVx3_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx5_ASAP7_75t_L g487 ( .A(n_405), .Y(n_487) );
BUFx12f_ASAP7_75t_L g424 ( .A(n_407), .Y(n_424) );
BUFx6f_ASAP7_75t_L g526 ( .A(n_407), .Y(n_526) );
BUFx2_ASAP7_75t_SL g524 ( .A(n_411), .Y(n_524) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
AO22x2_ASAP7_75t_SL g418 ( .A1(n_419), .A2(n_420), .B1(n_450), .B2(n_451), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
NAND4xp75_ASAP7_75t_SL g421 ( .A(n_422), .B(n_427), .C(n_432), .D(n_437), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_423), .B(n_426), .Y(n_422) );
AND2x2_ASAP7_75t_L g427 ( .A(n_428), .B(n_429), .Y(n_427) );
AND2x2_ASAP7_75t_L g432 ( .A(n_433), .B(n_435), .Y(n_432) );
HB1xp67_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx2_ASAP7_75t_L g491 ( .A(n_440), .Y(n_491) );
INVx2_ASAP7_75t_L g651 ( .A(n_440), .Y(n_651) );
BUFx6f_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx2_ASAP7_75t_L g473 ( .A(n_441), .Y(n_473) );
OAI22xp5_ASAP7_75t_L g442 ( .A1(n_443), .A2(n_444), .B1(n_447), .B2(n_448), .Y(n_442) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx4_ASAP7_75t_L g475 ( .A(n_446), .Y(n_475) );
INVx2_ASAP7_75t_SL g448 ( .A(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
AO21x2_ASAP7_75t_L g451 ( .A1(n_452), .A2(n_453), .B(n_476), .Y(n_451) );
NOR3xp33_ASAP7_75t_SL g476 ( .A(n_452), .B(n_455), .C(n_464), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_454), .B(n_463), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
NAND4xp25_ASAP7_75t_SL g455 ( .A(n_456), .B(n_457), .C(n_458), .D(n_461), .Y(n_455) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
NAND4xp25_ASAP7_75t_L g464 ( .A(n_465), .B(n_469), .C(n_471), .D(n_474), .Y(n_464) );
INVx2_ASAP7_75t_SL g466 ( .A(n_467), .Y(n_466) );
BUFx3_ASAP7_75t_L g541 ( .A(n_468), .Y(n_541) );
BUFx3_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
XNOR2xp5_ASAP7_75t_L g478 ( .A(n_479), .B(n_508), .Y(n_478) );
XOR2xp5_ASAP7_75t_L g580 ( .A(n_479), .B(n_508), .Y(n_580) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
NAND4xp75_ASAP7_75t_L g482 ( .A(n_483), .B(n_488), .C(n_498), .D(n_503), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_484), .B(n_486), .Y(n_483) );
BUFx3_ASAP7_75t_L g521 ( .A(n_485), .Y(n_521) );
OA21x2_ASAP7_75t_L g488 ( .A1(n_489), .A2(n_490), .B(n_492), .Y(n_488) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_495), .B(n_496), .Y(n_494) );
INVx3_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
AND2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_501), .Y(n_498) );
AND2x2_ASAP7_75t_L g503 ( .A(n_504), .B(n_506), .Y(n_503) );
BUFx2_ASAP7_75t_L g543 ( .A(n_505), .Y(n_543) );
OA22x2_ASAP7_75t_L g508 ( .A1(n_509), .A2(n_548), .B1(n_549), .B2(n_579), .Y(n_508) );
INVx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
OR2x2_ASAP7_75t_L g511 ( .A(n_512), .B(n_529), .Y(n_511) );
NAND4xp25_ASAP7_75t_SL g512 ( .A(n_513), .B(n_518), .C(n_522), .D(n_525), .Y(n_512) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
BUFx6f_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
BUFx2_ASAP7_75t_SL g527 ( .A(n_528), .Y(n_527) );
NAND3xp33_ASAP7_75t_L g529 ( .A(n_530), .B(n_538), .C(n_542), .Y(n_529) );
HB1xp67_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
BUFx3_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
OAI21xp33_ASAP7_75t_L g534 ( .A1(n_535), .A2(n_536), .B(n_537), .Y(n_534) );
BUFx3_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
OAI22xp5_ASAP7_75t_L g709 ( .A1(n_547), .A2(n_710), .B1(n_713), .B2(n_714), .Y(n_709) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
AO21x2_ASAP7_75t_L g551 ( .A1(n_552), .A2(n_564), .B(n_576), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_554), .B(n_555), .Y(n_553) );
NAND2xp5_ASAP7_75t_SL g558 ( .A(n_559), .B(n_562), .Y(n_558) );
NOR2xp33_ASAP7_75t_L g564 ( .A(n_565), .B(n_570), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_566), .B(n_567), .Y(n_565) );
INVx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
NAND2x1_ASAP7_75t_SL g570 ( .A(n_571), .B(n_574), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_577), .B(n_578), .Y(n_576) );
XNOR2xp5_ASAP7_75t_L g582 ( .A(n_583), .B(n_635), .Y(n_582) );
OAI22xp5_ASAP7_75t_L g583 ( .A1(n_584), .A2(n_614), .B1(n_633), .B2(n_634), .Y(n_583) );
INVx2_ASAP7_75t_L g633 ( .A(n_584), .Y(n_633) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
NOR2x1_ASAP7_75t_L g587 ( .A(n_588), .B(n_601), .Y(n_587) );
NAND4xp25_ASAP7_75t_L g588 ( .A(n_589), .B(n_592), .C(n_595), .D(n_596), .Y(n_588) );
NOR2xp33_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
INVx4_ASAP7_75t_L g630 ( .A(n_600), .Y(n_630) );
NOR2xp33_ASAP7_75t_L g647 ( .A(n_600), .B(n_648), .Y(n_647) );
NOR2xp33_ASAP7_75t_L g906 ( .A(n_600), .B(n_907), .Y(n_906) );
NAND4xp25_ASAP7_75t_L g601 ( .A(n_602), .B(n_605), .C(n_608), .D(n_611), .Y(n_601) );
INVx1_ASAP7_75t_L g634 ( .A(n_614), .Y(n_634) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx2_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
XNOR2x1_ASAP7_75t_L g616 ( .A(n_617), .B(n_618), .Y(n_616) );
NOR2x1_ASAP7_75t_L g618 ( .A(n_619), .B(n_624), .Y(n_618) );
NAND4xp25_ASAP7_75t_L g619 ( .A(n_620), .B(n_621), .C(n_622), .D(n_623), .Y(n_619) );
NAND3xp33_ASAP7_75t_L g624 ( .A(n_625), .B(n_631), .C(n_632), .Y(n_624) );
NOR2xp33_ASAP7_75t_L g627 ( .A(n_628), .B(n_629), .Y(n_627) );
INVx2_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx2_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
XNOR2x1_ASAP7_75t_L g636 ( .A(n_637), .B(n_657), .Y(n_636) );
NAND4xp25_ASAP7_75t_L g654 ( .A(n_639), .B(n_640), .C(n_642), .D(n_650), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_641), .B(n_652), .Y(n_656) );
NAND3xp33_ASAP7_75t_L g643 ( .A(n_644), .B(n_650), .C(n_652), .Y(n_643) );
INVxp67_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
OR2x2_ASAP7_75t_L g655 ( .A(n_645), .B(n_656), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_646), .B(n_649), .Y(n_645) );
NOR2x1_ASAP7_75t_L g653 ( .A(n_654), .B(n_655), .Y(n_653) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
XOR2x2_ASAP7_75t_L g658 ( .A(n_659), .B(n_673), .Y(n_658) );
NOR2xp67_ASAP7_75t_L g659 ( .A(n_660), .B(n_665), .Y(n_659) );
NAND4xp25_ASAP7_75t_L g660 ( .A(n_661), .B(n_662), .C(n_663), .D(n_664), .Y(n_660) );
NAND4xp25_ASAP7_75t_L g665 ( .A(n_666), .B(n_667), .C(n_668), .D(n_671), .Y(n_665) );
OAI221xp5_ASAP7_75t_L g674 ( .A1(n_675), .A2(n_892), .B1(n_894), .B2(n_914), .C(n_919), .Y(n_674) );
NOR3xp33_ASAP7_75t_L g675 ( .A(n_676), .B(n_797), .C(n_857), .Y(n_675) );
AOI31xp33_ASAP7_75t_L g676 ( .A1(n_677), .A2(n_765), .A3(n_783), .B(n_791), .Y(n_676) );
AOI211xp5_ASAP7_75t_L g677 ( .A1(n_678), .A2(n_697), .B(n_748), .C(n_756), .Y(n_677) );
INVx3_ASAP7_75t_L g872 ( .A(n_678), .Y(n_872) );
INVx3_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g808 ( .A(n_679), .B(n_809), .Y(n_808) );
AOI221xp5_ASAP7_75t_L g817 ( .A1(n_679), .A2(n_818), .B1(n_821), .B2(n_823), .C(n_825), .Y(n_817) );
NAND2xp5_ASAP7_75t_L g834 ( .A(n_679), .B(n_750), .Y(n_834) );
INVx3_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_680), .B(n_737), .Y(n_803) );
INVx2_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
NOR3xp33_ASAP7_75t_L g804 ( .A(n_681), .B(n_728), .C(n_805), .Y(n_804) );
NAND2xp5_ASAP7_75t_L g838 ( .A(n_681), .B(n_700), .Y(n_838) );
INVx3_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_682), .B(n_700), .Y(n_785) );
NAND2xp5_ASAP7_75t_L g822 ( .A(n_682), .B(n_775), .Y(n_822) );
OR2x2_ASAP7_75t_L g855 ( .A(n_682), .B(n_700), .Y(n_855) );
AND2x2_ASAP7_75t_L g859 ( .A(n_682), .B(n_819), .Y(n_859) );
AND2x2_ASAP7_75t_L g865 ( .A(n_682), .B(n_701), .Y(n_865) );
INVx1_ASAP7_75t_L g877 ( .A(n_682), .Y(n_877) );
NOR2xp33_ASAP7_75t_L g891 ( .A(n_682), .B(n_827), .Y(n_891) );
AND2x4_ASAP7_75t_L g682 ( .A(n_683), .B(n_690), .Y(n_682) );
AND2x2_ASAP7_75t_L g684 ( .A(n_685), .B(n_687), .Y(n_684) );
AND2x4_ASAP7_75t_L g691 ( .A(n_685), .B(n_692), .Y(n_691) );
AND2x4_ASAP7_75t_L g703 ( .A(n_685), .B(n_687), .Y(n_703) );
AND2x2_ASAP7_75t_L g721 ( .A(n_685), .B(n_687), .Y(n_721) );
AND2x4_ASAP7_75t_L g688 ( .A(n_687), .B(n_689), .Y(n_688) );
AND2x2_ASAP7_75t_L g704 ( .A(n_687), .B(n_689), .Y(n_704) );
AND2x2_ASAP7_75t_L g718 ( .A(n_687), .B(n_689), .Y(n_718) );
CKINVDCx5p33_ASAP7_75t_R g940 ( .A(n_687), .Y(n_940) );
INVx2_ASAP7_75t_L g747 ( .A(n_688), .Y(n_747) );
BUFx2_ASAP7_75t_L g893 ( .A(n_688), .Y(n_893) );
AND2x4_ASAP7_75t_L g696 ( .A(n_689), .B(n_692), .Y(n_696) );
AND2x4_ASAP7_75t_L g706 ( .A(n_689), .B(n_692), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_689), .B(n_692), .Y(n_714) );
INVx3_ASAP7_75t_L g740 ( .A(n_691), .Y(n_740) );
INVx2_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx2_ASAP7_75t_SL g695 ( .A(n_696), .Y(n_695) );
OAI22xp33_ASAP7_75t_L g697 ( .A1(n_698), .A2(n_722), .B1(n_733), .B2(n_735), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_699), .B(n_707), .Y(n_698) );
OAI211xp5_ASAP7_75t_SL g825 ( .A1(n_699), .A2(n_826), .B(n_830), .C(n_843), .Y(n_825) );
INVx3_ASAP7_75t_L g841 ( .A(n_699), .Y(n_841) );
INVx3_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
AND2x2_ASAP7_75t_L g809 ( .A(n_700), .B(n_738), .Y(n_809) );
INVx2_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
AND2x2_ASAP7_75t_L g736 ( .A(n_701), .B(n_737), .Y(n_736) );
AND2x2_ASAP7_75t_L g775 ( .A(n_701), .B(n_738), .Y(n_775) );
OR2x2_ASAP7_75t_L g782 ( .A(n_701), .B(n_738), .Y(n_782) );
AND2x2_ASAP7_75t_L g701 ( .A(n_702), .B(n_705), .Y(n_701) );
INVx3_ASAP7_75t_L g745 ( .A(n_703), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_707), .B(n_736), .Y(n_735) );
NOR2xp33_ASAP7_75t_L g750 ( .A(n_707), .B(n_737), .Y(n_750) );
AND2x2_ASAP7_75t_L g772 ( .A(n_707), .B(n_773), .Y(n_772) );
NOR2xp33_ASAP7_75t_L g781 ( .A(n_707), .B(n_782), .Y(n_781) );
NOR2xp33_ASAP7_75t_L g788 ( .A(n_707), .B(n_789), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g805 ( .A(n_707), .B(n_775), .Y(n_805) );
AND2x2_ASAP7_75t_L g814 ( .A(n_707), .B(n_764), .Y(n_814) );
A2O1A1Ixp33_ASAP7_75t_L g843 ( .A1(n_707), .A2(n_727), .B(n_819), .C(n_844), .Y(n_843) );
INVx1_ASAP7_75t_L g851 ( .A(n_707), .Y(n_851) );
CKINVDCx6p67_ASAP7_75t_R g707 ( .A(n_708), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_708), .B(n_764), .Y(n_763) );
AND2x2_ASAP7_75t_L g801 ( .A(n_708), .B(n_761), .Y(n_801) );
INVx1_ASAP7_75t_L g828 ( .A(n_708), .Y(n_828) );
NOR2xp33_ASAP7_75t_L g831 ( .A(n_708), .B(n_832), .Y(n_831) );
NOR2xp33_ASAP7_75t_L g840 ( .A(n_708), .B(n_737), .Y(n_840) );
AND2x2_ASAP7_75t_L g848 ( .A(n_708), .B(n_771), .Y(n_848) );
AOI22xp33_ASAP7_75t_L g849 ( .A1(n_708), .A2(n_751), .B1(n_850), .B2(n_852), .Y(n_849) );
OR2x6_ASAP7_75t_SL g708 ( .A(n_709), .B(n_715), .Y(n_708) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
OAI22xp5_ASAP7_75t_L g739 ( .A1(n_714), .A2(n_740), .B1(n_741), .B2(n_742), .Y(n_739) );
OAI221xp5_ASAP7_75t_L g793 ( .A1(n_714), .A2(n_740), .B1(n_794), .B2(n_795), .C(n_796), .Y(n_793) );
OAI22xp5_ASAP7_75t_L g715 ( .A1(n_716), .A2(n_717), .B1(n_719), .B2(n_720), .Y(n_715) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
OR2x2_ASAP7_75t_L g722 ( .A(n_723), .B(n_731), .Y(n_722) );
AND2x2_ASAP7_75t_L g752 ( .A(n_723), .B(n_753), .Y(n_752) );
AND2x2_ASAP7_75t_L g813 ( .A(n_723), .B(n_814), .Y(n_813) );
AND2x2_ASAP7_75t_SL g844 ( .A(n_723), .B(n_764), .Y(n_844) );
AND2x2_ASAP7_75t_L g723 ( .A(n_724), .B(n_727), .Y(n_723) );
INVx1_ASAP7_75t_L g732 ( .A(n_724), .Y(n_732) );
AND2x2_ASAP7_75t_L g761 ( .A(n_724), .B(n_728), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_725), .B(n_726), .Y(n_724) );
AND2x2_ASAP7_75t_L g771 ( .A(n_727), .B(n_732), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_727), .B(n_773), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g820 ( .A(n_727), .B(n_772), .Y(n_820) );
CKINVDCx5p33_ASAP7_75t_R g727 ( .A(n_728), .Y(n_727) );
AND2x2_ASAP7_75t_L g731 ( .A(n_728), .B(n_732), .Y(n_731) );
OR2x2_ASAP7_75t_L g824 ( .A(n_728), .B(n_753), .Y(n_824) );
AND2x4_ASAP7_75t_SL g728 ( .A(n_729), .B(n_730), .Y(n_728) );
AND2x2_ASAP7_75t_L g778 ( .A(n_731), .B(n_764), .Y(n_778) );
INVx1_ASAP7_75t_L g832 ( .A(n_731), .Y(n_832) );
AND2x2_ASAP7_75t_L g853 ( .A(n_731), .B(n_753), .Y(n_853) );
INVx1_ASAP7_75t_L g734 ( .A(n_732), .Y(n_734) );
AND2x2_ASAP7_75t_L g829 ( .A(n_732), .B(n_773), .Y(n_829) );
AND2x2_ASAP7_75t_L g835 ( .A(n_732), .B(n_764), .Y(n_835) );
NOR2xp33_ASAP7_75t_L g889 ( .A(n_732), .B(n_773), .Y(n_889) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
OAI211xp5_ASAP7_75t_L g875 ( .A1(n_736), .A2(n_856), .B(n_876), .C(n_878), .Y(n_875) );
INVx3_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx2_ASAP7_75t_L g759 ( .A(n_738), .Y(n_759) );
OR2x2_ASAP7_75t_L g738 ( .A(n_739), .B(n_743), .Y(n_738) );
OAI22xp5_ASAP7_75t_L g743 ( .A1(n_744), .A2(n_745), .B1(n_746), .B2(n_747), .Y(n_743) );
NOR2xp33_ASAP7_75t_L g748 ( .A(n_749), .B(n_751), .Y(n_748) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
AOI22xp5_ASAP7_75t_L g783 ( .A1(n_752), .A2(n_784), .B1(n_786), .B2(n_790), .Y(n_783) );
CKINVDCx6p67_ASAP7_75t_R g764 ( .A(n_753), .Y(n_764) );
INVx1_ASAP7_75t_L g774 ( .A(n_753), .Y(n_774) );
AND2x2_ASAP7_75t_L g862 ( .A(n_753), .B(n_801), .Y(n_862) );
AND2x2_ASAP7_75t_L g753 ( .A(n_754), .B(n_755), .Y(n_753) );
INVxp67_ASAP7_75t_SL g756 ( .A(n_757), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_758), .B(n_760), .Y(n_757) );
AND2x2_ASAP7_75t_L g790 ( .A(n_758), .B(n_784), .Y(n_790) );
OAI22xp5_ASAP7_75t_L g818 ( .A1(n_758), .A2(n_777), .B1(n_819), .B2(n_820), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g868 ( .A(n_758), .B(n_869), .Y(n_868) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
BUFx2_ASAP7_75t_L g812 ( .A(n_759), .Y(n_812) );
NOR2xp33_ASAP7_75t_L g876 ( .A(n_759), .B(n_877), .Y(n_876) );
O2A1O1Ixp33_ASAP7_75t_L g882 ( .A1(n_760), .A2(n_775), .B(n_869), .C(n_883), .Y(n_882) );
AND2x2_ASAP7_75t_L g760 ( .A(n_761), .B(n_762), .Y(n_760) );
INVx1_ASAP7_75t_L g769 ( .A(n_761), .Y(n_769) );
NAND3xp33_ASAP7_75t_L g839 ( .A(n_761), .B(n_840), .C(n_841), .Y(n_839) );
AND2x2_ASAP7_75t_L g869 ( .A(n_761), .B(n_772), .Y(n_869) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
NOR2xp33_ASAP7_75t_L g768 ( .A(n_764), .B(n_769), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_764), .B(n_771), .Y(n_800) );
NAND2xp5_ASAP7_75t_L g847 ( .A(n_764), .B(n_848), .Y(n_847) );
AOI21xp33_ASAP7_75t_L g765 ( .A1(n_766), .A2(n_775), .B(n_776), .Y(n_765) );
INVxp67_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
NOR2xp33_ASAP7_75t_L g767 ( .A(n_768), .B(n_770), .Y(n_767) );
INVx1_ASAP7_75t_L g779 ( .A(n_768), .Y(n_779) );
AOI21xp33_ASAP7_75t_SL g887 ( .A1(n_769), .A2(n_888), .B(n_890), .Y(n_887) );
AND2x2_ASAP7_75t_L g770 ( .A(n_771), .B(n_772), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g816 ( .A(n_771), .B(n_814), .Y(n_816) );
AOI211xp5_ASAP7_75t_L g806 ( .A1(n_773), .A2(n_807), .B(n_810), .C(n_815), .Y(n_806) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
AOI221xp5_ASAP7_75t_L g830 ( .A1(n_775), .A2(n_831), .B1(n_833), .B2(n_835), .C(n_836), .Y(n_830) );
AOI21xp33_ASAP7_75t_L g776 ( .A1(n_777), .A2(n_779), .B(n_780), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_777), .B(n_787), .Y(n_786) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
INVx1_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
INVx1_ASAP7_75t_L g819 ( .A(n_782), .Y(n_819) );
INVx1_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
A2O1A1Ixp33_ASAP7_75t_L g873 ( .A1(n_787), .A2(n_852), .B(n_874), .C(n_875), .Y(n_873) );
INVx1_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
INVx1_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
BUFx3_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
INVx2_ASAP7_75t_L g842 ( .A(n_793), .Y(n_842) );
AOI32xp33_ASAP7_75t_L g797 ( .A1(n_798), .A2(n_806), .A3(n_817), .B1(n_845), .B2(n_856), .Y(n_797) );
O2A1O1Ixp33_ASAP7_75t_L g798 ( .A1(n_799), .A2(n_801), .B(n_802), .C(n_804), .Y(n_798) );
INVx1_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
NOR2xp33_ASAP7_75t_L g883 ( .A(n_800), .B(n_822), .Y(n_883) );
OAI21xp5_ASAP7_75t_L g880 ( .A1(n_801), .A2(n_859), .B(n_881), .Y(n_880) );
INVx1_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
AOI221xp5_ASAP7_75t_SL g884 ( .A1(n_807), .A2(n_829), .B1(n_885), .B2(n_886), .C(n_887), .Y(n_884) );
INVx1_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
INVx1_ASAP7_75t_L g874 ( .A(n_809), .Y(n_874) );
AND2x2_ASAP7_75t_L g810 ( .A(n_811), .B(n_813), .Y(n_810) );
NOR2xp33_ASAP7_75t_L g815 ( .A(n_811), .B(n_816), .Y(n_815) );
INVx2_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
A2O1A1Ixp33_ASAP7_75t_SL g845 ( .A1(n_812), .A2(n_846), .B(n_849), .C(n_854), .Y(n_845) );
INVx1_ASAP7_75t_L g870 ( .A(n_816), .Y(n_870) );
NAND2xp5_ASAP7_75t_L g890 ( .A(n_819), .B(n_891), .Y(n_890) );
INVx1_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
INVx1_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
AOI31xp33_ASAP7_75t_L g860 ( .A1(n_824), .A2(n_861), .A3(n_863), .B(n_864), .Y(n_860) );
AOI21xp5_ASAP7_75t_L g881 ( .A1(n_824), .A2(n_861), .B(n_864), .Y(n_881) );
INVx1_ASAP7_75t_L g885 ( .A(n_826), .Y(n_885) );
NAND2xp5_ASAP7_75t_L g826 ( .A(n_827), .B(n_829), .Y(n_826) );
NAND2xp5_ASAP7_75t_L g879 ( .A(n_827), .B(n_853), .Y(n_879) );
INVx3_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
INVx1_ASAP7_75t_L g837 ( .A(n_829), .Y(n_837) );
INVxp67_ASAP7_75t_SL g833 ( .A(n_834), .Y(n_833) );
A2O1A1Ixp33_ASAP7_75t_L g858 ( .A1(n_835), .A2(n_850), .B(n_859), .C(n_860), .Y(n_858) );
OAI211xp5_ASAP7_75t_L g836 ( .A1(n_837), .A2(n_838), .B(n_839), .C(n_842), .Y(n_836) );
INVx1_ASAP7_75t_L g886 ( .A(n_838), .Y(n_886) );
CKINVDCx16_ASAP7_75t_R g856 ( .A(n_842), .Y(n_856) );
INVx1_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
CKINVDCx14_ASAP7_75t_R g850 ( .A(n_851), .Y(n_850) );
INVx1_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
INVx1_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
NAND5xp2_ASAP7_75t_L g857 ( .A(n_858), .B(n_866), .C(n_880), .D(n_882), .E(n_884), .Y(n_857) );
INVx1_ASAP7_75t_L g863 ( .A(n_859), .Y(n_863) );
INVx1_ASAP7_75t_L g861 ( .A(n_862), .Y(n_861) );
INVx1_ASAP7_75t_L g864 ( .A(n_865), .Y(n_864) );
O2A1O1Ixp33_ASAP7_75t_L g866 ( .A1(n_867), .A2(n_870), .B(n_871), .C(n_873), .Y(n_866) );
INVx1_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
INVx1_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
INVx1_ASAP7_75t_L g878 ( .A(n_879), .Y(n_878) );
INVx1_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
CKINVDCx5p33_ASAP7_75t_R g892 ( .A(n_893), .Y(n_892) );
INVx2_ASAP7_75t_L g894 ( .A(n_895), .Y(n_894) );
BUFx2_ASAP7_75t_SL g895 ( .A(n_896), .Y(n_895) );
INVx2_ASAP7_75t_L g896 ( .A(n_897), .Y(n_896) );
BUFx3_ASAP7_75t_L g897 ( .A(n_898), .Y(n_897) );
NAND2xp5_ASAP7_75t_L g899 ( .A(n_900), .B(n_908), .Y(n_899) );
AND4x1_ASAP7_75t_L g900 ( .A(n_901), .B(n_902), .C(n_904), .D(n_905), .Y(n_900) );
NOR4xp25_ASAP7_75t_L g908 ( .A(n_909), .B(n_911), .C(n_912), .D(n_913), .Y(n_908) );
INVx1_ASAP7_75t_L g909 ( .A(n_910), .Y(n_909) );
INVx1_ASAP7_75t_L g914 ( .A(n_915), .Y(n_914) );
HB1xp67_ASAP7_75t_L g915 ( .A(n_916), .Y(n_915) );
BUFx2_ASAP7_75t_SL g920 ( .A(n_921), .Y(n_920) );
INVx1_ASAP7_75t_L g924 ( .A(n_925), .Y(n_924) );
HB1xp67_ASAP7_75t_L g925 ( .A(n_926), .Y(n_925) );
INVx1_ASAP7_75t_L g926 ( .A(n_927), .Y(n_926) );
NAND3xp33_ASAP7_75t_L g927 ( .A(n_928), .B(n_933), .C(n_936), .Y(n_927) );
AND4x1_ASAP7_75t_L g928 ( .A(n_929), .B(n_930), .C(n_931), .D(n_932), .Y(n_928) );
BUFx2_ASAP7_75t_L g938 ( .A(n_939), .Y(n_938) );
endmodule