module fake_jpeg_29842_n_107 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_107);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_107;

wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx5p33_ASAP7_75t_R g35 ( 
.A(n_31),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_18),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_27),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_11),
.Y(n_42)
);

BUFx3_ASAP7_75t_SL g43 ( 
.A(n_23),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_25),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_37),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_50),
.B(n_51),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_52),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_41),
.B(n_0),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_35),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_49),
.A2(n_39),
.B1(n_43),
.B2(n_40),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_59),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_51),
.A2(n_44),
.B1(n_42),
.B2(n_45),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_60),
.B(n_64),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_47),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_63),
.B(n_4),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

MAJx2_ASAP7_75t_L g65 ( 
.A(n_48),
.B(n_40),
.C(n_14),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_65),
.A2(n_1),
.B(n_3),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_64),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_66),
.B(n_72),
.Y(n_90)
);

A2O1A1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_55),
.A2(n_40),
.B(n_2),
.C(n_3),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_68),
.Y(n_81)
);

O2A1O1Ixp33_ASAP7_75t_SL g69 ( 
.A1(n_65),
.A2(n_52),
.B(n_46),
.C(n_19),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_69),
.A2(n_75),
.B1(n_76),
.B2(n_79),
.Y(n_85)
);

NAND3xp33_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_16),
.C(n_33),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_61),
.A2(n_4),
.B(n_5),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_73),
.B(n_77),
.C(n_66),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_58),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_74),
.Y(n_82)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_57),
.B(n_5),
.Y(n_77)
);

OR2x2_ASAP7_75t_SL g84 ( 
.A(n_77),
.B(n_78),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_57),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_57),
.B(n_6),
.Y(n_80)
);

OAI32xp33_ASAP7_75t_L g87 ( 
.A1(n_80),
.A2(n_9),
.A3(n_12),
.B1(n_13),
.B2(n_20),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_71),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_83),
.B(n_86),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_69),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_87),
.B(n_89),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_67),
.A2(n_22),
.B1(n_24),
.B2(n_26),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_88),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_70),
.A2(n_28),
.B1(n_32),
.B2(n_34),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_91),
.B(n_72),
.C(n_81),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_93),
.B(n_95),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_91),
.B(n_81),
.C(n_84),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_94),
.A2(n_85),
.B(n_90),
.Y(n_97)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_97),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_96),
.Y(n_99)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_99),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_101),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_102),
.B(n_82),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_100),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g105 ( 
.A(n_104),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_105),
.A2(n_98),
.B(n_84),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_92),
.Y(n_107)
);


endmodule