module fake_jpeg_4977_n_190 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_190);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_190;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

INVx8_ASAP7_75t_SL g16 ( 
.A(n_5),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx8_ASAP7_75t_SL g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx9p33_ASAP7_75t_R g31 ( 
.A(n_16),
.Y(n_31)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_28),
.B(n_0),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_32),
.B(n_28),
.Y(n_55)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_35),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_0),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_37),
.Y(n_43)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_39),
.Y(n_47)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_53),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_36),
.A2(n_23),
.B1(n_24),
.B2(n_17),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_46),
.A2(n_50),
.B1(n_54),
.B2(n_38),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_32),
.B(n_30),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_48),
.B(n_52),
.Y(n_68)
);

NAND2x1_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_24),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_49),
.A2(n_33),
.B(n_37),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_36),
.A2(n_23),
.B1(n_24),
.B2(n_17),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_40),
.A2(n_23),
.B1(n_17),
.B2(n_25),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_51),
.A2(n_38),
.B1(n_37),
.B2(n_19),
.Y(n_73)
);

NAND2xp67_ASAP7_75t_SL g52 ( 
.A(n_32),
.B(n_28),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_36),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_43),
.Y(n_69)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_30),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_40),
.A2(n_27),
.B1(n_26),
.B2(n_22),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_58),
.A2(n_40),
.B1(n_22),
.B2(n_56),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_59),
.B(n_63),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_60),
.A2(n_62),
.B(n_50),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_49),
.A2(n_40),
.B1(n_38),
.B2(n_34),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_61),
.A2(n_64),
.B1(n_73),
.B2(n_58),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_49),
.A2(n_38),
.B1(n_34),
.B2(n_39),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_66),
.B(n_70),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_67),
.B(n_72),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_74),
.Y(n_79)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_35),
.Y(n_71)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_48),
.B(n_28),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_74),
.B(n_41),
.Y(n_76)
);

A2O1A1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_68),
.A2(n_52),
.B(n_41),
.C(n_43),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_75),
.B(n_85),
.Y(n_107)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_76),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_72),
.A2(n_51),
.B1(n_57),
.B2(n_53),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_77),
.A2(n_88),
.B1(n_89),
.B2(n_45),
.Y(n_101)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_82),
.Y(n_93)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_79),
.Y(n_104)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

AND2x2_ASAP7_75t_SL g83 ( 
.A(n_60),
.B(n_34),
.Y(n_83)
);

A2O1A1O1Ixp25_ASAP7_75t_L g95 ( 
.A1(n_83),
.A2(n_64),
.B(n_73),
.C(n_39),
.D(n_28),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_84),
.A2(n_19),
.B1(n_21),
.B2(n_29),
.Y(n_103)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_69),
.A2(n_57),
.B1(n_47),
.B2(n_42),
.Y(n_88)
);

OA22x2_ASAP7_75t_L g89 ( 
.A1(n_61),
.A2(n_45),
.B1(n_57),
.B2(n_47),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_90),
.A2(n_73),
.B1(n_45),
.B2(n_39),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_71),
.B(n_42),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_92),
.B(n_66),
.Y(n_109)
);

AOI32xp33_ASAP7_75t_L g94 ( 
.A1(n_83),
.A2(n_60),
.A3(n_68),
.B1(n_67),
.B2(n_62),
.Y(n_94)
);

NAND3xp33_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_89),
.C(n_79),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_SL g112 ( 
.A(n_95),
.B(n_77),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_91),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_97),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_101),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_29),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_100),
.B(n_103),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_83),
.A2(n_19),
.B(n_21),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_102),
.A2(n_92),
.B(n_89),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_105),
.B(n_109),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_89),
.A2(n_29),
.B1(n_21),
.B2(n_15),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_106),
.A2(n_89),
.B(n_86),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_76),
.C(n_88),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_108),
.B(n_104),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_112),
.B(n_114),
.C(n_102),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_113),
.B(n_124),
.Y(n_133)
);

XOR2x2_ASAP7_75t_L g128 ( 
.A(n_115),
.B(n_100),
.Y(n_128)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_93),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_119),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_118),
.A2(n_126),
.B(n_85),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_97),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_108),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_120),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_96),
.B(n_82),
.Y(n_121)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_121),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_96),
.B(n_78),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_122),
.B(n_123),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_107),
.B(n_80),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_80),
.Y(n_124)
);

AOI21xp33_ASAP7_75t_L g126 ( 
.A1(n_104),
.A2(n_79),
.B(n_75),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_127),
.B(n_129),
.C(n_139),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_128),
.A2(n_132),
.B(n_135),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_120),
.B(n_114),
.C(n_112),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_117),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_130),
.B(n_87),
.Y(n_145)
);

FAx1_ASAP7_75t_L g132 ( 
.A(n_113),
.B(n_105),
.CI(n_95),
.CON(n_132),
.SN(n_132)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_111),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_138),
.B(n_98),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_99),
.C(n_106),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_125),
.B(n_90),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_140),
.B(n_141),
.C(n_15),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_125),
.B(n_81),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_136),
.A2(n_119),
.B1(n_111),
.B2(n_116),
.Y(n_143)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_143),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_139),
.A2(n_110),
.B1(n_126),
.B2(n_98),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_144),
.A2(n_133),
.B1(n_132),
.B2(n_140),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_145),
.B(n_146),
.Y(n_154)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_134),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_147),
.B(n_148),
.Y(n_160)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_137),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_149),
.B(n_132),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_135),
.B(n_1),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_150),
.A2(n_153),
.B(n_131),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g151 ( 
.A(n_130),
.Y(n_151)
);

HB1xp67_ASAP7_75t_L g158 ( 
.A(n_151),
.Y(n_158)
);

HB1xp67_ASAP7_75t_L g153 ( 
.A(n_128),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_149),
.B(n_129),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_155),
.B(n_150),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_142),
.B(n_127),
.C(n_141),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_156),
.B(n_159),
.C(n_162),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_157),
.A2(n_14),
.B1(n_13),
.B2(n_4),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_161),
.A2(n_1),
.B(n_2),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_142),
.B(n_15),
.C(n_66),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_163),
.A2(n_152),
.B1(n_144),
.B2(n_157),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_164),
.A2(n_169),
.B1(n_171),
.B2(n_165),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_159),
.B(n_152),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_165),
.B(n_166),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_167),
.B(n_168),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_158),
.B(n_154),
.Y(n_168)
);

INVx11_ASAP7_75t_L g169 ( 
.A(n_160),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_169),
.B(n_156),
.Y(n_177)
);

OAI221xp5_ASAP7_75t_L g174 ( 
.A1(n_170),
.A2(n_14),
.B1(n_13),
.B2(n_4),
.C(n_5),
.Y(n_174)
);

OAI21x1_ASAP7_75t_L g172 ( 
.A1(n_166),
.A2(n_162),
.B(n_155),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_172),
.A2(n_174),
.B(n_175),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_177),
.B(n_1),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_175),
.A2(n_171),
.B1(n_164),
.B2(n_4),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_178),
.B(n_181),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_179),
.A2(n_182),
.B(n_7),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_176),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_173),
.A2(n_3),
.B(n_6),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_180),
.B(n_7),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_184),
.B(n_185),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_183),
.A2(n_7),
.B(n_9),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_187),
.B(n_9),
.C(n_10),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_188),
.A2(n_186),
.B(n_66),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_189),
.B(n_11),
.Y(n_190)
);


endmodule