module fake_jpeg_4001_n_141 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_141);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_141;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_4),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

HB1xp67_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_32),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_1),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_16),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_22),
.B(n_1),
.Y(n_35)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_36),
.A2(n_15),
.B1(n_21),
.B2(n_20),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_2),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_37),
.B(n_25),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_38),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_36),
.A2(n_26),
.B1(n_14),
.B2(n_25),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_40),
.A2(n_23),
.B1(n_19),
.B2(n_17),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_42),
.B(n_44),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_46),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_13),
.C(n_14),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_SL g56 ( 
.A1(n_48),
.A2(n_13),
.B(n_15),
.Y(n_56)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

BUFx2_ASAP7_75t_SL g54 ( 
.A(n_50),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_21),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_51),
.B(n_55),
.Y(n_78)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_52),
.B(n_56),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_53),
.B(n_61),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_20),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_16),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_57),
.B(n_60),
.Y(n_84)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_58),
.Y(n_83)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_47),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_62),
.A2(n_65),
.B1(n_67),
.B2(n_50),
.Y(n_76)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_39),
.Y(n_63)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_41),
.B(n_47),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_66),
.B(n_71),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_49),
.A2(n_23),
.B1(n_19),
.B2(n_5),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_47),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_68),
.B(n_72),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_24),
.Y(n_70)
);

NOR3xp33_ASAP7_75t_L g87 ( 
.A(n_70),
.B(n_8),
.C(n_10),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_34),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_48),
.Y(n_72)
);

OAI32xp33_ASAP7_75t_L g75 ( 
.A1(n_52),
.A2(n_38),
.A3(n_23),
.B1(n_30),
.B2(n_28),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_75),
.B(n_51),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_76),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_69),
.B(n_49),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_79),
.Y(n_89)
);

NOR3xp33_ASAP7_75t_SL g79 ( 
.A(n_70),
.B(n_49),
.C(n_29),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_87),
.B(n_9),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_72),
.A2(n_39),
.B1(n_28),
.B2(n_17),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_88),
.A2(n_80),
.B(n_57),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_90),
.B(n_78),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_85),
.B(n_60),
.Y(n_91)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_92),
.B(n_93),
.Y(n_105)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_84),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_75),
.B(n_54),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_94),
.A2(n_100),
.B(n_79),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_81),
.A2(n_62),
.B1(n_69),
.B2(n_56),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_95),
.B(n_101),
.Y(n_107)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_84),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_98),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_78),
.B(n_55),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_85),
.B(n_66),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_99),
.B(n_82),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_73),
.A2(n_71),
.B(n_68),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_88),
.B(n_54),
.C(n_34),
.Y(n_101)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_103),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_104),
.A2(n_108),
.B(n_112),
.Y(n_119)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_98),
.Y(n_110)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_110),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_99),
.B(n_34),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_111),
.B(n_112),
.Y(n_114)
);

AOI322xp5_ASAP7_75t_SL g113 ( 
.A1(n_104),
.A2(n_100),
.A3(n_93),
.B1(n_96),
.B2(n_95),
.C1(n_89),
.C2(n_92),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_SL g123 ( 
.A(n_113),
.B(n_119),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g116 ( 
.A(n_108),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g125 ( 
.A(n_116),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_105),
.A2(n_102),
.B1(n_97),
.B2(n_101),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_118),
.B(n_107),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_109),
.A2(n_94),
.B1(n_64),
.B2(n_82),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_120),
.B(n_94),
.C(n_111),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_113),
.A2(n_106),
.B(n_107),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_121),
.A2(n_86),
.B(n_74),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_122),
.B(n_29),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_124),
.B(n_126),
.C(n_86),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_114),
.B(n_117),
.C(n_115),
.Y(n_126)
);

A2O1A1Ixp33_ASAP7_75t_L g127 ( 
.A1(n_123),
.A2(n_116),
.B(n_83),
.C(n_7),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_127),
.B(n_10),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_128),
.B(n_131),
.C(n_29),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_129),
.A2(n_130),
.B(n_59),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_125),
.B(n_74),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_132),
.B(n_133),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_130),
.A2(n_58),
.B1(n_63),
.B2(n_12),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_134),
.A2(n_135),
.B1(n_63),
.B2(n_4),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_137),
.B(n_3),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_138),
.A2(n_136),
.B(n_137),
.Y(n_139)
);

MAJx2_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_6),
.C(n_24),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_6),
.Y(n_141)
);


endmodule