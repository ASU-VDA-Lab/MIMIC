module fake_jpeg_3629_n_232 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_232);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_232;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_11),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_35),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

BUFx8_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_6),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_5),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_37),
.Y(n_66)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_14),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_12),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_14),
.Y(n_69)
);

BUFx16f_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_24),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

BUFx10_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_10),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_32),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_18),
.B(n_9),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_11),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_48),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_79),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_70),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_78),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_0),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_81),
.B(n_85),
.Y(n_89)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_82),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_84),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_76),
.B(n_19),
.Y(n_85)
);

BUFx24_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_86),
.Y(n_94)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_84),
.Y(n_90)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_79),
.A2(n_69),
.B1(n_74),
.B2(n_75),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_91),
.A2(n_69),
.B1(n_74),
.B2(n_75),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_93),
.B(n_59),
.Y(n_101)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_95),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_83),
.A2(n_62),
.B1(n_67),
.B2(n_55),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_96),
.A2(n_86),
.B1(n_67),
.B2(n_55),
.Y(n_111)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_97),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_85),
.B(n_77),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_66),
.Y(n_117)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_86),
.Y(n_100)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_100),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_101),
.B(n_102),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_89),
.B(n_53),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_92),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_105),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_88),
.B(n_80),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_106),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_88),
.B(n_53),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_107),
.B(n_115),
.Y(n_129)
);

INVx4_ASAP7_75t_SL g108 ( 
.A(n_87),
.Y(n_108)
);

INVx4_ASAP7_75t_SL g128 ( 
.A(n_108),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_90),
.B(n_65),
.C(n_70),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_109),
.B(n_113),
.C(n_86),
.Y(n_126)
);

BUFx2_ASAP7_75t_SL g110 ( 
.A(n_97),
.Y(n_110)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_110),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_111),
.A2(n_118),
.B1(n_62),
.B2(n_98),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_92),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_112),
.B(n_117),
.Y(n_122)
);

MAJx2_ASAP7_75t_L g113 ( 
.A(n_87),
.B(n_70),
.C(n_58),
.Y(n_113)
);

INVx11_ASAP7_75t_L g114 ( 
.A(n_94),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_114),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_56),
.Y(n_115)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_94),
.Y(n_119)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_119),
.Y(n_130)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_116),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_121),
.B(n_50),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_118),
.A2(n_77),
.B1(n_56),
.B2(n_58),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_125),
.A2(n_141),
.B1(n_73),
.B2(n_63),
.Y(n_147)
);

XNOR2x1_ASAP7_75t_L g144 ( 
.A(n_126),
.B(n_137),
.Y(n_144)
);

AND2x6_ASAP7_75t_L g127 ( 
.A(n_113),
.B(n_27),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_29),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_109),
.B(n_71),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_131),
.B(n_132),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_71),
.Y(n_132)
);

AO22x1_ASAP7_75t_SL g134 ( 
.A1(n_103),
.A2(n_100),
.B1(n_98),
.B2(n_54),
.Y(n_134)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_134),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_108),
.B(n_57),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_135),
.B(n_51),
.Y(n_163)
);

INVx13_ASAP7_75t_L g136 ( 
.A(n_105),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_136),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_111),
.A2(n_72),
.B(n_60),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_137),
.A2(n_39),
.B(n_38),
.Y(n_167)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_104),
.Y(n_138)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_138),
.Y(n_150)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_120),
.Y(n_140)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_140),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_133),
.A2(n_120),
.B1(n_72),
.B2(n_60),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_143),
.A2(n_147),
.B1(n_34),
.B2(n_33),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_144),
.B(n_153),
.Y(n_185)
);

AO22x1_ASAP7_75t_L g145 ( 
.A1(n_129),
.A2(n_114),
.B1(n_116),
.B2(n_57),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_145),
.B(n_148),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g149 ( 
.A(n_126),
.B(n_73),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_149),
.B(n_165),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_123),
.B(n_122),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_151),
.B(n_154),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_130),
.B(n_142),
.C(n_127),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_128),
.B(n_139),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_134),
.A2(n_73),
.B1(n_63),
.B2(n_52),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_155),
.A2(n_30),
.B1(n_28),
.B2(n_25),
.Y(n_171)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_128),
.Y(n_157)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_157),
.Y(n_168)
);

AOI221xp5_ASAP7_75t_L g158 ( 
.A1(n_134),
.A2(n_73),
.B1(n_1),
.B2(n_2),
.C(n_3),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_158),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_121),
.B(n_0),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_159),
.A2(n_1),
.B(n_2),
.Y(n_169)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_124),
.Y(n_160)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_160),
.Y(n_176)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_124),
.Y(n_161)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_161),
.Y(n_178)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_163),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_164),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_136),
.B(n_46),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_138),
.Y(n_166)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_166),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_167),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_169),
.B(n_162),
.Y(n_190)
);

OAI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_170),
.A2(n_184),
.B1(n_186),
.B2(n_187),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_171),
.A2(n_155),
.B1(n_152),
.B2(n_150),
.Y(n_194)
);

CKINVDCx14_ASAP7_75t_R g174 ( 
.A(n_156),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_174),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_144),
.A2(n_22),
.B(n_21),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_175),
.A2(n_189),
.B(n_165),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_149),
.B(n_20),
.C(n_4),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_179),
.B(n_181),
.C(n_13),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_SL g181 ( 
.A(n_153),
.B(n_3),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_146),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_145),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_167),
.A2(n_7),
.B(n_8),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_190),
.B(n_194),
.Y(n_211)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_176),
.Y(n_191)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_191),
.Y(n_204)
);

AOI21x1_ASAP7_75t_L g205 ( 
.A1(n_193),
.A2(n_199),
.B(n_202),
.Y(n_205)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_195),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_172),
.B(n_10),
.Y(n_196)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_196),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_187),
.A2(n_158),
.B1(n_13),
.B2(n_15),
.Y(n_197)
);

INVxp67_ASAP7_75t_SL g206 ( 
.A(n_197),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_177),
.B(n_12),
.Y(n_198)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_198),
.Y(n_209)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_178),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_200),
.B(n_201),
.C(n_181),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_185),
.B(n_15),
.C(n_16),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_188),
.Y(n_202)
);

NOR3xp33_ASAP7_75t_L g203 ( 
.A(n_192),
.B(n_183),
.C(n_180),
.Y(n_203)
);

OR2x2_ASAP7_75t_L g217 ( 
.A(n_203),
.B(n_200),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_201),
.B(n_173),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_207),
.B(n_205),
.C(n_173),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_210),
.B(n_182),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_213),
.B(n_218),
.C(n_219),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_208),
.A2(n_183),
.B1(n_194),
.B2(n_197),
.Y(n_214)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_214),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_212),
.B(n_172),
.Y(n_215)
);

INVx11_ASAP7_75t_L g223 ( 
.A(n_215),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_211),
.A2(n_168),
.B1(n_174),
.B2(n_193),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_216),
.A2(n_217),
.B1(n_206),
.B2(n_203),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_204),
.B(n_16),
.C(n_17),
.Y(n_219)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_220),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_221),
.B(n_217),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_225),
.B(n_221),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_226),
.B(n_220),
.Y(n_227)
);

AO21x1_ASAP7_75t_L g228 ( 
.A1(n_227),
.A2(n_224),
.B(n_222),
.Y(n_228)
);

OAI21x1_ASAP7_75t_L g229 ( 
.A1(n_228),
.A2(n_222),
.B(n_206),
.Y(n_229)
);

NAND3xp33_ASAP7_75t_L g230 ( 
.A(n_229),
.B(n_223),
.C(n_209),
.Y(n_230)
);

OAI21x1_ASAP7_75t_L g231 ( 
.A1(n_230),
.A2(n_223),
.B(n_219),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_231),
.B(n_17),
.Y(n_232)
);


endmodule