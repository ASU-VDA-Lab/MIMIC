module fake_jpeg_25863_n_310 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_310);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_310;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx11_ASAP7_75t_SL g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_32),
.B(n_33),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_19),
.B(n_0),
.C(n_1),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_19),
.B(n_1),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_35),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_16),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_19),
.B(n_1),
.Y(n_37)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_21),
.A2(n_30),
.B1(n_23),
.B2(n_16),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_39),
.A2(n_21),
.B1(n_30),
.B2(n_17),
.Y(n_55)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_45),
.Y(n_63)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_47),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_55),
.A2(n_39),
.B1(n_37),
.B2(n_18),
.Y(n_81)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_56),
.B(n_57),
.Y(n_80)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_58),
.B(n_65),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_33),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_61),
.B(n_62),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_33),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_49),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_42),
.A2(n_48),
.B1(n_55),
.B2(n_21),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_66),
.A2(n_15),
.B1(n_20),
.B2(n_26),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_33),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_67),
.B(n_76),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_41),
.A2(n_37),
.B1(n_38),
.B2(n_21),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_69),
.A2(n_52),
.B1(n_43),
.B2(n_53),
.Y(n_88)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_70),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_41),
.A2(n_33),
.B1(n_34),
.B2(n_39),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_71),
.A2(n_81),
.B1(n_27),
.B2(n_31),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_57),
.A2(n_34),
.B1(n_30),
.B2(n_38),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_72),
.A2(n_18),
.B1(n_27),
.B2(n_22),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_49),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_73),
.Y(n_104)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_74),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_54),
.A2(n_25),
.B1(n_16),
.B2(n_24),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_75),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_44),
.B(n_34),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_44),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_82),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_56),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_45),
.B(n_37),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_84),
.B(n_38),
.C(n_46),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_85),
.B(n_101),
.Y(n_128)
);

INVx3_ASAP7_75t_SL g86 ( 
.A(n_59),
.Y(n_86)
);

INVx13_ASAP7_75t_L g119 ( 
.A(n_86),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_88),
.A2(n_96),
.B1(n_97),
.B2(n_77),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_62),
.A2(n_35),
.B(n_18),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_89),
.Y(n_127)
);

INVx2_ASAP7_75t_SL g90 ( 
.A(n_83),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_90),
.B(n_98),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_68),
.Y(n_92)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_92),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_94),
.B(n_110),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_66),
.A2(n_43),
.B1(n_35),
.B2(n_31),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_95),
.A2(n_108),
.B1(n_29),
.B2(n_22),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_67),
.A2(n_43),
.B1(n_35),
.B2(n_31),
.Y(n_96)
);

INVx1_ASAP7_75t_SL g98 ( 
.A(n_68),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_59),
.Y(n_99)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_99),
.Y(n_134)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_64),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_100),
.B(n_109),
.Y(n_136)
);

AO22x1_ASAP7_75t_L g101 ( 
.A1(n_78),
.A2(n_15),
.B1(n_20),
.B2(n_26),
.Y(n_101)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_101),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_106),
.A2(n_78),
.B1(n_77),
.B2(n_83),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_68),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_107),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_71),
.A2(n_29),
.B1(n_22),
.B2(n_27),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_64),
.Y(n_109)
);

OA22x2_ASAP7_75t_SL g110 ( 
.A1(n_61),
.A2(n_26),
.B1(n_20),
.B2(n_15),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_81),
.A2(n_2),
.B(n_3),
.Y(n_112)
);

OAI21xp33_ASAP7_75t_L g116 ( 
.A1(n_112),
.A2(n_14),
.B(n_3),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_105),
.B(n_58),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_113),
.B(n_123),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_114),
.A2(n_86),
.B1(n_60),
.B2(n_63),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_96),
.A2(n_76),
.B1(n_84),
.B2(n_70),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_115),
.A2(n_118),
.B1(n_125),
.B2(n_130),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_116),
.B(n_129),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_88),
.A2(n_72),
.B1(n_78),
.B2(n_80),
.Y(n_118)
);

AOI21xp33_ASAP7_75t_SL g120 ( 
.A1(n_110),
.A2(n_80),
.B(n_69),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_120),
.A2(n_93),
.B(n_103),
.Y(n_144)
);

BUFx24_ASAP7_75t_SL g121 ( 
.A(n_102),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_121),
.B(n_111),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_122),
.A2(n_126),
.B1(n_117),
.B2(n_131),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_105),
.B(n_82),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_91),
.A2(n_74),
.B1(n_83),
.B2(n_77),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_128),
.B(n_86),
.Y(n_162)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_87),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_94),
.A2(n_110),
.B1(n_97),
.B2(n_112),
.Y(n_130)
);

AND2x2_ASAP7_75t_SL g131 ( 
.A(n_110),
.B(n_79),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_131),
.B(n_140),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_89),
.B(n_25),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_133),
.B(n_137),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_95),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_85),
.A2(n_60),
.B1(n_65),
.B2(n_73),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_139),
.A2(n_92),
.B1(n_29),
.B2(n_28),
.Y(n_170)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_104),
.Y(n_140)
);

INVxp33_ASAP7_75t_L g141 ( 
.A(n_136),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_141),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_113),
.B(n_93),
.C(n_123),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_143),
.B(n_145),
.C(n_153),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_144),
.A2(n_132),
.B(n_133),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_128),
.B(n_103),
.C(n_108),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_146),
.A2(n_152),
.B1(n_119),
.B2(n_124),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_120),
.A2(n_104),
.B1(n_111),
.B2(n_90),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_147),
.A2(n_164),
.B1(n_170),
.B2(n_172),
.Y(n_177)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_136),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_148),
.B(n_149),
.Y(n_179)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_135),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_150),
.B(n_163),
.Y(n_174)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_135),
.Y(n_151)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_151),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_117),
.A2(n_90),
.B1(n_60),
.B2(n_98),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_139),
.B(n_109),
.C(n_100),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_125),
.B(n_63),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_155),
.A2(n_131),
.B(n_118),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_115),
.B(n_101),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_156),
.B(n_162),
.Y(n_196)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_140),
.Y(n_158)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_158),
.Y(n_175)
);

INVx3_ASAP7_75t_SL g160 ( 
.A(n_134),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_160),
.A2(n_124),
.B1(n_119),
.B2(n_5),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_127),
.B(n_99),
.Y(n_161)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_161),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_129),
.B(n_107),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_130),
.B(n_63),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_165),
.B(n_166),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_132),
.B(n_107),
.C(n_92),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_138),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_168),
.Y(n_178)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_122),
.Y(n_169)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_169),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_138),
.B(n_28),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_171),
.B(n_24),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_114),
.A2(n_28),
.B1(n_24),
.B2(n_4),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_176),
.B(n_185),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_183),
.B(n_186),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_159),
.A2(n_132),
.B1(n_131),
.B2(n_126),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_185),
.A2(n_199),
.B1(n_201),
.B2(n_7),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_168),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_167),
.B(n_154),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_187),
.B(n_189),
.Y(n_214)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_157),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_157),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_190),
.B(n_197),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_191),
.A2(n_192),
.B1(n_198),
.B2(n_7),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_169),
.A2(n_146),
.B1(n_166),
.B2(n_145),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_193),
.B(n_9),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_144),
.B(n_132),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_194),
.B(n_7),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_161),
.A2(n_134),
.B(n_3),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_195),
.A2(n_200),
.B(n_202),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_158),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_153),
.A2(n_151),
.B1(n_149),
.B2(n_159),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_160),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_147),
.A2(n_124),
.B1(n_119),
.B2(n_14),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_155),
.A2(n_2),
.B(n_4),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_170),
.Y(n_203)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_203),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_192),
.A2(n_165),
.B1(n_155),
.B2(n_148),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_204),
.A2(n_215),
.B1(n_225),
.B2(n_195),
.Y(n_234)
);

AOI21x1_ASAP7_75t_SL g205 ( 
.A1(n_193),
.A2(n_162),
.B(n_156),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_205),
.B(n_208),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_182),
.B(n_143),
.C(n_142),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_206),
.B(n_210),
.C(n_211),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_182),
.B(n_142),
.C(n_172),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_196),
.B(n_160),
.C(n_14),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_179),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_212),
.B(n_213),
.Y(n_228)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_179),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_188),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_196),
.B(n_4),
.C(n_5),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_216),
.B(n_217),
.C(n_227),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_180),
.B(n_5),
.C(n_6),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_201),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_218),
.B(n_202),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_219),
.A2(n_221),
.B(n_200),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_203),
.A2(n_188),
.B1(n_173),
.B2(n_181),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_223),
.B(n_226),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_224),
.B(n_177),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_184),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_180),
.B(n_9),
.C(n_10),
.Y(n_227)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_231),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_207),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_233),
.Y(n_261)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_234),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_205),
.B(n_194),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_236),
.B(n_237),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_204),
.B(n_176),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_208),
.A2(n_184),
.B(n_186),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_238),
.A2(n_241),
.B(n_246),
.Y(n_248)
);

NOR3xp33_ASAP7_75t_L g239 ( 
.A(n_222),
.B(n_178),
.C(n_173),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_239),
.B(n_243),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g240 ( 
.A(n_223),
.B(n_177),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_240),
.B(n_225),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_221),
.Y(n_241)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_242),
.Y(n_251)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_220),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_206),
.B(n_190),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_244),
.B(n_227),
.Y(n_255)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_214),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_245),
.B(n_234),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_244),
.B(n_174),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_252),
.B(n_235),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_232),
.B(n_210),
.C(n_211),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_254),
.B(n_259),
.C(n_240),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_255),
.B(n_260),
.Y(n_263)
);

BUFx12_ASAP7_75t_L g256 ( 
.A(n_238),
.Y(n_256)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_256),
.Y(n_265)
);

A2O1A1Ixp33_ASAP7_75t_SL g257 ( 
.A1(n_241),
.A2(n_178),
.B(n_209),
.C(n_189),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_257),
.A2(n_228),
.B(n_175),
.Y(n_271)
);

OA21x2_ASAP7_75t_SL g258 ( 
.A1(n_229),
.A2(n_216),
.B(n_226),
.Y(n_258)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_258),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_232),
.B(n_217),
.C(n_175),
.Y(n_259)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_262),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_255),
.B(n_237),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_264),
.B(n_250),
.Y(n_280)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_249),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_268),
.B(n_269),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_270),
.B(n_276),
.C(n_254),
.Y(n_277)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_271),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_261),
.B(n_215),
.Y(n_272)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_272),
.Y(n_285)
);

OR2x2_ASAP7_75t_L g273 ( 
.A(n_257),
.B(n_230),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_273),
.A2(n_248),
.B(n_257),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_253),
.A2(n_230),
.B1(n_260),
.B2(n_247),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_274),
.A2(n_256),
.B1(n_250),
.B2(n_229),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_251),
.B(n_235),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_275),
.B(n_263),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_259),
.B(n_230),
.C(n_236),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_277),
.B(n_283),
.C(n_284),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_278),
.B(n_280),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_282),
.B(n_267),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_270),
.B(n_253),
.C(n_248),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_276),
.B(n_257),
.C(n_256),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_286),
.B(n_287),
.C(n_266),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_263),
.B(n_264),
.C(n_274),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_289),
.B(n_291),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_290),
.B(n_292),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_277),
.B(n_265),
.C(n_273),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_283),
.B(n_271),
.C(n_11),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_279),
.B(n_10),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_294),
.B(n_285),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_287),
.B(n_10),
.C(n_11),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_295),
.B(n_296),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_284),
.B(n_11),
.C(n_12),
.Y(n_296)
);

BUFx24_ASAP7_75t_SL g297 ( 
.A(n_293),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_297),
.B(n_298),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_288),
.B(n_281),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_301),
.B(n_280),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_304),
.B(n_305),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_302),
.B(n_286),
.C(n_12),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_306),
.B(n_303),
.Y(n_307)
);

OAI321xp33_ASAP7_75t_L g308 ( 
.A1(n_307),
.A2(n_11),
.A3(n_13),
.B1(n_299),
.B2(n_300),
.C(n_306),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_308),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_309),
.B(n_13),
.Y(n_310)
);


endmodule