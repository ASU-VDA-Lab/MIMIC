module fake_netlist_6_4331_n_718 (n_16, n_1, n_9, n_8, n_18, n_10, n_21, n_24, n_6, n_15, n_27, n_3, n_14, n_0, n_4, n_22, n_26, n_13, n_11, n_28, n_17, n_23, n_12, n_20, n_7, n_2, n_5, n_19, n_25, n_718);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_6;
input n_15;
input n_27;
input n_3;
input n_14;
input n_0;
input n_4;
input n_22;
input n_26;
input n_13;
input n_11;
input n_28;
input n_17;
input n_23;
input n_12;
input n_20;
input n_7;
input n_2;
input n_5;
input n_19;
input n_25;

output n_718;

wire n_52;
wire n_591;
wire n_435;
wire n_91;
wire n_326;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_209;
wire n_465;
wire n_367;
wire n_680;
wire n_590;
wire n_625;
wire n_63;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_148;
wire n_226;
wire n_161;
wire n_208;
wire n_462;
wire n_68;
wire n_607;
wire n_671;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_50;
wire n_694;
wire n_578;
wire n_703;
wire n_144;
wire n_365;
wire n_125;
wire n_168;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_77;
wire n_106;
wire n_358;
wire n_160;
wire n_449;
wire n_131;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_575;
wire n_368;
wire n_677;
wire n_396;
wire n_495;
wire n_350;
wire n_78;
wire n_84;
wire n_585;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_142;
wire n_143;
wire n_382;
wire n_673;
wire n_180;
wire n_62;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_255;
wire n_284;
wire n_400;
wire n_140;
wire n_337;
wire n_214;
wire n_485;
wire n_67;
wire n_443;
wire n_246;
wire n_38;
wire n_471;
wire n_289;
wire n_421;
wire n_424;
wire n_615;
wire n_59;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_202;
wire n_320;
wire n_108;
wire n_639;
wire n_676;
wire n_327;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_65;
wire n_230;
wire n_605;
wire n_461;
wire n_141;
wire n_383;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_114;
wire n_86;
wire n_198;
wire n_104;
wire n_222;
wire n_179;
wire n_248;
wire n_300;
wire n_517;
wire n_667;
wire n_71;
wire n_74;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_72;
wire n_532;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_111;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_35;
wire n_183;
wire n_510;
wire n_79;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_506;
wire n_56;
wire n_360;
wire n_603;
wire n_119;
wire n_235;
wire n_536;
wire n_622;
wire n_147;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_39;
wire n_344;
wire n_73;
wire n_581;
wire n_428;
wire n_609;
wire n_432;
wire n_641;
wire n_693;
wire n_101;
wire n_167;
wire n_631;
wire n_174;
wire n_127;
wire n_516;
wire n_153;
wire n_525;
wire n_611;
wire n_156;
wire n_491;
wire n_145;
wire n_42;
wire n_133;
wire n_656;
wire n_96;
wire n_666;
wire n_371;
wire n_567;
wire n_189;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_129;
wire n_705;
wire n_647;
wire n_197;
wire n_137;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_155;
wire n_109;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_122;
wire n_45;
wire n_454;
wire n_34;
wire n_218;
wire n_638;
wire n_70;
wire n_234;
wire n_37;
wire n_486;
wire n_381;
wire n_82;
wire n_236;
wire n_653;
wire n_112;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_126;
wire n_414;
wire n_97;
wire n_563;
wire n_58;
wire n_490;
wire n_290;
wire n_220;
wire n_118;
wire n_224;
wire n_48;
wire n_93;
wire n_80;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_460;
wire n_107;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_89;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_407;
wire n_450;
wire n_103;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_69;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_31;
wire n_334;
wire n_559;
wire n_53;
wire n_370;
wire n_44;
wire n_458;
wire n_232;
wire n_650;
wire n_163;
wire n_717;
wire n_46;
wire n_330;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_154;
wire n_699;
wire n_456;
wire n_564;
wire n_98;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_686;
wire n_252;
wire n_228;
wire n_565;
wire n_594;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_83;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_716;
wire n_152;
wire n_623;
wire n_92;
wire n_599;
wire n_513;
wire n_321;
wire n_645;
wire n_331;
wire n_105;
wire n_227;
wire n_132;
wire n_570;
wire n_406;
wire n_483;
wire n_102;
wire n_204;
wire n_482;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_32;
wire n_66;
wire n_130;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_100;
wire n_121;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_150;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_325;
wire n_329;
wire n_464;
wire n_600;
wire n_561;
wire n_33;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_61;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_76;
wire n_243;
wire n_124;
wire n_548;
wire n_94;
wire n_282;
wire n_436;
wire n_116;
wire n_211;
wire n_523;
wire n_117;
wire n_175;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_40;
wire n_505;
wire n_240;
wire n_139;
wire n_319;
wire n_41;
wire n_134;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_95;
wire n_311;
wire n_403;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_123;
wire n_136;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_556;
wire n_159;
wire n_157;
wire n_162;
wire n_692;
wire n_115;
wire n_487;
wire n_550;
wire n_128;
wire n_241;
wire n_30;
wire n_275;
wire n_553;
wire n_43;
wire n_652;
wire n_560;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_146;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_88;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_113;
wire n_618;
wire n_582;
wire n_199;
wire n_138;
wire n_266;
wire n_296;
wire n_674;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_158;
wire n_217;
wire n_49;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_355;
wire n_426;
wire n_317;
wire n_149;
wire n_632;
wire n_702;
wire n_431;
wire n_90;
wire n_347;
wire n_459;
wire n_54;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_87;
wire n_195;
wire n_285;
wire n_497;
wire n_675;
wire n_85;
wire n_99;
wire n_257;
wire n_655;
wire n_706;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_47;
wire n_690;
wire n_29;
wire n_75;
wire n_401;
wire n_324;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_120;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_681;
wire n_110;
wire n_151;
wire n_412;
wire n_640;
wire n_81;
wire n_660;
wire n_36;
wire n_55;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_515;
wire n_64;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_135;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_457;
wire n_391;
wire n_687;
wire n_697;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_187;
wire n_501;
wire n_531;
wire n_60;
wire n_361;
wire n_508;
wire n_663;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_410;
wire n_398;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_171;
wire n_678;
wire n_192;
wire n_57;
wire n_169;
wire n_51;
wire n_649;
wire n_283;

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx5p33_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx5p33_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_28),
.Y(n_33)
);

CKINVDCx5p33_ASAP7_75t_R g34 ( 
.A(n_27),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_9),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

CKINVDCx5p33_ASAP7_75t_R g37 ( 
.A(n_18),
.Y(n_37)
);

CKINVDCx5p33_ASAP7_75t_R g38 ( 
.A(n_13),
.Y(n_38)
);

CKINVDCx5p33_ASAP7_75t_R g39 ( 
.A(n_6),
.Y(n_39)
);

CKINVDCx5p33_ASAP7_75t_R g40 ( 
.A(n_18),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_12),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

CKINVDCx5p33_ASAP7_75t_R g44 ( 
.A(n_6),
.Y(n_44)
);

CKINVDCx5p33_ASAP7_75t_R g45 ( 
.A(n_21),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_3),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_14),
.Y(n_49)
);

CKINVDCx5p33_ASAP7_75t_R g50 ( 
.A(n_22),
.Y(n_50)
);

CKINVDCx5p33_ASAP7_75t_R g51 ( 
.A(n_7),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_11),
.Y(n_52)
);

CKINVDCx5p33_ASAP7_75t_R g53 ( 
.A(n_25),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_10),
.Y(n_54)
);

CKINVDCx5p33_ASAP7_75t_R g55 ( 
.A(n_24),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_1),
.Y(n_56)
);

CKINVDCx5p33_ASAP7_75t_R g57 ( 
.A(n_10),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

HB1xp67_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

CKINVDCx5p33_ASAP7_75t_R g61 ( 
.A(n_30),
.Y(n_61)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

BUFx8_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

AND2x4_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_23),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_35),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_31),
.B(n_0),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_67),
.Y(n_72)
);

CKINVDCx5p33_ASAP7_75t_R g73 ( 
.A(n_61),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_61),
.Y(n_75)
);

CKINVDCx5p33_ASAP7_75t_R g76 ( 
.A(n_59),
.Y(n_76)
);

CKINVDCx5p33_ASAP7_75t_R g77 ( 
.A(n_59),
.Y(n_77)
);

CKINVDCx5p33_ASAP7_75t_R g78 ( 
.A(n_58),
.Y(n_78)
);

NOR2x1p5_ASAP7_75t_L g79 ( 
.A(n_58),
.B(n_56),
.Y(n_79)
);

CKINVDCx5p33_ASAP7_75t_R g80 ( 
.A(n_64),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

CKINVDCx5p33_ASAP7_75t_R g84 ( 
.A(n_64),
.Y(n_84)
);

CKINVDCx5p33_ASAP7_75t_R g85 ( 
.A(n_58),
.Y(n_85)
);

CKINVDCx5p33_ASAP7_75t_R g86 ( 
.A(n_58),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

CKINVDCx5p33_ASAP7_75t_R g88 ( 
.A(n_71),
.Y(n_88)
);

CKINVDCx5p33_ASAP7_75t_R g89 ( 
.A(n_71),
.Y(n_89)
);

CKINVDCx5p33_ASAP7_75t_R g90 ( 
.A(n_71),
.Y(n_90)
);

CKINVDCx5p33_ASAP7_75t_R g91 ( 
.A(n_71),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_71),
.Y(n_92)
);

CKINVDCx5p33_ASAP7_75t_R g93 ( 
.A(n_71),
.Y(n_93)
);

NAND2xp33_ASAP7_75t_R g94 ( 
.A(n_66),
.B(n_69),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_78),
.B(n_63),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_78),
.B(n_33),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_85),
.B(n_69),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_63),
.Y(n_98)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_88),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_76),
.B(n_66),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_77),
.B(n_80),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_66),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_73),
.B(n_66),
.Y(n_103)
);

NAND3xp33_ASAP7_75t_L g104 ( 
.A(n_94),
.B(n_68),
.C(n_44),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_92),
.Y(n_105)
);

OR2x6_ASAP7_75t_L g106 ( 
.A(n_79),
.B(n_47),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_63),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_81),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_90),
.B(n_63),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_74),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g111 ( 
.A(n_92),
.Y(n_111)
);

NOR2xp67_ASAP7_75t_L g112 ( 
.A(n_91),
.B(n_62),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_93),
.B(n_66),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_79),
.B(n_70),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_74),
.B(n_66),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_75),
.B(n_50),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_82),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_82),
.Y(n_118)
);

NAND3xp33_ASAP7_75t_L g119 ( 
.A(n_94),
.B(n_68),
.C(n_57),
.Y(n_119)
);

NAND2xp33_ASAP7_75t_L g120 ( 
.A(n_83),
.B(n_45),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_83),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_81),
.B(n_65),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_72),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_75),
.B(n_55),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g125 ( 
.A(n_81),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_87),
.B(n_70),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_72),
.B(n_34),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_72),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_81),
.B(n_65),
.Y(n_129)
);

NOR2xp67_ASAP7_75t_L g130 ( 
.A(n_87),
.B(n_62),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_87),
.B(n_53),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_85),
.B(n_65),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_78),
.B(n_63),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_92),
.Y(n_134)
);

NAND2xp33_ASAP7_75t_L g135 ( 
.A(n_78),
.B(n_65),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_97),
.B(n_39),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_132),
.B(n_63),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_126),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_132),
.B(n_65),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_113),
.A2(n_62),
.B(n_67),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_110),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_117),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_114),
.B(n_65),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_97),
.B(n_37),
.Y(n_144)
);

INVx2_ASAP7_75t_SL g145 ( 
.A(n_106),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_R g146 ( 
.A(n_135),
.B(n_41),
.Y(n_146)
);

INVx1_ASAP7_75t_SL g147 ( 
.A(n_101),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_101),
.B(n_52),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_99),
.B(n_65),
.Y(n_149)
);

INVx2_ASAP7_75t_SL g150 ( 
.A(n_106),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_104),
.A2(n_49),
.B1(n_46),
.B2(n_119),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_99),
.B(n_65),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_118),
.Y(n_153)
);

OR2x2_ASAP7_75t_L g154 ( 
.A(n_96),
.B(n_43),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_102),
.B(n_71),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_102),
.B(n_38),
.Y(n_156)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_108),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_103),
.B(n_40),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_106),
.A2(n_65),
.B1(n_71),
.B2(n_32),
.Y(n_159)
);

INVxp67_ASAP7_75t_SL g160 ( 
.A(n_108),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_121),
.B(n_71),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_111),
.B(n_62),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_108),
.Y(n_163)
);

INVx2_ASAP7_75t_SL g164 ( 
.A(n_100),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_116),
.Y(n_165)
);

AND2x4_ASAP7_75t_L g166 ( 
.A(n_127),
.B(n_131),
.Y(n_166)
);

OAI21xp33_ASAP7_75t_L g167 ( 
.A1(n_124),
.A2(n_47),
.B(n_42),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_115),
.A2(n_134),
.B1(n_105),
.B2(n_127),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_123),
.Y(n_169)
);

BUFx2_ASAP7_75t_L g170 ( 
.A(n_115),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_111),
.B(n_62),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_128),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_120),
.A2(n_51),
.B1(n_70),
.B2(n_56),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_111),
.B(n_62),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_108),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_111),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_111),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_95),
.B(n_43),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_111),
.Y(n_179)
);

O2A1O1Ixp33_ASAP7_75t_L g180 ( 
.A1(n_131),
.A2(n_42),
.B(n_32),
.C(n_70),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_125),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_125),
.B(n_62),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_98),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_133),
.A2(n_67),
.B1(n_70),
.B2(n_62),
.Y(n_184)
);

BUFx8_ASAP7_75t_L g185 ( 
.A(n_125),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_125),
.B(n_109),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_122),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_125),
.B(n_62),
.Y(n_188)
);

AND3x2_ASAP7_75t_SL g189 ( 
.A(n_122),
.B(n_2),
.C(n_4),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_125),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_112),
.B(n_70),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_129),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_129),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_107),
.B(n_8),
.Y(n_194)
);

BUFx2_ASAP7_75t_L g195 ( 
.A(n_130),
.Y(n_195)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_108),
.Y(n_196)
);

O2A1O1Ixp5_ASAP7_75t_L g197 ( 
.A1(n_194),
.A2(n_67),
.B(n_20),
.C(n_62),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_136),
.A2(n_67),
.B1(n_12),
.B2(n_13),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_163),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_147),
.B(n_8),
.Y(n_200)
);

O2A1O1Ixp33_ASAP7_75t_L g201 ( 
.A1(n_170),
.A2(n_178),
.B(n_144),
.C(n_154),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_165),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_148),
.B(n_15),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_143),
.A2(n_67),
.B(n_16),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_141),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_170),
.B(n_67),
.Y(n_206)
);

NOR3xp33_ASAP7_75t_L g207 ( 
.A(n_151),
.B(n_167),
.C(n_158),
.Y(n_207)
);

OAI22xp33_ASAP7_75t_L g208 ( 
.A1(n_164),
.A2(n_183),
.B1(n_154),
.B2(n_150),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_155),
.A2(n_149),
.B(n_152),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_153),
.B(n_15),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_183),
.A2(n_16),
.B1(n_17),
.B2(n_19),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_163),
.Y(n_212)
);

OR2x6_ASAP7_75t_L g213 ( 
.A(n_145),
.B(n_17),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_153),
.B(n_19),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_196),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_177),
.A2(n_190),
.B(n_160),
.Y(n_216)
);

AOI21x1_ASAP7_75t_L g217 ( 
.A1(n_162),
.A2(n_174),
.B(n_171),
.Y(n_217)
);

NOR3xp33_ASAP7_75t_SL g218 ( 
.A(n_156),
.B(n_189),
.C(n_180),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_155),
.A2(n_139),
.B(n_138),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_138),
.A2(n_166),
.B(n_187),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_141),
.B(n_142),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_142),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_166),
.A2(n_187),
.B(n_176),
.Y(n_223)
);

INVx8_ASAP7_75t_L g224 ( 
.A(n_166),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_169),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_187),
.B(n_164),
.Y(n_226)
);

O2A1O1Ixp5_ASAP7_75t_L g227 ( 
.A1(n_186),
.A2(n_137),
.B(n_193),
.C(n_192),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_145),
.B(n_150),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_187),
.B(n_193),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_165),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_146),
.B(n_173),
.Y(n_231)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_196),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_187),
.A2(n_176),
.B(n_179),
.Y(n_233)
);

NOR2xp67_ASAP7_75t_L g234 ( 
.A(n_172),
.B(n_161),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_179),
.A2(n_177),
.B(n_168),
.Y(n_235)
);

OR2x2_ASAP7_75t_L g236 ( 
.A(n_172),
.B(n_159),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_169),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_175),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_185),
.B(n_195),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_192),
.B(n_175),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_181),
.A2(n_191),
.B(n_190),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_181),
.A2(n_184),
.B(n_196),
.Y(n_242)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_157),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_195),
.Y(n_244)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_157),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_157),
.A2(n_140),
.B1(n_182),
.B2(n_188),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_185),
.A2(n_136),
.B1(n_183),
.B2(n_166),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_185),
.A2(n_189),
.B1(n_136),
.B2(n_183),
.Y(n_248)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_245),
.Y(n_249)
);

BUFx4f_ASAP7_75t_L g250 ( 
.A(n_224),
.Y(n_250)
);

BUFx2_ASAP7_75t_L g251 ( 
.A(n_202),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_225),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_230),
.Y(n_253)
);

AO21x2_ASAP7_75t_L g254 ( 
.A1(n_209),
.A2(n_189),
.B(n_235),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_227),
.A2(n_235),
.B(n_219),
.Y(n_255)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_224),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_219),
.A2(n_223),
.B(n_209),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_229),
.B(n_226),
.Y(n_258)
);

OAI21x1_ASAP7_75t_L g259 ( 
.A1(n_217),
.A2(n_233),
.B(n_223),
.Y(n_259)
);

BUFx3_ASAP7_75t_L g260 ( 
.A(n_224),
.Y(n_260)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_245),
.Y(n_261)
);

OAI21x1_ASAP7_75t_L g262 ( 
.A1(n_233),
.A2(n_246),
.B(n_220),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_215),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_244),
.Y(n_264)
);

NAND2x1p5_ASAP7_75t_L g265 ( 
.A(n_243),
.B(n_220),
.Y(n_265)
);

OAI21x1_ASAP7_75t_SL g266 ( 
.A1(n_240),
.A2(n_242),
.B(n_214),
.Y(n_266)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_199),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_248),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_208),
.B(n_200),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g270 ( 
.A(n_199),
.Y(n_270)
);

OAI21x1_ASAP7_75t_L g271 ( 
.A1(n_241),
.A2(n_216),
.B(n_197),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_237),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_215),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_205),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_L g275 ( 
.A1(n_207),
.A2(n_203),
.B1(n_231),
.B2(n_222),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_238),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_221),
.Y(n_277)
);

INVx1_ASAP7_75t_SL g278 ( 
.A(n_210),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_232),
.Y(n_279)
);

AOI21x1_ASAP7_75t_L g280 ( 
.A1(n_234),
.A2(n_206),
.B(n_241),
.Y(n_280)
);

BUFx10_ASAP7_75t_L g281 ( 
.A(n_228),
.Y(n_281)
);

OA21x2_ASAP7_75t_L g282 ( 
.A1(n_204),
.A2(n_218),
.B(n_198),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_201),
.B(n_236),
.Y(n_283)
);

BUFx8_ASAP7_75t_L g284 ( 
.A(n_199),
.Y(n_284)
);

INVx4_ASAP7_75t_L g285 ( 
.A(n_243),
.Y(n_285)
);

NOR2x1_ASAP7_75t_R g286 ( 
.A(n_239),
.B(n_212),
.Y(n_286)
);

BUFx12f_ASAP7_75t_L g287 ( 
.A(n_213),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_232),
.Y(n_288)
);

BUFx3_ASAP7_75t_L g289 ( 
.A(n_212),
.Y(n_289)
);

INVx1_ASAP7_75t_SL g290 ( 
.A(n_212),
.Y(n_290)
);

INVx6_ASAP7_75t_L g291 ( 
.A(n_215),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_204),
.Y(n_292)
);

INVxp33_ASAP7_75t_L g293 ( 
.A(n_247),
.Y(n_293)
);

INVx1_ASAP7_75t_SL g294 ( 
.A(n_213),
.Y(n_294)
);

NAND2x1p5_ASAP7_75t_L g295 ( 
.A(n_211),
.B(n_213),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_200),
.Y(n_296)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_245),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_227),
.A2(n_235),
.B(n_219),
.Y(n_298)
);

BUFx2_ASAP7_75t_L g299 ( 
.A(n_202),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_225),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_225),
.Y(n_301)
);

BUFx12f_ASAP7_75t_L g302 ( 
.A(n_202),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_225),
.Y(n_303)
);

BUFx3_ASAP7_75t_L g304 ( 
.A(n_224),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_245),
.A2(n_177),
.B(n_190),
.Y(n_305)
);

AND2x4_ASAP7_75t_L g306 ( 
.A(n_256),
.B(n_304),
.Y(n_306)
);

BUFx3_ASAP7_75t_L g307 ( 
.A(n_284),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_252),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_252),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_252),
.Y(n_310)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_285),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_L g312 ( 
.A1(n_269),
.A2(n_295),
.B1(n_275),
.B2(n_293),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_251),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_277),
.B(n_254),
.Y(n_314)
);

BUFx2_ASAP7_75t_L g315 ( 
.A(n_264),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_SL g316 ( 
.A1(n_268),
.A2(n_295),
.B1(n_254),
.B2(n_296),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_257),
.A2(n_298),
.B(n_255),
.Y(n_317)
);

NAND2x1_ASAP7_75t_L g318 ( 
.A(n_249),
.B(n_261),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_274),
.Y(n_319)
);

INVx1_ASAP7_75t_SL g320 ( 
.A(n_264),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_302),
.Y(n_321)
);

NOR2x1_ASAP7_75t_SL g322 ( 
.A(n_292),
.B(n_280),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_302),
.Y(n_323)
);

BUFx2_ASAP7_75t_L g324 ( 
.A(n_284),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_277),
.B(n_258),
.Y(n_325)
);

NAND2x1p5_ASAP7_75t_L g326 ( 
.A(n_262),
.B(n_259),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_302),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_L g328 ( 
.A1(n_295),
.A2(n_254),
.B1(n_278),
.B2(n_282),
.Y(n_328)
);

OAI21x1_ASAP7_75t_L g329 ( 
.A1(n_259),
.A2(n_271),
.B(n_262),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_SL g330 ( 
.A1(n_268),
.A2(n_254),
.B1(n_287),
.B2(n_282),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_251),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g332 ( 
.A(n_267),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_276),
.Y(n_333)
);

OAI21x1_ASAP7_75t_L g334 ( 
.A1(n_271),
.A2(n_257),
.B(n_280),
.Y(n_334)
);

AO21x2_ASAP7_75t_L g335 ( 
.A1(n_255),
.A2(n_298),
.B(n_266),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_276),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_283),
.B(n_278),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_276),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_250),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g340 ( 
.A(n_282),
.B(n_300),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_282),
.A2(n_250),
.B1(n_265),
.B2(n_292),
.Y(n_341)
);

AOI21x1_ASAP7_75t_L g342 ( 
.A1(n_266),
.A2(n_305),
.B(n_303),
.Y(n_342)
);

AOI22xp33_ASAP7_75t_L g343 ( 
.A1(n_294),
.A2(n_287),
.B1(n_272),
.B2(n_300),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_272),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_301),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_L g346 ( 
.A1(n_294),
.A2(n_287),
.B1(n_301),
.B2(n_303),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_279),
.Y(n_347)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_285),
.Y(n_348)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_267),
.Y(n_349)
);

INVx1_ASAP7_75t_SL g350 ( 
.A(n_299),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_279),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_253),
.B(n_299),
.Y(n_352)
);

CKINVDCx16_ASAP7_75t_R g353 ( 
.A(n_313),
.Y(n_353)
);

BUFx3_ASAP7_75t_L g354 ( 
.A(n_315),
.Y(n_354)
);

A2O1A1Ixp33_ASAP7_75t_L g355 ( 
.A1(n_317),
.A2(n_250),
.B(n_249),
.C(n_297),
.Y(n_355)
);

BUFx2_ASAP7_75t_L g356 ( 
.A(n_317),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_340),
.Y(n_357)
);

NOR3xp33_ASAP7_75t_SL g358 ( 
.A(n_331),
.B(n_286),
.C(n_288),
.Y(n_358)
);

NOR3xp33_ASAP7_75t_SL g359 ( 
.A(n_321),
.B(n_286),
.C(n_288),
.Y(n_359)
);

INVx3_ASAP7_75t_L g360 ( 
.A(n_326),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_340),
.Y(n_361)
);

NAND3xp33_ASAP7_75t_SL g362 ( 
.A(n_312),
.B(n_265),
.C(n_290),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_323),
.Y(n_363)
);

OR2x2_ASAP7_75t_L g364 ( 
.A(n_314),
.B(n_265),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_340),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_329),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_327),
.Y(n_367)
);

NOR2x1_ASAP7_75t_SL g368 ( 
.A(n_341),
.B(n_285),
.Y(n_368)
);

BUFx3_ASAP7_75t_L g369 ( 
.A(n_307),
.Y(n_369)
);

CKINVDCx8_ASAP7_75t_R g370 ( 
.A(n_339),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_314),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_329),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_325),
.B(n_249),
.Y(n_373)
);

OR2x2_ASAP7_75t_L g374 ( 
.A(n_335),
.B(n_261),
.Y(n_374)
);

CKINVDCx16_ASAP7_75t_R g375 ( 
.A(n_307),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_333),
.Y(n_376)
);

AND2x2_ASAP7_75t_L g377 ( 
.A(n_328),
.B(n_263),
.Y(n_377)
);

HB1xp67_ASAP7_75t_L g378 ( 
.A(n_341),
.Y(n_378)
);

OR2x6_ASAP7_75t_L g379 ( 
.A(n_326),
.B(n_304),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_333),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_334),
.Y(n_381)
);

HB1xp67_ASAP7_75t_L g382 ( 
.A(n_332),
.Y(n_382)
);

BUFx3_ASAP7_75t_L g383 ( 
.A(n_307),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_330),
.B(n_263),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_330),
.B(n_263),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_338),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_338),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_337),
.B(n_290),
.Y(n_388)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_316),
.B(n_273),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_357),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_366),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_357),
.Y(n_392)
);

HB1xp67_ASAP7_75t_L g393 ( 
.A(n_374),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_371),
.B(n_335),
.Y(n_394)
);

HB1xp67_ASAP7_75t_L g395 ( 
.A(n_374),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_379),
.Y(n_396)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_360),
.Y(n_397)
);

INVx5_ASAP7_75t_L g398 ( 
.A(n_379),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_366),
.Y(n_399)
);

AOI221xp5_ASAP7_75t_L g400 ( 
.A1(n_356),
.A2(n_337),
.B1(n_316),
.B2(n_320),
.C(n_315),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_366),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_372),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_371),
.B(n_357),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_361),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_361),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_356),
.B(n_335),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_356),
.B(n_335),
.Y(n_407)
);

INVx2_ASAP7_75t_SL g408 ( 
.A(n_379),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_370),
.A2(n_325),
.B1(n_350),
.B2(n_346),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_388),
.B(n_350),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_365),
.Y(n_411)
);

AND2x4_ASAP7_75t_L g412 ( 
.A(n_379),
.B(n_322),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_372),
.Y(n_413)
);

INVx3_ASAP7_75t_L g414 ( 
.A(n_360),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_365),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_388),
.B(n_336),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_376),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_384),
.B(n_334),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_384),
.B(n_334),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_376),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_384),
.B(n_326),
.Y(n_421)
);

NAND4xp25_ASAP7_75t_L g422 ( 
.A(n_373),
.B(n_343),
.C(n_352),
.D(n_320),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_372),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_385),
.B(n_326),
.Y(n_424)
);

OR2x2_ASAP7_75t_L g425 ( 
.A(n_378),
.B(n_347),
.Y(n_425)
);

INVx1_ASAP7_75t_SL g426 ( 
.A(n_354),
.Y(n_426)
);

NAND3xp33_ASAP7_75t_L g427 ( 
.A(n_358),
.B(n_344),
.C(n_345),
.Y(n_427)
);

OR2x2_ASAP7_75t_L g428 ( 
.A(n_393),
.B(n_378),
.Y(n_428)
);

INVx2_ASAP7_75t_SL g429 ( 
.A(n_396),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_418),
.B(n_385),
.Y(n_430)
);

AND2x2_ASAP7_75t_L g431 ( 
.A(n_418),
.B(n_385),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_417),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_403),
.B(n_382),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g434 ( 
.A(n_418),
.B(n_419),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_419),
.B(n_389),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_410),
.B(n_353),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_417),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_419),
.B(n_389),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_401),
.Y(n_439)
);

OR2x6_ASAP7_75t_SL g440 ( 
.A(n_427),
.B(n_364),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_420),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_409),
.B(n_353),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_401),
.Y(n_443)
);

OR2x2_ASAP7_75t_L g444 ( 
.A(n_393),
.B(n_395),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_421),
.B(n_389),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_403),
.B(n_382),
.Y(n_446)
);

AND2x2_ASAP7_75t_L g447 ( 
.A(n_421),
.B(n_364),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_420),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_404),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_403),
.B(n_394),
.Y(n_450)
);

OAI21xp33_ASAP7_75t_L g451 ( 
.A1(n_400),
.A2(n_358),
.B(n_359),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_404),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_401),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_394),
.B(n_364),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_405),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_401),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_394),
.B(n_374),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_423),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_423),
.Y(n_459)
);

NAND4xp25_ASAP7_75t_L g460 ( 
.A(n_410),
.B(n_354),
.C(n_373),
.D(n_362),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_405),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_395),
.B(n_354),
.Y(n_462)
);

INVxp67_ASAP7_75t_L g463 ( 
.A(n_425),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_423),
.Y(n_464)
);

AND2x4_ASAP7_75t_L g465 ( 
.A(n_396),
.B(n_379),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_411),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_434),
.B(n_421),
.Y(n_467)
);

OR2x2_ASAP7_75t_L g468 ( 
.A(n_444),
.B(n_406),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_436),
.B(n_422),
.Y(n_469)
);

AND2x2_ASAP7_75t_L g470 ( 
.A(n_434),
.B(n_430),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_462),
.B(n_426),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_462),
.B(n_426),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_447),
.B(n_400),
.Y(n_473)
);

OR2x2_ASAP7_75t_L g474 ( 
.A(n_444),
.B(n_406),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_432),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_430),
.B(n_424),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_451),
.B(n_422),
.Y(n_477)
);

AND2x4_ASAP7_75t_L g478 ( 
.A(n_465),
.B(n_396),
.Y(n_478)
);

OR2x2_ASAP7_75t_L g479 ( 
.A(n_450),
.B(n_457),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_439),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_439),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_447),
.B(n_406),
.Y(n_482)
);

INVxp67_ASAP7_75t_SL g483 ( 
.A(n_428),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_R g484 ( 
.A(n_433),
.B(n_363),
.Y(n_484)
);

AND2x4_ASAP7_75t_L g485 ( 
.A(n_465),
.B(n_396),
.Y(n_485)
);

AND2x4_ASAP7_75t_L g486 ( 
.A(n_465),
.B(n_396),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_431),
.B(n_424),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_432),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_439),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_437),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_454),
.B(n_407),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_437),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_441),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_431),
.B(n_424),
.Y(n_494)
);

NAND2x1p5_ASAP7_75t_L g495 ( 
.A(n_465),
.B(n_398),
.Y(n_495)
);

NAND4xp25_ASAP7_75t_L g496 ( 
.A(n_451),
.B(n_427),
.C(n_409),
.D(n_416),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_441),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_448),
.Y(n_498)
);

AND2x2_ASAP7_75t_L g499 ( 
.A(n_435),
.B(n_407),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_454),
.B(n_407),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_433),
.B(n_416),
.Y(n_501)
);

INVx1_ASAP7_75t_SL g502 ( 
.A(n_446),
.Y(n_502)
);

OR2x2_ASAP7_75t_L g503 ( 
.A(n_450),
.B(n_408),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_435),
.B(n_438),
.Y(n_504)
);

AND2x2_ASAP7_75t_L g505 ( 
.A(n_438),
.B(n_396),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_448),
.Y(n_506)
);

OR2x2_ASAP7_75t_L g507 ( 
.A(n_457),
.B(n_408),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_443),
.Y(n_508)
);

AND2x4_ASAP7_75t_L g509 ( 
.A(n_478),
.B(n_429),
.Y(n_509)
);

AND2x4_ASAP7_75t_L g510 ( 
.A(n_478),
.B(n_485),
.Y(n_510)
);

NAND4xp75_ASAP7_75t_SL g511 ( 
.A(n_477),
.B(n_440),
.C(n_377),
.D(n_342),
.Y(n_511)
);

NAND2xp67_ASAP7_75t_SL g512 ( 
.A(n_505),
.B(n_440),
.Y(n_512)
);

OR2x2_ASAP7_75t_L g513 ( 
.A(n_507),
.B(n_445),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_475),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_469),
.A2(n_442),
.B1(n_460),
.B2(n_396),
.Y(n_515)
);

AOI222xp33_ASAP7_75t_L g516 ( 
.A1(n_473),
.A2(n_463),
.B1(n_362),
.B2(n_445),
.C1(n_446),
.C2(n_396),
.Y(n_516)
);

OAI222xp33_ASAP7_75t_L g517 ( 
.A1(n_507),
.A2(n_429),
.B1(n_428),
.B2(n_463),
.C1(n_408),
.C2(n_370),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_475),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_488),
.Y(n_519)
);

OR2x2_ASAP7_75t_L g520 ( 
.A(n_503),
.B(n_443),
.Y(n_520)
);

OAI21xp5_ASAP7_75t_L g521 ( 
.A1(n_496),
.A2(n_460),
.B(n_359),
.Y(n_521)
);

NAND2x1_ASAP7_75t_L g522 ( 
.A(n_478),
.B(n_449),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_502),
.B(n_449),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_501),
.B(n_452),
.Y(n_524)
);

AND2x4_ASAP7_75t_L g525 ( 
.A(n_485),
.B(n_398),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_471),
.B(n_472),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_505),
.B(n_398),
.Y(n_527)
);

NOR2x1_ASAP7_75t_L g528 ( 
.A(n_488),
.B(n_452),
.Y(n_528)
);

OAI33xp33_ASAP7_75t_L g529 ( 
.A1(n_490),
.A2(n_461),
.A3(n_455),
.B1(n_466),
.B2(n_415),
.B3(n_411),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_490),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_483),
.B(n_455),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_492),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_492),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_L g534 ( 
.A1(n_485),
.A2(n_375),
.B1(n_281),
.B2(n_377),
.Y(n_534)
);

AND2x4_ASAP7_75t_L g535 ( 
.A(n_486),
.B(n_398),
.Y(n_535)
);

O2A1O1Ixp5_ASAP7_75t_R g536 ( 
.A1(n_491),
.A2(n_466),
.B(n_461),
.C(n_375),
.Y(n_536)
);

OR2x2_ASAP7_75t_L g537 ( 
.A(n_503),
.B(n_443),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_480),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_493),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_493),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_497),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_497),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_479),
.B(n_425),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_504),
.B(n_398),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_498),
.Y(n_545)
);

OR2x2_ASAP7_75t_L g546 ( 
.A(n_468),
.B(n_464),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_498),
.Y(n_547)
);

AOI32xp33_ASAP7_75t_L g548 ( 
.A1(n_504),
.A2(n_324),
.A3(n_383),
.B1(n_369),
.B2(n_377),
.Y(n_548)
);

OR2x2_ASAP7_75t_L g549 ( 
.A(n_468),
.B(n_453),
.Y(n_549)
);

INVx2_ASAP7_75t_SL g550 ( 
.A(n_470),
.Y(n_550)
);

XOR2x2_ASAP7_75t_L g551 ( 
.A(n_521),
.B(n_484),
.Y(n_551)
);

OAI211xp5_ASAP7_75t_SL g552 ( 
.A1(n_516),
.A2(n_479),
.B(n_500),
.C(n_506),
.Y(n_552)
);

AOI21xp33_ASAP7_75t_L g553 ( 
.A1(n_515),
.A2(n_506),
.B(n_425),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_528),
.Y(n_554)
);

XNOR2x2_ASAP7_75t_L g555 ( 
.A(n_536),
.B(n_470),
.Y(n_555)
);

OAI211xp5_ASAP7_75t_L g556 ( 
.A1(n_548),
.A2(n_474),
.B(n_482),
.C(n_355),
.Y(n_556)
);

OAI21xp33_ASAP7_75t_L g557 ( 
.A1(n_548),
.A2(n_495),
.B(n_486),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_526),
.B(n_367),
.Y(n_558)
);

OAI22xp5_ASAP7_75t_L g559 ( 
.A1(n_534),
.A2(n_370),
.B1(n_474),
.B2(n_398),
.Y(n_559)
);

AOI21xp5_ASAP7_75t_L g560 ( 
.A1(n_529),
.A2(n_517),
.B(n_524),
.Y(n_560)
);

AND2x2_ASAP7_75t_L g561 ( 
.A(n_510),
.B(n_476),
.Y(n_561)
);

AOI22xp33_ASAP7_75t_L g562 ( 
.A1(n_525),
.A2(n_486),
.B1(n_398),
.B2(n_495),
.Y(n_562)
);

XOR2x2_ASAP7_75t_L g563 ( 
.A(n_511),
.B(n_476),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_522),
.Y(n_564)
);

A2O1A1Ixp33_ASAP7_75t_L g565 ( 
.A1(n_534),
.A2(n_398),
.B(n_324),
.C(n_494),
.Y(n_565)
);

XNOR2x1_ASAP7_75t_L g566 ( 
.A(n_510),
.B(n_487),
.Y(n_566)
);

OAI22xp33_ASAP7_75t_L g567 ( 
.A1(n_550),
.A2(n_495),
.B1(n_369),
.B2(n_383),
.Y(n_567)
);

O2A1O1Ixp33_ASAP7_75t_L g568 ( 
.A1(n_531),
.A2(n_355),
.B(n_489),
.C(n_481),
.Y(n_568)
);

AOI21xp33_ASAP7_75t_L g569 ( 
.A1(n_523),
.A2(n_508),
.B(n_480),
.Y(n_569)
);

OR2x2_ASAP7_75t_L g570 ( 
.A(n_513),
.B(n_487),
.Y(n_570)
);

AOI22xp5_ASAP7_75t_SL g571 ( 
.A1(n_525),
.A2(n_494),
.B1(n_467),
.B2(n_499),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_528),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_514),
.Y(n_573)
);

INVx1_ASAP7_75t_SL g574 ( 
.A(n_509),
.Y(n_574)
);

INVx3_ASAP7_75t_L g575 ( 
.A(n_509),
.Y(n_575)
);

INVxp67_ASAP7_75t_L g576 ( 
.A(n_543),
.Y(n_576)
);

AOI21xp33_ASAP7_75t_SL g577 ( 
.A1(n_535),
.A2(n_499),
.B(n_467),
.Y(n_577)
);

AOI21xp33_ASAP7_75t_L g578 ( 
.A1(n_518),
.A2(n_532),
.B(n_547),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_519),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_530),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_533),
.Y(n_581)
);

AOI21xp33_ASAP7_75t_L g582 ( 
.A1(n_539),
.A2(n_412),
.B(n_489),
.Y(n_582)
);

OAI22xp33_ASAP7_75t_L g583 ( 
.A1(n_546),
.A2(n_369),
.B1(n_383),
.B2(n_379),
.Y(n_583)
);

NOR3xp33_ASAP7_75t_L g584 ( 
.A(n_540),
.B(n_414),
.C(n_397),
.Y(n_584)
);

INVx1_ASAP7_75t_SL g585 ( 
.A(n_551),
.Y(n_585)
);

AOI22xp5_ASAP7_75t_L g586 ( 
.A1(n_557),
.A2(n_535),
.B1(n_544),
.B2(n_527),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_560),
.B(n_541),
.Y(n_587)
);

AOI21xp5_ASAP7_75t_L g588 ( 
.A1(n_565),
.A2(n_553),
.B(n_552),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_573),
.Y(n_589)
);

HB1xp67_ASAP7_75t_L g590 ( 
.A(n_554),
.Y(n_590)
);

OAI221xp5_ASAP7_75t_L g591 ( 
.A1(n_562),
.A2(n_545),
.B1(n_542),
.B2(n_537),
.C(n_520),
.Y(n_591)
);

O2A1O1Ixp33_ASAP7_75t_L g592 ( 
.A1(n_553),
.A2(n_512),
.B(n_538),
.C(n_549),
.Y(n_592)
);

AOI22xp5_ASAP7_75t_L g593 ( 
.A1(n_563),
.A2(n_412),
.B1(n_369),
.B2(n_383),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_576),
.B(n_508),
.Y(n_594)
);

AOI211xp5_ASAP7_75t_SL g595 ( 
.A1(n_559),
.A2(n_412),
.B(n_414),
.C(n_397),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_579),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_580),
.Y(n_597)
);

HB1xp67_ASAP7_75t_L g598 ( 
.A(n_572),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_575),
.Y(n_599)
);

BUFx3_ASAP7_75t_L g600 ( 
.A(n_575),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_581),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_568),
.B(n_481),
.Y(n_602)
);

OR2x2_ASAP7_75t_L g603 ( 
.A(n_570),
.B(n_464),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_561),
.B(n_556),
.Y(n_604)
);

INVx2_ASAP7_75t_SL g605 ( 
.A(n_566),
.Y(n_605)
);

NAND2xp33_ASAP7_75t_SL g606 ( 
.A(n_564),
.B(n_339),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_574),
.Y(n_607)
);

O2A1O1Ixp33_ASAP7_75t_L g608 ( 
.A1(n_559),
.A2(n_412),
.B(n_397),
.C(n_414),
.Y(n_608)
);

OR2x2_ASAP7_75t_L g609 ( 
.A(n_555),
.B(n_464),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_574),
.B(n_415),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_578),
.Y(n_611)
);

OAI22xp33_ASAP7_75t_L g612 ( 
.A1(n_567),
.A2(n_379),
.B1(n_397),
.B2(n_414),
.Y(n_612)
);

INVx3_ASAP7_75t_L g613 ( 
.A(n_571),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_587),
.B(n_605),
.Y(n_614)
);

BUFx2_ASAP7_75t_L g615 ( 
.A(n_600),
.Y(n_615)
);

NAND3xp33_ASAP7_75t_SL g616 ( 
.A(n_588),
.B(n_577),
.C(n_558),
.Y(n_616)
);

NAND3xp33_ASAP7_75t_L g617 ( 
.A(n_611),
.B(n_584),
.C(n_582),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_604),
.B(n_569),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_589),
.Y(n_619)
);

OAI21xp33_ASAP7_75t_L g620 ( 
.A1(n_613),
.A2(n_569),
.B(n_583),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_607),
.B(n_412),
.Y(n_621)
);

HB1xp67_ASAP7_75t_L g622 ( 
.A(n_590),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_602),
.B(n_459),
.Y(n_623)
);

AOI211xp5_ASAP7_75t_L g624 ( 
.A1(n_585),
.A2(n_339),
.B(n_306),
.C(n_260),
.Y(n_624)
);

AOI221xp5_ASAP7_75t_L g625 ( 
.A1(n_592),
.A2(n_390),
.B1(n_392),
.B2(n_456),
.C(n_453),
.Y(n_625)
);

HB1xp67_ASAP7_75t_L g626 ( 
.A(n_590),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_596),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_597),
.Y(n_628)
);

NAND4xp25_ASAP7_75t_L g629 ( 
.A(n_613),
.B(n_414),
.C(n_397),
.D(n_306),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_601),
.Y(n_630)
);

AOI211xp5_ASAP7_75t_L g631 ( 
.A1(n_612),
.A2(n_339),
.B(n_306),
.C(n_260),
.Y(n_631)
);

CKINVDCx20_ASAP7_75t_R g632 ( 
.A(n_593),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_610),
.Y(n_633)
);

OAI21xp5_ASAP7_75t_L g634 ( 
.A1(n_614),
.A2(n_609),
.B(n_595),
.Y(n_634)
);

AOI22x1_ASAP7_75t_SL g635 ( 
.A1(n_632),
.A2(n_599),
.B1(n_600),
.B2(n_606),
.Y(n_635)
);

BUFx2_ASAP7_75t_L g636 ( 
.A(n_615),
.Y(n_636)
);

NOR4xp25_ASAP7_75t_L g637 ( 
.A(n_616),
.B(n_620),
.C(n_618),
.D(n_625),
.Y(n_637)
);

AOI221xp5_ASAP7_75t_L g638 ( 
.A1(n_617),
.A2(n_591),
.B1(n_608),
.B2(n_612),
.C(n_598),
.Y(n_638)
);

OR2x2_ASAP7_75t_L g639 ( 
.A(n_633),
.B(n_594),
.Y(n_639)
);

AOI22x1_ASAP7_75t_SL g640 ( 
.A1(n_629),
.A2(n_606),
.B1(n_586),
.B2(n_598),
.Y(n_640)
);

XNOR2x1_ASAP7_75t_SL g641 ( 
.A(n_619),
.B(n_284),
.Y(n_641)
);

AOI22xp5_ASAP7_75t_L g642 ( 
.A1(n_624),
.A2(n_603),
.B1(n_306),
.B2(n_339),
.Y(n_642)
);

INVx1_ASAP7_75t_SL g643 ( 
.A(n_622),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_622),
.Y(n_644)
);

NOR2x1p5_ASAP7_75t_SL g645 ( 
.A(n_627),
.B(n_630),
.Y(n_645)
);

NOR3xp33_ASAP7_75t_L g646 ( 
.A(n_628),
.B(n_345),
.C(n_344),
.Y(n_646)
);

AOI21xp5_ASAP7_75t_SL g647 ( 
.A1(n_626),
.A2(n_339),
.B(n_368),
.Y(n_647)
);

AOI22xp5_ASAP7_75t_L g648 ( 
.A1(n_631),
.A2(n_339),
.B1(n_390),
.B2(n_392),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_623),
.B(n_332),
.Y(n_649)
);

OAI21xp5_ASAP7_75t_L g650 ( 
.A1(n_626),
.A2(n_250),
.B(n_349),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_621),
.B(n_459),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_622),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_614),
.B(n_281),
.Y(n_653)
);

AOI21xp33_ASAP7_75t_SL g654 ( 
.A1(n_614),
.A2(n_349),
.B(n_284),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_614),
.B(n_281),
.Y(n_655)
);

OR2x2_ASAP7_75t_L g656 ( 
.A(n_636),
.B(n_459),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_637),
.B(n_281),
.Y(n_657)
);

AOI311xp33_ASAP7_75t_L g658 ( 
.A1(n_634),
.A2(n_347),
.A3(n_351),
.B(n_380),
.C(n_387),
.Y(n_658)
);

OA211x2_ASAP7_75t_L g659 ( 
.A1(n_638),
.A2(n_318),
.B(n_368),
.C(n_256),
.Y(n_659)
);

AOI21xp5_ASAP7_75t_L g660 ( 
.A1(n_634),
.A2(n_458),
.B(n_456),
.Y(n_660)
);

NOR4xp25_ASAP7_75t_L g661 ( 
.A(n_643),
.B(n_351),
.C(n_308),
.D(n_309),
.Y(n_661)
);

AOI21xp33_ASAP7_75t_L g662 ( 
.A1(n_653),
.A2(n_256),
.B(n_260),
.Y(n_662)
);

OAI211xp5_ASAP7_75t_L g663 ( 
.A1(n_643),
.A2(n_289),
.B(n_267),
.C(n_270),
.Y(n_663)
);

AOI221xp5_ASAP7_75t_L g664 ( 
.A1(n_652),
.A2(n_458),
.B1(n_456),
.B2(n_453),
.C(n_380),
.Y(n_664)
);

OAI21xp5_ASAP7_75t_SL g665 ( 
.A1(n_648),
.A2(n_458),
.B(n_360),
.Y(n_665)
);

OAI221xp5_ASAP7_75t_L g666 ( 
.A1(n_650),
.A2(n_304),
.B1(n_270),
.B2(n_289),
.C(n_360),
.Y(n_666)
);

NOR2x1_ASAP7_75t_L g667 ( 
.A(n_644),
.B(n_270),
.Y(n_667)
);

NAND3xp33_ASAP7_75t_L g668 ( 
.A(n_635),
.B(n_289),
.C(n_387),
.Y(n_668)
);

NAND4xp25_ASAP7_75t_L g669 ( 
.A(n_655),
.B(n_386),
.C(n_360),
.D(n_309),
.Y(n_669)
);

OAI21xp33_ASAP7_75t_L g670 ( 
.A1(n_645),
.A2(n_386),
.B(n_423),
.Y(n_670)
);

OAI211xp5_ASAP7_75t_SL g671 ( 
.A1(n_650),
.A2(n_310),
.B(n_319),
.C(n_308),
.Y(n_671)
);

NAND4xp25_ASAP7_75t_SL g672 ( 
.A(n_642),
.B(n_413),
.C(n_402),
.D(n_399),
.Y(n_672)
);

INVx1_ASAP7_75t_SL g673 ( 
.A(n_640),
.Y(n_673)
);

AOI222xp33_ASAP7_75t_L g674 ( 
.A1(n_649),
.A2(n_322),
.B1(n_402),
.B2(n_399),
.C1(n_391),
.C2(n_413),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_639),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_675),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_656),
.Y(n_677)
);

NOR2x1_ASAP7_75t_L g678 ( 
.A(n_668),
.B(n_673),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_667),
.Y(n_679)
);

NOR2xp67_ASAP7_75t_L g680 ( 
.A(n_663),
.B(n_654),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_669),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_670),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_666),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_671),
.Y(n_684)
);

AOI22xp5_ASAP7_75t_L g685 ( 
.A1(n_657),
.A2(n_646),
.B1(n_641),
.B2(n_651),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_659),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_658),
.B(n_647),
.Y(n_687)
);

NAND3xp33_ASAP7_75t_L g688 ( 
.A(n_678),
.B(n_662),
.C(n_674),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_682),
.B(n_660),
.Y(n_689)
);

AOI221xp5_ASAP7_75t_SL g690 ( 
.A1(n_686),
.A2(n_664),
.B1(n_672),
.B2(n_661),
.C(n_665),
.Y(n_690)
);

AOI222xp33_ASAP7_75t_L g691 ( 
.A1(n_676),
.A2(n_661),
.B1(n_381),
.B2(n_310),
.C1(n_319),
.C2(n_413),
.Y(n_691)
);

NAND5xp2_ASAP7_75t_L g692 ( 
.A(n_685),
.B(n_342),
.C(n_291),
.D(n_318),
.E(n_285),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_684),
.B(n_683),
.Y(n_693)
);

A2O1A1Ixp33_ASAP7_75t_L g694 ( 
.A1(n_680),
.A2(n_381),
.B(n_399),
.C(n_391),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_677),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_R g696 ( 
.A(n_695),
.B(n_679),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_689),
.Y(n_697)
);

HB1xp67_ASAP7_75t_L g698 ( 
.A(n_693),
.Y(n_698)
);

OR2x2_ASAP7_75t_L g699 ( 
.A(n_688),
.B(n_681),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_690),
.B(n_686),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_692),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_694),
.Y(n_702)
);

INVx1_ASAP7_75t_SL g703 ( 
.A(n_691),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_693),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_704),
.Y(n_705)
);

OAI22xp5_ASAP7_75t_L g706 ( 
.A1(n_700),
.A2(n_685),
.B1(n_687),
.B2(n_291),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_698),
.Y(n_707)
);

AOI22xp5_ASAP7_75t_L g708 ( 
.A1(n_701),
.A2(n_291),
.B1(n_263),
.B2(n_273),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_707),
.Y(n_709)
);

AO22x2_ASAP7_75t_L g710 ( 
.A1(n_706),
.A2(n_699),
.B1(n_697),
.B2(n_703),
.Y(n_710)
);

AOI22xp33_ASAP7_75t_SL g711 ( 
.A1(n_705),
.A2(n_698),
.B1(n_696),
.B2(n_702),
.Y(n_711)
);

OAI22xp5_ASAP7_75t_L g712 ( 
.A1(n_711),
.A2(n_708),
.B1(n_291),
.B2(n_402),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_709),
.B(n_291),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_713),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_714),
.B(n_710),
.Y(n_715)
);

OAI22xp5_ASAP7_75t_SL g716 ( 
.A1(n_715),
.A2(n_712),
.B1(n_263),
.B2(n_273),
.Y(n_716)
);

OR2x6_ASAP7_75t_L g717 ( 
.A(n_716),
.B(n_263),
.Y(n_717)
);

OAI22xp5_ASAP7_75t_L g718 ( 
.A1(n_717),
.A2(n_273),
.B1(n_348),
.B2(n_311),
.Y(n_718)
);


endmodule