module fake_jpeg_30239_n_39 (n_3, n_2, n_1, n_0, n_4, n_5, n_39);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_39;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx5_ASAP7_75t_L g6 ( 
.A(n_1),
.Y(n_6)
);

INVx2_ASAP7_75t_L g7 ( 
.A(n_3),
.Y(n_7)
);

NOR2xp33_ASAP7_75t_L g8 ( 
.A(n_2),
.B(n_3),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_4),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

INVx11_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

BUFx12_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

MAJIxp5_ASAP7_75t_L g13 ( 
.A(n_7),
.B(n_0),
.C(n_1),
.Y(n_13)
);

OAI21xp5_ASAP7_75t_L g24 ( 
.A1(n_13),
.A2(n_11),
.B(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_8),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g20 ( 
.A(n_14),
.B(n_19),
.Y(n_20)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_15),
.Y(n_22)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

OR2x2_ASAP7_75t_L g23 ( 
.A(n_16),
.B(n_17),
.Y(n_23)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_18),
.Y(n_21)
);

OR2x2_ASAP7_75t_L g19 ( 
.A(n_8),
.B(n_1),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_L g26 ( 
.A1(n_24),
.A2(n_13),
.B(n_19),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_22),
.A2(n_10),
.B1(n_18),
.B2(n_9),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_27),
.Y(n_30)
);

AOI221xp5_ASAP7_75t_L g32 ( 
.A1(n_26),
.A2(n_21),
.B1(n_2),
.B2(n_5),
.C(n_4),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_24),
.B(n_10),
.C(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

OA21x2_ASAP7_75t_SL g29 ( 
.A1(n_27),
.A2(n_20),
.B(n_23),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_29),
.B(n_32),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_30),
.Y(n_33)
);

AO21x1_ASAP7_75t_L g37 ( 
.A1(n_33),
.A2(n_35),
.B(n_31),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_2),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g36 ( 
.A1(n_35),
.A2(n_34),
.B(n_29),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_36),
.A2(n_37),
.B1(n_31),
.B2(n_12),
.Y(n_38)
);

O2A1O1Ixp33_ASAP7_75t_SL g39 ( 
.A1(n_38),
.A2(n_12),
.B(n_37),
.C(n_30),
.Y(n_39)
);


endmodule