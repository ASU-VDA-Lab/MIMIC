module fake_jpeg_10908_n_204 (n_13, n_21, n_57, n_53, n_33, n_54, n_1, n_45, n_10, n_23, n_27, n_55, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_56, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_204);

input n_13;
input n_21;
input n_57;
input n_53;
input n_33;
input n_54;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_55;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_56;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_204;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_54),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_33),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_12),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_27),
.Y(n_69)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

INVx6_ASAP7_75t_SL g71 ( 
.A(n_4),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_55),
.Y(n_72)
);

INVx11_ASAP7_75t_SL g73 ( 
.A(n_50),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_53),
.Y(n_74)
);

INVx11_ASAP7_75t_SL g75 ( 
.A(n_5),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_18),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_12),
.B(n_11),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_42),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_38),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_41),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_13),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_22),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_14),
.Y(n_83)
);

BUFx16f_ASAP7_75t_L g84 ( 
.A(n_17),
.Y(n_84)
);

INVx2_ASAP7_75t_SL g85 ( 
.A(n_21),
.Y(n_85)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_28),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_15),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_88),
.Y(n_102)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_84),
.Y(n_89)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_58),
.Y(n_90)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_90),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_91),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_68),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_92),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_77),
.B(n_0),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_93),
.B(n_85),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_0),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_94),
.B(n_69),
.Y(n_98)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_71),
.Y(n_95)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_95),
.Y(n_113)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_86),
.Y(n_96)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_96),
.Y(n_111)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_97),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_98),
.B(n_99),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_90),
.B(n_67),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_95),
.B(n_67),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_101),
.B(n_84),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_103),
.B(n_104),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_82),
.Y(n_104)
);

BUFx10_ASAP7_75t_L g106 ( 
.A(n_96),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_106),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_88),
.A2(n_59),
.B1(n_80),
.B2(n_85),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_110),
.A2(n_87),
.B1(n_76),
.B2(n_75),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_91),
.B(n_74),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_112),
.B(n_65),
.Y(n_118)
);

AND2x2_ASAP7_75t_SL g114 ( 
.A(n_100),
.B(n_63),
.Y(n_114)
);

INVx1_ASAP7_75t_SL g148 ( 
.A(n_114),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_106),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_115),
.B(n_57),
.Y(n_151)
);

A2O1A1Ixp33_ASAP7_75t_L g116 ( 
.A1(n_99),
.A2(n_62),
.B(n_64),
.C(n_81),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_116),
.B(n_120),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_118),
.B(n_127),
.Y(n_144)
);

OAI21xp33_ASAP7_75t_L g119 ( 
.A1(n_101),
.A2(n_66),
.B(n_79),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_119),
.A2(n_126),
.B(n_9),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_108),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_113),
.Y(n_121)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_121),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_102),
.A2(n_92),
.B1(n_75),
.B2(n_68),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_122),
.A2(n_73),
.B1(n_83),
.B2(n_26),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_106),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_123),
.B(n_128),
.Y(n_145)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_109),
.Y(n_125)
);

HB1xp67_ASAP7_75t_L g137 ( 
.A(n_125),
.Y(n_137)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_105),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_105),
.B(n_72),
.Y(n_128)
);

AND2x2_ASAP7_75t_SL g129 ( 
.A(n_111),
.B(n_70),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_129),
.B(n_73),
.Y(n_139)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_102),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_131),
.B(n_132),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_107),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_110),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_133),
.B(n_134),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_107),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_135),
.B(n_7),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_114),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_136),
.B(n_156),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_133),
.A2(n_87),
.B1(n_76),
.B2(n_78),
.Y(n_138)
);

A2O1A1Ixp33_ASAP7_75t_SL g173 ( 
.A1(n_138),
.A2(n_56),
.B(n_19),
.C(n_20),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_139),
.B(n_154),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_141),
.A2(n_143),
.B1(n_146),
.B2(n_149),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_126),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_142),
.A2(n_134),
.B1(n_130),
.B2(n_10),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_124),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_117),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_129),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_151),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_152),
.B(n_155),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_119),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_116),
.B(n_8),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_130),
.B(n_9),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_157),
.A2(n_16),
.B(n_23),
.Y(n_174)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_147),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_158),
.B(n_162),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_160),
.A2(n_165),
.B1(n_148),
.B2(n_159),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_140),
.B(n_10),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_142),
.A2(n_148),
.B1(n_150),
.B2(n_138),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_145),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_166),
.B(n_168),
.Y(n_175)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_153),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_137),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_169),
.B(n_170),
.Y(n_176)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_144),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_143),
.B(n_11),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_171),
.B(n_172),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_149),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_173),
.Y(n_182)
);

XNOR2x1_ASAP7_75t_L g178 ( 
.A(n_174),
.B(n_139),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_177),
.A2(n_161),
.B1(n_173),
.B2(n_47),
.Y(n_188)
);

OR2x2_ASAP7_75t_L g187 ( 
.A(n_178),
.B(n_164),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_165),
.A2(n_25),
.B1(n_30),
.B2(n_31),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_179),
.A2(n_183),
.B1(n_161),
.B2(n_173),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_163),
.Y(n_180)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_180),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_164),
.A2(n_32),
.B1(n_37),
.B2(n_39),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_167),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_184),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_SL g195 ( 
.A(n_187),
.B(n_192),
.C(n_181),
.Y(n_195)
);

CKINVDCx14_ASAP7_75t_R g194 ( 
.A(n_188),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_176),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_190),
.B(n_191),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_182),
.A2(n_173),
.B1(n_46),
.B2(n_48),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_195),
.A2(n_189),
.B(n_185),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_196),
.B(n_186),
.Y(n_197)
);

OAI21xp33_ASAP7_75t_L g198 ( 
.A1(n_197),
.A2(n_175),
.B(n_193),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_198),
.B(n_192),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_199),
.B(n_194),
.Y(n_200)
);

MAJx2_ASAP7_75t_L g201 ( 
.A(n_200),
.B(n_178),
.C(n_182),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_201),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_202),
.A2(n_43),
.B(n_49),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_203),
.B(n_51),
.Y(n_204)
);


endmodule