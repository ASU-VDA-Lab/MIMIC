module fake_jpeg_30368_n_126 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_126);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_126;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_15),
.B(n_13),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_12),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_9),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_3),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_2),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_29),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_31),
.Y(n_52)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_53),
.Y(n_55)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

OA22x2_ASAP7_75t_L g56 ( 
.A1(n_46),
.A2(n_19),
.B1(n_39),
.B2(n_38),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_60),
.Y(n_64)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_54),
.Y(n_57)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g59 ( 
.A1(n_41),
.A2(n_0),
.B(n_1),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_59),
.B(n_2),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_48),
.B(n_0),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_1),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_4),
.Y(n_72)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_63),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_70),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_56),
.B(n_51),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_3),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_10),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_4),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_56),
.B(n_44),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_5),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_61),
.A2(n_43),
.B1(n_50),
.B2(n_47),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_74),
.A2(n_45),
.B1(n_52),
.B2(n_42),
.Y(n_80)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_76),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_63),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_84),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_71),
.A2(n_50),
.B(n_47),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_78),
.Y(n_104)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_79),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_80),
.A2(n_89),
.B1(n_18),
.B2(n_21),
.Y(n_105)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_91),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_75),
.B(n_45),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_85),
.B(n_87),
.Y(n_95)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_86),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_74),
.A2(n_5),
.B(n_6),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_69),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_90),
.B(n_17),
.Y(n_103)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_65),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_92),
.B(n_11),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_69),
.C(n_16),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_94),
.B(n_106),
.C(n_107),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_88),
.B(n_40),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_98),
.B(n_100),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_84),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_102),
.B(n_103),
.Y(n_113)
);

AO22x1_ASAP7_75t_SL g111 ( 
.A1(n_105),
.A2(n_24),
.B1(n_26),
.B2(n_30),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_88),
.B(n_22),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_37),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_82),
.B(n_23),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_108),
.B(n_36),
.C(n_94),
.Y(n_116)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_97),
.Y(n_110)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_110),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_111),
.B(n_112),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_104),
.A2(n_32),
.B(n_34),
.Y(n_112)
);

XNOR2x1_ASAP7_75t_SL g115 ( 
.A(n_93),
.B(n_35),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_115),
.B(n_116),
.Y(n_119)
);

A2O1A1O1Ixp25_ASAP7_75t_L g120 ( 
.A1(n_118),
.A2(n_95),
.B(n_113),
.C(n_104),
.D(n_99),
.Y(n_120)
);

FAx1_ASAP7_75t_SL g122 ( 
.A(n_120),
.B(n_121),
.CI(n_96),
.CON(n_122),
.SN(n_122)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_119),
.B(n_114),
.C(n_109),
.Y(n_121)
);

INVx11_ASAP7_75t_L g123 ( 
.A(n_122),
.Y(n_123)
);

A2O1A1Ixp33_ASAP7_75t_SL g124 ( 
.A1(n_123),
.A2(n_122),
.B(n_117),
.C(n_96),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_123),
.C(n_110),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_125),
.B(n_101),
.Y(n_126)
);


endmodule