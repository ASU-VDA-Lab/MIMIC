module fake_netlist_5_1396_n_121 (n_16, n_0, n_12, n_9, n_25, n_18, n_27, n_22, n_1, n_8, n_10, n_24, n_21, n_4, n_11, n_17, n_19, n_7, n_15, n_26, n_20, n_5, n_14, n_2, n_23, n_13, n_3, n_6, n_121);

input n_16;
input n_0;
input n_12;
input n_9;
input n_25;
input n_18;
input n_27;
input n_22;
input n_1;
input n_8;
input n_10;
input n_24;
input n_21;
input n_4;
input n_11;
input n_17;
input n_19;
input n_7;
input n_15;
input n_26;
input n_20;
input n_5;
input n_14;
input n_2;
input n_23;
input n_13;
input n_3;
input n_6;

output n_121;

wire n_91;
wire n_82;
wire n_86;
wire n_83;
wire n_61;
wire n_90;
wire n_75;
wire n_101;
wire n_65;
wire n_78;
wire n_74;
wire n_114;
wire n_57;
wire n_96;
wire n_37;
wire n_111;
wire n_108;
wire n_31;
wire n_66;
wire n_98;
wire n_60;
wire n_43;
wire n_107;
wire n_58;
wire n_69;
wire n_116;
wire n_42;
wire n_45;
wire n_117;
wire n_46;
wire n_94;
wire n_113;
wire n_38;
wire n_105;
wire n_80;
wire n_35;
wire n_73;
wire n_92;
wire n_120;
wire n_30;
wire n_33;
wire n_84;
wire n_29;
wire n_79;
wire n_47;
wire n_53;
wire n_44;
wire n_40;
wire n_34;
wire n_100;
wire n_62;
wire n_71;
wire n_109;
wire n_112;
wire n_85;
wire n_95;
wire n_119;
wire n_59;
wire n_55;
wire n_99;
wire n_49;
wire n_39;
wire n_54;
wire n_67;
wire n_36;
wire n_76;
wire n_87;
wire n_64;
wire n_77;
wire n_102;
wire n_106;
wire n_81;
wire n_118;
wire n_28;
wire n_89;
wire n_70;
wire n_115;
wire n_68;
wire n_93;
wire n_72;
wire n_32;
wire n_41;
wire n_104;
wire n_103;
wire n_56;
wire n_51;
wire n_63;
wire n_97;
wire n_48;
wire n_50;
wire n_52;
wire n_88;
wire n_110;

HB1xp67_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_23),
.Y(n_29)
);

HB1xp67_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

CKINVDCx5p33_ASAP7_75t_R g33 ( 
.A(n_21),
.Y(n_33)
);

CKINVDCx5p33_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_11),
.Y(n_36)
);

HB1xp67_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

INVxp67_ASAP7_75t_SL g40 ( 
.A(n_8),
.Y(n_40)
);

CKINVDCx5p33_ASAP7_75t_R g41 ( 
.A(n_26),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_1),
.B(n_12),
.Y(n_42)
);

NOR2xp67_ASAP7_75t_L g43 ( 
.A(n_16),
.B(n_6),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

INVxp33_ASAP7_75t_SL g45 ( 
.A(n_2),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

CKINVDCx5p33_ASAP7_75t_R g48 ( 
.A(n_6),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

CKINVDCx5p33_ASAP7_75t_R g51 ( 
.A(n_3),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_28),
.B(n_0),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_50),
.B(n_3),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_50),
.Y(n_60)
);

AND2x6_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_15),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_49),
.B(n_4),
.Y(n_64)
);

AND2x4_ASAP7_75t_L g65 ( 
.A(n_38),
.B(n_46),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_60),
.B(n_34),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_53),
.B(n_43),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_53),
.B(n_43),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_65),
.B(n_30),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_57),
.B(n_45),
.Y(n_70)
);

NAND2xp33_ASAP7_75t_SL g71 ( 
.A(n_64),
.B(n_37),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_64),
.B(n_51),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_65),
.B(n_54),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_55),
.B(n_42),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_58),
.B(n_48),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_59),
.B(n_41),
.Y(n_76)
);

NAND2xp33_ASAP7_75t_SL g77 ( 
.A(n_63),
.B(n_36),
.Y(n_77)
);

OAI21x1_ASAP7_75t_L g78 ( 
.A1(n_73),
.A2(n_67),
.B(n_68),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_72),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_L g80 ( 
.A1(n_72),
.A2(n_40),
.B1(n_39),
.B2(n_31),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_77),
.B(n_29),
.Y(n_81)
);

OA21x2_ASAP7_75t_L g82 ( 
.A1(n_74),
.A2(n_63),
.B(n_56),
.Y(n_82)
);

NAND2x1p5_ASAP7_75t_L g83 ( 
.A(n_70),
.B(n_44),
.Y(n_83)
);

OAI21x1_ASAP7_75t_L g84 ( 
.A1(n_76),
.A2(n_56),
.B(n_52),
.Y(n_84)
);

OAI21x1_ASAP7_75t_L g85 ( 
.A1(n_69),
.A2(n_52),
.B(n_46),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

OAI21x1_ASAP7_75t_L g87 ( 
.A1(n_71),
.A2(n_44),
.B(n_62),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_67),
.A2(n_61),
.B1(n_31),
.B2(n_40),
.Y(n_88)
);

NAND2xp33_ASAP7_75t_SL g89 ( 
.A(n_79),
.B(n_33),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_86),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_82),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

NAND2xp33_ASAP7_75t_SL g93 ( 
.A(n_81),
.B(n_61),
.Y(n_93)
);

AND2x4_ASAP7_75t_L g94 ( 
.A(n_87),
.B(n_61),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_86),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_90),
.B(n_79),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_92),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_95),
.B(n_78),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_94),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_96),
.B(n_78),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_98),
.B(n_78),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_97),
.A2(n_89),
.B1(n_93),
.B2(n_80),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_97),
.A2(n_89),
.B1(n_88),
.B2(n_83),
.Y(n_103)
);

OAI222xp33_ASAP7_75t_L g104 ( 
.A1(n_102),
.A2(n_83),
.B1(n_39),
.B2(n_98),
.C1(n_97),
.C2(n_94),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_103),
.A2(n_99),
.B1(n_91),
.B2(n_94),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_100),
.A2(n_99),
.B1(n_87),
.B2(n_61),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_101),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_107),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_105),
.Y(n_109)
);

AOI221xp5_ASAP7_75t_L g110 ( 
.A1(n_109),
.A2(n_104),
.B1(n_106),
.B2(n_99),
.C(n_9),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_108),
.A2(n_61),
.B1(n_87),
.B2(n_82),
.Y(n_111)
);

AND2x4_ASAP7_75t_L g112 ( 
.A(n_108),
.B(n_85),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_R g113 ( 
.A(n_112),
.B(n_24),
.Y(n_113)
);

NAND2xp33_ASAP7_75t_SL g114 ( 
.A(n_110),
.B(n_4),
.Y(n_114)
);

INVx2_ASAP7_75t_SL g115 ( 
.A(n_113),
.Y(n_115)
);

NAND2x1p5_ASAP7_75t_L g116 ( 
.A(n_114),
.B(n_111),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_114),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_116),
.A2(n_82),
.B1(n_85),
.B2(n_84),
.Y(n_118)
);

AOI31xp33_ASAP7_75t_L g119 ( 
.A1(n_115),
.A2(n_5),
.A3(n_7),
.B(n_9),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_118),
.A2(n_117),
.B1(n_82),
.B2(n_84),
.Y(n_120)
);

AOI221xp5_ASAP7_75t_L g121 ( 
.A1(n_120),
.A2(n_119),
.B1(n_117),
.B2(n_7),
.C(n_22),
.Y(n_121)
);


endmodule